

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9706, n9707, n9708, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871;

  NOR2_X1 U11150 ( .A1(n17565), .A2(n16455), .ZN(n17881) );
  CLKBUF_X2 U11151 ( .A(n13703), .Z(n9716) );
  CLKBUF_X1 U11152 ( .A(n13683), .Z(n9717) );
  INV_X1 U11153 ( .A(n9756), .ZN(n9730) );
  INV_X1 U11154 ( .A(n17180), .ZN(n9728) );
  BUF_X1 U11155 ( .A(n10769), .Z(n12964) );
  CLKBUF_X1 U11156 ( .A(n13274), .Z(n15508) );
  INV_X1 U11157 ( .A(n17128), .ZN(n17085) );
  CLKBUF_X3 U11158 ( .A(n13278), .Z(n9725) );
  CLKBUF_X1 U11160 ( .A(n11239), .Z(n12963) );
  AND2_X1 U11161 ( .A1(n13118), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10728) );
  AND2_X1 U11162 ( .A1(n13131), .A2(n10470), .ZN(n10723) );
  AND2_X1 U11163 ( .A1(n13082), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12899) );
  AND2_X1 U11164 ( .A1(n10663), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10775) );
  AND2_X1 U11165 ( .A1(n9737), .A2(n10470), .ZN(n12971) );
  INV_X2 U11166 ( .A(n19283), .ZN(n11191) );
  NAND2_X1 U11167 ( .A1(n16351), .A2(n19283), .ZN(n11001) );
  CLKBUF_X2 U11168 ( .A(n11582), .Z(n12103) );
  INV_X1 U11169 ( .A(n19968), .ZN(n16351) );
  CLKBUF_X2 U11170 ( .A(n11542), .Z(n9713) );
  INV_X2 U11171 ( .A(n11196), .ZN(n19283) );
  INV_X1 U11172 ( .A(n11078), .ZN(n10544) );
  INV_X1 U11173 ( .A(n13854), .ZN(n20196) );
  NOR2_X1 U11174 ( .A1(n12212), .A2(n12278), .ZN(n13382) );
  CLKBUF_X3 U11175 ( .A(n10509), .Z(n13082) );
  INV_X2 U11176 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10470) );
  AND2_X1 U11177 ( .A1(n13654), .A2(n11390), .ZN(n11567) );
  AND2_X1 U11178 ( .A1(n11387), .A2(n13656), .ZN(n11582) );
  AND2_X1 U11179 ( .A1(n11391), .A2(n13647), .ZN(n11646) );
  AND2_X2 U11180 ( .A1(n11387), .A2(n11388), .ZN(n11542) );
  AND2_X1 U11181 ( .A1(n10000), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11391) );
  INV_X2 U11182 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16318) );
  CLKBUF_X1 U11183 ( .A(n18701), .Z(n9706) );
  NOR2_X1 U11184 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18803), .ZN(n18701) );
  CLKBUF_X1 U11185 ( .A(n19046), .Z(n9707) );
  NOR2_X1 U11186 ( .A1(n19081), .A2(n19533), .ZN(n19046) );
  AOI22_X1 U11187 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n19626), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10642) );
  AOI21_X1 U11188 ( .B1(n10012), .B2(n9913), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9911) );
  OR2_X1 U11189 ( .A1(n10830), .A2(n9881), .ZN(n9878) );
  INV_X1 U11190 ( .A(n11040), .ZN(n10568) );
  AND2_X1 U11191 ( .A1(n13656), .A2(n13647), .ZN(n11681) );
  AND2_X1 U11192 ( .A1(n11388), .A2(n13673), .ZN(n11584) );
  NAND3_X2 U11193 ( .A1(n15369), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13129) );
  XNOR2_X1 U11194 ( .A(n9863), .B(n13179), .ZN(n14312) );
  AND3_X1 U11195 ( .A1(n10586), .A2(n10585), .A3(n10584), .ZN(n9763) );
  INV_X1 U11196 ( .A(n10107), .ZN(n15511) );
  OR2_X1 U11197 ( .A1(n11557), .A2(n11556), .ZN(n12600) );
  OAI22_X2 U11198 ( .A1(n14312), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19969), 
        .B2(n13180), .ZN(n13703) );
  NAND2_X1 U11200 ( .A1(n15278), .A2(n15262), .ZN(n15261) );
  OR2_X1 U11201 ( .A1(n10640), .A2(n10633), .ZN(n19498) );
  NAND2_X1 U11202 ( .A1(n11629), .A2(n12209), .ZN(n11621) );
  AND2_X1 U11203 ( .A1(n12674), .A2(n12673), .ZN(n9757) );
  AND2_X1 U11205 ( .A1(n13600), .A2(n12853), .ZN(n13741) );
  NAND2_X2 U11206 ( .A1(n13741), .A2(n12855), .ZN(n13738) );
  OR2_X1 U11207 ( .A1(n10970), .A2(n10969), .ZN(n12440) );
  NOR2_X1 U11208 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15664), .ZN(
        n16382) );
  INV_X1 U11209 ( .A(n17565), .ZN(n18010) );
  AND2_X1 U11210 ( .A1(n14478), .A2(n14480), .ZN(n14467) );
  NAND2_X1 U11211 ( .A1(n9885), .A2(n9884), .ZN(n10932) );
  NAND4_X1 U11212 ( .A1(n9933), .A2(n9931), .A3(n14355), .A4(n9930), .ZN(
        n15042) );
  NAND3_X1 U11213 ( .A1(n10197), .A2(n10196), .A3(n10195), .ZN(n16398) );
  OAI21_X1 U11214 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18845), .A(n16555), 
        .ZN(n17872) );
  INV_X1 U11215 ( .A(n16121), .ZN(n16122) );
  XNOR2_X1 U11216 ( .A(n12387), .B(n12782), .ZN(n14784) );
  INV_X2 U11218 ( .A(n9757), .ZN(n15790) );
  OR2_X2 U11219 ( .A1(n10202), .A2(n13269), .ZN(n10203) );
  NAND4_X4 U11220 ( .A1(n11530), .A2(n9766), .A3(n11529), .A4(n11528), .ZN(
        n11536) );
  NOR2_X2 U11221 ( .A1(n17503), .A2(n17324), .ZN(n17316) );
  AND4_X2 U11222 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n11530) );
  OAI21_X2 U11223 ( .B1(n9718), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n16232), .ZN(n10843) );
  AND2_X4 U11224 ( .A1(n15378), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9708) );
  INV_X4 U11227 ( .A(n10543), .ZN(n11084) );
  MUX2_X2 U11228 ( .A(n10498), .B(n10497), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10543) );
  NAND2_X2 U11230 ( .A1(n9827), .A2(n10584), .ZN(n10612) );
  OR2_X2 U11231 ( .A1(n13356), .A2(n11346), .ZN(n11199) );
  BUF_X4 U11232 ( .A(n15790), .Z(n9711) );
  NAND2_X2 U11234 ( .A1(n12624), .A2(n12623), .ZN(n12628) );
  NOR2_X2 U11237 ( .A1(n10101), .A2(n9869), .ZN(n10098) );
  OR2_X4 U11238 ( .A1(n10648), .A2(n12824), .ZN(n10659) );
  AND2_X4 U11239 ( .A1(n11391), .A2(n11389), .ZN(n12096) );
  CLKBUF_X1 U11240 ( .A(n13703), .Z(n9714) );
  OAI21_X2 U11241 ( .B1(n14299), .B2(n14300), .A(n12498), .ZN(n12502) );
  BUF_X2 U11242 ( .A(n16234), .Z(n9718) );
  NOR2_X2 U11243 ( .A1(n10175), .A2(n10174), .ZN(n18217) );
  NOR2_X2 U11244 ( .A1(n18810), .A2(n17868), .ZN(n17729) );
  AND3_X1 U11245 ( .A1(n9887), .A2(n9749), .A3(n9886), .ZN(n15054) );
  INV_X1 U11247 ( .A(n15308), .ZN(n9719) );
  AND2_X1 U11248 ( .A1(n14467), .A2(n9788), .ZN(n14442) );
  NAND2_X1 U11249 ( .A1(n15146), .A2(n15147), .ZN(n10881) );
  NOR2_X1 U11250 ( .A1(n11055), .A2(n14095), .ZN(n14089) );
  NAND2_X1 U11251 ( .A1(n10787), .A2(n11065), .ZN(n11055) );
  AND2_X1 U11252 ( .A1(n13227), .A2(n9818), .ZN(n13158) );
  OR2_X1 U11253 ( .A1(n12459), .A2(n12458), .ZN(n15083) );
  NAND2_X2 U11254 ( .A1(n12861), .A2(n12860), .ZN(n14007) );
  NOR2_X1 U11255 ( .A1(n19505), .A2(n19419), .ZN(n19521) );
  NAND2_X1 U11256 ( .A1(n9929), .A2(n10676), .ZN(n10827) );
  AND2_X1 U11257 ( .A1(n16279), .A2(n9799), .ZN(n14070) );
  NAND2_X1 U11258 ( .A1(n16295), .A2(n16294), .ZN(n16293) );
  INV_X4 U11259 ( .A(n9716), .ZN(n19069) );
  NAND2_X1 U11260 ( .A1(n10911), .A2(n10910), .ZN(n10920) );
  AND2_X1 U11261 ( .A1(n17198), .A2(P3_EBX_REG_7__SCAN_IN), .ZN(n17201) );
  BUF_X2 U11262 ( .A(n16791), .Z(n16843) );
  AOI21_X1 U11263 ( .B1(n18646), .B2(n10201), .A(n10200), .ZN(n13266) );
  AND2_X1 U11264 ( .A1(n11076), .A2(n10569), .ZN(n13728) );
  AND2_X1 U11265 ( .A1(n13172), .A2(n9800), .ZN(n13186) );
  AND2_X1 U11266 ( .A1(n13189), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13172) );
  CLKBUF_X1 U11267 ( .A(n12336), .Z(n13546) );
  INV_X2 U11268 ( .A(n17387), .ZN(n18191) );
  NAND2_X1 U11269 ( .A1(n9940), .A2(n19305), .ZN(n11201) );
  NAND2_X2 U11271 ( .A1(n19968), .A2(n11196), .ZN(n11040) );
  INV_X1 U11272 ( .A(n10549), .ZN(n19305) );
  INV_X2 U11273 ( .A(n18213), .ZN(n17238) );
  NOR2_X2 U11274 ( .A1(n13854), .A2(n13860), .ZN(n13852) );
  CLKBUF_X2 U11275 ( .A(n11617), .Z(n20221) );
  INV_X2 U11276 ( .A(n12209), .ZN(n11608) );
  CLKBUF_X2 U11277 ( .A(n11589), .Z(n12023) );
  AND4_X1 U11278 ( .A1(n11503), .A2(n11502), .A3(n11501), .A4(n11500), .ZN(
        n11509) );
  AND4_X1 U11279 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n11508) );
  BUF_X2 U11280 ( .A(n11583), .Z(n12115) );
  BUF_X2 U11281 ( .A(n11584), .Z(n12102) );
  BUF_X2 U11282 ( .A(n11537), .Z(n12125) );
  BUF_X2 U11283 ( .A(n11646), .Z(n12123) );
  INV_X2 U11284 ( .A(n13276), .ZN(n10125) );
  NOR2_X4 U11285 ( .A1(n16903), .A2(n10113), .ZN(n13276) );
  INV_X4 U11286 ( .A(n9761), .ZN(n17163) );
  CLKBUF_X2 U11287 ( .A(n11567), .Z(n12118) );
  CLKBUF_X2 U11288 ( .A(n11599), .Z(n12097) );
  CLKBUF_X2 U11289 ( .A(n11681), .Z(n11660) );
  AND2_X1 U11290 ( .A1(n9906), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11387) );
  NOR2_X4 U11292 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13673) );
  INV_X4 U11293 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15369) );
  AOI21_X1 U11294 ( .B1(n14357), .B2(n14356), .A(n15054), .ZN(n14360) );
  AOI211_X1 U11295 ( .C1(n14374), .C2(n19263), .A(n14373), .B(n14372), .ZN(
        n14375) );
  AOI21_X1 U11296 ( .B1(n14315), .B2(n19260), .A(n9840), .ZN(n14316) );
  AOI21_X1 U11297 ( .B1(n12396), .B2(n14258), .A(n12395), .ZN(n12418) );
  XNOR2_X1 U11298 ( .A(n12593), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14315) );
  NOR2_X1 U11299 ( .A1(n14694), .A2(n14710), .ZN(n14700) );
  INV_X1 U11300 ( .A(n14318), .ZN(n9934) );
  NOR2_X1 U11301 ( .A1(n15045), .A2(n15046), .ZN(n15044) );
  INV_X1 U11302 ( .A(n15276), .ZN(n16159) );
  NOR2_X1 U11303 ( .A1(n15276), .A2(n15242), .ZN(n16142) );
  NAND2_X1 U11304 ( .A1(n15053), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15045) );
  NAND2_X1 U11305 ( .A1(n15085), .A2(n12462), .ZN(n15076) );
  NOR2_X1 U11306 ( .A1(n15114), .A2(n15212), .ZN(n15207) );
  AOI21_X1 U11307 ( .B1(n9719), .B2(n9752), .A(n9795), .ZN(n15260) );
  NAND2_X2 U11308 ( .A1(n9858), .A2(n11072), .ZN(n12591) );
  NAND2_X1 U11309 ( .A1(n14901), .A2(n14900), .ZN(n14899) );
  XNOR2_X1 U11310 ( .A(n12721), .B(n12720), .ZN(n14411) );
  AOI21_X1 U11311 ( .B1(n12208), .B2(n12207), .A(n12721), .ZN(n14690) );
  NAND2_X1 U11312 ( .A1(n10881), .A2(n9773), .ZN(n15134) );
  AOI211_X1 U11313 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15160), .A(
        n15159), .B(n15158), .ZN(n15163) );
  NAND2_X1 U11314 ( .A1(n14927), .A2(n10042), .ZN(n10043) );
  AND2_X1 U11315 ( .A1(n13165), .A2(n13164), .ZN(n13166) );
  NAND3_X1 U11316 ( .A1(n10033), .A2(n10032), .A3(n10031), .ZN(n14090) );
  NAND2_X1 U11317 ( .A1(n11053), .A2(n14037), .ZN(n10033) );
  AND2_X1 U11318 ( .A1(n10088), .A2(n10082), .ZN(n10042) );
  AOI21_X1 U11319 ( .B1(n9974), .B2(n12589), .A(n12588), .ZN(n12595) );
  NOR2_X1 U11320 ( .A1(n14195), .A2(n14531), .ZN(n14519) );
  AND2_X1 U11321 ( .A1(n9936), .A2(n14357), .ZN(n9935) );
  XNOR2_X1 U11322 ( .A(n11069), .B(n12494), .ZN(n15132) );
  INV_X1 U11323 ( .A(n11069), .ZN(n11071) );
  NAND2_X1 U11324 ( .A1(n12499), .A2(n12478), .ZN(n12484) );
  OR2_X1 U11325 ( .A1(n16073), .A2(n12494), .ZN(n12487) );
  INV_X1 U11326 ( .A(n14049), .ZN(n9720) );
  OR2_X1 U11327 ( .A1(n15791), .A2(n12690), .ZN(n12691) );
  AND2_X1 U11328 ( .A1(n15792), .A2(n12695), .ZN(n14224) );
  INV_X1 U11329 ( .A(n12477), .ZN(n12499) );
  OR2_X1 U11330 ( .A1(n16101), .A2(n12494), .ZN(n12467) );
  AND2_X1 U11331 ( .A1(n14771), .A2(n15804), .ZN(n15792) );
  NOR3_X1 U11332 ( .A1(n17567), .A2(n17574), .A3(n17917), .ZN(n17546) );
  NOR2_X1 U11333 ( .A1(n10827), .A2(n11222), .ZN(n9928) );
  AND2_X1 U11334 ( .A1(n15793), .A2(n12686), .ZN(n14776) );
  NOR2_X1 U11335 ( .A1(n12474), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12479) );
  AND2_X1 U11336 ( .A1(n10784), .A2(n10783), .ZN(n10786) );
  NOR2_X1 U11337 ( .A1(n17568), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17567) );
  NOR2_X1 U11338 ( .A1(n14121), .A2(n11169), .ZN(n14237) );
  NAND2_X1 U11339 ( .A1(n12468), .A2(n14912), .ZN(n12474) );
  INV_X1 U11340 ( .A(n14264), .ZN(n9954) );
  NOR2_X1 U11341 ( .A1(n13812), .A2(n13874), .ZN(n13953) );
  OR2_X1 U11342 ( .A1(n15601), .A2(n12494), .ZN(n12450) );
  NAND2_X1 U11343 ( .A1(n17656), .A2(n17610), .ZN(n17622) );
  AND2_X1 U11344 ( .A1(n12657), .A2(n12656), .ZN(n12658) );
  NOR2_X1 U11345 ( .A1(n9882), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U11346 ( .A1(n13945), .A2(n9792), .ZN(n14146) );
  AND3_X1 U11347 ( .A1(n9845), .A2(n9839), .A3(n9838), .ZN(n9837) );
  NOR2_X1 U11348 ( .A1(n14561), .A2(n14482), .ZN(n14481) );
  AND2_X1 U11349 ( .A1(n9771), .A2(n11864), .ZN(n12641) );
  INV_X1 U11350 ( .A(n10677), .ZN(n19276) );
  AND2_X1 U11351 ( .A1(n9836), .A2(n9835), .ZN(n9839) );
  AOI22_X1 U11352 ( .A1(n19321), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10749), .ZN(n9838) );
  NOR2_X1 U11353 ( .A1(n13745), .A2(n13777), .ZN(n13787) );
  NAND2_X1 U11354 ( .A1(n10632), .A2(n10631), .ZN(n19326) );
  OR2_X1 U11355 ( .A1(n10640), .A2(n10637), .ZN(n19381) );
  NAND2_X1 U11356 ( .A1(n12854), .A2(n12850), .ZN(n13740) );
  AND2_X1 U11357 ( .A1(n10041), .A2(n9796), .ZN(n12854) );
  NOR2_X1 U11358 ( .A1(n10651), .A2(n10649), .ZN(n10757) );
  INV_X1 U11359 ( .A(n17824), .ZN(n17877) );
  NOR2_X1 U11360 ( .A1(n15580), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17785) );
  CLKBUF_X1 U11361 ( .A(n12749), .Z(n14675) );
  NAND2_X1 U11362 ( .A1(n9853), .A2(n10636), .ZN(n10637) );
  XNOR2_X1 U11363 ( .A(n15375), .B(n12835), .ZN(n13584) );
  NAND2_X2 U11364 ( .A1(n14670), .A2(n13748), .ZN(n14679) );
  NAND2_X1 U11365 ( .A1(n18846), .A2(n18687), .ZN(n16555) );
  NAND2_X1 U11366 ( .A1(n9883), .A2(n9789), .ZN(n10943) );
  NOR2_X1 U11367 ( .A1(n9770), .A2(n10629), .ZN(n10636) );
  NAND2_X1 U11368 ( .A1(n12834), .A2(n12833), .ZN(n15375) );
  INV_X1 U11369 ( .A(n16391), .ZN(n18687) );
  INV_X1 U11370 ( .A(n10932), .ZN(n9883) );
  OR2_X1 U11371 ( .A1(n11707), .A2(n11706), .ZN(n11708) );
  XNOR2_X1 U11372 ( .A(n11707), .B(n11705), .ZN(n11822) );
  NAND2_X1 U11373 ( .A1(n14611), .A2(n20234), .ZN(n14612) );
  INV_X1 U11374 ( .A(n18639), .ZN(n16380) );
  NAND2_X1 U11375 ( .A1(n13272), .A2(n18076), .ZN(n18639) );
  NAND2_X1 U11376 ( .A1(n10616), .A2(n10615), .ZN(n11101) );
  INV_X1 U11377 ( .A(n10920), .ZN(n9885) );
  NAND2_X1 U11378 ( .A1(n10606), .A2(n10604), .ZN(n10626) );
  CLKBUF_X1 U11379 ( .A(n12616), .Z(n20579) );
  NOR2_X2 U11380 ( .A1(n16398), .A2(n18091), .ZN(n18633) );
  INV_X1 U11381 ( .A(n18091), .ZN(n18076) );
  NAND2_X1 U11382 ( .A1(n10912), .A2(n12473), .ZN(n10911) );
  AND2_X1 U11383 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17202), .ZN(n17198) );
  NOR2_X2 U11384 ( .A1(n19300), .A2(n19310), .ZN(n19301) );
  NAND3_X1 U11385 ( .A1(n10609), .A2(n10611), .A3(n9758), .ZN(n10617) );
  AND2_X1 U11386 ( .A1(n11698), .A2(n11697), .ZN(n11701) );
  OAI211_X1 U11387 ( .C1(n10588), .C2(n19969), .A(n9763), .B(n10587), .ZN(
        n10620) );
  AOI21_X1 U11388 ( .B1(n11714), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11718), .ZN(n11723) );
  INV_X2 U11389 ( .A(n17502), .ZN(n17495) );
  INV_X2 U11390 ( .A(n17228), .ZN(n17225) );
  INV_X2 U11391 ( .A(n11102), .ZN(n12538) );
  NAND2_X1 U11392 ( .A1(n10888), .A2(n11235), .ZN(n12473) );
  NOR2_X1 U11393 ( .A1(n10599), .A2(n10598), .ZN(n10601) );
  NOR2_X2 U11394 ( .A1(n9878), .A2(n10844), .ZN(n10888) );
  OR2_X1 U11395 ( .A1(n15692), .A2(n9926), .ZN(n17227) );
  NAND3_X1 U11396 ( .A1(n10049), .A2(n10591), .A3(n10048), .ZN(n10607) );
  NAND2_X1 U11397 ( .A1(n14244), .A2(n14245), .ZN(n18631) );
  NAND2_X1 U11398 ( .A1(n13728), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10610) );
  NOR2_X2 U11399 ( .A1(n17349), .A2(n16447), .ZN(n17786) );
  NAND2_X1 U11400 ( .A1(n11081), .A2(n9828), .ZN(n10580) );
  AND2_X1 U11401 ( .A1(n9941), .A2(n13535), .ZN(n13534) );
  BUF_X4 U11402 ( .A(n10608), .Z(n12543) );
  OR2_X1 U11403 ( .A1(n11185), .A2(n19967), .ZN(n10584) );
  AND2_X2 U11404 ( .A1(n10565), .A2(n13023), .ZN(n10608) );
  NAND2_X1 U11405 ( .A1(n11199), .A2(n11198), .ZN(n9941) );
  NAND2_X1 U11406 ( .A1(n10542), .A2(n10541), .ZN(n11081) );
  NAND2_X1 U11407 ( .A1(n10567), .A2(n10528), .ZN(n10055) );
  NAND2_X1 U11408 ( .A1(n13211), .A2(n16353), .ZN(n11186) );
  NAND2_X1 U11409 ( .A1(n10805), .A2(n10804), .ZN(n10840) );
  INV_X1 U11410 ( .A(n10567), .ZN(n11076) );
  NAND2_X1 U11411 ( .A1(n10554), .A2(n16351), .ZN(n16353) );
  INV_X1 U11412 ( .A(n10919), .ZN(n9884) );
  OR2_X1 U11413 ( .A1(n12764), .A2(n12284), .ZN(n12734) );
  AND2_X1 U11414 ( .A1(n10502), .A2(n10501), .ZN(n10529) );
  INV_X1 U11415 ( .A(n12356), .ZN(n12380) );
  AND3_X1 U11416 ( .A1(n9747), .A2(n10543), .A3(n9848), .ZN(n10554) );
  INV_X1 U11417 ( .A(n11610), .ZN(n11790) );
  NAND3_X1 U11418 ( .A1(n13382), .A2(n11558), .A3(n11619), .ZN(n12764) );
  NAND2_X1 U11419 ( .A1(n12301), .A2(n12329), .ZN(n12371) );
  AND2_X1 U11420 ( .A1(n11612), .A2(n11628), .ZN(n11615) );
  INV_X2 U11421 ( .A(n17321), .ZN(n18226) );
  INV_X2 U11422 ( .A(n16398), .ZN(n18850) );
  OR2_X1 U11423 ( .A1(n10548), .A2(n9940), .ZN(n11190) );
  NAND2_X1 U11424 ( .A1(n9765), .A2(n9987), .ZN(n17376) );
  OR2_X1 U11425 ( .A1(n11621), .A2(n11611), .ZN(n14829) );
  OR2_X1 U11426 ( .A1(n10675), .A2(n10674), .ZN(n10814) );
  OR2_X2 U11427 ( .A1(n10797), .A2(n10796), .ZN(n12496) );
  NOR2_X1 U11428 ( .A1(n12278), .A2(n20764), .ZN(n11994) );
  INV_X1 U11429 ( .A(n12284), .ZN(n12301) );
  INV_X1 U11430 ( .A(n18199), .ZN(n13269) );
  AND2_X1 U11431 ( .A1(n11620), .A2(n11619), .ZN(n11630) );
  INV_X2 U11432 ( .A(n11019), .ZN(n10499) );
  NAND2_X1 U11433 ( .A1(n9727), .A2(n13854), .ZN(n11631) );
  CLKBUF_X1 U11434 ( .A(n11629), .Z(n20228) );
  INV_X1 U11435 ( .A(n11609), .ZN(n11629) );
  AND4_X1 U11436 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10498) );
  AND4_X1 U11437 ( .A1(n10496), .A2(n10495), .A3(n10494), .A4(n10493), .ZN(
        n10497) );
  AND4_X1 U11438 ( .A1(n11566), .A2(n11565), .A3(n11564), .A4(n11563), .ZN(
        n11578) );
  AND4_X1 U11439 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11576) );
  AND2_X2 U11440 ( .A1(n9731), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10704) );
  INV_X4 U11441 ( .A(n15511), .ZN(n17175) );
  AND4_X1 U11442 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11579) );
  AND4_X1 U11443 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11577) );
  INV_X4 U11444 ( .A(n15522), .ZN(n17174) );
  AND4_X1 U11445 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(
        n11511) );
  AND4_X1 U11446 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11510) );
  INV_X2 U11447 ( .A(n17128), .ZN(n17184) );
  AND4_X1 U11448 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11607) );
  AND2_X1 U11449 ( .A1(n13193), .A2(n12410), .ZN(n13201) );
  AND4_X1 U11450 ( .A1(n11598), .A2(n11597), .A3(n11596), .A4(n11595), .ZN(
        n11605) );
  AND2_X1 U11451 ( .A1(n10465), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10468) );
  AND4_X1 U11452 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n11606) );
  INV_X2 U11453 ( .A(n16540), .ZN(U215) );
  INV_X2 U11454 ( .A(n9756), .ZN(n17116) );
  NAND2_X2 U11455 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19985), .ZN(n19898) );
  NAND2_X2 U11456 ( .A1(n19985), .A2(n19852), .ZN(n19901) );
  NOR2_X1 U11457 ( .A1(n17697), .A2(n9874), .ZN(n9873) );
  INV_X2 U11459 ( .A(n17180), .ZN(n17125) );
  NAND2_X1 U11460 ( .A1(n9997), .A2(n9996), .ZN(n15522) );
  INV_X2 U11461 ( .A(n12404), .ZN(n9722) );
  AND2_X2 U11462 ( .A1(n11387), .A2(n11391), .ZN(n11583) );
  INV_X2 U11463 ( .A(n13117), .ZN(n9723) );
  INV_X2 U11464 ( .A(n16542), .ZN(n16544) );
  INV_X2 U11465 ( .A(n18162), .ZN(n9724) );
  AND2_X1 U11466 ( .A1(n9866), .A2(n9865), .ZN(n13198) );
  CLKBUF_X1 U11467 ( .A(n12116), .Z(n12080) );
  NOR2_X1 U11468 ( .A1(n10115), .A2(n10111), .ZN(n13274) );
  AND2_X2 U11469 ( .A1(n11388), .A2(n13647), .ZN(n11647) );
  AND2_X2 U11470 ( .A1(n9708), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12965) );
  NAND2_X1 U11471 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18825), .ZN(
        n10110) );
  NAND2_X1 U11472 ( .A1(n18825), .A2(n18831), .ZN(n16903) );
  INV_X2 U11473 ( .A(n20133), .ZN(n9726) );
  AND2_X1 U11474 ( .A1(n11381), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11388) );
  NOR2_X1 U11475 ( .A1(n11382), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11389) );
  AND2_X1 U11476 ( .A1(n13656), .A2(n13647), .ZN(n9741) );
  AND2_X2 U11477 ( .A1(n13673), .A2(n13656), .ZN(n12124) );
  INV_X2 U11478 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18817) );
  AND2_X1 U11479 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13647) );
  AND2_X1 U11480 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13656) );
  NOR2_X2 U11481 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13655) );
  AND2_X2 U11482 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13654) );
  INV_X1 U11483 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13473) );
  NAND2_X1 U11484 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13195) );
  NOR2_X2 U11485 ( .A1(n14007), .A2(n12862), .ZN(n14015) );
  OR2_X1 U11486 ( .A1(n14282), .A2(n12704), .ZN(n14682) );
  AND2_X2 U11487 ( .A1(n14709), .A2(n14282), .ZN(n9744) );
  INV_X1 U11488 ( .A(n13860), .ZN(n9727) );
  OR2_X1 U11489 ( .A1(n10110), .A2(n10112), .ZN(n17180) );
  NAND2_X1 U11490 ( .A1(n10043), .A2(n10044), .ZN(n13027) );
  NOR2_X1 U11491 ( .A1(n10115), .A2(n10110), .ZN(n13273) );
  OR2_X1 U11492 ( .A1(n12791), .A2(n11536), .ZN(n11637) );
  NOR2_X1 U11493 ( .A1(n16052), .A2(n19069), .ZN(n16035) );
  OR2_X1 U11494 ( .A1(n18657), .A2(n10114), .ZN(n9756) );
  AND2_X2 U11495 ( .A1(n12591), .A2(n9857), .ZN(n16192) );
  AND2_X2 U11496 ( .A1(n14153), .A2(n10052), .ZN(n12980) );
  INV_X4 U11497 ( .A(n17144), .ZN(n17080) );
  OR2_X2 U11498 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n14252), .ZN(
        n17144) );
  OAI21_X2 U11499 ( .B1(n10737), .B2(n10736), .A(n10735), .ZN(n10828) );
  NAND2_X1 U11500 ( .A1(n12698), .A2(n14761), .ZN(n14744) );
  AND2_X1 U11501 ( .A1(n14761), .A2(n10003), .ZN(n10002) );
  OR2_X1 U11502 ( .A1(n11065), .A2(n11064), .ZN(n11069) );
  NAND2_X2 U11503 ( .A1(n9831), .A2(n10786), .ZN(n11065) );
  INV_X4 U11504 ( .A(n13117), .ZN(n9731) );
  INV_X4 U11505 ( .A(n13117), .ZN(n9732) );
  NAND2_X4 U11506 ( .A1(n10442), .A2(n15369), .ZN(n13117) );
  INV_X1 U11507 ( .A(n12544), .ZN(n9733) );
  INV_X2 U11508 ( .A(n12544), .ZN(n12542) );
  NOR2_X4 U11509 ( .A1(n10659), .A2(n13995), .ZN(n10764) );
  OR2_X2 U11510 ( .A1(n11186), .A2(n10557), .ZN(n11180) );
  INV_X1 U11511 ( .A(n19094), .ZN(n10622) );
  NAND2_X1 U11512 ( .A1(n9905), .A2(n11694), .ZN(n11713) );
  NAND3_X1 U11513 ( .A1(n10049), .A2(n10591), .A3(n10048), .ZN(n9734) );
  NAND3_X1 U11514 ( .A1(n10049), .A2(n10591), .A3(n10048), .ZN(n9735) );
  INV_X1 U11515 ( .A(n12283), .ZN(n9736) );
  AND2_X1 U11516 ( .A1(n12600), .A2(n13860), .ZN(n12283) );
  INV_X1 U11517 ( .A(n9856), .ZN(n10627) );
  NOR2_X4 U11518 ( .A1(n18657), .A2(n10113), .ZN(n10107) );
  NAND2_X1 U11519 ( .A1(n10621), .A2(n10620), .ZN(n9856) );
  INV_X2 U11521 ( .A(n13129), .ZN(n9738) );
  AND2_X4 U11523 ( .A1(n10665), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11244) );
  AND2_X1 U11524 ( .A1(n11747), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12232) );
  INV_X1 U11525 ( .A(n12270), .ZN(n12259) );
  OR2_X1 U11526 ( .A1(n10874), .A2(n10873), .ZN(n10877) );
  NAND2_X1 U11527 ( .A1(n11184), .A2(n10050), .ZN(n10591) );
  NOR2_X1 U11528 ( .A1(n10051), .A2(n19969), .ZN(n10050) );
  NAND2_X1 U11529 ( .A1(n10055), .A2(n16351), .ZN(n9828) );
  INV_X1 U11530 ( .A(n14444), .ZN(n10026) );
  NAND2_X1 U11531 ( .A1(n11867), .A2(n11866), .ZN(n12674) );
  INV_X1 U11532 ( .A(n11865), .ZN(n11866) );
  OR2_X1 U11533 ( .A1(n11666), .A2(n11665), .ZN(n12676) );
  AOI21_X1 U11534 ( .B1(n12615), .B2(n12627), .A(n20172), .ZN(n9916) );
  NAND2_X1 U11535 ( .A1(n12616), .A2(n12615), .ZN(n9917) );
  AND2_X1 U11536 ( .A1(n20760), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12276) );
  NAND2_X1 U11537 ( .A1(n13051), .A2(n13053), .ZN(n13054) );
  INV_X1 U11538 ( .A(n10618), .ZN(n10615) );
  INV_X1 U11539 ( .A(n10617), .ZN(n10616) );
  NOR2_X1 U11540 ( .A1(n12509), .A2(n9978), .ZN(n9977) );
  INV_X1 U11541 ( .A(n14151), .ZN(n9978) );
  OR2_X1 U11542 ( .A1(n14940), .A2(n12508), .ZN(n12509) );
  AND2_X1 U11543 ( .A1(n9751), .A2(n10067), .ZN(n10066) );
  INV_X1 U11544 ( .A(n12455), .ZN(n10067) );
  OAI21_X1 U11545 ( .B1(n9750), .B2(n10070), .A(n15272), .ZN(n10069) );
  INV_X1 U11546 ( .A(n12436), .ZN(n10070) );
  INV_X1 U11547 ( .A(n15315), .ZN(n9959) );
  NOR2_X1 U11548 ( .A1(n9786), .A2(n10060), .ZN(n10059) );
  NAND2_X1 U11549 ( .A1(n15134), .A2(n10062), .ZN(n9832) );
  NOR2_X1 U11550 ( .A1(n16187), .A2(n10061), .ZN(n10060) );
  NAND2_X1 U11551 ( .A1(n18831), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10111) );
  AND2_X1 U11552 ( .A1(n15675), .A2(n12699), .ZN(n14751) );
  NAND2_X1 U11553 ( .A1(n14759), .A2(n9711), .ZN(n14761) );
  NAND2_X1 U11554 ( .A1(n14182), .A2(n10012), .ZN(n14759) );
  AND2_X1 U11555 ( .A1(n12276), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13460) );
  AOI21_X1 U11556 ( .B1(n12271), .B2(n12270), .A(n12269), .ZN(n12274) );
  NAND2_X1 U11557 ( .A1(n12261), .A2(n12260), .ZN(n12275) );
  OR2_X1 U11558 ( .A1(n14146), .A2(n11156), .ZN(n14121) );
  OR2_X1 U11559 ( .A1(n11155), .A2(n14145), .ZN(n11156) );
  OR2_X1 U11560 ( .A1(n14920), .A2(n14321), .ZN(n14903) );
  AND2_X1 U11561 ( .A1(n19969), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12848) );
  NAND2_X1 U11562 ( .A1(n11020), .A2(n11017), .ZN(n16344) );
  NAND2_X1 U11563 ( .A1(n13398), .A2(n11016), .ZN(n11017) );
  AND2_X1 U11564 ( .A1(n10976), .A2(n10975), .ZN(n11011) );
  OR2_X1 U11565 ( .A1(n16661), .A2(n16791), .ZN(n9875) );
  AND2_X1 U11566 ( .A1(n19988), .A2(n19986), .ZN(n13847) );
  XOR2_X1 U11567 ( .A(n14304), .B(n14303), .Z(n16047) );
  OAI21_X1 U11568 ( .B1(n19381), .B2(n10687), .A(n11191), .ZN(n10688) );
  NAND2_X1 U11569 ( .A1(n9846), .A2(n10647), .ZN(n9836) );
  AOI21_X1 U11570 ( .B1(n12115), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n9897), .ZN(n11765) );
  AND2_X1 U11571 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n9897)
         );
  NAND2_X1 U11572 ( .A1(n9743), .A2(n9760), .ZN(n11636) );
  OR2_X1 U11573 ( .A1(n12209), .A2(n11629), .ZN(n11620) );
  AND2_X1 U11574 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n9898)
         );
  BUF_X1 U11575 ( .A(n12096), .Z(n12024) );
  BUF_X1 U11576 ( .A(n12124), .Z(n12064) );
  INV_X1 U11577 ( .A(n12684), .ZN(n9913) );
  INV_X1 U11578 ( .A(n10012), .ZN(n9914) );
  INV_X1 U11579 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10000) );
  INV_X1 U11580 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9906) );
  AOI21_X1 U11581 ( .B1(n12115), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n9896), .ZN(n11752) );
  AND2_X1 U11582 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n9896)
         );
  NAND2_X1 U11583 ( .A1(n13860), .A2(n13854), .ZN(n12284) );
  AOI21_X1 U11584 ( .B1(n12097), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A(n9903), .ZN(n11677) );
  AND2_X1 U11585 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n9903)
         );
  BUF_X1 U11586 ( .A(n12004), .Z(n12117) );
  AND2_X1 U11587 ( .A1(n10876), .A2(n10875), .ZN(n11061) );
  NAND2_X1 U11588 ( .A1(n9856), .A2(n10578), .ZN(n9939) );
  OAI21_X1 U11589 ( .B1(n10610), .B2(n19090), .A(n10582), .ZN(n10583) );
  NOR2_X1 U11590 ( .A1(n15374), .A2(n19077), .ZN(n10581) );
  OAI211_X1 U11591 ( .C1(n10499), .C2(n11029), .A(n10056), .B(n10547), .ZN(
        n11082) );
  NAND2_X1 U11592 ( .A1(n10499), .A2(n11201), .ZN(n10056) );
  NOR2_X1 U11593 ( .A1(n10554), .A2(n19968), .ZN(n10541) );
  AND2_X1 U11594 ( .A1(n10561), .A2(n10544), .ZN(n10540) );
  NOR2_X1 U11595 ( .A1(n10651), .A2(n15387), .ZN(n10658) );
  INV_X1 U11596 ( .A(n10637), .ZN(n10641) );
  NAND2_X1 U11597 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18817), .ZN(
        n10114) );
  AOI21_X1 U11598 ( .B1(n15394), .B2(n18213), .A(n10203), .ZN(n13243) );
  NOR2_X1 U11599 ( .A1(n17871), .A2(n13329), .ZN(n13330) );
  NOR2_X1 U11600 ( .A1(n18217), .A2(n17238), .ZN(n10202) );
  NAND2_X1 U11601 ( .A1(n13243), .A2(n13240), .ZN(n13237) );
  NAND2_X1 U11602 ( .A1(n11609), .A2(n11619), .ZN(n11610) );
  AND2_X1 U11603 ( .A1(n12138), .A2(n14596), .ZN(n10029) );
  AND2_X1 U11604 ( .A1(n14570), .A2(n14493), .ZN(n12138) );
  NOR2_X1 U11605 ( .A1(n14765), .A2(n12032), .ZN(n12033) );
  INV_X1 U11606 ( .A(n12195), .ZN(n12201) );
  NAND2_X1 U11607 ( .A1(n9767), .A2(n14142), .ZN(n10024) );
  AND2_X1 U11608 ( .A1(n9802), .A2(n14129), .ZN(n10023) );
  NAND2_X1 U11609 ( .A1(n11892), .A2(n10021), .ZN(n10020) );
  INV_X1 U11610 ( .A(n14021), .ZN(n10021) );
  AOI21_X1 U11611 ( .B1(n12123), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n9899), .ZN(n11880) );
  INV_X1 U11612 ( .A(n12718), .ZN(n12035) );
  NAND2_X1 U11613 ( .A1(n20234), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12112) );
  NAND2_X1 U11614 ( .A1(n12703), .A2(n9712), .ZN(n14718) );
  NAND2_X1 U11615 ( .A1(n15768), .A2(n12703), .ZN(n14692) );
  NOR2_X1 U11616 ( .A1(n9973), .A2(n14567), .ZN(n9972) );
  INV_X1 U11617 ( .A(n14573), .ZN(n9973) );
  NOR2_X2 U11618 ( .A1(n9736), .A2(n12284), .ZN(n12356) );
  INV_X1 U11619 ( .A(n12283), .ZN(n9907) );
  INV_X1 U11620 ( .A(n14030), .ZN(n9969) );
  XNOR2_X1 U11621 ( .A(n12674), .B(n11870), .ZN(n10016) );
  NAND2_X1 U11622 ( .A1(n9736), .A2(n12296), .ZN(n12336) );
  AND2_X1 U11623 ( .A1(n12209), .A2(n13860), .ZN(n12670) );
  OAI21_X1 U11624 ( .B1(n12259), .B2(n11674), .A(n11673), .ZN(n11829) );
  AND2_X1 U11625 ( .A1(n11690), .A2(n11689), .ZN(n11705) );
  NAND2_X1 U11626 ( .A1(n9826), .A2(n10552), .ZN(n11185) );
  INV_X1 U11627 ( .A(n10553), .ZN(n9826) );
  NAND2_X1 U11628 ( .A1(n11186), .A2(n10564), .ZN(n10049) );
  NAND2_X1 U11629 ( .A1(n10557), .A2(n10564), .ZN(n10048) );
  NAND2_X1 U11630 ( .A1(n12443), .A2(n9754), .ZN(n9882) );
  INV_X1 U11631 ( .A(n9881), .ZN(n9876) );
  INV_X1 U11632 ( .A(n10830), .ZN(n9877) );
  NAND2_X1 U11633 ( .A1(n10082), .A2(n14916), .ZN(n10044) );
  NOR2_X1 U11634 ( .A1(n11361), .A2(n9955), .ZN(n9953) );
  AND2_X1 U11635 ( .A1(n12934), .A2(n14154), .ZN(n10054) );
  INV_X1 U11636 ( .A(n14008), .ZN(n9981) );
  NOR2_X1 U11637 ( .A1(n14950), .A2(n9958), .ZN(n9957) );
  INV_X1 U11638 ( .A(n13228), .ZN(n9958) );
  NOR2_X1 U11639 ( .A1(n15173), .A2(n10038), .ZN(n10037) );
  AND2_X1 U11640 ( .A1(n12590), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10034) );
  AND2_X1 U11641 ( .A1(n10918), .A2(n15311), .ZN(n12455) );
  INV_X1 U11642 ( .A(n16267), .ZN(n9961) );
  AND2_X1 U11643 ( .A1(n10892), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16209) );
  NAND2_X1 U11644 ( .A1(n9850), .A2(n11068), .ZN(n16204) );
  INV_X1 U11645 ( .A(n15136), .ZN(n10886) );
  NAND2_X1 U11646 ( .A1(n10058), .A2(n10057), .ZN(n9844) );
  NAND2_X1 U11647 ( .A1(n11101), .A2(n10619), .ZN(n10030) );
  NAND2_X1 U11648 ( .A1(n9939), .A2(n10594), .ZN(n10624) );
  AND2_X1 U11649 ( .A1(n10561), .A2(n11023), .ZN(n10562) );
  NOR2_X1 U11650 ( .A1(n12824), .A2(n10628), .ZN(n10631) );
  INV_X1 U11651 ( .A(n13293), .ZN(n13277) );
  INV_X1 U11652 ( .A(n13288), .ZN(n17128) );
  NOR2_X1 U11653 ( .A1(n16903), .A2(n10114), .ZN(n13278) );
  NOR2_X1 U11654 ( .A1(n17356), .A2(n15556), .ZN(n15555) );
  NAND2_X1 U11655 ( .A1(n15582), .A2(n17610), .ZN(n15588) );
  NOR2_X1 U11656 ( .A1(n10110), .A2(n10113), .ZN(n13289) );
  NAND2_X1 U11657 ( .A1(n9986), .A2(n9985), .ZN(n9984) );
  NAND2_X1 U11658 ( .A1(n15541), .A2(n18129), .ZN(n9985) );
  INV_X1 U11659 ( .A(n17819), .ZN(n9986) );
  NAND2_X1 U11660 ( .A1(n15536), .A2(n15537), .ZN(n15539) );
  INV_X1 U11661 ( .A(n17376), .ZN(n13329) );
  NAND2_X1 U11662 ( .A1(n18217), .A2(n15394), .ZN(n18646) );
  AOI22_X1 U11663 ( .A1(n18638), .A2(n16380), .B1(n18635), .B2(n18633), .ZN(
        n16391) );
  INV_X2 U11664 ( .A(n12112), .ZN(n12719) );
  AND2_X1 U11665 ( .A1(n9788), .A2(n12709), .ZN(n10025) );
  NAND2_X1 U11666 ( .A1(n11378), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12189) );
  INV_X1 U11667 ( .A(n12184), .ZN(n11378) );
  OR2_X1 U11668 ( .A1(n14598), .A2(n14492), .ZN(n14586) );
  OR2_X1 U11669 ( .A1(n14598), .A2(n14507), .ZN(n14584) );
  NOR2_X1 U11670 ( .A1(n11985), .A2(n14201), .ZN(n12002) );
  NAND2_X1 U11671 ( .A1(n12002), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12032) );
  NAND2_X1 U11672 ( .A1(n9910), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9909) );
  INV_X1 U11673 ( .A(n12757), .ZN(n9910) );
  AND2_X1 U11674 ( .A1(n14761), .A2(n9745), .ZN(n10001) );
  NAND2_X1 U11675 ( .A1(n13957), .A2(n9762), .ZN(n14033) );
  NAND2_X1 U11676 ( .A1(n13957), .A2(n12315), .ZN(n14031) );
  NOR2_X1 U11677 ( .A1(n15685), .A2(n15928), .ZN(n15966) );
  AND2_X1 U11678 ( .A1(n12776), .A2(n13460), .ZN(n12807) );
  XNOR2_X1 U11679 ( .A(n11830), .B(n11829), .ZN(n12616) );
  CLKBUF_X1 U11680 ( .A(n12722), .Z(n12723) );
  INV_X1 U11681 ( .A(n20342), .ZN(n20238) );
  NOR2_X1 U11682 ( .A1(n20521), .A2(n20342), .ZN(n20666) );
  AND2_X1 U11683 ( .A1(n12484), .A2(n12482), .ZN(n16059) );
  INV_X1 U11684 ( .A(n19300), .ZN(n10803) );
  AND2_X1 U11685 ( .A1(n11168), .A2(n11167), .ZN(n12402) );
  AND2_X1 U11686 ( .A1(n13794), .A2(n13792), .ZN(n13793) );
  NAND2_X1 U11687 ( .A1(n9768), .A2(n14899), .ZN(n10045) );
  AND2_X1 U11688 ( .A1(n9806), .A2(n9951), .ZN(n9950) );
  INV_X1 U11689 ( .A(n14977), .ZN(n9951) );
  NAND2_X1 U11690 ( .A1(n14995), .A2(n9806), .ZN(n14978) );
  NAND2_X1 U11691 ( .A1(n13175), .A2(n9753), .ZN(n9863) );
  NOR2_X1 U11692 ( .A1(n14903), .A2(n14902), .ZN(n14904) );
  NAND2_X1 U11693 ( .A1(n11055), .A2(n14095), .ZN(n10031) );
  AND2_X1 U11694 ( .A1(n9849), .A2(n11101), .ZN(n13744) );
  OAI21_X1 U11695 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n14358), .ZN(n9930) );
  NAND2_X1 U11696 ( .A1(n9932), .A2(n9934), .ZN(n9931) );
  AND2_X1 U11697 ( .A1(n16059), .A2(n12496), .ZN(n14357) );
  INV_X1 U11698 ( .A(n14922), .ZN(n9975) );
  NAND2_X1 U11699 ( .A1(n14237), .A2(n9976), .ZN(n14933) );
  NAND2_X1 U11700 ( .A1(n15202), .A2(n15296), .ZN(n10068) );
  NAND2_X1 U11701 ( .A1(n10923), .A2(n15296), .ZN(n10071) );
  NAND2_X1 U11702 ( .A1(n13786), .A2(n9772), .ZN(n13946) );
  AND2_X1 U11703 ( .A1(n10900), .A2(n10896), .ZN(n10064) );
  OR2_X1 U11704 ( .A1(n15134), .A2(n16209), .ZN(n10065) );
  AND2_X1 U11705 ( .A1(n11235), .A2(n13431), .ZN(n11236) );
  AND3_X1 U11706 ( .A1(n13579), .A2(n11094), .A3(n14380), .ZN(n11096) );
  NAND2_X1 U11707 ( .A1(n12825), .A2(n19533), .ZN(n12845) );
  NAND2_X1 U11708 ( .A1(n12838), .A2(n12837), .ZN(n13700) );
  NAND2_X1 U11709 ( .A1(n13583), .A2(n13584), .ZN(n12838) );
  INV_X1 U11710 ( .A(n19505), .ZN(n19763) );
  AOI21_X2 U11711 ( .B1(n15390), .B2(n13980), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19768) );
  NAND2_X1 U11712 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19768), .ZN(n19310) );
  AND2_X1 U11713 ( .A1(n10988), .A2(n10987), .ZN(n16339) );
  NOR2_X1 U11714 ( .A1(n18199), .A2(n18647), .ZN(n16546) );
  NAND3_X1 U11715 ( .A1(n10098), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10095) );
  NOR2_X1 U11716 ( .A1(n16791), .A2(n10106), .ZN(n16662) );
  NAND2_X1 U11717 ( .A1(n15523), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n9989) );
  NAND2_X1 U11718 ( .A1(n17778), .A2(n15551), .ZN(n17747) );
  XNOR2_X1 U11719 ( .A(n9984), .B(n15544), .ZN(n17809) );
  NAND2_X1 U11720 ( .A1(n17809), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17808) );
  NAND2_X1 U11721 ( .A1(n17747), .A2(n9998), .ZN(n18037) );
  INV_X1 U11722 ( .A(n18043), .ZN(n9998) );
  NOR2_X1 U11723 ( .A1(n17798), .A2(n17797), .ZN(n17796) );
  OR2_X1 U11724 ( .A1(n15565), .A2(n15564), .ZN(n17816) );
  XOR2_X1 U11725 ( .A(n13329), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17865) );
  INV_X1 U11726 ( .A(n18208), .ZN(n15394) );
  NOR2_X1 U11727 ( .A1(n18213), .A2(n18217), .ZN(n13261) );
  AND2_X1 U11728 ( .A1(n14458), .A2(n13851), .ZN(n20051) );
  INV_X1 U11729 ( .A(n20024), .ZN(n20093) );
  AND2_X1 U11730 ( .A1(n14458), .A2(n13868), .ZN(n20102) );
  AND2_X1 U11731 ( .A1(n12282), .A2(n12281), .ZN(n14568) );
  INV_X1 U11732 ( .A(n14595), .ZN(n13760) );
  INV_X2 U11733 ( .A(n14568), .ZN(n14611) );
  INV_X1 U11734 ( .A(n15775), .ZN(n14655) );
  INV_X1 U11735 ( .A(n14670), .ZN(n14666) );
  NOR2_X1 U11737 ( .A1(n16035), .A2(n16034), .ZN(n16036) );
  XNOR2_X1 U11738 ( .A(n13158), .B(n12573), .ZN(n19101) );
  NAND2_X1 U11739 ( .A1(n9974), .A2(n19263), .ZN(n9841) );
  INV_X1 U11740 ( .A(n16220), .ZN(n19264) );
  OAI21_X1 U11741 ( .B1(n16047), .B2(n16283), .A(n9946), .ZN(n9945) );
  NOR2_X1 U11742 ( .A1(n9947), .A2(n15034), .ZN(n9946) );
  INV_X1 U11743 ( .A(n14309), .ZN(n9947) );
  XNOR2_X1 U11744 ( .A(n15205), .B(n15206), .ZN(n16138) );
  NAND2_X1 U11745 ( .A1(n9830), .A2(n9782), .ZN(n15204) );
  AOI21_X1 U11746 ( .B1(n15107), .B2(n12452), .A(n10963), .ZN(n10972) );
  INV_X1 U11747 ( .A(n16307), .ZN(n16274) );
  OR2_X1 U11748 ( .A1(n15375), .A2(n13433), .ZN(n19945) );
  INV_X1 U11749 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19943) );
  INV_X1 U11750 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15374) );
  NAND2_X1 U11751 ( .A1(n16344), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15390) );
  OAI21_X1 U11752 ( .B1(n16966), .B2(n9919), .A(n9811), .ZN(n16960) );
  OR2_X1 U11753 ( .A1(n9922), .A2(n16956), .ZN(n9919) );
  OR2_X1 U11754 ( .A1(n16381), .A2(n18191), .ZN(n9926) );
  NAND2_X1 U11755 ( .A1(n9995), .A2(n9994), .ZN(n9993) );
  AOI21_X1 U11756 ( .B1(n16433), .B2(n18099), .A(n9784), .ZN(n9994) );
  NAND2_X1 U11757 ( .A1(n16434), .A2(n18633), .ZN(n9995) );
  NAND2_X1 U11758 ( .A1(n13328), .A2(n18159), .ZN(n18133) );
  NAND2_X1 U11759 ( .A1(n19723), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10654) );
  AOI21_X1 U11760 ( .B1(n12115), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n9895), .ZN(n11729) );
  AND2_X1 U11761 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n9895)
         );
  NAND2_X1 U11762 ( .A1(n11621), .A2(n12600), .ZN(n11628) );
  NAND2_X1 U11763 ( .A1(n10757), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10693) );
  INV_X1 U11764 ( .A(n10580), .ZN(n9825) );
  NOR2_X1 U11765 ( .A1(n10571), .A2(n10570), .ZN(n10572) );
  NOR2_X1 U11766 ( .A1(n10610), .A2(n13585), .ZN(n10570) );
  NAND2_X1 U11767 ( .A1(n10547), .A2(n10499), .ZN(n10560) );
  AOI21_X1 U11768 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18677), .A(
        n10207), .ZN(n10208) );
  AOI21_X1 U11769 ( .B1(n12103), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A(n9900), .ZN(n11477) );
  AND2_X1 U11770 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n9900)
         );
  AOI21_X1 U11771 ( .B1(n12080), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A(n9902), .ZN(n11899) );
  AND2_X1 U11772 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n9902)
         );
  AND2_X1 U11773 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n9899)
         );
  OAI21_X1 U11774 ( .B1(n12259), .B2(n11463), .A(n11782), .ZN(n11783) );
  AOI21_X1 U11775 ( .B1(n12102), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A(n9901), .ZN(n11656) );
  AND2_X1 U11776 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n9901)
         );
  OR2_X1 U11777 ( .A1(n11771), .A2(n11770), .ZN(n12642) );
  INV_X1 U11778 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11382) );
  NOR2_X1 U11779 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11390) );
  AND2_X1 U11780 ( .A1(n9894), .A2(n9893), .ZN(n11652) );
  NAND2_X1 U11781 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n9894) );
  NAND2_X1 U11782 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n9893) );
  INV_X1 U11783 ( .A(n12613), .ZN(n11671) );
  NAND2_X1 U11784 ( .A1(n9904), .A2(n11627), .ZN(n11698) );
  NAND2_X1 U11785 ( .A1(n11713), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9904) );
  NAND2_X1 U11786 ( .A1(n12797), .A2(n12283), .ZN(n9962) );
  BUF_X1 U11787 ( .A(n11618), .Z(n12792) );
  CLKBUF_X1 U11788 ( .A(n12764), .Z(n13464) );
  AND2_X1 U11789 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U11790 ( .A1(n11630), .A2(n11623), .ZN(n12791) );
  INV_X1 U11791 ( .A(n12232), .ZN(n12268) );
  NAND2_X1 U11792 ( .A1(n10825), .A2(n10882), .ZN(n9881) );
  NAND2_X1 U11793 ( .A1(n10064), .A2(n16209), .ZN(n10061) );
  NOR2_X1 U11794 ( .A1(n10063), .A2(n16187), .ZN(n10062) );
  INV_X1 U11795 ( .A(n10064), .ZN(n10063) );
  NAND2_X1 U11796 ( .A1(n11201), .A2(n11084), .ZN(n10561) );
  AND3_X2 U11797 ( .A1(n15369), .A2(n9855), .A3(n16318), .ZN(n10509) );
  NAND2_X1 U11798 ( .A1(n9938), .A2(n10594), .ZN(n10629) );
  INV_X1 U11799 ( .A(n9939), .ZN(n9938) );
  AND2_X2 U11800 ( .A1(n9834), .A2(n16318), .ZN(n10488) );
  NOR2_X1 U11801 ( .A1(n17364), .A2(n15552), .ZN(n15557) );
  NOR2_X1 U11802 ( .A1(n13330), .A2(n17370), .ZN(n15507) );
  AOI21_X1 U11803 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18672), .A(
        n10206), .ZN(n10214) );
  AND2_X1 U11804 ( .A1(n13260), .A2(n13256), .ZN(n10206) );
  NAND2_X1 U11805 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11561) );
  INV_X1 U11806 ( .A(n14292), .ZN(n10027) );
  AOI21_X1 U11807 ( .B1(n12115), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n9898), .ZN(n12122) );
  AND2_X1 U11808 ( .A1(n14521), .A2(n14596), .ZN(n14494) );
  NAND2_X1 U11809 ( .A1(n12692), .A2(n12685), .ZN(n10013) );
  NOR2_X1 U11810 ( .A1(n15784), .A2(n15781), .ZN(n12692) );
  NOR2_X1 U11811 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  AND2_X1 U11812 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11374), .ZN(
        n11794) );
  NAND2_X1 U11813 ( .A1(n12620), .A2(n12619), .ZN(n12622) );
  INV_X1 U11814 ( .A(n14025), .ZN(n9968) );
  AND2_X1 U11815 ( .A1(n13956), .A2(n13955), .ZN(n12315) );
  NAND2_X1 U11816 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11587) );
  OR2_X1 U11817 ( .A1(n11758), .A2(n11757), .ZN(n12632) );
  INV_X1 U11818 ( .A(n12671), .ZN(n11702) );
  OR2_X1 U11819 ( .A1(n11687), .A2(n11686), .ZN(n12606) );
  AND2_X1 U11820 ( .A1(n13387), .A2(n12772), .ZN(n13456) );
  INV_X1 U11821 ( .A(n11536), .ZN(n11617) );
  INV_X1 U11822 ( .A(n20579), .ZN(n20194) );
  OAI21_X1 U11823 ( .B1(n20867), .B2(n16019), .A(n14848), .ZN(n20195) );
  INV_X1 U11824 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13669) );
  AND2_X1 U11825 ( .A1(n11746), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U11826 ( .A1(n12270), .A2(n12670), .ZN(n12272) );
  OR2_X1 U11827 ( .A1(n10954), .A2(n10952), .ZN(n10957) );
  NOR2_X1 U11828 ( .A1(n10943), .A2(n10942), .ZN(n10945) );
  NAND2_X1 U11829 ( .A1(n10945), .A2(n10944), .ZN(n10954) );
  NAND2_X1 U11830 ( .A1(n9890), .A2(n9889), .ZN(n10912) );
  NOR2_X1 U11831 ( .A1(n9891), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n9889) );
  INV_X1 U11832 ( .A(n10898), .ZN(n9890) );
  NAND2_X1 U11833 ( .A1(n18991), .A2(n9892), .ZN(n9891) );
  NOR2_X1 U11834 ( .A1(n10898), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U11835 ( .A1(n9949), .A2(n10884), .ZN(n10887) );
  OR2_X1 U11836 ( .A1(n10830), .A2(n9880), .ZN(n9879) );
  NAND2_X1 U11837 ( .A1(n19300), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10804) );
  NAND2_X1 U11838 ( .A1(n10973), .A2(n10803), .ZN(n10805) );
  INV_X1 U11839 ( .A(n14323), .ZN(n9952) );
  NAND2_X1 U11840 ( .A1(n13030), .A2(n13029), .ZN(n13031) );
  INV_X1 U11841 ( .A(n16343), .ZN(n13143) );
  NOR2_X1 U11842 ( .A1(n15048), .A2(n9862), .ZN(n9861) );
  AND2_X1 U11843 ( .A1(n13223), .A2(n14877), .ZN(n9982) );
  AND2_X1 U11844 ( .A1(n13192), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13191) );
  NAND2_X1 U11845 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9867) );
  NOR2_X1 U11846 ( .A1(n10547), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11200) );
  AND2_X1 U11847 ( .A1(n9977), .A2(n14931), .ZN(n9976) );
  AND2_X1 U11848 ( .A1(n9787), .A2(n14014), .ZN(n9980) );
  AND2_X1 U11849 ( .A1(n9785), .A2(n15335), .ZN(n9960) );
  AND2_X1 U11850 ( .A1(n13817), .A2(n13801), .ZN(n9983) );
  INV_X1 U11851 ( .A(n11061), .ZN(n11064) );
  OAI21_X1 U11852 ( .B1(n11055), .B2(n12496), .A(n19048), .ZN(n10848) );
  NAND2_X1 U11853 ( .A1(n10057), .A2(n9928), .ZN(n11052) );
  NAND2_X1 U11854 ( .A1(n9844), .A2(n10829), .ZN(n11041) );
  AND4_X1 U11855 ( .A1(n10556), .A2(n11077), .A3(n19300), .A4(n9848), .ZN(
        n10557) );
  OR2_X1 U11856 ( .A1(n13071), .A2(n19287), .ZN(n12835) );
  AND2_X1 U11857 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13725) );
  NAND3_X1 U11858 ( .A1(n19934), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19768), 
        .ZN(n13983) );
  AND3_X1 U11859 ( .A1(n10544), .A2(n11019), .A3(n11084), .ZN(n10550) );
  NAND2_X1 U11860 ( .A1(n10447), .A2(n10470), .ZN(n9859) );
  NAND2_X1 U11861 ( .A1(n10452), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9860) );
  NAND2_X1 U11862 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18807), .ZN(
        n10115) );
  INV_X1 U11863 ( .A(n10114), .ZN(n9997) );
  INV_X1 U11864 ( .A(n10111), .ZN(n9996) );
  NOR2_X1 U11865 ( .A1(n10112), .A2(n16903), .ZN(n13288) );
  NAND2_X1 U11866 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n10092), .ZN(
        n9871) );
  NOR2_X1 U11867 ( .A1(n18226), .A2(n18204), .ZN(n13240) );
  NOR2_X1 U11868 ( .A1(n17796), .A2(n18107), .ZN(n15546) );
  INV_X1 U11869 ( .A(n13266), .ZN(n13247) );
  OAI22_X1 U11870 ( .A1(n18825), .A2(n18672), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13260) );
  NAND2_X1 U11871 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10112) );
  NOR2_X1 U11872 ( .A1(n13237), .A2(n18646), .ZN(n15396) );
  AND2_X1 U11873 ( .A1(n12730), .A2(n12729), .ZN(n13386) );
  AND2_X1 U11874 ( .A1(n20091), .A2(n14458), .ZN(n20060) );
  NAND2_X1 U11875 ( .A1(n13547), .A2(n12301), .ZN(n9970) );
  INV_X1 U11876 ( .A(n13608), .ZN(n11840) );
  AND2_X1 U11877 ( .A1(n11821), .A2(n11841), .ZN(n10075) );
  OAI21_X1 U11878 ( .B1(n20192), .B2(n11982), .A(n11820), .ZN(n11821) );
  NAND2_X1 U11879 ( .A1(n10075), .A2(n11840), .ZN(n13609) );
  INV_X1 U11880 ( .A(n20189), .ZN(n20190) );
  NOR2_X2 U11881 ( .A1(n12207), .A2(n12208), .ZN(n12721) );
  NAND2_X1 U11882 ( .A1(n11379), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12204) );
  INV_X1 U11883 ( .A(n12189), .ZN(n11379) );
  NAND2_X1 U11884 ( .A1(n14467), .A2(n9781), .ZN(n14443) );
  AND2_X1 U11885 ( .A1(n12162), .A2(n14722), .ZN(n12163) );
  NOR2_X1 U11886 ( .A1(n12145), .A2(n15713), .ZN(n12148) );
  NAND2_X1 U11887 ( .A1(n12148), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12161) );
  AND2_X1 U11888 ( .A1(n10074), .A2(n10029), .ZN(n10028) );
  NOR2_X1 U11889 ( .A1(n12135), .A2(n14514), .ZN(n12093) );
  NAND2_X1 U11890 ( .A1(n12093), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12094) );
  CLKBUF_X1 U11891 ( .A(n14519), .Z(n14520) );
  NAND2_X1 U11892 ( .A1(n11970), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11985) );
  AND2_X1 U11893 ( .A1(n10023), .A2(n12001), .ZN(n10022) );
  NOR2_X1 U11894 ( .A1(n11939), .A2(n15740), .ZN(n11970) );
  AND2_X1 U11895 ( .A1(n11919), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11934) );
  NOR2_X1 U11896 ( .A1(n11893), .A2(n20016), .ZN(n11919) );
  AOI21_X1 U11897 ( .B1(n11908), .B2(n12162), .A(n11907), .ZN(n14021) );
  AND3_X1 U11898 ( .A1(n11891), .A2(n11890), .A3(n11889), .ZN(n13973) );
  NAND2_X1 U11899 ( .A1(n11871), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11887) );
  NAND2_X1 U11900 ( .A1(n11876), .A2(n11875), .ZN(n13952) );
  INV_X1 U11901 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11857) );
  NOR2_X1 U11902 ( .A1(n11858), .A2(n11857), .ZN(n11871) );
  NAND2_X1 U11903 ( .A1(n11793), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11858) );
  NAND2_X1 U11904 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11803) );
  XNOR2_X1 U11905 ( .A(n12622), .B(n12621), .ZN(n13690) );
  NAND2_X1 U11906 ( .A1(n14481), .A2(n14470), .ZN(n14469) );
  OR2_X1 U11907 ( .A1(n14469), .A2(n14285), .ZN(n14453) );
  NAND2_X1 U11908 ( .A1(n14574), .A2(n9809), .ZN(n14561) );
  INV_X1 U11909 ( .A(n14559), .ZN(n9971) );
  NAND2_X1 U11910 ( .A1(n14574), .A2(n9972), .ZN(n14565) );
  NAND2_X1 U11911 ( .A1(n14574), .A2(n14573), .ZN(n14576) );
  AND2_X1 U11912 ( .A1(n9745), .A2(n9822), .ZN(n10003) );
  AND2_X1 U11913 ( .A1(n12700), .A2(n12701), .ZN(n9918) );
  AND2_X1 U11914 ( .A1(n14589), .A2(n14496), .ZN(n14574) );
  AND3_X1 U11915 ( .A1(n12352), .A2(n12351), .A3(n12350), .ZN(n14587) );
  NOR2_X1 U11916 ( .A1(n14588), .A2(n14587), .ZN(n14589) );
  NAND2_X1 U11917 ( .A1(n14600), .A2(n14599), .ZN(n14602) );
  OR2_X1 U11918 ( .A1(n14602), .A2(n14511), .ZN(n14588) );
  NAND2_X1 U11919 ( .A1(n9907), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12341) );
  NOR2_X1 U11920 ( .A1(n14540), .A2(n14525), .ZN(n14600) );
  NAND2_X1 U11921 ( .A1(n9967), .A2(n9966), .ZN(n14540) );
  INV_X1 U11922 ( .A(n14537), .ZN(n9966) );
  AND2_X1 U11923 ( .A1(n9712), .A2(n15898), .ZN(n15781) );
  NAND2_X1 U11924 ( .A1(n14182), .A2(n10014), .ZN(n15783) );
  NOR2_X1 U11925 ( .A1(n12691), .A2(n10015), .ZN(n10014) );
  INV_X1 U11926 ( .A(n15914), .ZN(n15685) );
  NOR2_X1 U11927 ( .A1(n14169), .A2(n14165), .ZN(n14164) );
  NOR2_X1 U11928 ( .A1(n12621), .A2(n20186), .ZN(n15948) );
  OR2_X1 U11929 ( .A1(n14175), .A2(n14167), .ZN(n14169) );
  AND2_X1 U11930 ( .A1(n12326), .A2(n12325), .ZN(n14176) );
  NAND2_X1 U11931 ( .A1(n9742), .A2(n14176), .ZN(n14175) );
  AND3_X1 U11933 ( .A1(n12317), .A2(n12351), .A3(n12316), .ZN(n14030) );
  NOR2_X1 U11934 ( .A1(n13893), .A2(n12308), .ZN(n13957) );
  NAND2_X1 U11935 ( .A1(n12295), .A2(n12294), .ZN(n13755) );
  INV_X1 U11936 ( .A(n13610), .ZN(n12294) );
  INV_X1 U11937 ( .A(n13611), .ZN(n12295) );
  OR2_X1 U11938 ( .A1(n13755), .A2(n13754), .ZN(n13893) );
  NOR2_X1 U11939 ( .A1(n20175), .A2(n15948), .ZN(n15939) );
  CLKBUF_X1 U11940 ( .A(n11832), .Z(n11833) );
  BUF_X1 U11941 ( .A(n11742), .Z(n13675) );
  INV_X1 U11942 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14831) );
  CLKBUF_X1 U11943 ( .A(n13647), .Z(n14834) );
  OR2_X1 U11944 ( .A1(n20192), .A2(n14824), .ZN(n20427) );
  INV_X1 U11945 ( .A(n20368), .ZN(n20627) );
  INV_X1 U11946 ( .A(n12600), .ZN(n20217) );
  AND2_X1 U11947 ( .A1(n9717), .A2(n20579), .ZN(n20657) );
  INV_X1 U11948 ( .A(n20704), .ZN(n20658) );
  AND2_X1 U11949 ( .A1(n9717), .A2(n20194), .ZN(n20548) );
  AOI21_X1 U11950 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20628), .A(n20342), 
        .ZN(n20705) );
  NAND3_X1 U11951 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20761), .A3(n20195), 
        .ZN(n20235) );
  NAND2_X1 U11952 ( .A1(n19968), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19967) );
  AND2_X1 U11953 ( .A1(n10980), .A2(n10979), .ZN(n11016) );
  OR2_X1 U11954 ( .A1(n10978), .A2(n10977), .ZN(n10980) );
  NAND2_X1 U11955 ( .A1(n12491), .A2(n12490), .ZN(n16023) );
  INV_X1 U11956 ( .A(n9882), .ZN(n12465) );
  NOR2_X1 U11957 ( .A1(n14853), .A2(n19069), .ZN(n15604) );
  NOR2_X1 U11958 ( .A1(n15604), .A2(n15605), .ZN(n15603) );
  NOR2_X1 U11959 ( .A1(n14865), .A2(n15099), .ZN(n14853) );
  NOR2_X1 U11960 ( .A1(n18895), .A2(n18897), .ZN(n14866) );
  AND2_X1 U11961 ( .A1(n9868), .A2(n9714), .ZN(n14865) );
  NAND2_X1 U11962 ( .A1(n14866), .A2(n15117), .ZN(n9868) );
  NAND2_X1 U11963 ( .A1(n18907), .A2(n18908), .ZN(n18895) );
  NOR2_X1 U11964 ( .A1(n18918), .A2(n18920), .ZN(n18907) );
  AND2_X1 U11965 ( .A1(n10939), .A2(n10938), .ZN(n18930) );
  NAND2_X1 U11966 ( .A1(n18957), .A2(n18962), .ZN(n18948) );
  NOR2_X1 U11967 ( .A1(n14069), .A2(n16163), .ZN(n18957) );
  NAND2_X1 U11968 ( .A1(n18971), .A2(n18972), .ZN(n14069) );
  NOR2_X1 U11969 ( .A1(n18982), .A2(n18984), .ZN(n18971) );
  NAND2_X1 U11970 ( .A1(n19016), .A2(n19017), .ZN(n19005) );
  NOR2_X1 U11971 ( .A1(n19024), .A2(n19025), .ZN(n19016) );
  NOR2_X1 U11972 ( .A1(n19050), .A2(n19052), .ZN(n19039) );
  AND2_X1 U11973 ( .A1(n12858), .A2(n13793), .ZN(n13877) );
  AND2_X1 U11974 ( .A1(n12857), .A2(n13804), .ZN(n13792) );
  INV_X1 U11975 ( .A(n11211), .ZN(n12572) );
  XNOR2_X1 U11976 ( .A(n13051), .B(n13052), .ZN(n14901) );
  XNOR2_X1 U11977 ( .A(n13027), .B(n13029), .ZN(n14911) );
  NAND2_X1 U11978 ( .A1(n14911), .A2(n14910), .ZN(n14909) );
  NAND2_X1 U11979 ( .A1(n14927), .A2(n10088), .ZN(n14915) );
  NAND2_X1 U11980 ( .A1(n9954), .A2(n9810), .ZN(n15219) );
  NAND2_X1 U11981 ( .A1(n9954), .A2(n9953), .ZN(n15217) );
  AND2_X1 U11982 ( .A1(n10054), .A2(n10053), .ZN(n10052) );
  INV_X1 U11983 ( .A(n14938), .ZN(n10053) );
  NAND2_X1 U11984 ( .A1(n14153), .A2(n10054), .ZN(n14937) );
  AND3_X1 U11985 ( .A1(n11309), .A2(n11308), .A3(n11307), .ZN(n15315) );
  CLKBUF_X1 U11986 ( .A(n14070), .Z(n15314) );
  INV_X1 U11987 ( .A(n19967), .ZN(n13398) );
  NOR2_X1 U11988 ( .A1(n13349), .A2(n13225), .ZN(n19231) );
  INV_X1 U11989 ( .A(n13157), .ZN(n16121) );
  NAND2_X1 U11990 ( .A1(n13175), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15047) );
  AND2_X1 U11992 ( .A1(n12529), .A2(n12528), .ZN(n14902) );
  NOR2_X2 U11993 ( .A1(n13181), .A2(n16085), .ZN(n13182) );
  NAND2_X1 U11994 ( .A1(n13186), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13184) );
  AND2_X1 U11995 ( .A1(n11178), .A2(n11177), .ZN(n12508) );
  NAND2_X1 U11996 ( .A1(n13945), .A2(n9980), .ZN(n14065) );
  NAND2_X1 U11997 ( .A1(n13192), .A2(n9793), .ZN(n13203) );
  AND2_X1 U11998 ( .A1(n11134), .A2(n11133), .ZN(n14008) );
  INV_X1 U11999 ( .A(n13191), .ZN(n13202) );
  NAND2_X1 U12000 ( .A1(n13945), .A2(n14341), .ZN(n14342) );
  NAND2_X1 U12001 ( .A1(n13201), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13200) );
  NAND2_X1 U12002 ( .A1(n9865), .A2(n9864), .ZN(n13196) );
  INV_X1 U12003 ( .A(n9867), .ZN(n9864) );
  INV_X1 U12004 ( .A(n11041), .ZN(n16230) );
  INV_X1 U12005 ( .A(n13159), .ZN(n9956) );
  INV_X1 U12006 ( .A(n14357), .ZN(n9888) );
  AND2_X1 U12007 ( .A1(n12591), .A2(n9819), .ZN(n12592) );
  OR3_X1 U12008 ( .A1(n16086), .A2(n12494), .A3(n14329), .ZN(n15063) );
  NAND2_X1 U12009 ( .A1(n12591), .A2(n12590), .ZN(n15089) );
  NOR2_X1 U12010 ( .A1(n12457), .A2(n12456), .ZN(n12458) );
  INV_X1 U12011 ( .A(n15202), .ZN(n9830) );
  OR2_X1 U12012 ( .A1(n14235), .A2(n12402), .ZN(n11169) );
  AND2_X1 U12013 ( .A1(n11154), .A2(n11153), .ZN(n14145) );
  NOR2_X1 U12014 ( .A1(n14146), .A2(n14145), .ZN(n14147) );
  NAND2_X1 U12015 ( .A1(n14070), .A2(n14071), .ZN(n16253) );
  OR3_X1 U12016 ( .A1(n18967), .A2(n12494), .A3(n15320), .ZN(n15310) );
  CLKBUF_X1 U12017 ( .A(n15308), .Z(n15329) );
  NAND2_X1 U12018 ( .A1(n16279), .A2(n9960), .ZN(n15334) );
  NOR2_X1 U12019 ( .A1(n16270), .A2(n15350), .ZN(n9857) );
  AND3_X1 U12020 ( .A1(n11280), .A2(n11279), .A3(n11278), .ZN(n16267) );
  NAND2_X1 U12021 ( .A1(n16279), .A2(n15352), .ZN(n16266) );
  NAND2_X1 U12022 ( .A1(n12591), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16190) );
  NOR2_X1 U12023 ( .A1(n16288), .A2(n16287), .ZN(n15351) );
  OR2_X1 U12024 ( .A1(n11102), .A2(n15350), .ZN(n11119) );
  NAND2_X1 U12025 ( .A1(n13786), .A2(n9983), .ZN(n13802) );
  AND2_X1 U12026 ( .A1(n19027), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15136) );
  NAND2_X1 U12027 ( .A1(n14096), .A2(n11231), .ZN(n15359) );
  NAND2_X1 U12028 ( .A1(n14089), .A2(n11064), .ZN(n11062) );
  INV_X1 U12029 ( .A(n14089), .ZN(n11060) );
  NAND2_X1 U12030 ( .A1(n16228), .A2(n11050), .ZN(n11054) );
  OAI21_X1 U12031 ( .B1(n11041), .B2(n12496), .A(n13713), .ZN(n16234) );
  NAND2_X1 U12032 ( .A1(n10623), .A2(n10606), .ZN(n9842) );
  INV_X1 U12033 ( .A(n10030), .ZN(n9843) );
  NAND2_X1 U12034 ( .A1(n10625), .A2(n10626), .ZN(n9854) );
  AND2_X1 U12035 ( .A1(n11184), .A2(n11077), .ZN(n13729) );
  NAND2_X1 U12036 ( .A1(n15245), .A2(n15249), .ZN(n15247) );
  NOR2_X1 U12037 ( .A1(n10549), .A2(n19969), .ZN(n13429) );
  NOR2_X1 U12038 ( .A1(n11196), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13431) );
  AOI21_X1 U12039 ( .B1(n13995), .B2(n12848), .A(n12832), .ZN(n13583) );
  NAND2_X1 U12040 ( .A1(n19323), .A2(n19945), .ZN(n19419) );
  NAND2_X1 U12041 ( .A1(n19929), .A2(n19917), .ZN(n19915) );
  OR2_X1 U12042 ( .A1(n19929), .A2(n19917), .ZN(n19676) );
  INV_X1 U12043 ( .A(n11084), .ZN(n19291) );
  NOR2_X2 U12044 ( .A1(n16122), .A2(n13983), .ZN(n19315) );
  OR2_X1 U12045 ( .A1(n19929), .A2(n19937), .ZN(n19505) );
  OR2_X1 U12046 ( .A1(n19323), .A2(n19945), .ZN(n19675) );
  INV_X1 U12047 ( .A(n19768), .ZN(n19357) );
  INV_X1 U12048 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19973) );
  NOR2_X1 U12049 ( .A1(n16843), .A2(n16580), .ZN(n16572) );
  NOR2_X1 U12050 ( .A1(n16591), .A2(n17505), .ZN(n16590) );
  NOR2_X1 U12051 ( .A1(n16620), .A2(n16843), .ZN(n16609) );
  NOR2_X1 U12052 ( .A1(n16609), .A2(n17540), .ZN(n16608) );
  NOR2_X1 U12053 ( .A1(n16629), .A2(n16843), .ZN(n16621) );
  NOR2_X1 U12054 ( .A1(n16621), .A2(n16622), .ZN(n16620) );
  NOR2_X1 U12055 ( .A1(n16652), .A2(n16843), .ZN(n16641) );
  NOR2_X1 U12056 ( .A1(n17591), .A2(n16641), .ZN(n16640) );
  NOR2_X1 U12057 ( .A1(n16662), .A2(n17620), .ZN(n16661) );
  OR2_X1 U12058 ( .A1(n10112), .A2(n18657), .ZN(n9761) );
  NOR2_X1 U12059 ( .A1(n18191), .A2(n18859), .ZN(n10221) );
  NAND2_X1 U12060 ( .A1(n17022), .A2(n9816), .ZN(n16981) );
  NOR2_X1 U12061 ( .A1(n9925), .A2(n16644), .ZN(n9923) );
  NOR2_X1 U12062 ( .A1(n17321), .A2(n16667), .ZN(n9924) );
  NAND2_X1 U12063 ( .A1(n17022), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n16998) );
  XOR2_X1 U12064 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n10093), .Z(
        n16791) );
  NOR2_X1 U12065 ( .A1(n10095), .A2(n16392), .ZN(n10094) );
  NAND2_X1 U12066 ( .A1(n17579), .A2(n9870), .ZN(n9869) );
  NOR2_X1 U12067 ( .A1(n9871), .A2(n17537), .ZN(n9870) );
  NOR3_X1 U12068 ( .A1(n10101), .A2(n17600), .A3(n9872), .ZN(n17549) );
  INV_X1 U12069 ( .A(n17549), .ZN(n10100) );
  OR2_X1 U12070 ( .A1(n18012), .A2(n18011), .ZN(n17565) );
  NOR3_X1 U12071 ( .A1(n16698), .A2(n17646), .A3(n16678), .ZN(n17588) );
  AND2_X1 U12072 ( .A1(n17655), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16699) );
  NAND2_X1 U12073 ( .A1(n16699), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16698) );
  INV_X1 U12074 ( .A(n16699), .ZN(n16710) );
  NAND3_X1 U12075 ( .A1(n17803), .A2(n9873), .A3(n10087), .ZN(n17679) );
  NOR2_X1 U12076 ( .A1(n18037), .A2(n17719), .ZN(n17696) );
  NOR2_X1 U12077 ( .A1(n17713), .A2(n17724), .ZN(n17708) );
  AND2_X1 U12078 ( .A1(n9873), .A2(n17803), .ZN(n17709) );
  NOR2_X1 U12079 ( .A1(n17754), .A2(n18092), .ZN(n17749) );
  INV_X1 U12080 ( .A(n16828), .ZN(n17803) );
  AOI22_X1 U12081 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U12082 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9725), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10197) );
  AOI211_X1 U12083 ( .C1(n17163), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n10194), .B(n10193), .ZN(n10195) );
  INV_X1 U12084 ( .A(n17833), .ZN(n16858) );
  AND2_X1 U12085 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17833) );
  OR2_X1 U12086 ( .A1(n15594), .A2(n9807), .ZN(n15595) );
  NAND2_X1 U12087 ( .A1(n15596), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17521) );
  NAND2_X1 U12088 ( .A1(n17622), .A2(n15591), .ZN(n17568) );
  NAND2_X1 U12089 ( .A1(n15590), .A2(n10086), .ZN(n15591) );
  NAND2_X1 U12090 ( .A1(n17665), .A2(n17912), .ZN(n15590) );
  INV_X1 U12091 ( .A(n17786), .ZN(n17610) );
  NAND2_X1 U12092 ( .A1(n17696), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18012) );
  INV_X1 U12093 ( .A(n18648), .ZN(n13250) );
  NOR2_X1 U12094 ( .A1(n17786), .A2(n15580), .ZN(n17754) );
  INV_X1 U12095 ( .A(n17747), .ZN(n18063) );
  NAND2_X1 U12096 ( .A1(n17808), .A2(n15545), .ZN(n17797) );
  INV_X1 U12097 ( .A(n9984), .ZN(n15543) );
  NAND2_X1 U12098 ( .A1(n17834), .A2(n15540), .ZN(n17820) );
  XNOR2_X1 U12099 ( .A(n15539), .B(n18139), .ZN(n17835) );
  NAND2_X1 U12100 ( .A1(n17835), .A2(n17836), .ZN(n17834) );
  XNOR2_X1 U12101 ( .A(n15559), .B(n13326), .ZN(n13327) );
  INV_X1 U12102 ( .A(n15560), .ZN(n13326) );
  NAND2_X1 U12103 ( .A1(n18858), .A2(n15396), .ZN(n18144) );
  XNOR2_X1 U12104 ( .A(n13303), .B(n13302), .ZN(n17852) );
  OR2_X1 U12105 ( .A1(n18647), .A2(n13247), .ZN(n13238) );
  NOR2_X1 U12106 ( .A1(n13313), .A2(n13312), .ZN(n17871) );
  NAND2_X2 U12107 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18657) );
  NAND2_X1 U12108 ( .A1(n10108), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14252) );
  INV_X1 U12109 ( .A(n10112), .ZN(n10108) );
  INV_X1 U12110 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18672) );
  NOR2_X1 U12111 ( .A1(n10135), .A2(n10134), .ZN(n18208) );
  NOR2_X1 U12112 ( .A1(n10165), .A2(n10164), .ZN(n18213) );
  INV_X1 U12113 ( .A(n18231), .ZN(n18487) );
  NOR2_X1 U12114 ( .A1(n10186), .A2(n10185), .ZN(n18199) );
  INV_X1 U12115 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18643) );
  NOR2_X1 U12116 ( .A1(n18700), .A2(n18862), .ZN(n18846) );
  NOR2_X1 U12117 ( .A1(n20091), .A2(n14414), .ZN(n20067) );
  OR2_X1 U12118 ( .A1(n20051), .A2(n13853), .ZN(n20104) );
  INV_X1 U12119 ( .A(n20081), .ZN(n20099) );
  INV_X1 U12120 ( .A(n20102), .ZN(n20088) );
  OR2_X1 U12121 ( .A1(n13865), .A2(n13859), .ZN(n20091) );
  OR3_X1 U12122 ( .A1(n13865), .A2(n13862), .A3(n13861), .ZN(n20024) );
  INV_X1 U12123 ( .A(n14612), .ZN(n14607) );
  INV_X1 U12124 ( .A(n15733), .ZN(n14665) );
  INV_X1 U12125 ( .A(n14218), .ZN(n14173) );
  NAND2_X1 U12126 ( .A1(n13454), .A2(n13460), .ZN(n12738) );
  OR2_X1 U12127 ( .A1(n14666), .A2(n13748), .ZN(n14218) );
  AND2_X1 U12128 ( .A1(n13618), .A2(n15638), .ZN(n20120) );
  OR2_X2 U12129 ( .A1(n19988), .A2(n13438), .ZN(n20152) );
  XNOR2_X1 U12130 ( .A(n13850), .B(n13849), .ZN(n14351) );
  NAND2_X1 U12131 ( .A1(n12207), .A2(n12710), .ZN(n14400) );
  AND2_X1 U12132 ( .A1(n12189), .A2(n12185), .ZN(n14460) );
  NAND2_X1 U12133 ( .A1(n14744), .A2(n12700), .ZN(n14736) );
  AND2_X1 U12134 ( .A1(n14586), .A2(n14585), .ZN(n15775) );
  AND2_X1 U12135 ( .A1(n12034), .A2(n12053), .ZN(n14769) );
  INV_X1 U12136 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14765) );
  NAND2_X1 U12137 ( .A1(n20158), .A2(n12712), .ZN(n15837) );
  OR3_X1 U12138 ( .A1(n12732), .A2(n15627), .A3(n19992), .ZN(n20158) );
  INV_X1 U12139 ( .A(n15837), .ZN(n20165) );
  XNOR2_X1 U12140 ( .A(n12784), .B(n12783), .ZN(n14546) );
  MUX2_X1 U12141 ( .A(n12782), .B(n13375), .S(n14406), .Z(n12784) );
  XNOR2_X1 U12142 ( .A(n9908), .B(n12760), .ZN(n14354) );
  XNOR2_X1 U12143 ( .A(n14703), .B(n14702), .ZN(n14809) );
  NAND2_X1 U12144 ( .A1(n10085), .A2(n14701), .ZN(n14703) );
  XNOR2_X1 U12145 ( .A(n14719), .B(n12813), .ZN(n15840) );
  OAI21_X1 U12146 ( .B1(n14731), .B2(n10080), .A(n9764), .ZN(n14719) );
  NAND2_X1 U12147 ( .A1(n15852), .A2(n9820), .ZN(n10007) );
  XNOR2_X1 U12148 ( .A(n10009), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15849) );
  AOI21_X1 U12149 ( .B1(n15761), .B2(n15760), .A(n10010), .ZN(n10009) );
  NOR2_X1 U12150 ( .A1(n15760), .A2(n10011), .ZN(n10010) );
  NOR2_X1 U12151 ( .A1(n15939), .A2(n15682), .ZN(n15875) );
  CLKBUF_X1 U12152 ( .A(n15820), .Z(n15823) );
  CLKBUF_X1 U12153 ( .A(n15826), .Z(n15827) );
  CLKBUF_X1 U12154 ( .A(n13886), .Z(n13887) );
  CLKBUF_X1 U12155 ( .A(n13822), .Z(n13823) );
  AND2_X1 U12156 ( .A1(n12807), .A2(n12787), .ZN(n15999) );
  CLKBUF_X1 U12157 ( .A(n13764), .Z(n13765) );
  INV_X1 U12158 ( .A(n15916), .ZN(n20175) );
  CLKBUF_X1 U12159 ( .A(n13587), .Z(n13588) );
  AND2_X1 U12160 ( .A1(n15916), .A2(n15966), .ZN(n13892) );
  OR2_X1 U12161 ( .A1(n12616), .A2(n12627), .ZN(n9915) );
  INV_X1 U12162 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20628) );
  CLKBUF_X1 U12163 ( .A(n12596), .Z(n20192) );
  CLKBUF_X1 U12164 ( .A(n13642), .Z(n13643) );
  INV_X1 U12165 ( .A(n20636), .ZN(n20698) );
  AND2_X1 U12166 ( .A1(n12723), .A2(n12804), .ZN(n15612) );
  NOR2_X1 U12167 ( .A1(n15646), .A2(n20593), .ZN(n14840) );
  NOR2_X1 U12168 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16008) );
  OAI21_X1 U12169 ( .B1(n20276), .B2(n20275), .A(n20274), .ZN(n20293) );
  AND2_X1 U12170 ( .A1(n20270), .A2(n20627), .ZN(n20292) );
  OAI21_X1 U12171 ( .B1(n20359), .B2(n20343), .A(n20666), .ZN(n20361) );
  NOR2_X2 U12172 ( .A1(n20427), .A2(n20368), .ZN(n20414) );
  NOR2_X2 U12173 ( .A1(n20427), .A2(n20426), .ZN(n20483) );
  INV_X1 U12174 ( .A(n20515), .ZN(n20482) );
  INV_X1 U12175 ( .A(n20527), .ZN(n20544) );
  AND2_X1 U12176 ( .A1(n20553), .A2(n20657), .ZN(n20575) );
  OAI211_X1 U12177 ( .C1(n20619), .C2(n20593), .A(n20666), .B(n20592), .ZN(
        n20622) );
  OAI211_X1 U12178 ( .C1(n20691), .C2(n20667), .A(n20666), .B(n20665), .ZN(
        n20693) );
  INV_X1 U12179 ( .A(n20600), .ZN(n20711) );
  INV_X1 U12180 ( .A(n20758), .ZN(n20732) );
  INV_X1 U12181 ( .A(n20735), .ZN(n20754) );
  NAND2_X1 U12182 ( .A1(n20658), .A2(n20548), .ZN(n20758) );
  INV_X1 U12183 ( .A(n20625), .ZN(n20750) );
  INV_X1 U12184 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20761) );
  NOR2_X1 U12185 ( .A1(n16053), .A2(n16054), .ZN(n16052) );
  INV_X1 U12186 ( .A(n12491), .ZN(n12486) );
  NOR2_X1 U12187 ( .A1(n9852), .A2(n19069), .ZN(n13209) );
  NOR2_X1 U12188 ( .A1(n13209), .A2(n13210), .ZN(n16029) );
  NOR2_X1 U12189 ( .A1(n16106), .A2(n19069), .ZN(n16098) );
  NOR2_X1 U12190 ( .A1(n16107), .A2(n16108), .ZN(n16106) );
  INV_X1 U12191 ( .A(n19086), .ZN(n19063) );
  AND2_X1 U12192 ( .A1(n18870), .A2(n16369), .ZN(n19019) );
  NAND2_X1 U12193 ( .A1(n19039), .A2(n19040), .ZN(n19024) );
  INV_X1 U12194 ( .A(n19034), .ZN(n19081) );
  INV_X1 U12195 ( .A(n9707), .ZN(n19079) );
  OR2_X1 U12196 ( .A1(n13222), .A2(n14897), .ZN(n16068) );
  OR2_X1 U12197 ( .A1(n11331), .A2(n11330), .ZN(n14017) );
  OR2_X1 U12198 ( .A1(n11305), .A2(n11304), .ZN(n14345) );
  AND2_X1 U12199 ( .A1(n13738), .A2(n12859), .ZN(n14346) );
  OR2_X1 U12200 ( .A1(n11290), .A2(n11289), .ZN(n13943) );
  INV_X1 U12201 ( .A(n14926), .ZN(n14939) );
  OAI21_X1 U12202 ( .B1(n13598), .B2(n13599), .A(n13600), .ZN(n19323) );
  AND2_X1 U12203 ( .A1(n14887), .A2(n10045), .ZN(n14895) );
  INV_X1 U12204 ( .A(n19105), .ZN(n14999) );
  AND2_X1 U12205 ( .A1(n19132), .A2(n13147), .ZN(n19105) );
  NOR2_X1 U12206 ( .A1(n19146), .A2(n19158), .ZN(n19142) );
  INV_X1 U12207 ( .A(n19162), .ZN(n19146) );
  INV_X1 U12208 ( .A(n16124), .ZN(n19158) );
  INV_X1 U12209 ( .A(n19134), .ZN(n19166) );
  AND2_X1 U12210 ( .A1(n13397), .A2(n19970), .ZN(n19203) );
  NOR2_X2 U12211 ( .A1(n19203), .A2(n13399), .ZN(n19211) );
  OR2_X1 U12212 ( .A1(n19231), .A2(n19245), .ZN(n13444) );
  NAND2_X1 U12213 ( .A1(n14303), .A2(n14878), .ZN(n16058) );
  INV_X1 U12214 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18941) );
  OAI21_X1 U12215 ( .B1(n15202), .B2(n10923), .A(n15296), .ZN(n16158) );
  INV_X1 U12216 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16225) );
  NAND2_X1 U12217 ( .A1(n10033), .A2(n10032), .ZN(n14086) );
  INV_X1 U12218 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16240) );
  NAND2_X1 U12219 ( .A1(n18875), .A2(n12403), .ZN(n16239) );
  AND2_X1 U12220 ( .A1(n16239), .A2(n13360), .ZN(n16227) );
  INV_X1 U12221 ( .A(n16239), .ZN(n19258) );
  NAND2_X1 U12222 ( .A1(n15037), .A2(n16274), .ZN(n9948) );
  NAND2_X1 U12223 ( .A1(n15045), .A2(n10035), .ZN(n14371) );
  OR2_X1 U12224 ( .A1(n13221), .A2(n13224), .ZN(n14890) );
  AND2_X1 U12225 ( .A1(n15184), .A2(n12583), .ZN(n15167) );
  NAND2_X1 U12226 ( .A1(n10068), .A2(n9750), .ZN(n15273) );
  NAND2_X1 U12227 ( .A1(n10065), .A2(n10064), .ZN(n16186) );
  INV_X1 U12228 ( .A(n19917), .ZN(n19937) );
  INV_X1 U12229 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19933) );
  INV_X1 U12230 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19926) );
  INV_X1 U12231 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16336) );
  NAND2_X1 U12232 ( .A1(n19094), .A2(n12848), .ZN(n12834) );
  XNOR2_X1 U12233 ( .A(n13699), .B(n13700), .ZN(n19929) );
  INV_X1 U12234 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16358) );
  NOR2_X1 U12235 ( .A1(n19506), .A2(n19676), .ZN(n19486) );
  OR2_X1 U12236 ( .A1(n19500), .A2(n19499), .ZN(n19527) );
  INV_X1 U12237 ( .A(n19561), .ZN(n19553) );
  NOR2_X1 U12238 ( .A1(n19675), .A2(n19562), .ZN(n19614) );
  INV_X1 U12239 ( .A(n19773), .ZN(n19715) );
  INV_X1 U12240 ( .A(n19785), .ZN(n19732) );
  INV_X1 U12241 ( .A(n19808), .ZN(n19746) );
  OAI21_X1 U12242 ( .B1(n19726), .B2(n19725), .A(n19724), .ZN(n19753) );
  INV_X1 U12243 ( .A(n19745), .ZN(n19751) );
  INV_X1 U12244 ( .A(n19729), .ZN(n19770) );
  INV_X1 U12245 ( .A(n19692), .ZN(n19776) );
  INV_X1 U12246 ( .A(n19735), .ZN(n19782) );
  INV_X1 U12247 ( .A(n19739), .ZN(n19788) );
  INV_X1 U12248 ( .A(n19704), .ZN(n19799) );
  NOR2_X2 U12249 ( .A1(n19675), .A2(n19505), .ZN(n19814) );
  INV_X1 U12250 ( .A(n19757), .ZN(n19813) );
  AND2_X1 U12251 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11038), .ZN(n16367) );
  AND2_X1 U12252 ( .A1(n10994), .A2(n10993), .ZN(n19956) );
  INV_X1 U12253 ( .A(n19055), .ZN(n19825) );
  OAI21_X1 U12254 ( .B1(n18632), .B2(n18631), .A(n17453), .ZN(n18859) );
  NOR2_X1 U12255 ( .A1(n16554), .A2(n18697), .ZN(n17453) );
  NOR2_X1 U12256 ( .A1(n16573), .A2(n16572), .ZN(n16571) );
  NOR2_X1 U12257 ( .A1(n16590), .A2(n16843), .ZN(n16581) );
  NOR2_X1 U12258 ( .A1(n16581), .A2(n16582), .ZN(n16580) );
  NOR2_X1 U12259 ( .A1(n16608), .A2(n16843), .ZN(n16600) );
  AND2_X1 U12260 ( .A1(n10218), .A2(n16888), .ZN(n16617) );
  NOR2_X1 U12261 ( .A1(n13341), .A2(n16843), .ZN(n16630) );
  NOR2_X1 U12262 ( .A1(n17559), .A2(n16630), .ZN(n16629) );
  NOR2_X1 U12263 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16643), .ZN(n16634) );
  NOR2_X1 U12264 ( .A1(n16640), .A2(n16843), .ZN(n13342) );
  NOR2_X1 U12265 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16666), .ZN(n16651) );
  AND2_X1 U12266 ( .A1(n9875), .A2(n17604), .ZN(n16652) );
  INV_X1 U12267 ( .A(n9875), .ZN(n16653) );
  INV_X1 U12268 ( .A(n16902), .ZN(n16888) );
  INV_X1 U12269 ( .A(n16898), .ZN(n16891) );
  INV_X1 U12270 ( .A(n16914), .ZN(n16894) );
  NOR2_X2 U12271 ( .A1(n16894), .A2(n18803), .ZN(n16898) );
  INV_X1 U12272 ( .A(n16871), .ZN(n16910) );
  NOR2_X1 U12273 ( .A1(n16925), .A2(n16924), .ZN(n16950) );
  NOR3_X1 U12274 ( .A1(n16981), .A2(n16919), .A3(n16975), .ZN(n16980) );
  NOR2_X1 U12275 ( .A1(n17038), .A2(n17035), .ZN(n17022) );
  NAND3_X1 U12276 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(n17079), .ZN(n17035) );
  NOR2_X1 U12277 ( .A1(n17039), .A2(n17092), .ZN(n17079) );
  NOR2_X1 U12278 ( .A1(n17095), .A2(n9927), .ZN(n17093) );
  NAND2_X1 U12279 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .ZN(n9927) );
  NAND2_X1 U12280 ( .A1(n17093), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n17092) );
  NAND2_X1 U12281 ( .A1(n17142), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n17095) );
  NAND2_X1 U12282 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17154), .ZN(n17139) );
  INV_X1 U12283 ( .A(n17170), .ZN(n17154) );
  NAND2_X1 U12284 ( .A1(n17171), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n17170) );
  AND2_X1 U12285 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17206), .ZN(n17202) );
  INV_X1 U12286 ( .A(n17209), .ZN(n17206) );
  NOR2_X1 U12287 ( .A1(n17227), .A2(n17215), .ZN(n17210) );
  NAND2_X1 U12288 ( .A1(n17210), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n17209) );
  NOR2_X1 U12289 ( .A1(n17394), .A2(n17259), .ZN(n17255) );
  NAND2_X1 U12290 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17263), .ZN(n17259) );
  NOR2_X1 U12291 ( .A1(n17408), .A2(n17294), .ZN(n17288) );
  NOR2_X1 U12292 ( .A1(n15506), .A2(n15505), .ZN(n17356) );
  INV_X1 U12293 ( .A(n17317), .ZN(n17363) );
  INV_X1 U12294 ( .A(n17378), .ZN(n17375) );
  NOR2_X1 U12295 ( .A1(n9990), .A2(n9988), .ZN(n9987) );
  INV_X1 U12296 ( .A(n13300), .ZN(n9990) );
  NOR2_X1 U12297 ( .A1(n17363), .A2(n18667), .ZN(n17378) );
  INV_X1 U12298 ( .A(n17372), .ZN(n17377) );
  INV_X1 U12299 ( .A(n17451), .ZN(n17440) );
  NOR2_X1 U12300 ( .A1(n17449), .A2(n17440), .ZN(n17446) );
  INV_X1 U12301 ( .A(n17442), .ZN(n17448) );
  BUF_X1 U12302 ( .A(n17469), .Z(n17499) );
  NOR2_X1 U12303 ( .A1(n18850), .A2(n17499), .ZN(n17500) );
  NOR2_X1 U12304 ( .A1(n17679), .A2(n17671), .ZN(n17655) );
  INV_X1 U12305 ( .A(n18037), .ZN(n17717) );
  NOR2_X1 U12306 ( .A1(n17794), .A2(n16816), .ZN(n17781) );
  NOR2_X1 U12307 ( .A1(n16401), .A2(n17876), .ZN(n17788) );
  INV_X1 U12308 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17794) );
  AND2_X1 U12309 ( .A1(n17833), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17814) );
  INV_X1 U12310 ( .A(n18221), .ZN(n18577) );
  INV_X1 U12311 ( .A(n16400), .ZN(n17876) );
  INV_X1 U12312 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18862) );
  INV_X1 U12313 ( .A(n18080), .ZN(n18096) );
  NOR2_X1 U12314 ( .A1(n18639), .A2(n16401), .ZN(n18099) );
  INV_X1 U12315 ( .A(n18144), .ZN(n18664) );
  INV_X1 U12316 ( .A(n18633), .ZN(n18153) );
  NAND2_X1 U12317 ( .A1(n18648), .A2(n13238), .ZN(n18658) );
  CLKBUF_X1 U12318 ( .A(n13328), .Z(n18162) );
  INV_X1 U12319 ( .A(n18133), .ZN(n18164) );
  INV_X1 U12320 ( .A(n18658), .ZN(n18668) );
  INV_X1 U12321 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18677) );
  INV_X1 U12322 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18680) );
  INV_X1 U12323 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18803) );
  CLKBUF_X1 U12324 ( .A(n18795), .Z(n18786) );
  OAI21_X1 U12326 ( .B1(n14784), .B2(n14612), .A(n12389), .ZN(n12390) );
  OAI211_X1 U12327 ( .C1(n14354), .C2(n15988), .A(n9964), .B(n9963), .ZN(
        P1_U3000) );
  NOR2_X1 U12328 ( .A1(n12818), .A2(n9965), .ZN(n9964) );
  NAND2_X1 U12329 ( .A1(n14546), .A2(n15999), .ZN(n9963) );
  INV_X1 U12330 ( .A(n12823), .ZN(n9965) );
  INV_X1 U12331 ( .A(n10005), .ZN(P1_U3007) );
  AOI211_X1 U12332 ( .C1(n15849), .C2(n20182), .A(n10008), .B(n10006), .ZN(
        n10005) );
  NOR2_X1 U12333 ( .A1(n15853), .A2(n20179), .ZN(n10008) );
  OR2_X1 U12334 ( .A1(n15848), .A2(n10007), .ZN(n10006) );
  INV_X1 U12335 ( .A(n16036), .ZN(n16044) );
  NAND2_X1 U12336 ( .A1(n9841), .A2(n14314), .ZN(n9840) );
  OAI21_X1 U12337 ( .B1(n12431), .B2(n16219), .A(n12414), .ZN(n12415) );
  NAND2_X1 U12338 ( .A1(n14315), .A2(n16274), .ZN(n12594) );
  OAI21_X1 U12339 ( .B1(n15039), .B2(n16315), .A(n9942), .ZN(P2_U3016) );
  AOI21_X1 U12340 ( .B1(n16281), .B2(n16041), .A(n9943), .ZN(n9942) );
  NAND2_X1 U12341 ( .A1(n9948), .A2(n9944), .ZN(n9943) );
  INV_X1 U12342 ( .A(n9945), .ZN(n9944) );
  NAND2_X1 U12343 ( .A1(n9829), .A2(n15225), .ZN(P2_U3024) );
  NAND2_X1 U12344 ( .A1(n16138), .A2(n16301), .ZN(n9829) );
  INV_X1 U12345 ( .A(n11371), .ZN(n11372) );
  INV_X1 U12346 ( .A(n12432), .ZN(n12433) );
  OAI21_X1 U12347 ( .B1(n12431), .B2(n16307), .A(n12430), .ZN(n12432) );
  NOR2_X1 U12348 ( .A1(n9921), .A2(n9803), .ZN(n9920) );
  NOR2_X1 U12349 ( .A1(n16971), .A2(n17228), .ZN(n16963) );
  INV_X1 U12350 ( .A(n17171), .ZN(n17195) );
  OAI211_X1 U12351 ( .C1(n16439), .C2(n18080), .A(n9992), .B(n9991), .ZN(
        P3_U2831) );
  AOI21_X1 U12352 ( .B1(n16438), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n16437), .ZN(n9991) );
  NAND2_X1 U12353 ( .A1(n9993), .A2(n18169), .ZN(n9992) );
  CLKBUF_X1 U12354 ( .A(n13274), .Z(n17173) );
  INV_X1 U12355 ( .A(n11619), .ZN(n20234) );
  OR2_X2 U12356 ( .A1(n11521), .A2(n11520), .ZN(n11619) );
  AND3_X1 U12357 ( .A1(n13957), .A2(n9746), .A3(n14053), .ZN(n9742) );
  INV_X1 U12358 ( .A(n13277), .ZN(n17176) );
  NAND2_X1 U12359 ( .A1(n14182), .A2(n12685), .ZN(n14183) );
  INV_X1 U12360 ( .A(n12592), .ZN(n14331) );
  AND2_X1 U12361 ( .A1(n9962), .A2(n12801), .ZN(n9743) );
  AND2_X1 U12362 ( .A1(n10024), .A2(n9802), .ZN(n14128) );
  NOR2_X1 U12363 ( .A1(n15874), .A2(n14751), .ZN(n9745) );
  XNOR2_X1 U12364 ( .A(n12549), .B(n12548), .ZN(n16033) );
  INV_X1 U12365 ( .A(n16033), .ZN(n9974) );
  OR2_X1 U12366 ( .A1(n10115), .A2(n16903), .ZN(n13299) );
  NOR2_X1 U12367 ( .A1(n16063), .A2(n16064), .ZN(n9852) );
  NAND2_X2 U12368 ( .A1(n9854), .A2(n10623), .ZN(n12824) );
  INV_X1 U12369 ( .A(n12824), .ZN(n9853) );
  AND2_X1 U12370 ( .A1(n9762), .A2(n9968), .ZN(n9746) );
  AND3_X1 U12371 ( .A1(n11078), .A2(n9940), .A3(n11019), .ZN(n9747) );
  AND2_X1 U12372 ( .A1(n9983), .A2(n11120), .ZN(n9748) );
  AND2_X1 U12373 ( .A1(n14355), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9749) );
  INV_X1 U12374 ( .A(n10824), .ZN(n10844) );
  NAND2_X1 U12375 ( .A1(n13183), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13181) );
  NAND2_X1 U12376 ( .A1(n13190), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13188) );
  AND2_X1 U12377 ( .A1(n13945), .A2(n9787), .ZN(n14009) );
  AND2_X1 U12378 ( .A1(n16279), .A2(n9785), .ZN(n15333) );
  AND2_X1 U12379 ( .A1(n16156), .A2(n10071), .ZN(n9750) );
  OAI21_X1 U12380 ( .B1(n20193), .B2(n11982), .A(n11810), .ZN(n13752) );
  AND2_X1 U12381 ( .A1(n12436), .A2(n15296), .ZN(n9751) );
  AND2_X1 U12382 ( .A1(n9751), .A2(n10072), .ZN(n9752) );
  OR2_X1 U12383 ( .A1(n15326), .A2(n10916), .ZN(n12441) );
  INV_X1 U12384 ( .A(n10664), .ZN(n13727) );
  INV_X2 U12385 ( .A(n13727), .ZN(n10665) );
  NOR2_X1 U12386 ( .A1(n13177), .A2(n15056), .ZN(n13175) );
  AND2_X1 U12387 ( .A1(n9861), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9753) );
  AND2_X1 U12388 ( .A1(n12442), .A2(n9815), .ZN(n9754) );
  NAND2_X2 U12389 ( .A1(n13147), .A2(n13431), .ZN(n11211) );
  NAND2_X1 U12390 ( .A1(n10594), .A2(n10578), .ZN(n9755) );
  INV_X1 U12391 ( .A(n12283), .ZN(n12329) );
  NAND2_X1 U12392 ( .A1(n14237), .A2(n14151), .ZN(n12510) );
  INV_X1 U12393 ( .A(n9949), .ZN(n11235) );
  AND2_X1 U12394 ( .A1(n14995), .A2(n9950), .ZN(n14966) );
  INV_X1 U12395 ( .A(n9711), .ZN(n10011) );
  NAND2_X1 U12396 ( .A1(n14467), .A2(n14468), .ZN(n14290) );
  NOR2_X1 U12397 ( .A1(n14556), .A2(n14557), .ZN(n14478) );
  NAND2_X1 U12398 ( .A1(n20217), .A2(n13854), .ZN(n12296) );
  AND3_X1 U12399 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13194) );
  NAND2_X1 U12400 ( .A1(n14467), .A2(n10025), .ZN(n12207) );
  OR2_X1 U12401 ( .A1(n9733), .A2(n13712), .ZN(n9758) );
  AND2_X1 U12402 ( .A1(n12592), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9759) );
  OR2_X1 U12403 ( .A1(n11631), .A2(n20221), .ZN(n9760) );
  NOR2_X1 U12404 ( .A1(n10110), .A2(n10114), .ZN(n13293) );
  AND2_X1 U12405 ( .A1(n12315), .A2(n9969), .ZN(n9762) );
  AND2_X1 U12406 ( .A1(n14519), .A2(n14523), .ZN(n14521) );
  OR3_X1 U12407 ( .A1(n15760), .A2(n15762), .A3(n10011), .ZN(n9764) );
  AND4_X1 U12408 ( .A1(n13297), .A2(n13296), .A3(n13295), .A4(n13294), .ZN(
        n9765) );
  AND2_X1 U12409 ( .A1(n11527), .A2(n11526), .ZN(n9766) );
  OR2_X1 U12410 ( .A1(n14049), .A2(n14172), .ZN(n9767) );
  AND2_X1 U12411 ( .A1(n13054), .A2(n10047), .ZN(n9768) );
  NAND2_X1 U12412 ( .A1(n10065), .A2(n10896), .ZN(n15346) );
  NAND2_X1 U12413 ( .A1(n10046), .A2(n13073), .ZN(n14887) );
  NOR3_X1 U12414 ( .A1(n16039), .A2(n12494), .A3(n12576), .ZN(n9769) );
  NAND2_X1 U12415 ( .A1(n10881), .A2(n10880), .ZN(n15135) );
  NAND2_X1 U12416 ( .A1(n10004), .A2(n9712), .ZN(n15767) );
  NOR2_X1 U12417 ( .A1(n10621), .A2(n10620), .ZN(n9770) );
  OR2_X1 U12418 ( .A1(n11784), .A2(n11783), .ZN(n9771) );
  AND2_X1 U12419 ( .A1(n9748), .A2(n13881), .ZN(n9772) );
  AND2_X1 U12420 ( .A1(n10880), .A2(n10886), .ZN(n9773) );
  INV_X1 U12421 ( .A(n12685), .ZN(n10015) );
  NAND2_X1 U12422 ( .A1(n13989), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9774) );
  NOR2_X1 U12423 ( .A1(n15219), .A2(n15004), .ZN(n14995) );
  AND2_X1 U12424 ( .A1(n12698), .A2(n10001), .ZN(n9775) );
  INV_X1 U12425 ( .A(n10607), .ZN(n11102) );
  AND2_X1 U12426 ( .A1(n14915), .A2(n13001), .ZN(n9776) );
  AND2_X1 U12427 ( .A1(n9755), .A2(n19094), .ZN(n9777) );
  OR2_X1 U12428 ( .A1(n14318), .A2(n12476), .ZN(n9778) );
  AND2_X1 U12429 ( .A1(n14904), .A2(n14896), .ZN(n13222) );
  NAND2_X1 U12430 ( .A1(n14995), .A2(n14996), .ZN(n14322) );
  NAND2_X1 U12431 ( .A1(n10504), .A2(n10503), .ZN(n10579) );
  INV_X1 U12432 ( .A(n12778), .ZN(n15627) );
  NAND2_X1 U12433 ( .A1(n14909), .A2(n13031), .ZN(n13051) );
  NAND2_X1 U12434 ( .A1(n14521), .A2(n10029), .ZN(n14563) );
  NOR2_X1 U12435 ( .A1(n14282), .A2(n14693), .ZN(n9779) );
  NAND2_X1 U12436 ( .A1(n10547), .A2(n10549), .ZN(n10555) );
  INV_X1 U12437 ( .A(n10555), .ZN(n9848) );
  XNOR2_X1 U12438 ( .A(n11065), .B(n11061), .ZN(n11056) );
  AND2_X1 U12439 ( .A1(n12592), .A2(n10037), .ZN(n15053) );
  INV_X1 U12440 ( .A(n15053), .ZN(n10036) );
  AND2_X1 U12441 ( .A1(n15063), .A2(n12489), .ZN(n14355) );
  XNOR2_X1 U12442 ( .A(n11823), .B(n11704), .ZN(n13683) );
  NOR2_X1 U12443 ( .A1(n9879), .A2(n10844), .ZN(n10883) );
  NOR2_X1 U12444 ( .A1(n13203), .A2(n18941), .ZN(n13190) );
  NOR2_X1 U12445 ( .A1(n13200), .A2(n18978), .ZN(n13192) );
  AND2_X1 U12446 ( .A1(n17022), .A2(n9924), .ZN(n9780) );
  AND2_X1 U12447 ( .A1(n10027), .A2(n14468), .ZN(n9781) );
  NAND2_X1 U12448 ( .A1(n14153), .A2(n14154), .ZN(n14155) );
  NAND2_X1 U12449 ( .A1(n10024), .A2(n10023), .ZN(n14127) );
  NOR2_X1 U12450 ( .A1(n13951), .A2(n10020), .ZN(n14022) );
  NOR2_X1 U12451 ( .A1(n13946), .A2(n13947), .ZN(n13945) );
  AND2_X1 U12452 ( .A1(n13786), .A2(n9748), .ZN(n13796) );
  NAND2_X1 U12453 ( .A1(n13609), .A2(n11841), .ZN(n13751) );
  AND4_X1 U12454 ( .A1(n12454), .A2(n15259), .A3(n12453), .A4(n12452), .ZN(
        n9782) );
  AND2_X1 U12455 ( .A1(n14237), .A2(n9977), .ZN(n9783) );
  NAND2_X1 U12456 ( .A1(n9740), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10101) );
  AND4_X1 U12457 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16436), .A3(
        n16435), .A4(n18808), .ZN(n9784) );
  AND2_X1 U12458 ( .A1(n13198), .A2(n12409), .ZN(n13193) );
  NOR2_X1 U12459 ( .A1(n16253), .A2(n16254), .ZN(n15280) );
  AND2_X1 U12460 ( .A1(n9961), .A2(n15352), .ZN(n9785) );
  OR2_X1 U12461 ( .A1(n10084), .A2(n10906), .ZN(n9786) );
  AND2_X1 U12462 ( .A1(n9981), .A2(n14341), .ZN(n9787) );
  NOR2_X1 U12463 ( .A1(n16097), .A2(n19069), .ZN(n16082) );
  AND2_X1 U12464 ( .A1(n13172), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13185) );
  NOR2_X2 U12465 ( .A1(n11084), .A2(n11078), .ZN(n11077) );
  INV_X1 U12466 ( .A(n11077), .ZN(n10051) );
  NOR2_X1 U12467 ( .A1(n16098), .A2(n16099), .ZN(n16097) );
  AND2_X1 U12468 ( .A1(n9781), .A2(n10026), .ZN(n9788) );
  OR2_X1 U12469 ( .A1(n9940), .A2(n10931), .ZN(n9789) );
  AND2_X1 U12470 ( .A1(n12859), .A2(n14345), .ZN(n9790) );
  OR2_X1 U12471 ( .A1(n10898), .A2(n9891), .ZN(n9791) );
  AND2_X1 U12472 ( .A1(n9980), .A2(n9979), .ZN(n9792) );
  AND2_X1 U12473 ( .A1(n12411), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9793) );
  NAND2_X1 U12474 ( .A1(n10017), .A2(n11892), .ZN(n13971) );
  XOR2_X1 U12475 ( .A(n13989), .B(n15992), .Z(n9794) );
  INV_X1 U12476 ( .A(n12441), .ZN(n10072) );
  INV_X2 U12477 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19969) );
  OR2_X1 U12478 ( .A1(n10066), .A2(n10069), .ZN(n9795) );
  OR2_X1 U12479 ( .A1(n12849), .A2(n12848), .ZN(n9796) );
  NOR2_X1 U12480 ( .A1(n10830), .A2(n10844), .ZN(n9797) );
  AND2_X1 U12481 ( .A1(n11050), .A2(n14094), .ZN(n9798) );
  AND2_X1 U12482 ( .A1(n9960), .A2(n9959), .ZN(n9799) );
  AND2_X1 U12483 ( .A1(n13173), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9800) );
  AND2_X1 U12484 ( .A1(n9976), .A2(n9975), .ZN(n9801) );
  INV_X1 U12485 ( .A(n11200), .ZN(n11350) );
  AND2_X1 U12486 ( .A1(n11189), .A2(n19955), .ZN(n16301) );
  INV_X1 U12487 ( .A(n9853), .ZN(n15387) );
  NOR2_X1 U12488 ( .A1(n13184), .A2(n13174), .ZN(n13183) );
  AND2_X1 U12489 ( .A1(n14159), .A2(n14160), .ZN(n9802) );
  AND2_X1 U12490 ( .A1(n17228), .A2(n17249), .ZN(n9803) );
  AND2_X1 U12491 ( .A1(n13787), .A2(n13788), .ZN(n13786) );
  AND2_X1 U12492 ( .A1(n13957), .A2(n9746), .ZN(n9804) );
  OR3_X1 U12493 ( .A1(n10101), .A2(n17600), .A3(n9871), .ZN(n9805) );
  INV_X1 U12494 ( .A(n19263), .ZN(n16214) );
  AND2_X1 U12495 ( .A1(n16239), .A2(n19936), .ZN(n19263) );
  AND2_X1 U12496 ( .A1(n14996), .A2(n9952), .ZN(n9806) );
  AND2_X1 U12497 ( .A1(n13786), .A2(n13817), .ZN(n13800) );
  AND2_X1 U12498 ( .A1(n17786), .A2(n15593), .ZN(n9807) );
  AND2_X2 U12499 ( .A1(n13125), .A2(n10470), .ZN(n12898) );
  OR2_X1 U12500 ( .A1(n19269), .A2(n18962), .ZN(n9808) );
  AND2_X1 U12501 ( .A1(n9972), .A2(n9971), .ZN(n9809) );
  AND2_X1 U12502 ( .A1(n9953), .A2(n15216), .ZN(n9810) );
  INV_X1 U12503 ( .A(n9967), .ZN(n14538) );
  NOR2_X1 U12504 ( .A1(n14198), .A2(n14199), .ZN(n9967) );
  NAND2_X1 U12505 ( .A1(n13738), .A2(n9790), .ZN(n14344) );
  OR2_X1 U12506 ( .A1(n10747), .A2(n10746), .ZN(n10821) );
  OR2_X1 U12507 ( .A1(n17225), .A2(n9922), .ZN(n9811) );
  AND2_X1 U12508 ( .A1(n13175), .A2(n9861), .ZN(n9812) );
  AND2_X1 U12509 ( .A1(n9982), .A2(n14304), .ZN(n9813) );
  AND2_X1 U12510 ( .A1(n17803), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9814) );
  INV_X1 U12511 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n9892) );
  XNOR2_X1 U12512 ( .A(n12290), .B(n13547), .ZN(n13590) );
  INV_X1 U12513 ( .A(n14048), .ZN(n10019) );
  OR2_X1 U12514 ( .A1(n9940), .A2(n12513), .ZN(n9815) );
  AND2_X1 U12515 ( .A1(n9924), .A2(n9923), .ZN(n9816) );
  AND2_X1 U12516 ( .A1(n9915), .A2(n12615), .ZN(n9817) );
  AND2_X1 U12517 ( .A1(n9957), .A2(n9956), .ZN(n9818) );
  AND2_X1 U12518 ( .A1(n10034), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9819) );
  INV_X1 U12519 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9862) );
  OR2_X1 U12520 ( .A1(n20177), .A2(n20824), .ZN(n9820) );
  NOR2_X2 U12521 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15378) );
  OR2_X1 U12522 ( .A1(n14695), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9821) );
  AND2_X1 U12523 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9822) );
  INV_X1 U12524 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9855) );
  INV_X1 U12525 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10038) );
  INV_X1 U12526 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9874) );
  INV_X1 U12527 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n9925) );
  INV_X1 U12528 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n9847) );
  NOR3_X2 U12529 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9706), .A3(
        n18316), .ZN(n18246) );
  NOR3_X2 U12530 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n9706), .A3(
        n18407), .ZN(n18379) );
  NOR3_X2 U12531 ( .A1(n9706), .A2(n18672), .A3(n18316), .ZN(n18288) );
  NOR3_X2 U12532 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9706), .A3(
        n18363), .ZN(n18334) );
  AOI22_X2 U12533 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19314), .ZN(n19779) );
  NOR2_X2 U12534 ( .A1(n16121), .A2(n13983), .ZN(n19314) );
  NOR3_X2 U12535 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9706), .A3(
        n18457), .ZN(n18425) );
  NOR2_X2 U12536 ( .A1(n18222), .A2(n18221), .ZN(n18622) );
  NAND2_X1 U12537 ( .A1(n10579), .A2(n10568), .ZN(n9824) );
  NAND2_X1 U12538 ( .A1(n9823), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U12539 ( .A1(n9825), .A2(n9824), .ZN(n9823) );
  AND2_X2 U12540 ( .A1(n9855), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10442) );
  XNOR2_X1 U12541 ( .A(n15202), .B(n15298), .ZN(n16164) );
  NOR2_X2 U12542 ( .A1(n10627), .A2(n9770), .ZN(n19094) );
  INV_X1 U12543 ( .A(n11052), .ZN(n9831) );
  INV_X1 U12544 ( .A(n10828), .ZN(n10057) );
  NAND2_X2 U12545 ( .A1(n9832), .A2(n10059), .ZN(n15308) );
  NOR2_X2 U12546 ( .A1(n10639), .A2(n10640), .ZN(n10749) );
  AND2_X2 U12547 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9834) );
  INV_X2 U12548 ( .A(n9833), .ZN(n10664) );
  NAND2_X1 U12549 ( .A1(n9834), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9833) );
  NOR2_X1 U12550 ( .A1(n9834), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15381) );
  NAND2_X1 U12551 ( .A1(n10756), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n9835) );
  NAND3_X1 U12552 ( .A1(n10686), .A2(n10685), .A3(n9837), .ZN(n10737) );
  NAND3_X1 U12553 ( .A1(n12846), .A2(n9849), .A3(n10622), .ZN(n10651) );
  NAND2_X2 U12554 ( .A1(n9843), .A2(n9842), .ZN(n9849) );
  NAND2_X1 U12555 ( .A1(n16230), .A2(n16229), .ZN(n16228) );
  NAND2_X1 U12556 ( .A1(n9844), .A2(n11222), .ZN(n11051) );
  NOR2_X1 U12557 ( .A1(n10650), .A2(n10648), .ZN(n14109) );
  NAND2_X1 U12558 ( .A1(n19723), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9845) );
  NOR2_X1 U12559 ( .A1(n10648), .A2(n9847), .ZN(n9846) );
  INV_X1 U12560 ( .A(n19723), .ZN(n19720) );
  NAND2_X1 U12561 ( .A1(n16228), .A2(n9798), .ZN(n10032) );
  INV_X1 U12562 ( .A(n11054), .ZN(n14039) );
  NAND2_X2 U12563 ( .A1(n9859), .A2(n9860), .ZN(n10549) );
  NAND2_X4 U12564 ( .A1(n9849), .A2(n12846), .ZN(n10640) );
  NAND3_X1 U12565 ( .A1(n9849), .A2(n12846), .A3(n12847), .ZN(n10041) );
  XNOR2_X1 U12566 ( .A(n15044), .B(n12576), .ZN(n15037) );
  NAND2_X1 U12567 ( .A1(n15131), .A2(n11066), .ZN(n9850) );
  NAND2_X1 U12568 ( .A1(n9851), .A2(n11063), .ZN(n15131) );
  NAND2_X1 U12569 ( .A1(n11057), .A2(n11056), .ZN(n11063) );
  OAI21_X1 U12570 ( .B1(n10039), .B2(n11059), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U12571 ( .A1(n16204), .A2(n16202), .ZN(n9858) );
  NAND3_X1 U12572 ( .A1(n16161), .A2(n16162), .A3(n9808), .ZN(P2_U3000) );
  INV_X1 U12573 ( .A(n13195), .ZN(n9865) );
  NOR2_X1 U12574 ( .A1(n9867), .A2(n16225), .ZN(n9866) );
  NOR2_X1 U12575 ( .A1(n10101), .A2(n17600), .ZN(n17578) );
  INV_X1 U12576 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9872) );
  NAND4_X1 U12577 ( .A1(n10824), .A2(n9877), .A3(n10887), .A4(n9876), .ZN(
        n10890) );
  INV_X1 U12578 ( .A(n10825), .ZN(n9880) );
  NAND2_X1 U12579 ( .A1(n12443), .A2(n12442), .ZN(n12463) );
  NAND2_X2 U12580 ( .A1(n12445), .A2(n12473), .ZN(n12443) );
  NAND2_X1 U12581 ( .A1(n9935), .A2(n9934), .ZN(n9886) );
  NAND2_X1 U12582 ( .A1(n9778), .A2(n9888), .ZN(n9887) );
  NAND3_X1 U12583 ( .A1(n9887), .A2(n14355), .A3(n9886), .ZN(n15055) );
  NAND2_X1 U12584 ( .A1(n12277), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9905) );
  NAND3_X1 U12585 ( .A1(n9909), .A2(n12759), .A3(n12758), .ZN(n9908) );
  NAND2_X2 U12586 ( .A1(n12705), .A2(n14682), .ZN(n12757) );
  OAI21_X1 U12587 ( .B1(n9914), .B2(n14080), .A(n9911), .ZN(n9912) );
  NAND2_X1 U12588 ( .A1(n9912), .A2(n10011), .ZN(n12697) );
  NAND2_X2 U12589 ( .A1(n14080), .A2(n12684), .ZN(n14182) );
  NAND2_X2 U12590 ( .A1(n9744), .A2(n14800), .ZN(n14681) );
  NOR2_X2 U12591 ( .A1(n14692), .A2(n9821), .ZN(n14709) );
  XNOR2_X1 U12592 ( .A(n12680), .B(n9794), .ZN(n15987) );
  AND2_X2 U12593 ( .A1(n12669), .A2(n12668), .ZN(n12680) );
  NAND2_X1 U12594 ( .A1(n9917), .A2(n9916), .ZN(n13544) );
  NAND2_X1 U12595 ( .A1(n14744), .A2(n9918), .ZN(n12702) );
  AND2_X2 U12596 ( .A1(n17201), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17171) );
  NAND2_X2 U12597 ( .A1(n18817), .A2(n18807), .ZN(n10113) );
  INV_X2 U12598 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18807) );
  NOR2_X1 U12599 ( .A1(n16960), .A2(n16593), .ZN(n9921) );
  NOR2_X2 U12600 ( .A1(n16966), .A2(n16956), .ZN(n16971) );
  OAI21_X1 U12601 ( .B1(n15468), .B2(P3_EBX_REG_28__SCAN_IN), .A(n9920), .ZN(
        P3_U2675) );
  AND2_X1 U12602 ( .A1(n17223), .A2(n16955), .ZN(n9922) );
  NOR2_X2 U12603 ( .A1(n17139), .A2(n17138), .ZN(n17142) );
  NAND3_X1 U12604 ( .A1(n10661), .A2(n10662), .A3(n10660), .ZN(n9929) );
  AND2_X1 U12605 ( .A1(n9937), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9932) );
  NAND3_X1 U12606 ( .A1(n9935), .A2(n9934), .A3(n14358), .ZN(n9933) );
  INV_X1 U12607 ( .A(n12476), .ZN(n9936) );
  NOR2_X1 U12608 ( .A1(n12476), .A2(n15173), .ZN(n9937) );
  NAND2_X2 U12609 ( .A1(n10624), .A2(n10605), .ZN(n10623) );
  NAND2_X4 U12610 ( .A1(n10463), .A2(n10464), .ZN(n9940) );
  NOR2_X1 U12611 ( .A1(n9940), .A2(n14149), .ZN(n10942) );
  NOR2_X1 U12612 ( .A1(n9940), .A2(n11165), .ZN(n10952) );
  NOR2_X1 U12613 ( .A1(n9940), .A2(n11159), .ZN(n10956) );
  NOR2_X1 U12614 ( .A1(n9940), .A2(n11172), .ZN(n10958) );
  NOR2_X1 U12615 ( .A1(n9940), .A2(n14945), .ZN(n12444) );
  NAND2_X1 U12616 ( .A1(n10549), .A2(n9940), .ZN(n10501) );
  INV_X4 U12617 ( .A(n9940), .ZN(n19300) );
  NAND2_X1 U12618 ( .A1(n13431), .A2(n9940), .ZN(n11346) );
  XNOR2_X1 U12619 ( .A(n10549), .B(n9940), .ZN(n11029) );
  NAND2_X1 U12620 ( .A1(n12496), .A2(n9940), .ZN(n9949) );
  INV_X1 U12621 ( .A(n9941), .ZN(n13537) );
  NOR2_X1 U12622 ( .A1(n14264), .A2(n11361), .ZN(n14864) );
  INV_X1 U12623 ( .A(n11364), .ZN(n9955) );
  NAND2_X1 U12624 ( .A1(n13227), .A2(n9957), .ZN(n14952) );
  NAND2_X1 U12625 ( .A1(n13227), .A2(n13228), .ZN(n13226) );
  NAND2_X1 U12626 ( .A1(n9970), .A2(n12290), .ZN(n13611) );
  NAND2_X1 U12627 ( .A1(n14237), .A2(n9801), .ZN(n14920) );
  INV_X1 U12628 ( .A(n14064), .ZN(n9979) );
  NAND2_X1 U12629 ( .A1(n13222), .A2(n9982), .ZN(n14303) );
  NAND2_X1 U12630 ( .A1(n13222), .A2(n9813), .ZN(n12549) );
  AND2_X1 U12631 ( .A1(n13222), .A2(n13223), .ZN(n13221) );
  NAND3_X1 U12632 ( .A1(n13298), .A2(n13301), .A3(n9989), .ZN(n9988) );
  INV_X2 U12633 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18831) );
  NAND4_X1 U12634 ( .A1(n11626), .A2(n11625), .A3(n9999), .A4(n11624), .ZN(
        n12277) );
  INV_X1 U12635 ( .A(n12798), .ZN(n9999) );
  NAND2_X1 U12636 ( .A1(n12796), .A2(n13857), .ZN(n12798) );
  AND2_X2 U12637 ( .A1(n13673), .A2(n11391), .ZN(n11589) );
  NAND2_X1 U12638 ( .A1(n12698), .A2(n10002), .ZN(n10004) );
  NOR2_X2 U12639 ( .A1(n12691), .A2(n10013), .ZN(n10012) );
  NAND2_X1 U12640 ( .A1(n10016), .A2(n11994), .ZN(n11876) );
  AOI21_X1 U12641 ( .B1(n10016), .B2(n12670), .A(n12665), .ZN(n15821) );
  INV_X1 U12642 ( .A(n13951), .ZN(n10017) );
  NAND2_X1 U12643 ( .A1(n10017), .A2(n10018), .ZN(n14049) );
  NAND2_X1 U12644 ( .A1(n10024), .A2(n10022), .ZN(n14195) );
  NAND2_X1 U12645 ( .A1(n14521), .A2(n10028), .ZN(n14556) );
  NOR2_X2 U12646 ( .A1(n10648), .A2(n10649), .ZN(n19723) );
  NAND2_X2 U12647 ( .A1(n10640), .A2(n10622), .ZN(n10648) );
  NAND3_X2 U12648 ( .A1(n10030), .A2(n10606), .A3(n10623), .ZN(n12846) );
  NAND2_X1 U12649 ( .A1(n14090), .A2(n11060), .ZN(n11057) );
  INV_X1 U12650 ( .A(n10031), .ZN(n14087) );
  AND2_X1 U12651 ( .A1(n12591), .A2(n10034), .ZN(n14328) );
  NAND2_X1 U12652 ( .A1(n10036), .A2(n12575), .ZN(n10035) );
  INV_X1 U12653 ( .A(n11062), .ZN(n10039) );
  NAND2_X1 U12654 ( .A1(n10040), .A2(n11062), .ZN(n15145) );
  NAND2_X1 U12655 ( .A1(n11063), .A2(n11059), .ZN(n10040) );
  NAND2_X1 U12656 ( .A1(n14899), .A2(n13054), .ZN(n10046) );
  NAND3_X1 U12657 ( .A1(n14887), .A2(n14894), .A3(n10045), .ZN(n14893) );
  INV_X1 U12658 ( .A(n13073), .ZN(n10047) );
  INV_X1 U12659 ( .A(n14344), .ZN(n12861) );
  AND2_X1 U12660 ( .A1(n10055), .A2(n11077), .ZN(n11089) );
  AOI21_X1 U12661 ( .B1(n10579), .B2(n10055), .A(n10580), .ZN(n10588) );
  INV_X1 U12662 ( .A(n11201), .ZN(n13146) );
  INV_X1 U12663 ( .A(n10827), .ZN(n10058) );
  OAI21_X1 U12664 ( .B1(n15308), .B2(n12441), .A(n12455), .ZN(n15202) );
  OR2_X1 U12665 ( .A1(n14121), .A2(n12402), .ZN(n14236) );
  NAND2_X1 U12666 ( .A1(n11802), .A2(n11801), .ZN(n20193) );
  NAND2_X1 U12667 ( .A1(n14090), .A2(n11058), .ZN(n11059) );
  NAND2_X1 U12668 ( .A1(n12680), .A2(n9774), .ZN(n12683) );
  NAND2_X1 U12669 ( .A1(n15767), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12703) );
  AOI211_X2 U12670 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15160), .A(
        n14366), .B(n14365), .ZN(n14367) );
  CLKBUF_X1 U12671 ( .A(n15134), .Z(n16206) );
  XNOR2_X1 U12672 ( .A(n14262), .B(n10089), .ZN(n14278) );
  NAND2_X1 U12673 ( .A1(n14259), .A2(n14258), .ZN(n14262) );
  OR2_X1 U12674 ( .A1(n14442), .A2(n12709), .ZN(n12710) );
  INV_X1 U12675 ( .A(n13814), .ZN(n11843) );
  OR2_X1 U12676 ( .A1(n18875), .A2(n19283), .ZN(n16220) );
  NAND2_X1 U12677 ( .A1(n10553), .A2(n19968), .ZN(n13211) );
  NAND2_X1 U12678 ( .A1(n9720), .A2(n11938), .ZN(n14142) );
  AND2_X1 U12679 ( .A1(n13130), .A2(n10470), .ZN(n10722) );
  INV_X1 U12680 ( .A(n10695), .ZN(n19352) );
  INV_X1 U12681 ( .A(n11864), .ZN(n11867) );
  NOR2_X1 U12682 ( .A1(n20519), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10073) );
  AND2_X1 U12683 ( .A1(n12147), .A2(n12146), .ZN(n10074) );
  INV_X1 U12684 ( .A(n12198), .ZN(n12162) );
  NAND2_X1 U12685 ( .A1(n11189), .A2(n11183), .ZN(n16283) );
  AND3_X1 U12686 ( .A1(n14306), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14099), .ZN(n10076) );
  AND2_X2 U12687 ( .A1(n13436), .A2(n16367), .ZN(n14936) );
  INV_X1 U12688 ( .A(n14936), .ZN(n14907) );
  NOR2_X1 U12689 ( .A1(n12449), .A2(n12448), .ZN(n10077) );
  AND2_X1 U12690 ( .A1(n15103), .A2(n16274), .ZN(n10078) );
  NOR2_X1 U12691 ( .A1(n12586), .A2(n10076), .ZN(n10079) );
  INV_X1 U12692 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20016) );
  OR2_X1 U12693 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10080) );
  AND3_X1 U12694 ( .A1(n19283), .A2(n19305), .A3(n19300), .ZN(n10081) );
  OR3_X1 U12695 ( .A1(n13005), .A2(n13004), .A3(n14919), .ZN(n10082) );
  OR2_X1 U12696 ( .A1(n14400), .A2(n20191), .ZN(n10083) );
  NOR3_X1 U12697 ( .A1(n10904), .A2(n12494), .A3(n16270), .ZN(n10084) );
  NAND2_X1 U12698 ( .A1(n17712), .A2(n17872), .ZN(n17618) );
  OR2_X1 U12699 ( .A1(n14700), .A2(n14696), .ZN(n10085) );
  OR3_X1 U12700 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17593), .ZN(n10086) );
  AND2_X1 U12701 ( .A1(n17708), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10087) );
  INV_X1 U12702 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12760) );
  INV_X1 U12703 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12756) );
  INV_X1 U12704 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13174) );
  AND2_X1 U12705 ( .A1(n12711), .A2(n20636), .ZN(n15799) );
  INV_X1 U12706 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11816) );
  INV_X1 U12707 ( .A(n14006), .ZN(n12860) );
  NAND2_X1 U12708 ( .A1(n12980), .A2(n13002), .ZN(n10088) );
  AND2_X1 U12709 ( .A1(n14261), .A2(n14260), .ZN(n10089) );
  AND4_X1 U12710 ( .A1(n11541), .A2(n11540), .A3(n11539), .A4(n11538), .ZN(
        n10090) );
  INV_X1 U12711 ( .A(n12329), .ZN(n13375) );
  AND4_X1 U12712 ( .A1(n11546), .A2(n11545), .A3(n11544), .A4(n11543), .ZN(
        n10091) );
  AOI22_X1 U12713 ( .A1(n10608), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10566) );
  OR2_X1 U12714 ( .A1(n12228), .A2(n12227), .ZN(n12230) );
  NOR2_X1 U12715 ( .A1(n10610), .A2(n13701), .ZN(n10598) );
  NOR2_X1 U12716 ( .A1(n19963), .A2(n10581), .ZN(n10582) );
  INV_X1 U12717 ( .A(n10688), .ZN(n10692) );
  NOR2_X1 U12718 ( .A1(n11191), .A2(n19969), .ZN(n10564) );
  INV_X1 U12719 ( .A(n11746), .ZN(n11747) );
  AND2_X1 U12720 ( .A1(n12223), .A2(n12222), .ZN(n12225) );
  OR2_X1 U12721 ( .A1(n11853), .A2(n11852), .ZN(n12662) );
  NAND2_X1 U12722 ( .A1(n9782), .A2(n12455), .ZN(n12456) );
  AND3_X1 U12723 ( .A1(n10693), .A2(n10692), .A3(n10691), .ZN(n10699) );
  NAND2_X1 U12724 ( .A1(n10567), .A2(n19291), .ZN(n10503) );
  AND2_X1 U12725 ( .A1(n19950), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10833) );
  NOR2_X1 U12726 ( .A1(n10214), .A2(n10213), .ZN(n10207) );
  NAND2_X1 U12727 ( .A1(n20221), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12671) );
  OR2_X1 U12728 ( .A1(n11781), .A2(n11780), .ZN(n12653) );
  OR2_X1 U12729 ( .A1(n11654), .A2(n11653), .ZN(n12613) );
  INV_X1 U12730 ( .A(n13211), .ZN(n10565) );
  INV_X1 U12731 ( .A(n13052), .ZN(n13053) );
  INV_X1 U12732 ( .A(n12479), .ZN(n12480) );
  INV_X1 U12733 ( .A(n16185), .ZN(n10906) );
  AND2_X1 U12734 ( .A1(n11536), .A2(n13854), .ZN(n11746) );
  INV_X1 U12735 ( .A(n13973), .ZN(n11892) );
  AND2_X1 U12736 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n11377), .ZN(
        n12171) );
  NAND2_X1 U12737 ( .A1(n11531), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12195) );
  INV_X1 U12738 ( .A(n14141), .ZN(n11938) );
  NOR2_X1 U12739 ( .A1(n11735), .A2(n11734), .ZN(n12599) );
  INV_X1 U12740 ( .A(n10560), .ZN(n11023) );
  AND2_X1 U12741 ( .A1(n11077), .A2(n10568), .ZN(n10569) );
  INV_X1 U12742 ( .A(n13028), .ZN(n13029) );
  INV_X1 U12743 ( .A(n14916), .ZN(n13001) );
  OR2_X1 U12744 ( .A1(n14861), .A2(n14263), .ZN(n11361) );
  OR2_X1 U12745 ( .A1(n10734), .A2(n10733), .ZN(n10802) );
  INV_X1 U12746 ( .A(n14017), .ZN(n12862) );
  OR2_X1 U12747 ( .A1(n10978), .A2(n10979), .ZN(n10976) );
  INV_X1 U12748 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15438) );
  INV_X1 U12749 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17127) );
  INV_X1 U12750 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15584) );
  INV_X1 U12751 ( .A(n11964), .ZN(n11376) );
  INV_X1 U12752 ( .A(n11629), .ZN(n12278) );
  AND2_X1 U12753 ( .A1(n20764), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12718) );
  AND2_X1 U12754 ( .A1(n11380), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13848) );
  NAND2_X1 U12755 ( .A1(n12171), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12184) );
  OR2_X1 U12756 ( .A1(n14583), .A2(n14507), .ZN(n14492) );
  AND2_X1 U12757 ( .A1(n12057), .A2(n12056), .ZN(n14596) );
  NOR2_X1 U12758 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13843) );
  INV_X1 U12759 ( .A(n11887), .ZN(n11375) );
  AOI21_X1 U12760 ( .B1(n12651), .B2(n11994), .A(n11863), .ZN(n13874) );
  INV_X1 U12761 ( .A(n13843), .ZN(n12198) );
  NAND2_X1 U12762 ( .A1(n12702), .A2(n10011), .ZN(n15768) );
  OR2_X1 U12763 ( .A1(n12373), .A2(n12301), .ZN(n12351) );
  INV_X1 U12764 ( .A(n15612), .ZN(n13666) );
  NAND2_X1 U12765 ( .A1(n11745), .A2(n11744), .ZN(n20336) );
  INV_X1 U12766 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12247) );
  INV_X1 U12767 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20587) );
  AND2_X1 U12768 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12829) );
  OR2_X1 U12769 ( .A1(n11355), .A2(n15026), .ZN(n11356) );
  OR2_X1 U12770 ( .A1(n10781), .A2(n10780), .ZN(n11226) );
  AND2_X1 U12771 ( .A1(n11146), .A2(n11145), .ZN(n14064) );
  INV_X1 U12772 ( .A(n10802), .ZN(n11210) );
  OR2_X1 U12773 ( .A1(n18922), .A2(n12494), .ZN(n10948) );
  AND2_X1 U12774 ( .A1(n10925), .A2(n10930), .ZN(n18955) );
  OR2_X1 U12775 ( .A1(n16299), .A2(n11098), .ZN(n15349) );
  INV_X1 U12776 ( .A(n12496), .ZN(n12494) );
  NOR2_X1 U12777 ( .A1(n18831), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13256) );
  NAND2_X1 U12778 ( .A1(n17520), .A2(n15597), .ZN(n15664) );
  OAI211_X1 U12779 ( .C1(n15585), .C2(n15584), .A(n15588), .B(n15583), .ZN(
        n15586) );
  NAND2_X1 U12780 ( .A1(n17791), .A2(n15572), .ZN(n15580) );
  NOR2_X1 U12781 ( .A1(n12272), .A2(n12729), .ZN(n12273) );
  INV_X1 U12782 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15740) );
  NAND2_X1 U12783 ( .A1(n11376), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11939) );
  INV_X1 U12784 ( .A(n13860), .ZN(n12214) );
  AND2_X1 U12785 ( .A1(n14351), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U12786 ( .A1(n13847), .A2(n13846), .ZN(n14458) );
  NAND2_X1 U12787 ( .A1(n13451), .A2(n12735), .ZN(n13454) );
  NOR2_X1 U12788 ( .A1(n12094), .A2(n12087), .ZN(n12058) );
  NAND2_X1 U12789 ( .A1(n12033), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12135) );
  NAND2_X1 U12790 ( .A1(n11375), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11893) );
  AND2_X2 U12791 ( .A1(n11617), .A2(n12209), .ZN(n12778) );
  NAND2_X1 U12792 ( .A1(n12757), .A2(n12756), .ZN(n12759) );
  AOI21_X1 U12793 ( .B1(n14700), .B2(n14699), .A(n14698), .ZN(n14701) );
  AND3_X1 U12794 ( .A1(n12340), .A2(n12351), .A3(n12339), .ZN(n14537) );
  AND3_X1 U12795 ( .A1(n12328), .A2(n12351), .A3(n12327), .ZN(n14167) );
  NAND2_X1 U12796 ( .A1(n12807), .A2(n13646), .ZN(n15916) );
  INV_X1 U12797 ( .A(n20270), .ZN(n20307) );
  INV_X1 U12798 ( .A(n20548), .ZN(n20426) );
  INV_X1 U12799 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20549) );
  INV_X1 U12800 ( .A(n12276), .ZN(n15640) );
  OR2_X1 U12801 ( .A1(n11092), .A2(n11091), .ZN(n16343) );
  OR2_X1 U12802 ( .A1(n18870), .A2(n13216), .ZN(n19034) );
  AND2_X1 U12803 ( .A1(n12518), .A2(n12517), .ZN(n14922) );
  AND2_X1 U12804 ( .A1(n13943), .A2(n13877), .ZN(n12859) );
  AND3_X1 U12805 ( .A1(n11225), .A2(n11224), .A3(n11223), .ZN(n14041) );
  NOR2_X1 U12806 ( .A1(n13220), .A2(n12494), .ZN(n14358) );
  AND2_X1 U12807 ( .A1(n16155), .A2(n15271), .ZN(n12436) );
  OR2_X1 U12808 ( .A1(n14078), .A2(n10922), .ZN(n15296) );
  NAND2_X1 U12809 ( .A1(n11096), .A2(n15253), .ZN(n14099) );
  OR2_X1 U12810 ( .A1(n12398), .A2(n11037), .ZN(n11039) );
  XNOR2_X1 U12811 ( .A(n13534), .B(n11205), .ZN(n13906) );
  INV_X1 U12812 ( .A(n19945), .ZN(n14106) );
  NAND2_X1 U12813 ( .A1(n19929), .A2(n19937), .ZN(n19562) );
  OR2_X1 U12814 ( .A1(n19323), .A2(n14106), .ZN(n19713) );
  NOR2_X1 U12815 ( .A1(n18850), .A2(n17387), .ZN(n13236) );
  NOR2_X1 U12816 ( .A1(n16599), .A2(n16843), .ZN(n16591) );
  NOR2_X1 U12817 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16713), .ZN(n16703) );
  NOR2_X1 U12818 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16741), .ZN(n16724) );
  NOR2_X1 U12819 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16854), .ZN(n16847) );
  AOI211_X1 U12820 ( .C1(n17116), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n10152), .B(n10151), .ZN(n10153) );
  AOI211_X1 U12821 ( .C1(n10107), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n10121), .B(n10120), .ZN(n10122) );
  AOI21_X1 U12822 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(n16554) );
  INV_X1 U12823 ( .A(n17788), .ZN(n17748) );
  NOR2_X1 U12824 ( .A1(n17533), .A2(n15595), .ZN(n15596) );
  NAND2_X1 U12825 ( .A1(n15555), .A2(n15554), .ZN(n16447) );
  NOR2_X1 U12826 ( .A1(n18658), .A2(n18666), .ZN(n18145) );
  INV_X1 U12827 ( .A(n18099), .ZN(n18039) );
  AND2_X1 U12828 ( .A1(n15580), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17784) );
  INV_X1 U12829 ( .A(n15571), .ZN(n15569) );
  NAND2_X1 U12830 ( .A1(n13327), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15561) );
  INV_X1 U12831 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13302) );
  NAND2_X1 U12832 ( .A1(n18487), .A2(n18543), .ZN(n18221) );
  AOI21_X2 U12833 ( .B1(n12275), .B2(n12274), .A(n12273), .ZN(n15646) );
  AND2_X1 U12834 ( .A1(n14458), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20092) );
  AND2_X1 U12835 ( .A1(n11794), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11793) );
  INV_X1 U12836 ( .A(n20060), .ZN(n15737) );
  INV_X1 U12837 ( .A(n14673), .ZN(n14667) );
  OR2_X1 U12838 ( .A1(n12736), .A2(n13644), .ZN(n12737) );
  INV_X1 U12839 ( .A(n13475), .ZN(n13524) );
  NAND2_X1 U12840 ( .A1(n12058), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12145) );
  AND2_X1 U12841 ( .A1(n14598), .A2(n14597), .ZN(n15733) );
  NAND2_X1 U12842 ( .A1(n11934), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11964) );
  NAND2_X1 U12843 ( .A1(n12683), .A2(n12682), .ZN(n14080) );
  AND2_X1 U12844 ( .A1(n15837), .A2(n20164), .ZN(n15809) );
  INV_X1 U12845 ( .A(n20158), .ZN(n20167) );
  INV_X1 U12846 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14702) );
  NOR2_X1 U12847 ( .A1(n15863), .A2(n15862), .ZN(n15846) );
  AND2_X1 U12848 ( .A1(n12807), .A2(n15612), .ZN(n15928) );
  INV_X1 U12849 ( .A(n13892), .ZN(n15985) );
  INV_X1 U12850 ( .A(n15988), .ZN(n20182) );
  NAND2_X1 U12851 ( .A1(n20761), .A2(n20195), .ZN(n20342) );
  INV_X1 U12852 ( .A(n14840), .ZN(n14848) );
  AND2_X1 U12853 ( .A1(n20193), .A2(n20192), .ZN(n20270) );
  AND2_X1 U12854 ( .A1(n20270), .A2(n20657), .ZN(n20330) );
  NOR2_X2 U12855 ( .A1(n20307), .A2(n20426), .ZN(n20360) );
  INV_X1 U12856 ( .A(n20447), .ZN(n20415) );
  INV_X1 U12857 ( .A(n20427), .ZN(n20389) );
  NOR2_X1 U12858 ( .A1(n9717), .A2(n20194), .ZN(n20448) );
  AND2_X1 U12859 ( .A1(n20553), .A2(n20627), .ZN(n20543) );
  NOR2_X1 U12860 ( .A1(n20193), .A2(n12597), .ZN(n20553) );
  INV_X1 U12861 ( .A(n20594), .ZN(n20621) );
  AND2_X1 U12862 ( .A1(n20580), .A2(n20579), .ZN(n20653) );
  INV_X1 U12863 ( .A(n20662), .ZN(n20692) );
  INV_X1 U12864 ( .A(n20597), .ZN(n20700) );
  INV_X1 U12865 ( .A(n20607), .ZN(n20723) );
  INV_X1 U12866 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20760) );
  INV_X1 U12867 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20772) );
  AND2_X1 U12868 ( .A1(n13219), .A2(n13218), .ZN(n19086) );
  AND2_X1 U12869 ( .A1(n19231), .A2(n19914), .ZN(n19093) );
  AND2_X1 U12870 ( .A1(n14015), .A2(n14063), .ZN(n14207) );
  OR2_X1 U12871 ( .A1(n11250), .A2(n11249), .ZN(n13808) );
  AND2_X1 U12872 ( .A1(n14862), .A2(n14265), .ZN(n18902) );
  INV_X1 U12873 ( .A(n19132), .ZN(n19157) );
  INV_X1 U12874 ( .A(n13449), .ZN(n19245) );
  NOR2_X1 U12875 ( .A1(n13349), .A2(n11191), .ZN(n19229) );
  INV_X1 U12876 ( .A(n15222), .ZN(n16137) );
  AND2_X1 U12877 ( .A1(n14011), .A2(n14010), .ZN(n16167) );
  INV_X1 U12878 ( .A(n16219), .ZN(n19260) );
  AND2_X1 U12879 ( .A1(n12437), .A2(n12451), .ZN(n15122) );
  INV_X1 U12880 ( .A(n15319), .ZN(n16260) );
  AND2_X1 U12881 ( .A1(n11097), .A2(n14099), .ZN(n16299) );
  AND2_X1 U12882 ( .A1(n11039), .A2(n16367), .ZN(n11189) );
  XNOR2_X1 U12883 ( .A(n13584), .B(n13583), .ZN(n19917) );
  OAI21_X1 U12884 ( .B1(n19279), .B2(n19278), .A(n19277), .ZN(n19316) );
  OR2_X1 U12885 ( .A1(n19358), .A2(n19357), .ZN(n19376) );
  INV_X1 U12886 ( .A(n19410), .ZN(n19402) );
  INV_X1 U12887 ( .A(n19445), .ZN(n19437) );
  NOR2_X1 U12888 ( .A1(n19419), .A2(n19676), .ZN(n19470) );
  AND2_X1 U12889 ( .A1(n19504), .A2(n19503), .ZN(n19526) );
  INV_X1 U12890 ( .A(n19603), .ZN(n19620) );
  NOR2_X1 U12891 ( .A1(n19713), .A2(n19915), .ZN(n19619) );
  INV_X1 U12892 ( .A(n19818), .ZN(n19742) );
  INV_X1 U12893 ( .A(n19700), .ZN(n19794) );
  INV_X1 U12894 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19852) );
  AOI21_X1 U12895 ( .B1(n13260), .B2(n13259), .A(n13258), .ZN(n18635) );
  NOR2_X1 U12896 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16619), .ZN(n16618) );
  NAND2_X1 U12897 ( .A1(n10221), .A2(n18689), .ZN(n16902) );
  NOR2_X1 U12898 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16691), .ZN(n16682) );
  NOR2_X1 U12899 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16764), .ZN(n16749) );
  NOR2_X1 U12900 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n16787), .ZN(n16768) );
  NOR2_X1 U12901 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16812), .ZN(n16794) );
  NOR2_X1 U12902 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16833), .ZN(n16818) );
  INV_X1 U12903 ( .A(n16911), .ZN(n16906) );
  NOR2_X1 U12904 ( .A1(n17472), .A2(n17250), .ZN(n17243) );
  NAND2_X1 U12905 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17269), .ZN(n17268) );
  NAND2_X1 U12906 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17316), .ZN(n17312) );
  NAND2_X1 U12907 ( .A1(n17231), .A2(n17321), .ZN(n17369) );
  NAND3_X1 U12908 ( .A1(n10124), .A2(n10123), .A3(n10122), .ZN(n17387) );
  INV_X1 U12909 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18810) );
  OAI211_X1 U12910 ( .C1(n18850), .C2(n18851), .A(n17454), .B(n17453), .ZN(
        n17469) );
  INV_X1 U12911 ( .A(n14244), .ZN(n17454) );
  INV_X1 U12912 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17646) );
  INV_X1 U12913 ( .A(n17756), .ZN(n17787) );
  NAND2_X1 U12914 ( .A1(n17846), .A2(n17872), .ZN(n17868) );
  NAND2_X1 U12915 ( .A1(n18145), .A2(n18144), .ZN(n18091) );
  OAI21_X2 U12916 ( .B1(n18645), .B2(n13250), .A(n18644), .ZN(n18666) );
  NAND3_X1 U12917 ( .A1(n15496), .A2(n15495), .A3(n15494), .ZN(n16401) );
  NAND2_X1 U12918 ( .A1(n14253), .A2(n18189), .ZN(n18231) );
  INV_X1 U12919 ( .A(U212), .ZN(n16508) );
  OR3_X1 U12920 ( .A1(n15646), .A2(n19992), .A3(n12785), .ZN(n19988) );
  INV_X1 U12921 ( .A(n20092), .ZN(n20064) );
  INV_X1 U12922 ( .A(n20051), .ZN(n20029) );
  OR3_X1 U12923 ( .A1(n13865), .A2(n12214), .A3(n13864), .ZN(n20081) );
  INV_X1 U12924 ( .A(n12390), .ZN(n12391) );
  INV_X1 U12925 ( .A(n13760), .ZN(n14609) );
  NAND2_X1 U12926 ( .A1(n14611), .A2(n11619), .ZN(n14595) );
  INV_X1 U12927 ( .A(n15770), .ZN(n15714) );
  INV_X1 U12928 ( .A(n15800), .ZN(n14180) );
  NAND2_X1 U12929 ( .A1(n12738), .A2(n12737), .ZN(n14670) );
  INV_X1 U12930 ( .A(n20120), .ZN(n20146) );
  INV_X1 U12931 ( .A(n20152), .ZN(n20151) );
  INV_X1 U12932 ( .A(n15809), .ZN(n20157) );
  INV_X1 U12933 ( .A(n15799), .ZN(n20191) );
  INV_X1 U12934 ( .A(n15999), .ZN(n20179) );
  NAND2_X1 U12935 ( .A1(n12807), .A2(n12781), .ZN(n15988) );
  INV_X1 U12936 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20188) );
  NAND2_X1 U12937 ( .A1(n20270), .A2(n20448), .ZN(n20268) );
  AOI22_X1 U12938 ( .A1(n20272), .A2(n20275), .B1(n10073), .B2(n20521), .ZN(
        n20296) );
  AOI21_X1 U12939 ( .B1(n20698), .B2(n20304), .A(n20303), .ZN(n20335) );
  NAND2_X1 U12940 ( .A1(n20389), .A2(n20448), .ZN(n20388) );
  AOI22_X1 U12941 ( .A1(n20397), .A2(n20394), .B1(n10073), .B2(n20586), .ZN(
        n20419) );
  NAND2_X1 U12942 ( .A1(n20389), .A2(n20657), .ZN(n20447) );
  NAND2_X1 U12943 ( .A1(n20553), .A2(n20448), .ZN(n20515) );
  AOI22_X1 U12944 ( .A1(n20526), .A2(n20522), .B1(n20521), .B2(n20520), .ZN(
        n20547) );
  NAND2_X1 U12945 ( .A1(n20553), .A2(n20548), .ZN(n20594) );
  AOI22_X1 U12946 ( .A1(n20591), .A2(n20588), .B1(n20586), .B2(n20585), .ZN(
        n20626) );
  NAND2_X1 U12947 ( .A1(n20658), .A2(n20627), .ZN(n20662) );
  NAND2_X1 U12948 ( .A1(n20658), .A2(n20657), .ZN(n20735) );
  INV_X1 U12949 ( .A(n13460), .ZN(n19992) );
  INV_X1 U12950 ( .A(n20851), .ZN(n20847) );
  INV_X1 U12951 ( .A(n20837), .ZN(n20830) );
  AND2_X1 U12952 ( .A1(n16348), .A2(n16367), .ZN(n18870) );
  AOI22_X1 U12953 ( .A1(n16036), .A2(n16030), .B1(n19019), .B2(n19101), .ZN(
        n16031) );
  OR2_X1 U12954 ( .A1(n14148), .A2(n14147), .ZN(n18939) );
  INV_X1 U12955 ( .A(n19019), .ZN(n19083) );
  INV_X1 U12956 ( .A(n19093), .ZN(n19075) );
  INV_X1 U12957 ( .A(n14936), .ZN(n14884) );
  AND2_X1 U12958 ( .A1(n13145), .A2(n16367), .ZN(n19132) );
  NAND2_X1 U12959 ( .A1(n13146), .A2(n19132), .ZN(n19162) );
  INV_X1 U12960 ( .A(n19211), .ZN(n19205) );
  INV_X1 U12961 ( .A(n19231), .ZN(n19254) );
  INV_X1 U12962 ( .A(n19229), .ZN(n13449) );
  INV_X1 U12963 ( .A(n12415), .ZN(n12416) );
  INV_X1 U12964 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18978) );
  OR2_X1 U12965 ( .A1(n18875), .A2(n11191), .ZN(n16219) );
  INV_X1 U12966 ( .A(n16227), .ZN(n19269) );
  NOR2_X1 U12967 ( .A1(n10078), .A2(n11372), .ZN(n11373) );
  INV_X1 U12968 ( .A(n16301), .ZN(n16315) );
  INV_X1 U12969 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19950) );
  AOI211_X2 U12970 ( .C1(n19275), .C2(n19278), .A(n19274), .B(n19357), .ZN(
        n19320) );
  INV_X1 U12971 ( .A(n19371), .ZN(n19379) );
  OR2_X1 U12972 ( .A1(n19419), .A2(n19915), .ZN(n19410) );
  OR2_X1 U12973 ( .A1(n19506), .A2(n19915), .ZN(n19445) );
  INV_X1 U12974 ( .A(n19470), .ZN(n19466) );
  INV_X1 U12975 ( .A(n19486), .ZN(n19494) );
  INV_X1 U12976 ( .A(n19527), .ZN(n19525) );
  OR2_X1 U12977 ( .A1(n19506), .A2(n19505), .ZN(n19561) );
  INV_X1 U12978 ( .A(n19614), .ZN(n19623) );
  INV_X1 U12979 ( .A(n19619), .ZN(n19653) );
  AOI211_X2 U12980 ( .C1(n14112), .C2(n14111), .A(n14113), .B(n14110), .ZN(
        n19674) );
  NAND2_X1 U12981 ( .A1(n19677), .A2(n19682), .ZN(n19745) );
  NAND2_X1 U12982 ( .A1(n19714), .A2(n19763), .ZN(n19818) );
  INV_X1 U12983 ( .A(n19911), .ZN(n19834) );
  XNOR2_X1 U12984 ( .A(n10438), .B(n10437), .ZN(n10439) );
  INV_X1 U12985 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17724) );
  INV_X1 U12986 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16816) );
  INV_X1 U12987 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17213) );
  INV_X1 U12988 ( .A(n17369), .ZN(n17317) );
  INV_X1 U12989 ( .A(n16401), .ZN(n17349) );
  NOR2_X1 U12990 ( .A1(n13325), .A2(n13324), .ZN(n17364) );
  INV_X1 U12991 ( .A(n17446), .ZN(n17442) );
  NAND2_X1 U12992 ( .A1(n17453), .A2(n17385), .ZN(n17451) );
  INV_X1 U12993 ( .A(n17500), .ZN(n17497) );
  INV_X1 U12994 ( .A(n17729), .ZN(n17682) );
  NOR2_X1 U12995 ( .A1(n17729), .A2(n17539), .ZN(n17857) );
  INV_X1 U12996 ( .A(n18169), .ZN(n18159) );
  INV_X1 U12997 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18086) );
  INV_X1 U12998 ( .A(n18126), .ZN(n18175) );
  INV_X1 U12999 ( .A(n18846), .ZN(n18697) );
  INV_X1 U13000 ( .A(n18800), .ZN(n18713) );
  INV_X1 U13001 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18728) );
  CLKBUF_X1 U13002 ( .A(n18790), .Z(n18791) );
  AND2_X1 U13003 ( .A1(n12748), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20189)
         );
  INV_X1 U13004 ( .A(n16502), .ZN(n16511) );
  OAI21_X1 U13005 ( .B1(n14616), .B2(n14609), .A(n12391), .ZN(P1_U2842) );
  OAI211_X1 U13006 ( .C1(n14799), .C2(n20158), .A(n10083), .B(n12717), .ZN(
        P1_U2970) );
  XNOR2_X1 U13007 ( .A(n10440), .B(n10439), .ZN(P3_U2640) );
  NAND4_X1 U13008 ( .A1(n17781), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17697) );
  NAND2_X1 U13009 ( .A1(n17814), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16828) );
  INV_X1 U13010 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17713) );
  NAND2_X1 U13011 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17671) );
  INV_X1 U13012 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16678) );
  INV_X1 U13013 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10103) );
  INV_X1 U13014 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17607) );
  NOR2_X1 U13015 ( .A1(n10103), .A2(n17607), .ZN(n17579) );
  INV_X1 U13016 ( .A(n17579), .ZN(n17600) );
  NAND2_X1 U13017 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17551) );
  INV_X1 U13018 ( .A(n17551), .ZN(n10092) );
  INV_X1 U13019 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17537) );
  INV_X1 U13020 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16392) );
  NAND2_X1 U13021 ( .A1(n10094), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10093) );
  NOR3_X1 U13022 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18708) );
  NAND2_X1 U13023 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18708), .ZN(n18704) );
  INV_X1 U13024 ( .A(n18704), .ZN(n16830) );
  INV_X1 U13025 ( .A(n16830), .ZN(n16808) );
  NOR2_X1 U13026 ( .A1(n16791), .A2(n16808), .ZN(n16899) );
  XOR2_X1 U13027 ( .A(n10094), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16573) );
  AOI21_X1 U13028 ( .B1(n10095), .B2(n16392), .A(n10094), .ZN(n16582) );
  INV_X1 U13029 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U13030 ( .A1(n10098), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10097) );
  INV_X1 U13031 ( .A(n10095), .ZN(n16394) );
  AOI21_X1 U13032 ( .B1(n10096), .B2(n10097), .A(n16394), .ZN(n17505) );
  OAI21_X1 U13033 ( .B1(n10098), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n10097), .ZN(n17524) );
  INV_X1 U13034 ( .A(n17524), .ZN(n16601) );
  AOI21_X1 U13035 ( .B1(n9805), .B2(n17537), .A(n10098), .ZN(n17540) );
  INV_X1 U13036 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17562) );
  NOR2_X1 U13037 ( .A1(n10100), .A2(n17562), .ZN(n10099) );
  OAI21_X1 U13038 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n10099), .A(
        n9805), .ZN(n17553) );
  INV_X1 U13039 ( .A(n17553), .ZN(n16622) );
  AOI21_X1 U13040 ( .B1(n10100), .B2(n17562), .A(n10099), .ZN(n17559) );
  OAI21_X1 U13041 ( .B1(n17578), .B2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n10100), .ZN(n17581) );
  INV_X1 U13042 ( .A(n17581), .ZN(n13343) );
  INV_X1 U13043 ( .A(n10101), .ZN(n10104) );
  NAND2_X1 U13044 ( .A1(n10104), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10102) );
  AOI21_X1 U13045 ( .B1(n10103), .B2(n10102), .A(n17578), .ZN(n17591) );
  OAI22_X1 U13046 ( .A1(n10101), .A2(n17607), .B1(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n10104), .ZN(n17604) );
  INV_X1 U13047 ( .A(n17604), .ZN(n16654) );
  OAI21_X1 U13048 ( .B1(n9740), .B2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n10101), .ZN(n10105) );
  INV_X1 U13049 ( .A(n10105), .ZN(n17620) );
  INV_X1 U13050 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17685) );
  INV_X1 U13051 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16883) );
  NAND2_X1 U13052 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16883), .ZN(
        n16757) );
  NOR3_X1 U13053 ( .A1(n17685), .A2(n17679), .A3(n16757), .ZN(n16709) );
  AND2_X1 U13054 ( .A1(n9740), .A2(n16709), .ZN(n10106) );
  NOR2_X1 U13055 ( .A1(n13343), .A2(n13342), .ZN(n13341) );
  NOR2_X1 U13056 ( .A1(n16601), .A2(n16600), .ZN(n16599) );
  INV_X1 U13057 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18787) );
  INV_X1 U13058 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18780) );
  INV_X1 U13059 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18776) );
  INV_X1 U13060 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18774) );
  INV_X1 U13061 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18766) );
  NAND2_X1 U13062 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16887) );
  INV_X1 U13063 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18735) );
  NOR2_X1 U13064 ( .A1(n16887), .A2(n18735), .ZN(n16860) );
  NAND2_X1 U13065 ( .A1(n16860), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n16846) );
  INV_X1 U13066 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18739) );
  NOR2_X1 U13067 ( .A1(n16846), .A2(n18739), .ZN(n16821) );
  NAND2_X1 U13068 ( .A1(n16821), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n16822) );
  INV_X1 U13069 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18743) );
  NOR2_X1 U13070 ( .A1(n16822), .A2(n18743), .ZN(n16803) );
  NAND2_X1 U13071 ( .A1(n16803), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n16778) );
  NAND2_X1 U13072 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16786) );
  INV_X1 U13073 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18751) );
  NOR3_X1 U13074 ( .A1(n16778), .A2(n16786), .A3(n18751), .ZN(n16760) );
  NAND2_X1 U13075 ( .A1(n16760), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n16748) );
  INV_X1 U13076 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18755) );
  NOR2_X1 U13077 ( .A1(n16748), .A2(n18755), .ZN(n16736) );
  NAND2_X1 U13078 ( .A1(n16736), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n16673) );
  NAND2_X1 U13079 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16702) );
  INV_X1 U13080 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18763) );
  NOR2_X1 U13081 ( .A1(n16702), .A2(n18763), .ZN(n16672) );
  NAND2_X1 U13082 ( .A1(n16672), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n16676) );
  NOR3_X1 U13083 ( .A1(n18766), .A2(n16673), .A3(n16676), .ZN(n16660) );
  NAND2_X1 U13084 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16660), .ZN(n16639) );
  INV_X1 U13085 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18771) );
  NOR2_X1 U13086 ( .A1(n16639), .A2(n18771), .ZN(n16645) );
  NAND2_X1 U13087 ( .A1(n16645), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n13340) );
  OR2_X1 U13088 ( .A1(n18774), .A2(n13340), .ZN(n16631) );
  NOR2_X1 U13089 ( .A1(n18776), .A2(n16631), .ZN(n10218) );
  NOR2_X2 U13090 ( .A1(n10115), .A2(n18657), .ZN(n13290) );
  BUF_X4 U13091 ( .A(n13290), .Z(n17191) );
  AOI22_X1 U13092 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10124) );
  INV_X2 U13093 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18825) );
  AOI22_X1 U13094 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10123) );
  INV_X1 U13095 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13096 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10109) );
  OAI21_X1 U13097 ( .B1(n17144), .B2(n10394), .A(n10109), .ZN(n10121) );
  AOI22_X1 U13098 ( .A1(n13274), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10119) );
  NOR2_X2 U13099 ( .A1(n10113), .A2(n10111), .ZN(n10188) );
  AOI22_X1 U13100 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10118) );
  INV_X2 U13101 ( .A(n10125), .ZN(n17041) );
  AOI22_X1 U13102 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10117) );
  INV_X2 U13103 ( .A(n13299), .ZN(n15523) );
  AOI22_X1 U13104 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10116) );
  NAND4_X1 U13105 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n10120) );
  CLKBUF_X3 U13106 ( .A(n10188), .Z(n17182) );
  AOI22_X1 U13107 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13289), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10129) );
  INV_X2 U13108 ( .A(n10125), .ZN(n17177) );
  AOI22_X1 U13109 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U13110 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U13111 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10126) );
  NAND4_X1 U13112 ( .A1(n10129), .A2(n10128), .A3(n10127), .A4(n10126), .ZN(
        n10135) );
  AOI22_X1 U13113 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U13114 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U13115 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15508), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U13116 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10130) );
  NAND4_X1 U13117 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10134) );
  AOI22_X1 U13118 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U13119 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10144) );
  AOI22_X1 U13120 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10136) );
  OAI21_X1 U13121 ( .B1(n17144), .B2(n17127), .A(n10136), .ZN(n10142) );
  AOI22_X1 U13122 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U13123 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15508), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U13124 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10138) );
  AOI22_X1 U13125 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10137) );
  NAND4_X1 U13126 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10141) );
  AOI211_X1 U13127 ( .C1(n17175), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n10142), .B(n10141), .ZN(n10143) );
  NAND3_X1 U13128 ( .A1(n10145), .A2(n10144), .A3(n10143), .ZN(n10204) );
  BUF_X4 U13129 ( .A(n13289), .Z(n17181) );
  AOI22_X1 U13130 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U13131 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10154) );
  INV_X1 U13132 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17199) );
  INV_X2 U13133 ( .A(n13277), .ZN(n17162) );
  AOI22_X1 U13134 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10146) );
  OAI21_X1 U13135 ( .B1(n10125), .B2(n17199), .A(n10146), .ZN(n10152) );
  AOI22_X1 U13136 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13274), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10150) );
  INV_X2 U13137 ( .A(n13299), .ZN(n17183) );
  AOI22_X1 U13138 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13139 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U13140 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10147) );
  NAND4_X1 U13141 ( .A1(n10150), .A2(n10149), .A3(n10148), .A4(n10147), .ZN(
        n10151) );
  NAND3_X2 U13142 ( .A1(n10155), .A2(n10154), .A3(n10153), .ZN(n17321) );
  NAND2_X1 U13143 ( .A1(n18191), .A2(n17321), .ZN(n13245) );
  NOR2_X1 U13144 ( .A1(n10204), .A2(n13245), .ZN(n10176) );
  AOI22_X1 U13145 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13146 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13274), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U13147 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U13148 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10156) );
  NAND4_X1 U13149 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10165) );
  AOI22_X1 U13150 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U13151 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U13152 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13153 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10160) );
  NAND4_X1 U13154 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n10164) );
  AOI22_X1 U13155 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U13156 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U13157 ( .A1(n15508), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U13158 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9725), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10166) );
  NAND4_X1 U13159 ( .A1(n10169), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n10175) );
  AOI22_X1 U13160 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U13161 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U13162 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U13163 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10170) );
  NAND4_X1 U13164 ( .A1(n10173), .A2(n10172), .A3(n10171), .A4(n10170), .ZN(
        n10174) );
  NAND3_X1 U13165 ( .A1(n18208), .A2(n10176), .A3(n13261), .ZN(n18647) );
  AOI22_X1 U13166 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13167 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13168 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U13169 ( .A1(n15508), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10177) );
  NAND4_X1 U13170 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10186) );
  AOI22_X1 U13171 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U13172 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U13173 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13174 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10181) );
  NAND4_X1 U13175 ( .A1(n10184), .A2(n10183), .A3(n10182), .A4(n10181), .ZN(
        n10185) );
  NAND2_X1 U13176 ( .A1(n18217), .A2(n17238), .ZN(n13241) );
  OAI21_X1 U13177 ( .B1(n10203), .B2(n17387), .A(n13241), .ZN(n10201) );
  NOR2_X1 U13178 ( .A1(n18226), .A2(n13261), .ZN(n10199) );
  AOI22_X1 U13179 ( .A1(n13274), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10187) );
  OAI21_X1 U13180 ( .B1(n13299), .B2(n15438), .A(n10187), .ZN(n10194) );
  AOI22_X1 U13181 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U13182 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10188), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13183 ( .A1(n17177), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13184 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10189) );
  NAND4_X1 U13185 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10193) );
  NOR2_X1 U13186 ( .A1(n13236), .A2(n13269), .ZN(n10198) );
  OAI22_X1 U13187 ( .A1(n18208), .A2(n10199), .B1(n13261), .B2(n10198), .ZN(
        n10200) );
  NOR2_X1 U13188 ( .A1(n13269), .A2(n10204), .ZN(n13239) );
  NAND2_X1 U13189 ( .A1(n10202), .A2(n13239), .ZN(n15393) );
  NOR2_X1 U13190 ( .A1(n13245), .A2(n15393), .ZN(n10205) );
  INV_X1 U13191 ( .A(n10204), .ZN(n18204) );
  INV_X1 U13192 ( .A(n13237), .ZN(n13267) );
  NAND3_X1 U13193 ( .A1(n18213), .A2(n13267), .A3(n17387), .ZN(n14244) );
  NAND2_X1 U13194 ( .A1(n13236), .A2(n16546), .ZN(n14245) );
  AOI21_X2 U13195 ( .B1(n10205), .B2(n18850), .A(n18631), .ZN(n18648) );
  NOR2_X4 U13196 ( .A1(n13238), .A2(n13250), .ZN(n18632) );
  XNOR2_X1 U13197 ( .A(n13256), .B(n13260), .ZN(n10217) );
  INV_X1 U13198 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18681) );
  OAI22_X1 U13199 ( .A1(n18817), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18677), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U13200 ( .A1(n10208), .A2(n18807), .ZN(n10211) );
  OR2_X1 U13201 ( .A1(n10211), .A2(n18680), .ZN(n10209) );
  AOI22_X1 U13202 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18643), .B1(
        n10208), .B2(n18807), .ZN(n10212) );
  AOI22_X1 U13203 ( .A1(n18681), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n10209), .B2(n10212), .ZN(n10216) );
  NAND2_X1 U13204 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18643), .ZN(
        n10210) );
  OAI22_X1 U13205 ( .A1(n10212), .A2(n18680), .B1(n10211), .B2(n10210), .ZN(
        n13255) );
  XNOR2_X1 U13206 ( .A(n10214), .B(n10213), .ZN(n13254) );
  OAI21_X1 U13207 ( .B1(n13255), .B2(n13254), .A(n10216), .ZN(n13258) );
  INV_X1 U13208 ( .A(n13258), .ZN(n10215) );
  NAND2_X1 U13209 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18810), .ZN(n18700) );
  NAND2_X1 U13210 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18728), .ZN(n18841) );
  INV_X2 U13211 ( .A(n18841), .ZN(n18788) );
  NAND2_X1 U13212 ( .A1(n18788), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18795) );
  INV_X1 U13213 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18716) );
  INV_X1 U13214 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18730) );
  NAND2_X1 U13215 ( .A1(n18716), .A2(n18730), .ZN(n16551) );
  NAND3_X1 U13216 ( .A1(n18728), .A2(n18786), .A3(n16551), .ZN(n18848) );
  NAND2_X1 U13217 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18851) );
  INV_X1 U13218 ( .A(n18851), .ZN(n18722) );
  AOI211_X1 U13219 ( .C1(n18850), .C2(n18848), .A(n18722), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18689) );
  NAND2_X1 U13220 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16617), .ZN(n16616) );
  NOR2_X1 U13221 ( .A1(n18780), .A2(n16616), .ZN(n16605) );
  NAND3_X1 U13222 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16605), .ZN(n16585) );
  NOR2_X1 U13223 ( .A1(n18787), .A2(n16585), .ZN(n10222) );
  INV_X1 U13224 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18794) );
  NAND2_X1 U13225 ( .A1(n10222), .A2(n18794), .ZN(n16576) );
  NOR2_X1 U13226 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18863) );
  INV_X1 U13227 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n14253) );
  NAND3_X1 U13228 ( .A1(n18863), .A2(n14253), .A3(n18862), .ZN(n13328) );
  INV_X1 U13229 ( .A(n18700), .ZN(n17873) );
  NAND2_X1 U13230 ( .A1(n17873), .A2(n9706), .ZN(n18695) );
  NAND4_X1 U13231 ( .A1(n13328), .A2(n18859), .A3(n18695), .A4(n16808), .ZN(
        n16914) );
  NAND4_X1 U13232 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(P3_REIP_REG_26__SCAN_IN), 
        .A3(n10218), .A4(n16914), .ZN(n16592) );
  NAND3_X1 U13233 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U13234 ( .A1(n16902), .A2(n16914), .ZN(n16912) );
  OAI21_X1 U13235 ( .B1(n16592), .B2(n10219), .A(n16912), .ZN(n16584) );
  INV_X1 U13236 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18792) );
  AOI21_X1 U13237 ( .B1(n16576), .B2(n16584), .A(n18792), .ZN(n10226) );
  NOR2_X1 U13238 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16900) );
  NAND2_X1 U13239 ( .A1(n16900), .A2(n17213), .ZN(n16895) );
  NOR2_X1 U13240 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16895), .ZN(n16873) );
  INV_X1 U13241 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16857) );
  NAND2_X1 U13242 ( .A1(n16873), .A2(n16857), .ZN(n16854) );
  INV_X1 U13243 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16836) );
  NAND2_X1 U13244 ( .A1(n16847), .A2(n16836), .ZN(n16833) );
  INV_X1 U13245 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16813) );
  NAND2_X1 U13246 ( .A1(n16818), .A2(n16813), .ZN(n16812) );
  INV_X1 U13247 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17155) );
  NAND2_X1 U13248 ( .A1(n16794), .A2(n17155), .ZN(n16787) );
  INV_X1 U13249 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16765) );
  NAND2_X1 U13250 ( .A1(n16768), .A2(n16765), .ZN(n16764) );
  INV_X1 U13251 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17111) );
  NAND2_X1 U13252 ( .A1(n16749), .A2(n17111), .ZN(n16741) );
  INV_X1 U13253 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17039) );
  NAND2_X1 U13254 ( .A1(n16724), .A2(n17039), .ZN(n16713) );
  INV_X1 U13255 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17053) );
  NAND2_X1 U13256 ( .A1(n16703), .A2(n17053), .ZN(n16691) );
  INV_X1 U13257 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16667) );
  NAND2_X1 U13258 ( .A1(n16682), .A2(n16667), .ZN(n16666) );
  INV_X1 U13259 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16644) );
  NAND2_X1 U13260 ( .A1(n16651), .A2(n16644), .ZN(n16643) );
  INV_X1 U13261 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16919) );
  NAND2_X1 U13262 ( .A1(n16634), .A2(n16919), .ZN(n16619) );
  INV_X1 U13263 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16956) );
  NAND2_X1 U13264 ( .A1(n16618), .A2(n16956), .ZN(n16613) );
  NOR2_X1 U13265 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16613), .ZN(n16602) );
  INV_X1 U13266 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16593) );
  NAND2_X1 U13267 ( .A1(n16602), .A2(n16593), .ZN(n16589) );
  NOR2_X1 U13268 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16589), .ZN(n16579) );
  INV_X1 U13269 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16925) );
  NAND2_X1 U13270 ( .A1(n16579), .A2(n16925), .ZN(n16570) );
  INV_X1 U13271 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18849) );
  NAND2_X1 U13272 ( .A1(n18849), .A2(n18851), .ZN(n10220) );
  NAND4_X1 U13273 ( .A1(n10221), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n16398), 
        .A4(n10220), .ZN(n16911) );
  INV_X1 U13274 ( .A(n10221), .ZN(n18864) );
  AOI211_X4 U13275 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16398), .A(n18689), .B(
        n18864), .ZN(n16871) );
  AOI22_X1 U13276 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16898), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16871), .ZN(n10224) );
  NAND3_X1 U13277 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n10222), .A3(n18792), 
        .ZN(n10223) );
  OAI211_X1 U13278 ( .C1(n16570), .C2(n16911), .A(n10224), .B(n10223), .ZN(
        n10225) );
  AOI211_X1 U13279 ( .C1(n16899), .C2(n16571), .A(n10226), .B(n10225), .ZN(
        n10440) );
  INV_X1 U13280 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16507) );
  AOI22_X1 U13281 ( .A1(n18817), .A2(keyinput68), .B1(n16507), .B2(keyinput92), 
        .ZN(n10227) );
  OAI221_X1 U13282 ( .B1(n18817), .B2(keyinput68), .C1(n16507), .C2(keyinput92), .A(n10227), .ZN(n10236) );
  INV_X1 U13283 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19872) );
  INV_X1 U13284 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U13285 ( .A1(n19872), .A2(keyinput65), .B1(keyinput79), .B2(n10229), 
        .ZN(n10228) );
  OAI221_X1 U13286 ( .B1(n19872), .B2(keyinput65), .C1(n10229), .C2(keyinput79), .A(n10228), .ZN(n10235) );
  INV_X1 U13287 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10424) );
  INV_X1 U13288 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U13289 ( .A1(n10424), .A2(keyinput100), .B1(n10231), .B2(
        keyinput110), .ZN(n10230) );
  OAI221_X1 U13290 ( .B1(n10424), .B2(keyinput100), .C1(n10231), .C2(
        keyinput110), .A(n10230), .ZN(n10234) );
  INV_X1 U13291 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17402) );
  INV_X1 U13292 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U13293 ( .A1(n17402), .A2(keyinput52), .B1(n19866), .B2(keyinput44), 
        .ZN(n10232) );
  OAI221_X1 U13294 ( .B1(n17402), .B2(keyinput52), .C1(n19866), .C2(keyinput44), .A(n10232), .ZN(n10233) );
  NOR4_X1 U13295 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10267) );
  INV_X1 U13296 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20842) );
  AOI22_X1 U13297 ( .A1(n20842), .A2(keyinput54), .B1(n10394), .B2(keyinput25), 
        .ZN(n10237) );
  OAI221_X1 U13298 ( .B1(n20842), .B2(keyinput54), .C1(n10394), .C2(keyinput25), .A(n10237), .ZN(n10247) );
  INV_X1 U13299 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n19524) );
  INV_X1 U13300 ( .A(P2_DATAWIDTH_REG_29__SCAN_IN), .ZN(n19830) );
  AOI22_X1 U13301 ( .A1(n19524), .A2(keyinput95), .B1(keyinput12), .B2(n19830), 
        .ZN(n10238) );
  OAI221_X1 U13302 ( .B1(n19524), .B2(keyinput95), .C1(n19830), .C2(keyinput12), .A(n10238), .ZN(n10246) );
  INV_X1 U13303 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17097) );
  INV_X1 U13304 ( .A(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U13305 ( .A1(n17097), .A2(keyinput70), .B1(n10240), .B2(keyinput40), 
        .ZN(n10239) );
  OAI221_X1 U13306 ( .B1(n17097), .B2(keyinput70), .C1(n10240), .C2(keyinput40), .A(n10239), .ZN(n10245) );
  INV_X1 U13307 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10241) );
  XOR2_X1 U13308 ( .A(n10241), .B(keyinput124), .Z(n10243) );
  XNOR2_X1 U13309 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput50), 
        .ZN(n10242) );
  NAND2_X1 U13310 ( .A1(n10243), .A2(n10242), .ZN(n10244) );
  NOR4_X1 U13311 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10266) );
  INV_X1 U13312 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11804) );
  INV_X1 U13313 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19509) );
  AOI22_X1 U13314 ( .A1(n11804), .A2(keyinput23), .B1(n19509), .B2(keyinput66), 
        .ZN(n10248) );
  OAI221_X1 U13315 ( .B1(n11804), .B2(keyinput23), .C1(n19509), .C2(keyinput66), .A(n10248), .ZN(n10255) );
  INV_X1 U13316 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15510) );
  AOI22_X1 U13317 ( .A1(n15510), .A2(keyinput98), .B1(n15438), .B2(keyinput82), 
        .ZN(n10249) );
  OAI221_X1 U13318 ( .B1(n15510), .B2(keyinput98), .C1(n15438), .C2(keyinput82), .A(n10249), .ZN(n10254) );
  INV_X1 U13319 ( .A(P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19831) );
  INV_X1 U13320 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13321 ( .A1(n19831), .A2(keyinput34), .B1(n10694), .B2(keyinput56), 
        .ZN(n10250) );
  OAI221_X1 U13322 ( .B1(n19831), .B2(keyinput34), .C1(n10694), .C2(keyinput56), .A(n10250), .ZN(n10253) );
  INV_X1 U13323 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14295) );
  AOI22_X1 U13324 ( .A1(n14295), .A2(keyinput73), .B1(n18941), .B2(keyinput105), .ZN(n10251) );
  OAI221_X1 U13325 ( .B1(n14295), .B2(keyinput73), .C1(n18941), .C2(
        keyinput105), .A(n10251), .ZN(n10252) );
  NOR4_X1 U13326 ( .A1(n10255), .A2(n10254), .A3(n10253), .A4(n10252), .ZN(
        n10265) );
  INV_X1 U13327 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20113) );
  INV_X1 U13328 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17654) );
  AOI22_X1 U13329 ( .A1(n20113), .A2(keyinput125), .B1(n17654), .B2(keyinput96), .ZN(n10256) );
  OAI221_X1 U13330 ( .B1(n20113), .B2(keyinput125), .C1(n17654), .C2(
        keyinput96), .A(n10256), .ZN(n10263) );
  INV_X1 U13331 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18122) );
  AOI22_X1 U13332 ( .A1(n18122), .A2(keyinput114), .B1(n18643), .B2(keyinput11), .ZN(n10257) );
  OAI221_X1 U13333 ( .B1(n18122), .B2(keyinput114), .C1(n18643), .C2(
        keyinput11), .A(n10257), .ZN(n10262) );
  INV_X1 U13334 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n20134) );
  INV_X1 U13335 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U13336 ( .A1(n20134), .A2(keyinput43), .B1(n17443), .B2(keyinput5), 
        .ZN(n10258) );
  OAI221_X1 U13337 ( .B1(n20134), .B2(keyinput43), .C1(n17443), .C2(keyinput5), 
        .A(n10258), .ZN(n10261) );
  INV_X1 U13338 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19998) );
  INV_X1 U13339 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U13340 ( .A1(n19998), .A2(keyinput91), .B1(keyinput93), .B2(n17396), 
        .ZN(n10259) );
  OAI221_X1 U13341 ( .B1(n19998), .B2(keyinput91), .C1(n17396), .C2(keyinput93), .A(n10259), .ZN(n10260) );
  NOR4_X1 U13342 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10264) );
  NAND4_X1 U13343 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10392) );
  INV_X1 U13344 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16537) );
  INV_X1 U13345 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U13346 ( .A1(n16537), .A2(keyinput19), .B1(n10269), .B2(keyinput60), 
        .ZN(n10268) );
  OAI221_X1 U13347 ( .B1(n16537), .B2(keyinput19), .C1(n10269), .C2(keyinput60), .A(n10268), .ZN(n10277) );
  INV_X1 U13348 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11737) );
  INV_X1 U13349 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n20150) );
  AOI22_X1 U13350 ( .A1(n11737), .A2(keyinput51), .B1(keyinput47), .B2(n20150), 
        .ZN(n10270) );
  OAI221_X1 U13351 ( .B1(n11737), .B2(keyinput51), .C1(n20150), .C2(keyinput47), .A(n10270), .ZN(n10276) );
  INV_X1 U13352 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18180) );
  INV_X1 U13353 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U13354 ( .A1(n18180), .A2(keyinput31), .B1(n17179), .B2(keyinput49), 
        .ZN(n10271) );
  OAI221_X1 U13355 ( .B1(n18180), .B2(keyinput31), .C1(n17179), .C2(keyinput49), .A(n10271), .ZN(n10275) );
  INV_X1 U13356 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10273) );
  INV_X1 U13357 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16413) );
  AOI22_X1 U13358 ( .A1(n10273), .A2(keyinput46), .B1(keyinput27), .B2(n16413), 
        .ZN(n10272) );
  OAI221_X1 U13359 ( .B1(n10273), .B2(keyinput46), .C1(n16413), .C2(keyinput27), .A(n10272), .ZN(n10274) );
  NOR4_X1 U13360 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n10308) );
  INV_X1 U13361 ( .A(P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19829) );
  AOI22_X1 U13362 ( .A1(n15374), .A2(keyinput18), .B1(keyinput9), .B2(n19829), 
        .ZN(n10278) );
  OAI221_X1 U13363 ( .B1(n15374), .B2(keyinput18), .C1(n19829), .C2(keyinput9), 
        .A(n10278), .ZN(n10285) );
  INV_X1 U13364 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20854) );
  AOI22_X1 U13365 ( .A1(n14215), .A2(keyinput108), .B1(keyinput21), .B2(n20854), .ZN(n10279) );
  OAI221_X1 U13366 ( .B1(n14215), .B2(keyinput108), .C1(n20854), .C2(
        keyinput21), .A(n10279), .ZN(n10284) );
  INV_X1 U13367 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15986) );
  INV_X1 U13368 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U13369 ( .A1(n15986), .A2(keyinput126), .B1(n12422), .B2(keyinput58), .ZN(n10280) );
  OAI221_X1 U13370 ( .B1(n15986), .B2(keyinput126), .C1(n12422), .C2(
        keyinput58), .A(n10280), .ZN(n10283) );
  INV_X1 U13371 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18222) );
  INV_X1 U13372 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U13373 ( .A1(n18222), .A2(keyinput28), .B1(keyinput17), .B2(n17138), 
        .ZN(n10281) );
  OAI221_X1 U13374 ( .B1(n18222), .B2(keyinput28), .C1(n17138), .C2(keyinput17), .A(n10281), .ZN(n10282) );
  NOR4_X1 U13375 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10307) );
  INV_X1 U13376 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10287) );
  INV_X1 U13377 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n20464) );
  AOI22_X1 U13378 ( .A1(n10287), .A2(keyinput13), .B1(keyinput35), .B2(n20464), 
        .ZN(n10286) );
  OAI221_X1 U13379 ( .B1(n10287), .B2(keyinput13), .C1(n20464), .C2(keyinput35), .A(n10286), .ZN(n10295) );
  INV_X1 U13380 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13381 ( .A1(n17127), .A2(keyinput74), .B1(n10289), .B2(keyinput32), 
        .ZN(n10288) );
  OAI221_X1 U13382 ( .B1(n17127), .B2(keyinput74), .C1(n10289), .C2(keyinput32), .A(n10288), .ZN(n10294) );
  INV_X1 U13383 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20633) );
  INV_X1 U13384 ( .A(P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n20766) );
  AOI22_X1 U13385 ( .A1(n20633), .A2(keyinput24), .B1(keyinput39), .B2(n20766), 
        .ZN(n10290) );
  OAI221_X1 U13386 ( .B1(n20633), .B2(keyinput24), .C1(n20766), .C2(keyinput39), .A(n10290), .ZN(n10293) );
  INV_X1 U13387 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17000) );
  INV_X1 U13388 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U13389 ( .A1(n17000), .A2(keyinput113), .B1(n17488), .B2(keyinput94), .ZN(n10291) );
  OAI221_X1 U13390 ( .B1(n17000), .B2(keyinput113), .C1(n17488), .C2(
        keyinput94), .A(n10291), .ZN(n10292) );
  NOR4_X1 U13391 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10306) );
  AOI22_X1 U13392 ( .A1(n14765), .A2(keyinput41), .B1(keyinput122), .B2(n16667), .ZN(n10296) );
  OAI221_X1 U13393 ( .B1(n14765), .B2(keyinput41), .C1(n16667), .C2(
        keyinput122), .A(n10296), .ZN(n10304) );
  INV_X1 U13394 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10298) );
  INV_X1 U13395 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U13396 ( .A1(n10298), .A2(keyinput81), .B1(keyinput10), .B2(n11748), 
        .ZN(n10297) );
  OAI221_X1 U13397 ( .B1(n10298), .B2(keyinput81), .C1(n11748), .C2(keyinput10), .A(n10297), .ZN(n10303) );
  INV_X1 U13398 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14425) );
  INV_X1 U13399 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13572) );
  AOI22_X1 U13400 ( .A1(n14425), .A2(keyinput26), .B1(n13572), .B2(keyinput63), 
        .ZN(n10299) );
  OAI221_X1 U13401 ( .B1(n14425), .B2(keyinput26), .C1(n13572), .C2(keyinput63), .A(n10299), .ZN(n10302) );
  INV_X1 U13402 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16532) );
  INV_X1 U13403 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n20334) );
  AOI22_X1 U13404 ( .A1(n16532), .A2(keyinput97), .B1(n20334), .B2(keyinput29), 
        .ZN(n10300) );
  OAI221_X1 U13405 ( .B1(n16532), .B2(keyinput97), .C1(n20334), .C2(keyinput29), .A(n10300), .ZN(n10301) );
  NOR4_X1 U13406 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10305) );
  NAND4_X1 U13407 ( .A1(n10308), .A2(n10307), .A3(n10306), .A4(n10305), .ZN(
        n10391) );
  INV_X1 U13408 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U13409 ( .A1(n16593), .A2(keyinput88), .B1(keyinput2), .B2(n17424), 
        .ZN(n10309) );
  OAI221_X1 U13410 ( .B1(n16593), .B2(keyinput88), .C1(n17424), .C2(keyinput2), 
        .A(n10309), .ZN(n10317) );
  INV_X1 U13411 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15997) );
  INV_X1 U13412 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13413 ( .A1(n15997), .A2(keyinput76), .B1(n10311), .B2(keyinput107), .ZN(n10310) );
  OAI221_X1 U13414 ( .B1(n15997), .B2(keyinput76), .C1(n10311), .C2(
        keyinput107), .A(n10310), .ZN(n10316) );
  INV_X1 U13415 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16566) );
  INV_X1 U13416 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13417 ( .A1(n16566), .A2(keyinput115), .B1(n10774), .B2(keyinput85), .ZN(n10312) );
  OAI221_X1 U13418 ( .B1(n16566), .B2(keyinput115), .C1(n10774), .C2(
        keyinput85), .A(n10312), .ZN(n10315) );
  INV_X1 U13419 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n20310) );
  INV_X1 U13420 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18732) );
  AOI22_X1 U13421 ( .A1(n20310), .A2(keyinput53), .B1(keyinput119), .B2(n18732), .ZN(n10313) );
  OAI221_X1 U13422 ( .B1(n20310), .B2(keyinput53), .C1(n18732), .C2(
        keyinput119), .A(n10313), .ZN(n10314) );
  NOR4_X1 U13423 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10348) );
  INV_X1 U13424 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18785) );
  INV_X1 U13425 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15898) );
  AOI22_X1 U13426 ( .A1(n18785), .A2(keyinput3), .B1(n15898), .B2(keyinput4), 
        .ZN(n10318) );
  OAI221_X1 U13427 ( .B1(n18785), .B2(keyinput3), .C1(n15898), .C2(keyinput4), 
        .A(n10318), .ZN(n10325) );
  INV_X1 U13428 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17490) );
  AOI22_X1 U13429 ( .A1(n18849), .A2(keyinput75), .B1(n17490), .B2(keyinput80), 
        .ZN(n10319) );
  OAI221_X1 U13430 ( .B1(n18849), .B2(keyinput75), .C1(n17490), .C2(keyinput80), .A(n10319), .ZN(n10324) );
  INV_X1 U13431 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20843) );
  INV_X1 U13432 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n19188) );
  AOI22_X1 U13433 ( .A1(n20843), .A2(keyinput57), .B1(n19188), .B2(keyinput102), .ZN(n10320) );
  OAI221_X1 U13434 ( .B1(n20843), .B2(keyinput57), .C1(n19188), .C2(
        keyinput102), .A(n10320), .ZN(n10323) );
  INV_X1 U13435 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14775) );
  INV_X1 U13436 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15874) );
  AOI22_X1 U13437 ( .A1(n14775), .A2(keyinput103), .B1(n15874), .B2(keyinput78), .ZN(n10321) );
  OAI221_X1 U13438 ( .B1(n14775), .B2(keyinput103), .C1(n15874), .C2(
        keyinput78), .A(n10321), .ZN(n10322) );
  NOR4_X1 U13439 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10347) );
  INV_X1 U13440 ( .A(P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19833) );
  AOI22_X1 U13441 ( .A1(n19833), .A2(keyinput90), .B1(n19926), .B2(keyinput33), 
        .ZN(n10326) );
  OAI221_X1 U13442 ( .B1(n19833), .B2(keyinput90), .C1(n19926), .C2(keyinput33), .A(n10326), .ZN(n10334) );
  INV_X1 U13443 ( .A(P3_LWORD_REG_5__SCAN_IN), .ZN(n17437) );
  INV_X1 U13444 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U13445 ( .A1(n17437), .A2(keyinput69), .B1(n16469), .B2(keyinput14), 
        .ZN(n10327) );
  OAI221_X1 U13446 ( .B1(n17437), .B2(keyinput69), .C1(n16469), .C2(keyinput14), .A(n10327), .ZN(n10333) );
  INV_X1 U13447 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14699) );
  INV_X1 U13448 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18223) );
  AOI22_X1 U13449 ( .A1(n14699), .A2(keyinput0), .B1(keyinput83), .B2(n18223), 
        .ZN(n10328) );
  OAI221_X1 U13450 ( .B1(n14699), .B2(keyinput0), .C1(n18223), .C2(keyinput83), 
        .A(n10328), .ZN(n10332) );
  INV_X1 U13451 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n19172) );
  INV_X1 U13452 ( .A(P3_LWORD_REG_6__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13453 ( .A1(n19172), .A2(keyinput106), .B1(n10330), .B2(keyinput87), .ZN(n10329) );
  OAI221_X1 U13454 ( .B1(n19172), .B2(keyinput106), .C1(n10330), .C2(
        keyinput87), .A(n10329), .ZN(n10331) );
  NOR4_X1 U13455 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10346) );
  INV_X1 U13456 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n17432) );
  INV_X1 U13457 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20826) );
  AOI22_X1 U13458 ( .A1(n17432), .A2(keyinput55), .B1(n20826), .B2(keyinput48), 
        .ZN(n10335) );
  OAI221_X1 U13459 ( .B1(n17432), .B2(keyinput55), .C1(n20826), .C2(keyinput48), .A(n10335), .ZN(n10344) );
  INV_X1 U13460 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10338) );
  INV_X1 U13461 ( .A(DATAI_28_), .ZN(n10337) );
  AOI22_X1 U13462 ( .A1(n10338), .A2(keyinput20), .B1(keyinput64), .B2(n10337), 
        .ZN(n10336) );
  OAI221_X1 U13463 ( .B1(n10338), .B2(keyinput20), .C1(n10337), .C2(keyinput64), .A(n10336), .ZN(n10343) );
  INV_X1 U13464 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18779) );
  INV_X1 U13465 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U13466 ( .A1(n18779), .A2(keyinput61), .B1(n18202), .B2(keyinput36), 
        .ZN(n10339) );
  OAI221_X1 U13467 ( .B1(n18779), .B2(keyinput61), .C1(n18202), .C2(keyinput36), .A(n10339), .ZN(n10342) );
  INV_X1 U13468 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16530) );
  INV_X1 U13469 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n19190) );
  AOI22_X1 U13470 ( .A1(n16530), .A2(keyinput1), .B1(keyinput45), .B2(n19190), 
        .ZN(n10340) );
  OAI221_X1 U13471 ( .B1(n16530), .B2(keyinput1), .C1(n19190), .C2(keyinput45), 
        .A(n10340), .ZN(n10341) );
  NOR4_X1 U13472 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10345) );
  NAND4_X1 U13473 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10390) );
  INV_X1 U13474 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17486) );
  INV_X1 U13475 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13476 ( .A1(n17486), .A2(keyinput67), .B1(n10822), .B2(keyinput71), 
        .ZN(n10349) );
  OAI221_X1 U13477 ( .B1(n17486), .B2(keyinput67), .C1(n10822), .C2(keyinput71), .A(n10349), .ZN(n10356) );
  INV_X1 U13478 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n20461) );
  INV_X1 U13479 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n19178) );
  AOI22_X1 U13480 ( .A1(n20461), .A2(keyinput117), .B1(keyinput6), .B2(n19178), 
        .ZN(n10350) );
  OAI221_X1 U13481 ( .B1(n20461), .B2(keyinput117), .C1(n19178), .C2(keyinput6), .A(n10350), .ZN(n10355) );
  INV_X1 U13482 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13446) );
  INV_X1 U13483 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18768) );
  AOI22_X1 U13484 ( .A1(n13446), .A2(keyinput116), .B1(keyinput99), .B2(n18768), .ZN(n10351) );
  OAI221_X1 U13485 ( .B1(n13446), .B2(keyinput116), .C1(n18768), .C2(
        keyinput99), .A(n10351), .ZN(n10354) );
  INV_X1 U13486 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n20122) );
  INV_X1 U13487 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13935) );
  AOI22_X1 U13488 ( .A1(n20122), .A2(keyinput42), .B1(n13935), .B2(keyinput112), .ZN(n10352) );
  OAI221_X1 U13489 ( .B1(n20122), .B2(keyinput42), .C1(n13935), .C2(
        keyinput112), .A(n10352), .ZN(n10353) );
  NOR4_X1 U13490 ( .A1(n10356), .A2(n10355), .A3(n10354), .A4(n10353), .ZN(
        n10388) );
  INV_X1 U13491 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n10358) );
  INV_X1 U13492 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19863) );
  AOI22_X1 U13493 ( .A1(n10358), .A2(keyinput89), .B1(n19863), .B2(keyinput38), 
        .ZN(n10357) );
  OAI221_X1 U13494 ( .B1(n10358), .B2(keyinput89), .C1(n19863), .C2(keyinput38), .A(n10357), .ZN(n10365) );
  INV_X1 U13495 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n17400) );
  INV_X1 U13496 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20861) );
  AOI22_X1 U13497 ( .A1(n17400), .A2(keyinput37), .B1(n20861), .B2(keyinput123), .ZN(n10359) );
  OAI221_X1 U13498 ( .B1(n17400), .B2(keyinput37), .C1(n20861), .C2(
        keyinput123), .A(n10359), .ZN(n10364) );
  INV_X1 U13499 ( .A(P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19832) );
  INV_X1 U13500 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19902) );
  AOI22_X1 U13501 ( .A1(n19832), .A2(keyinput121), .B1(keyinput16), .B2(n19902), .ZN(n10360) );
  OAI221_X1 U13502 ( .B1(n19832), .B2(keyinput121), .C1(n19902), .C2(
        keyinput16), .A(n10360), .ZN(n10363) );
  INV_X1 U13503 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n19180) );
  INV_X1 U13504 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U13505 ( .A1(n19180), .A2(keyinput15), .B1(n10926), .B2(keyinput30), 
        .ZN(n10361) );
  OAI221_X1 U13506 ( .B1(n19180), .B2(keyinput15), .C1(n10926), .C2(keyinput30), .A(n10361), .ZN(n10362) );
  NOR4_X1 U13507 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10387) );
  INV_X1 U13508 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U13509 ( .A1(n9862), .A2(keyinput127), .B1(keyinput8), .B2(n11448), 
        .ZN(n10366) );
  OAI221_X1 U13510 ( .B1(n9862), .B2(keyinput127), .C1(n11448), .C2(keyinput8), 
        .A(n10366), .ZN(n10374) );
  INV_X1 U13511 ( .A(P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(n18709) );
  INV_X1 U13512 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n19175) );
  AOI22_X1 U13513 ( .A1(n18709), .A2(keyinput62), .B1(n19175), .B2(keyinput111), .ZN(n10367) );
  OAI221_X1 U13514 ( .B1(n18709), .B2(keyinput62), .C1(n19175), .C2(
        keyinput111), .A(n10367), .ZN(n10373) );
  INV_X1 U13515 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n19206) );
  INV_X1 U13516 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13517 ( .A1(n19206), .A2(keyinput7), .B1(n10369), .B2(keyinput86), 
        .ZN(n10368) );
  OAI221_X1 U13518 ( .B1(n19206), .B2(keyinput7), .C1(n10369), .C2(keyinput86), 
        .A(n10368), .ZN(n10372) );
  INV_X1 U13519 ( .A(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n18710) );
  INV_X1 U13520 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13521 ( .A1(n18710), .A2(keyinput120), .B1(n10393), .B2(keyinput22), .ZN(n10370) );
  OAI221_X1 U13522 ( .B1(n18710), .B2(keyinput120), .C1(n10393), .C2(
        keyinput22), .A(n10370), .ZN(n10371) );
  NOR4_X1 U13523 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10386) );
  INV_X1 U13524 ( .A(P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n18712) );
  INV_X1 U13525 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U13526 ( .A1(n18712), .A2(keyinput109), .B1(keyinput72), .B2(n17413), .ZN(n10375) );
  OAI221_X1 U13527 ( .B1(n18712), .B2(keyinput109), .C1(n17413), .C2(
        keyinput72), .A(n10375), .ZN(n10380) );
  INV_X1 U13528 ( .A(DATAI_13_), .ZN(n10377) );
  INV_X1 U13529 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19319) );
  AOI22_X1 U13530 ( .A1(n10377), .A2(keyinput59), .B1(n19319), .B2(keyinput118), .ZN(n10376) );
  OAI221_X1 U13531 ( .B1(n10377), .B2(keyinput59), .C1(n19319), .C2(
        keyinput118), .A(n10376), .ZN(n10379) );
  XOR2_X1 U13532 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B(keyinput77), .Z(
        n10378) );
  OR3_X1 U13533 ( .A1(n10380), .A2(n10379), .A3(n10378), .ZN(n10384) );
  INV_X1 U13534 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12575) );
  INV_X1 U13535 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20784) );
  AOI22_X1 U13536 ( .A1(n12575), .A2(keyinput104), .B1(keyinput101), .B2(
        n20784), .ZN(n10381) );
  OAI221_X1 U13537 ( .B1(n12575), .B2(keyinput104), .C1(n20784), .C2(
        keyinput101), .A(n10381), .ZN(n10383) );
  INV_X1 U13538 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n19187) );
  XNOR2_X1 U13539 ( .A(n19187), .B(keyinput84), .ZN(n10382) );
  NOR3_X1 U13540 ( .A1(n10384), .A2(n10383), .A3(n10382), .ZN(n10385) );
  NAND4_X1 U13541 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10389) );
  NOR4_X1 U13542 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10438) );
  NOR2_X1 U13543 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18878) );
  NOR4_X1 U13544 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_11__6__SCAN_IN), .A3(n18817), .A4(n10393), .ZN(n10395) );
  NAND4_X1 U13545 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18878), .A3(
        n10395), .A4(n10394), .ZN(n10403) );
  NAND4_X1 U13546 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(P3_EBX_REG_20__SCAN_IN), 
        .A3(P3_EBX_REG_15__SCAN_IN), .A4(n16593), .ZN(n10402) );
  NAND4_X1 U13547 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_14__3__SCAN_IN), .A3(n15510), .A4(n18643), .ZN(n10401) );
  NOR4_X1 U13548 ( .A1(DATAI_13_), .A2(P1_UWORD_REG_13__SCAN_IN), .A3(
        P1_LWORD_REG_15__SCAN_IN), .A4(P3_DATAO_REG_7__SCAN_IN), .ZN(n10399)
         );
  NOR4_X1 U13549 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_ADDRESS_REG_1__SCAN_IN), .A4(n18785), .ZN(n10398) );
  NOR4_X1 U13550 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(BUF1_REG_1__SCAN_IN), .A4(P2_LWORD_REG_10__SCAN_IN), .ZN(n10397)
         );
  NOR4_X1 U13551 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAO_REG_18__SCAN_IN), .A3(P1_BE_N_REG_2__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n10396) );
  NAND4_X1 U13552 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10400) );
  NOR4_X1 U13553 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n10436) );
  NAND4_X1 U13554 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(
        P2_BE_N_REG_3__SCAN_IN), .A3(P2_LWORD_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(n10407) );
  NAND4_X1 U13555 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(P2_DATAO_REG_10__SCAN_IN), 
        .A3(P3_ADDRESS_REG_19__SCAN_IN), .A4(P2_DATAWIDTH_REG_9__SCAN_IN), 
        .ZN(n10406) );
  NAND4_X1 U13556 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(
        P2_DATAO_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAO_REG_18__SCAN_IN), .ZN(n10405) );
  NAND4_X1 U13557 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(P2_DATAO_REG_3__SCAN_IN), 
        .A4(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n10404) );
  NOR4_X1 U13558 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        n10435) );
  NAND4_X1 U13559 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .A3(P1_INSTQUEUE_REG_3__0__SCAN_IN), 
        .A4(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10411) );
  NAND4_X1 U13560 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_3__7__SCAN_IN), .A3(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10410) );
  NAND4_X1 U13561 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        BUF1_REG_27__SCAN_IN), .A3(P2_DATAO_REG_26__SCAN_IN), .A4(
        P3_ADDRESS_REG_24__SCAN_IN), .ZN(n10409) );
  NAND4_X1 U13562 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        BUF2_REG_11__SCAN_IN), .A3(P1_BE_N_REG_1__SCAN_IN), .A4(
        P3_LWORD_REG_5__SCAN_IN), .ZN(n10408) );
  NOR4_X1 U13563 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10434) );
  NOR4_X1 U13564 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_7__6__SCAN_IN), .A3(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A4(P2_EAX_REG_24__SCAN_IN), .ZN(n10415) );
  NOR4_X1 U13565 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_REIP_REG_7__SCAN_IN), .A3(P2_EBX_REG_27__SCAN_IN), .A4(
        BUF2_REG_19__SCAN_IN), .ZN(n10414) );
  NOR4_X1 U13566 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_1__3__SCAN_IN), .A3(P1_INSTQUEUE_REG_13__3__SCAN_IN), 
        .A4(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10413) );
  NOR4_X1 U13567 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_12__4__SCAN_IN), .A3(P1_INSTQUEUE_REG_8__0__SCAN_IN), 
        .A4(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10412) );
  NAND4_X1 U13568 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10432) );
  NOR4_X1 U13569 ( .A1(BUF2_REG_10__SCAN_IN), .A2(P3_DATAO_REG_3__SCAN_IN), 
        .A3(P3_DATAO_REG_23__SCAN_IN), .A4(P3_DATAO_REG_24__SCAN_IN), .ZN(
        n10419) );
  NOR4_X1 U13570 ( .A1(BUF2_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(P3_LWORD_REG_6__SCAN_IN), 
        .ZN(n10418) );
  NOR4_X1 U13571 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(P2_DATAO_REG_21__SCAN_IN), .A3(P2_DATAO_REG_23__SCAN_IN), .A4(P2_DATAO_REG_28__SCAN_IN), .ZN(n10417) );
  NOR4_X1 U13572 ( .A1(BUF2_REG_7__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), .A3(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A4(P2_DATAO_REG_15__SCAN_IN), .ZN(
        n10416) );
  NAND4_X1 U13573 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(
        n10431) );
  NAND4_X1 U13574 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(
        P1_FLUSH_REG_SCAN_IN), .A3(P3_DATAO_REG_26__SCAN_IN), .A4(
        P3_FLUSH_REG_SCAN_IN), .ZN(n10423) );
  NAND4_X1 U13575 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(P1_DATAO_REG_5__SCAN_IN), .ZN(
        n10422) );
  NAND4_X1 U13576 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_14__2__SCAN_IN), .A3(P1_STATEBS16_REG_SCAN_IN), .A4(
        BUF2_REG_23__SCAN_IN), .ZN(n10421) );
  NAND4_X1 U13577 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_EBX_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n10420) );
  OR4_X1 U13578 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n10430) );
  NOR4_X1 U13579 ( .A1(n19872), .A2(n19866), .A3(n10424), .A4(n17402), .ZN(
        n10428) );
  NOR4_X1 U13580 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A4(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10426) );
  NOR4_X1 U13581 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_6__7__SCAN_IN), .A3(P1_REIP_REG_25__SCAN_IN), .A4(
        DATAI_28_), .ZN(n10425) );
  AND4_X1 U13582 ( .A1(n16413), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n10426), .A4(n10425), .ZN(n10427) );
  NAND4_X1 U13583 ( .A1(n10428), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A3(
        n10427), .A4(n14775), .ZN(n10429) );
  NOR4_X1 U13584 ( .A1(n10432), .A2(n10431), .A3(n10430), .A4(n10429), .ZN(
        n10433) );
  NAND4_X1 U13585 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n10437) );
  AND2_X4 U13586 ( .A1(n15378), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13130) );
  AOI22_X1 U13587 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13130), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10446) );
  AND2_X4 U13588 ( .A1(n10442), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13125) );
  AND2_X4 U13589 ( .A1(n10441), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13131) );
  AOI22_X1 U13590 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13591 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10444) );
  BUF_X4 U13592 ( .A(n10488), .Z(n13123) );
  INV_X2 U13593 ( .A(n13129), .ZN(n10663) );
  AOI22_X1 U13594 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10443) );
  NAND4_X1 U13595 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10447) );
  AOI22_X1 U13597 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13130), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13598 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U13599 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U13600 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10448) );
  NAND4_X1 U13601 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10452) );
  AOI22_X1 U13602 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13130), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13603 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13604 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U13605 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10453) );
  NAND4_X1 U13606 ( .A1(n10456), .A2(n10455), .A3(n10454), .A4(n10453), .ZN(
        n10457) );
  NAND2_X1 U13607 ( .A1(n10457), .A2(n10470), .ZN(n10464) );
  AOI22_X1 U13608 ( .A1(n10509), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U13609 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13610 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13611 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10458) );
  NAND4_X1 U13612 ( .A1(n10461), .A2(n10460), .A3(n10459), .A4(n10458), .ZN(
        n10462) );
  NAND2_X1 U13613 ( .A1(n10462), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10463) );
  AOI22_X1 U13614 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13615 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9737), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13616 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13617 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10466) );
  NAND4_X1 U13618 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n10477) );
  AOI22_X1 U13619 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13130), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13620 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9737), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10471) );
  AND2_X1 U13621 ( .A1(n10471), .A2(n10470), .ZN(n10474) );
  AOI22_X1 U13622 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13623 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10472) );
  NAND4_X1 U13624 ( .A1(n10475), .A2(n10474), .A3(n10473), .A4(n10472), .ZN(
        n10476) );
  NAND2_X2 U13625 ( .A1(n10477), .A2(n10476), .ZN(n11019) );
  AOI22_X1 U13626 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13130), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13627 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13628 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13629 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9738), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10478) );
  NAND4_X1 U13630 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10487) );
  AOI22_X1 U13631 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13632 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13633 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10483) );
  AOI22_X1 U13634 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10482) );
  NAND4_X1 U13635 ( .A1(n10485), .A2(n10484), .A3(n10483), .A4(n10482), .ZN(
        n10486) );
  MUX2_X2 U13636 ( .A(n10487), .B(n10486), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10547) );
  AOI22_X1 U13637 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13638 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13639 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10490) );
  BUF_X4 U13640 ( .A(n10488), .Z(n13118) );
  AOI22_X1 U13641 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13642 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13643 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13644 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13645 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10493) );
  NAND2_X1 U13646 ( .A1(n11082), .A2(n11084), .ZN(n10504) );
  NAND2_X1 U13647 ( .A1(n11019), .A2(n10549), .ZN(n10500) );
  NAND2_X1 U13648 ( .A1(n10560), .A2(n10500), .ZN(n10502) );
  INV_X1 U13649 ( .A(n10547), .ZN(n13160) );
  NAND2_X2 U13650 ( .A1(n10529), .A2(n13160), .ZN(n10567) );
  AOI22_X1 U13651 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13130), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13652 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13653 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13654 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10505) );
  NAND4_X1 U13655 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10515) );
  AOI22_X1 U13656 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13657 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9708), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13658 ( .A1(n10664), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13659 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10510) );
  NAND4_X1 U13660 ( .A1(n10513), .A2(n10512), .A3(n10511), .A4(n10510), .ZN(
        n10514) );
  MUX2_X2 U13661 ( .A(n10515), .B(n10514), .S(n10470), .Z(n19968) );
  AOI22_X1 U13662 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13663 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13664 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13665 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10516) );
  NAND4_X1 U13666 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(
        n10520) );
  NAND2_X1 U13667 ( .A1(n10520), .A2(n10470), .ZN(n10527) );
  AOI22_X1 U13668 ( .A1(n13082), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13669 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13670 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U13671 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10521) );
  NAND4_X1 U13672 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10525) );
  NAND2_X1 U13673 ( .A1(n10525), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10526) );
  NAND2_X2 U13674 ( .A1(n10527), .A2(n10526), .ZN(n11196) );
  AND2_X1 U13675 ( .A1(n11201), .A2(n19283), .ZN(n10528) );
  AOI22_X1 U13676 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13677 ( .A1(n13125), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13678 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13679 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9737), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10530) );
  NAND4_X1 U13680 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10539) );
  AOI22_X1 U13681 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13125), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13682 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13683 ( .A1(n13130), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10664), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13684 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10534) );
  NAND4_X1 U13685 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10538) );
  MUX2_X2 U13686 ( .A(n10539), .B(n10538), .S(n10470), .Z(n11078) );
  NAND2_X1 U13687 ( .A1(n10529), .A2(n10540), .ZN(n10542) );
  NOR2_X1 U13688 ( .A1(n10555), .A2(n19300), .ZN(n10545) );
  NAND2_X1 U13689 ( .A1(n10550), .A2(n10545), .ZN(n10982) );
  NOR2_X1 U13690 ( .A1(n19283), .A2(n11078), .ZN(n10546) );
  NAND2_X1 U13691 ( .A1(n10982), .A2(n10546), .ZN(n10552) );
  INV_X1 U13692 ( .A(n10547), .ZN(n10548) );
  NOR2_X1 U13693 ( .A1(n11190), .A2(n10549), .ZN(n10551) );
  AND2_X2 U13694 ( .A1(n10551), .A2(n10550), .ZN(n10553) );
  NAND2_X1 U13695 ( .A1(n10612), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10559) );
  INV_X1 U13696 ( .A(n11001), .ZN(n10556) );
  NOR2_X1 U13697 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19963) );
  AOI22_X1 U13698 ( .A1(n11180), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19963), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10558) );
  NAND2_X1 U13699 ( .A1(n10559), .A2(n10558), .ZN(n10577) );
  INV_X1 U13700 ( .A(n10577), .ZN(n10575) );
  NAND2_X1 U13701 ( .A1(n11001), .A2(n11040), .ZN(n13142) );
  OAI211_X1 U13702 ( .C1(n10081), .C2(n11084), .A(n10562), .B(n13142), .ZN(
        n10563) );
  INV_X1 U13703 ( .A(n10563), .ZN(n11184) );
  NAND2_X1 U13704 ( .A1(n10607), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10573) );
  AND2_X1 U13705 ( .A1(n13429), .A2(n11196), .ZN(n13023) );
  INV_X1 U13706 ( .A(n10566), .ZN(n10571) );
  INV_X1 U13707 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13585) );
  NAND2_X1 U13708 ( .A1(n10573), .A2(n10572), .ZN(n10576) );
  INV_X1 U13709 ( .A(n10576), .ZN(n10574) );
  NAND2_X1 U13710 ( .A1(n10575), .A2(n10574), .ZN(n10594) );
  NAND2_X1 U13711 ( .A1(n10577), .A2(n10576), .ZN(n10578) );
  INV_X1 U13712 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n19090) );
  INV_X1 U13713 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19077) );
  INV_X1 U13714 ( .A(n10583), .ZN(n10586) );
  NAND2_X1 U13715 ( .A1(n10608), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13716 ( .A1(n9734), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10587) );
  AND3_X1 U13717 ( .A1(n11077), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10568), 
        .ZN(n10589) );
  INV_X1 U13718 ( .A(n10610), .ZN(n12544) );
  OAI22_X1 U13719 ( .A1(n10612), .A2(n10589), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12544), .ZN(n10593) );
  NAND2_X1 U13720 ( .A1(n19963), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10590) );
  AND2_X1 U13721 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  NAND2_X1 U13722 ( .A1(n10593), .A2(n10592), .ZN(n10621) );
  NAND2_X1 U13723 ( .A1(n10612), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10596) );
  AOI21_X1 U13724 ( .B1(n19969), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U13725 ( .A1(n10596), .A2(n10595), .ZN(n10603) );
  AOI22_X1 U13726 ( .A1(n10608), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10597) );
  INV_X1 U13727 ( .A(n10597), .ZN(n10599) );
  INV_X1 U13728 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13701) );
  NAND2_X1 U13729 ( .A1(n9735), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10600) );
  NAND2_X1 U13730 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  OR2_X2 U13731 ( .A1(n10603), .A2(n10602), .ZN(n10606) );
  NAND2_X1 U13732 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  INV_X1 U13733 ( .A(n10626), .ZN(n10605) );
  NAND2_X1 U13734 ( .A1(n10607), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10611) );
  AOI22_X1 U13735 ( .A1(n12543), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10609) );
  INV_X1 U13736 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13712) );
  NAND2_X1 U13737 ( .A1(n10612), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10614) );
  NAND2_X1 U13738 ( .A1(n19963), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10613) );
  NAND2_X1 U13739 ( .A1(n10614), .A2(n10613), .ZN(n10618) );
  NAND2_X1 U13740 ( .A1(n10618), .A2(n10617), .ZN(n10619) );
  INV_X1 U13741 ( .A(n10624), .ZN(n10625) );
  XNOR2_X2 U13742 ( .A(n9755), .B(n10627), .ZN(n13995) );
  NAND2_X1 U13743 ( .A1(n10658), .A2(n13995), .ZN(n10695) );
  INV_X1 U13744 ( .A(n13995), .ZN(n10646) );
  NOR2_X4 U13745 ( .A1(n10659), .A2(n14399), .ZN(n19597) );
  AOI22_X1 U13746 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19352), .B1(
        n19597), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10662) );
  INV_X1 U13747 ( .A(n9777), .ZN(n10628) );
  NAND2_X1 U13748 ( .A1(n10631), .A2(n10640), .ZN(n19564) );
  INV_X1 U13749 ( .A(n19564), .ZN(n19567) );
  NAND2_X1 U13750 ( .A1(n12824), .A2(n10636), .ZN(n10633) );
  INV_X1 U13751 ( .A(n10633), .ZN(n10630) );
  NAND2_X1 U13752 ( .A1(n10640), .A2(n10630), .ZN(n10682) );
  INV_X1 U13753 ( .A(n10682), .ZN(n19758) );
  AOI22_X1 U13754 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19567), .B1(
        n19758), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10645) );
  INV_X1 U13755 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13033) );
  INV_X1 U13756 ( .A(n10640), .ZN(n10632) );
  INV_X1 U13757 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10634) );
  OAI22_X1 U13758 ( .A1(n13033), .A2(n19326), .B1(n19498), .B2(n10634), .ZN(
        n10635) );
  INV_X1 U13759 ( .A(n10635), .ZN(n10644) );
  INV_X1 U13760 ( .A(n19381), .ZN(n19386) );
  AND2_X1 U13761 ( .A1(n12824), .A2(n9777), .ZN(n10638) );
  NAND2_X1 U13762 ( .A1(n10640), .A2(n10638), .ZN(n10679) );
  INV_X1 U13763 ( .A(n10679), .ZN(n19680) );
  AOI22_X1 U13764 ( .A1(n19386), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n19680), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10643) );
  INV_X1 U13765 ( .A(n10638), .ZN(n10639) );
  NAND2_X1 U13766 ( .A1(n10641), .A2(n10640), .ZN(n10690) );
  INV_X1 U13767 ( .A(n10690), .ZN(n19626) );
  NAND4_X1 U13768 ( .A1(n10645), .A2(n10644), .A3(n10643), .A4(n10642), .ZN(
        n10657) );
  NAND2_X1 U13769 ( .A1(n12824), .A2(n10646), .ZN(n10650) );
  INV_X1 U13770 ( .A(n10650), .ZN(n10647) );
  NAND2_X1 U13771 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10655) );
  NAND2_X1 U13772 ( .A1(n12824), .A2(n13995), .ZN(n10649) );
  NAND2_X1 U13773 ( .A1(n10757), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10653) );
  NOR2_X2 U13774 ( .A1(n10651), .A2(n10650), .ZN(n10756) );
  NAND2_X1 U13775 ( .A1(n10756), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10652) );
  NAND4_X1 U13776 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(
        n10656) );
  NOR2_X1 U13777 ( .A1(n10657), .A2(n10656), .ZN(n10661) );
  NAND2_X1 U13778 ( .A1(n10658), .A2(n14399), .ZN(n10677) );
  AOI22_X1 U13779 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19276), .B1(
        n10764), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10660) );
  AND2_X2 U13780 ( .A1(n13125), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10768) );
  AOI22_X1 U13781 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10669) );
  NOR4_X2 U13782 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U13783 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10668) );
  AND2_X2 U13784 ( .A1(n13118), .A2(n10470), .ZN(n12970) );
  AOI22_X1 U13785 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12970), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10667) );
  AND2_X2 U13786 ( .A1(n10665), .A2(n10470), .ZN(n12972) );
  AOI22_X1 U13787 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10666) );
  NAND4_X1 U13788 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10675) );
  AND2_X2 U13789 ( .A1(n9723), .A2(n10470), .ZN(n12962) );
  AOI22_X1 U13790 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13791 ( .A1(n12899), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13792 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10671) );
  AND2_X1 U13793 ( .A1(n13131), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10769) );
  AOI22_X1 U13794 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10769), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10670) );
  NAND4_X1 U13795 ( .A1(n10673), .A2(n10672), .A3(n10671), .A4(n10670), .ZN(
        n10674) );
  INV_X1 U13796 ( .A(n10814), .ZN(n11219) );
  NAND2_X1 U13797 ( .A1(n11219), .A2(n19283), .ZN(n10676) );
  INV_X1 U13798 ( .A(n19326), .ZN(n19321) );
  INV_X1 U13799 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19287) );
  OR2_X1 U13800 ( .A1(n10677), .A2(n19287), .ZN(n10686) );
  INV_X1 U13801 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10680) );
  INV_X1 U13802 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10678) );
  OAI22_X1 U13803 ( .A1(n10680), .A2(n19498), .B1(n10679), .B2(n10678), .ZN(
        n10684) );
  INV_X1 U13804 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12989) );
  INV_X1 U13805 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10681) );
  OAI22_X1 U13806 ( .A1(n12989), .A2(n19564), .B1(n10682), .B2(n10681), .ZN(
        n10683) );
  NOR2_X1 U13807 ( .A1(n10684), .A2(n10683), .ZN(n10685) );
  INV_X1 U13808 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10687) );
  INV_X1 U13809 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10689) );
  OR2_X1 U13810 ( .A1(n10690), .A2(n10689), .ZN(n10691) );
  NAND2_X1 U13811 ( .A1(n19597), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10698) );
  OR2_X1 U13812 ( .A1(n10695), .A2(n10694), .ZN(n10697) );
  NAND2_X1 U13813 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10696) );
  NAND4_X1 U13814 ( .A1(n10699), .A2(n10698), .A3(n10697), .A4(n10696), .ZN(
        n10736) );
  AOI22_X1 U13815 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13816 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13817 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10769), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13818 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10700) );
  NAND4_X1 U13819 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n10710) );
  AOI22_X1 U13820 ( .A1(n12899), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10775), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13821 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13822 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13823 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10705) );
  NAND4_X1 U13824 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n10709) );
  NOR2_X1 U13825 ( .A1(n10710), .A2(n10709), .ZN(n13356) );
  OR2_X1 U13826 ( .A1(n13356), .A2(n11191), .ZN(n11043) );
  INV_X1 U13827 ( .A(n11043), .ZN(n10721) );
  AOI22_X1 U13828 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12962), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13829 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n11239), .ZN(n10713) );
  AOI22_X1 U13830 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13831 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10711) );
  NAND4_X1 U13832 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n10720) );
  AOI22_X1 U13833 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13834 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12970), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13835 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12971), .B1(
        n10775), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13836 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11244), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10715) );
  NAND4_X1 U13837 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10719) );
  OR2_X2 U13838 ( .A1(n10720), .A2(n10719), .ZN(n11044) );
  NAND2_X1 U13839 ( .A1(n10721), .A2(n11044), .ZN(n11042) );
  AOI22_X1 U13840 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13841 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11239), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13842 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10769), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13843 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10724) );
  NAND4_X1 U13844 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n10734) );
  AOI22_X1 U13845 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13846 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13847 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13848 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10729) );
  NAND4_X1 U13849 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        n10733) );
  NAND2_X1 U13850 ( .A1(n11042), .A2(n11210), .ZN(n10735) );
  AOI22_X1 U13851 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13852 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13853 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U13854 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10738) );
  NAND4_X1 U13855 ( .A1(n10741), .A2(n10740), .A3(n10739), .A4(n10738), .ZN(
        n10747) );
  AOI22_X1 U13856 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13857 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10775), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13858 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13859 ( .A1(n12971), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10742) );
  NAND4_X1 U13860 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(
        n10746) );
  INV_X1 U13861 ( .A(n10821), .ZN(n11222) );
  INV_X1 U13862 ( .A(n19498), .ZN(n10748) );
  AOI22_X1 U13863 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n19626), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10755) );
  INV_X1 U13864 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13076) );
  INV_X1 U13865 ( .A(n10749), .ZN(n19448) );
  INV_X1 U13866 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10750) );
  OAI22_X1 U13867 ( .A1(n13076), .A2(n19326), .B1(n19448), .B2(n10750), .ZN(
        n10751) );
  INV_X1 U13868 ( .A(n10751), .ZN(n10754) );
  AOI22_X1 U13869 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19567), .B1(
        n19758), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13870 ( .A1(n19386), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n19680), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10752) );
  NAND4_X1 U13871 ( .A1(n10755), .A2(n10754), .A3(n10753), .A4(n10752), .ZN(
        n10763) );
  NAND2_X1 U13872 ( .A1(n10756), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10761) );
  NAND2_X1 U13873 ( .A1(n10757), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10760) );
  NAND2_X1 U13874 ( .A1(n19723), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10759) );
  NAND2_X1 U13875 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10758) );
  NAND4_X1 U13876 ( .A1(n10761), .A2(n10760), .A3(n10759), .A4(n10758), .ZN(
        n10762) );
  NOR2_X1 U13877 ( .A1(n10763), .A2(n10762), .ZN(n10767) );
  AOI22_X1 U13878 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19352), .B1(
        n10764), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13879 ( .A1(n19276), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n19597), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10765) );
  NAND3_X1 U13880 ( .A1(n10767), .A2(n10766), .A3(n10765), .ZN(n10784) );
  AOI22_X1 U13881 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13882 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11239), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13883 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13884 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10770) );
  NAND4_X1 U13885 ( .A1(n10773), .A2(n10772), .A3(n10771), .A4(n10770), .ZN(
        n10781) );
  AOI22_X1 U13886 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U13887 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13888 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13889 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10776) );
  NAND4_X1 U13890 ( .A1(n10779), .A2(n10778), .A3(n10777), .A4(n10776), .ZN(
        n10780) );
  INV_X1 U13891 ( .A(n11226), .ZN(n10782) );
  NAND2_X1 U13892 ( .A1(n10782), .A2(n19283), .ZN(n10783) );
  INV_X1 U13893 ( .A(n10786), .ZN(n10785) );
  NAND2_X1 U13894 ( .A1(n11052), .A2(n10785), .ZN(n10787) );
  AOI22_X1 U13895 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13896 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n12964), .ZN(n10790) );
  AOI22_X1 U13897 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n10723), .ZN(n10789) );
  AOI22_X1 U13898 ( .A1(n12899), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12963), .ZN(n10788) );
  NAND4_X1 U13899 ( .A1(n10791), .A2(n10790), .A3(n10789), .A4(n10788), .ZN(
        n10797) );
  AOI22_X1 U13900 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13901 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12970), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13902 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12971), .B1(
        n10775), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13903 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11244), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10792) );
  NAND4_X1 U13904 ( .A1(n10795), .A2(n10794), .A3(n10793), .A4(n10792), .ZN(
        n10796) );
  INV_X1 U13905 ( .A(n11044), .ZN(n11204) );
  NAND2_X1 U13906 ( .A1(n13585), .A2(n19090), .ZN(n10798) );
  MUX2_X2 U13907 ( .A(n11204), .B(n10798), .S(n19300), .Z(n10838) );
  XNOR2_X1 U13908 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U13909 ( .A1(n10985), .A2(n10833), .ZN(n10800) );
  NAND2_X1 U13910 ( .A1(n19943), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10799) );
  NAND2_X1 U13911 ( .A1(n10800), .A2(n10799), .ZN(n10808) );
  XNOR2_X1 U13912 ( .A(n16318), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10806) );
  XNOR2_X1 U13913 ( .A(n10808), .B(n10806), .ZN(n10999) );
  INV_X1 U13914 ( .A(n10999), .ZN(n11008) );
  NAND2_X1 U13915 ( .A1(n11040), .A2(n11008), .ZN(n10801) );
  OAI21_X1 U13916 ( .B1(n10802), .B2(n11040), .A(n10801), .ZN(n10973) );
  NOR2_X2 U13917 ( .A1(n10838), .A2(n10840), .ZN(n10832) );
  INV_X1 U13918 ( .A(n10806), .ZN(n10807) );
  NAND2_X1 U13919 ( .A1(n10808), .A2(n10807), .ZN(n10810) );
  NAND2_X1 U13920 ( .A1(n19933), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10809) );
  NAND2_X1 U13921 ( .A1(n10810), .A2(n10809), .ZN(n10818) );
  XNOR2_X1 U13922 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10817) );
  INV_X1 U13923 ( .A(n10817), .ZN(n10811) );
  XNOR2_X1 U13924 ( .A(n10818), .B(n10811), .ZN(n10975) );
  INV_X1 U13925 ( .A(n10975), .ZN(n10812) );
  NAND2_X1 U13926 ( .A1(n11040), .A2(n10812), .ZN(n10813) );
  OAI21_X1 U13927 ( .B1(n11040), .B2(n10814), .A(n10813), .ZN(n10815) );
  INV_X1 U13928 ( .A(n10815), .ZN(n10816) );
  MUX2_X1 U13929 ( .A(n10816), .B(n13712), .S(n19300), .Z(n10831) );
  NAND2_X1 U13930 ( .A1(n10832), .A2(n10831), .ZN(n10830) );
  NAND2_X1 U13931 ( .A1(n10818), .A2(n10817), .ZN(n10820) );
  NAND2_X1 U13932 ( .A1(n19926), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10819) );
  NAND2_X1 U13933 ( .A1(n10820), .A2(n10819), .ZN(n10978) );
  NAND2_X1 U13934 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16358), .ZN(
        n10979) );
  MUX2_X1 U13935 ( .A(n10821), .B(n10976), .S(n11040), .Z(n10823) );
  MUX2_X1 U13936 ( .A(n10823), .B(n10822), .S(n19300), .Z(n10824) );
  INV_X1 U13937 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13778) );
  MUX2_X1 U13938 ( .A(n11226), .B(n13778), .S(n19300), .Z(n10825) );
  NOR2_X1 U13939 ( .A1(n9797), .A2(n10825), .ZN(n10826) );
  OR2_X1 U13940 ( .A1(n10883), .A2(n10826), .ZN(n19048) );
  INV_X1 U13941 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14095) );
  XNOR2_X1 U13942 ( .A(n10848), .B(n14095), .ZN(n14084) );
  NAND2_X1 U13943 ( .A1(n10827), .A2(n10828), .ZN(n10829) );
  OAI21_X1 U13944 ( .B1(n10832), .B2(n10831), .A(n10830), .ZN(n13713) );
  INV_X1 U13945 ( .A(n10833), .ZN(n10984) );
  NAND2_X1 U13946 ( .A1(n15369), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10834) );
  NAND2_X1 U13947 ( .A1(n10984), .A2(n10834), .ZN(n11004) );
  MUX2_X1 U13948 ( .A(n13356), .B(n11004), .S(n11040), .Z(n10974) );
  MUX2_X1 U13949 ( .A(n10974), .B(n19090), .S(n19300), .Z(n13353) );
  INV_X1 U13950 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10835) );
  NOR2_X1 U13951 ( .A1(n13353), .A2(n10835), .ZN(n13355) );
  INV_X1 U13952 ( .A(n13355), .ZN(n14382) );
  NAND3_X1 U13953 ( .A1(n19300), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U13954 ( .A1(n10838), .A2(n10836), .ZN(n14383) );
  NOR2_X1 U13955 ( .A1(n14382), .A2(n14383), .ZN(n10837) );
  NAND2_X1 U13956 ( .A1(n14382), .A2(n14383), .ZN(n14381) );
  OAI21_X1 U13957 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10837), .A(
        n14381), .ZN(n13424) );
  INV_X1 U13958 ( .A(n10838), .ZN(n10839) );
  XNOR2_X1 U13959 ( .A(n10840), .B(n10839), .ZN(n13834) );
  XNOR2_X1 U13960 ( .A(n13834), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13423) );
  OR2_X1 U13961 ( .A1(n13424), .A2(n13423), .ZN(n13566) );
  NAND2_X1 U13962 ( .A1(n13834), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10841) );
  NAND2_X1 U13963 ( .A1(n13566), .A2(n10841), .ZN(n16232) );
  NAND2_X1 U13964 ( .A1(n9718), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10842) );
  NAND2_X1 U13965 ( .A1(n10843), .A2(n10842), .ZN(n14035) );
  XNOR2_X1 U13966 ( .A(n10830), .B(n10844), .ZN(n19064) );
  XNOR2_X1 U13967 ( .A(n19064), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14036) );
  NAND2_X1 U13968 ( .A1(n14035), .A2(n14036), .ZN(n10847) );
  INV_X1 U13969 ( .A(n19064), .ZN(n10845) );
  NAND2_X1 U13970 ( .A1(n10845), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10846) );
  NAND2_X1 U13971 ( .A1(n10847), .A2(n10846), .ZN(n14085) );
  NAND2_X1 U13972 ( .A1(n14084), .A2(n14085), .ZN(n10850) );
  NAND2_X1 U13973 ( .A1(n10848), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10849) );
  NAND2_X1 U13974 ( .A1(n10850), .A2(n10849), .ZN(n15146) );
  AOI22_X1 U13975 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n19626), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10855) );
  INV_X1 U13976 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13093) );
  OAI22_X1 U13977 ( .A1(n13093), .A2(n19326), .B1(n19498), .B2(n19524), .ZN(
        n10851) );
  INV_X1 U13978 ( .A(n10851), .ZN(n10854) );
  AOI22_X1 U13979 ( .A1(n19386), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n19680), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13980 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19567), .B1(
        n19758), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10852) );
  NAND4_X1 U13981 ( .A1(n10855), .A2(n10854), .A3(n10853), .A4(n10852), .ZN(
        n10861) );
  NAND2_X1 U13982 ( .A1(n10756), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10859) );
  NAND2_X1 U13983 ( .A1(n10757), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10858) );
  NAND2_X1 U13984 ( .A1(n14109), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10857) );
  NAND2_X1 U13985 ( .A1(n19723), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10856) );
  NAND4_X1 U13986 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(
        n10860) );
  NOR2_X1 U13987 ( .A1(n10861), .A2(n10860), .ZN(n10864) );
  AOI22_X1 U13988 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19276), .B1(
        n10764), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U13989 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19352), .B1(
        n19597), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10862) );
  NAND3_X1 U13990 ( .A1(n10864), .A2(n10863), .A3(n10862), .ZN(n10876) );
  AOI22_X1 U13991 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12962), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13992 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12963), .ZN(n10867) );
  AOI22_X1 U13993 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13994 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10865) );
  NAND4_X1 U13995 ( .A1(n10868), .A2(n10867), .A3(n10866), .A4(n10865), .ZN(
        n10874) );
  AOI22_X1 U13996 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U13997 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12970), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13998 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12971), .B1(
        n10775), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13999 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11244), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10869) );
  NAND4_X1 U14000 ( .A1(n10872), .A2(n10871), .A3(n10870), .A4(n10869), .ZN(
        n10873) );
  INV_X1 U14001 ( .A(n10877), .ZN(n11230) );
  NAND2_X1 U14002 ( .A1(n11230), .A2(n19283), .ZN(n10875) );
  NAND2_X1 U14003 ( .A1(n11056), .A2(n12494), .ZN(n10878) );
  INV_X1 U14004 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19035) );
  MUX2_X1 U14005 ( .A(n10877), .B(n19035), .S(n19300), .Z(n10882) );
  XNOR2_X1 U14006 ( .A(n10883), .B(n10882), .ZN(n19036) );
  NAND2_X1 U14007 ( .A1(n10878), .A2(n19036), .ZN(n10879) );
  INV_X1 U14008 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15361) );
  XNOR2_X1 U14009 ( .A(n10879), .B(n15361), .ZN(n15147) );
  NAND2_X1 U14010 ( .A1(n10879), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10880) );
  INV_X1 U14011 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13819) );
  NAND2_X1 U14012 ( .A1(n19300), .A2(n13819), .ZN(n10884) );
  INV_X1 U14013 ( .A(n10887), .ZN(n10885) );
  XNOR2_X1 U14014 ( .A(n10888), .B(n10885), .ZN(n19027) );
  INV_X1 U14015 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11117) );
  NOR2_X1 U14016 ( .A1(n10803), .A2(n11117), .ZN(n10889) );
  OR2_X2 U14017 ( .A1(n10890), .A2(n10889), .ZN(n10898) );
  NAND2_X1 U14018 ( .A1(n10890), .A2(n10889), .ZN(n10891) );
  AND2_X1 U14019 ( .A1(n10898), .A2(n10891), .ZN(n19012) );
  NAND2_X1 U14020 ( .A1(n19012), .A2(n12496), .ZN(n10894) );
  INV_X1 U14021 ( .A(n10894), .ZN(n10892) );
  INV_X1 U14022 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U14023 ( .A1(n10894), .A2(n10893), .ZN(n16207) );
  INV_X1 U14024 ( .A(n19027), .ZN(n10895) );
  INV_X1 U14025 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16297) );
  NAND2_X1 U14026 ( .A1(n10895), .A2(n16297), .ZN(n16205) );
  AND2_X1 U14027 ( .A1(n16207), .A2(n16205), .ZN(n10896) );
  NOR2_X1 U14028 ( .A1(n10803), .A2(n9892), .ZN(n10897) );
  MUX2_X1 U14029 ( .A(n10803), .B(n10897), .S(n10898), .Z(n10899) );
  NOR2_X1 U14030 ( .A1(n10899), .A2(n10907), .ZN(n19000) );
  AOI21_X1 U14031 ( .B1(n19000), .B2(n12496), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15345) );
  INV_X1 U14032 ( .A(n15345), .ZN(n10900) );
  INV_X1 U14033 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n18991) );
  NOR2_X1 U14034 ( .A1(n10907), .A2(n18991), .ZN(n10901) );
  NAND2_X1 U14035 ( .A1(n19300), .A2(n10901), .ZN(n10902) );
  NAND2_X1 U14036 ( .A1(n12473), .A2(n10902), .ZN(n10903) );
  AOI21_X1 U14037 ( .B1(n10907), .B2(n18991), .A(n10903), .ZN(n18989) );
  AOI21_X1 U14038 ( .B1(n18989), .B2(n12496), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16187) );
  INV_X1 U14039 ( .A(n18989), .ZN(n10904) );
  INV_X1 U14040 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16270) );
  AND2_X1 U14041 ( .A1(n12496), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10905) );
  NAND2_X1 U14042 ( .A1(n19000), .A2(n10905), .ZN(n16185) );
  INV_X1 U14043 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U14044 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n9791), .ZN(n10908) );
  NOR2_X1 U14045 ( .A1(n10803), .A2(n10908), .ZN(n10909) );
  OR2_X1 U14046 ( .A1(n10911), .A2(n10909), .ZN(n18979) );
  NOR2_X1 U14047 ( .A1(n18979), .A2(n12494), .ZN(n10914) );
  AND2_X1 U14048 ( .A1(n10914), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15326) );
  NAND2_X1 U14049 ( .A1(n19300), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10910) );
  NAND3_X1 U14050 ( .A1(n19300), .A2(n10912), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n10913) );
  NAND2_X1 U14051 ( .A1(n10920), .A2(n10913), .ZN(n18967) );
  INV_X1 U14052 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15320) );
  INV_X1 U14053 ( .A(n15310), .ZN(n10916) );
  INV_X1 U14054 ( .A(n10914), .ZN(n10915) );
  INV_X1 U14055 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15337) );
  NAND2_X1 U14056 ( .A1(n10915), .A2(n15337), .ZN(n15325) );
  OR2_X1 U14057 ( .A1(n10916), .A2(n15325), .ZN(n10918) );
  OR2_X1 U14058 ( .A1(n18967), .A2(n12494), .ZN(n10917) );
  NAND2_X1 U14059 ( .A1(n10917), .A2(n15320), .ZN(n15311) );
  INV_X1 U14060 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11131) );
  NOR2_X1 U14061 ( .A1(n10803), .A2(n11131), .ZN(n10919) );
  NAND2_X1 U14062 ( .A1(n10920), .A2(n10919), .ZN(n10921) );
  NAND2_X1 U14063 ( .A1(n10932), .A2(n10921), .ZN(n14078) );
  INV_X1 U14064 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15299) );
  OAI21_X1 U14065 ( .B1(n14078), .B2(n12494), .A(n15299), .ZN(n15297) );
  INV_X1 U14066 ( .A(n15297), .ZN(n10923) );
  NAND2_X1 U14067 ( .A1(n12496), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10922) );
  NAND2_X1 U14068 ( .A1(n19300), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10924) );
  MUX2_X1 U14069 ( .A(n19300), .B(n10924), .S(n10932), .Z(n10925) );
  OR2_X1 U14070 ( .A1(n10932), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10930) );
  NAND2_X1 U14071 ( .A1(n18955), .A2(n12496), .ZN(n10927) );
  NAND2_X1 U14072 ( .A1(n10927), .A2(n10926), .ZN(n16156) );
  AND2_X1 U14073 ( .A1(n12496), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10928) );
  NAND2_X1 U14074 ( .A1(n18955), .A2(n10928), .ZN(n16155) );
  INV_X1 U14075 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11143) );
  NOR2_X1 U14076 ( .A1(n10803), .A2(n11143), .ZN(n10929) );
  NAND2_X1 U14077 ( .A1(n10930), .A2(n10929), .ZN(n10933) );
  NOR2_X1 U14078 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n10931) );
  NAND2_X1 U14079 ( .A1(n10933), .A2(n10943), .ZN(n10935) );
  INV_X1 U14080 ( .A(n10935), .ZN(n18944) );
  AND2_X1 U14081 ( .A1(n12496), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10934) );
  NAND2_X1 U14082 ( .A1(n18944), .A2(n10934), .ZN(n15271) );
  INV_X1 U14083 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15287) );
  OAI21_X1 U14084 ( .B1(n10935), .B2(n12494), .A(n15287), .ZN(n15272) );
  INV_X1 U14085 ( .A(n10943), .ZN(n10936) );
  INV_X1 U14086 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14149) );
  NAND2_X1 U14087 ( .A1(n10936), .A2(n14149), .ZN(n10939) );
  INV_X1 U14088 ( .A(n12473), .ZN(n10937) );
  AOI21_X1 U14089 ( .B1(n10943), .B2(n10942), .A(n10937), .ZN(n10938) );
  NAND2_X1 U14090 ( .A1(n18930), .A2(n12496), .ZN(n10940) );
  XNOR2_X1 U14091 ( .A(n10940), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15259) );
  NAND2_X1 U14092 ( .A1(n15260), .A2(n15259), .ZN(n15258) );
  AND2_X1 U14093 ( .A1(n12496), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10941) );
  NAND2_X1 U14094 ( .A1(n18930), .A2(n10941), .ZN(n12435) );
  NAND2_X1 U14095 ( .A1(n15258), .A2(n12435), .ZN(n15123) );
  NAND2_X1 U14096 ( .A1(n19300), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10944) );
  OAI21_X1 U14097 ( .B1(n10945), .B2(n10944), .A(n10954), .ZN(n18922) );
  INV_X1 U14098 ( .A(n10948), .ZN(n10946) );
  NAND2_X1 U14099 ( .A1(n10946), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12437) );
  INV_X1 U14100 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10947) );
  NAND2_X1 U14101 ( .A1(n10948), .A2(n10947), .ZN(n12451) );
  INV_X1 U14102 ( .A(n12437), .ZN(n10949) );
  AOI21_X1 U14103 ( .B1(n15123), .B2(n15122), .A(n10949), .ZN(n12392) );
  INV_X1 U14104 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11165) );
  INV_X1 U14105 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11159) );
  INV_X1 U14106 ( .A(n10956), .ZN(n10950) );
  XNOR2_X1 U14107 ( .A(n10957), .B(n10950), .ZN(n18898) );
  NAND2_X1 U14108 ( .A1(n18898), .A2(n12496), .ZN(n10960) );
  INV_X1 U14109 ( .A(n10960), .ZN(n10951) );
  NAND2_X1 U14110 ( .A1(n10951), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14261) );
  INV_X1 U14111 ( .A(n10952), .ZN(n10953) );
  XNOR2_X1 U14112 ( .A(n10954), .B(n10953), .ZN(n18910) );
  AND2_X1 U14113 ( .A1(n12496), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10955) );
  NAND2_X1 U14114 ( .A1(n18910), .A2(n10955), .ZN(n14258) );
  AND2_X1 U14115 ( .A1(n14261), .A2(n14258), .ZN(n12439) );
  NAND2_X1 U14116 ( .A1(n12392), .A2(n12439), .ZN(n15107) );
  NOR2_X2 U14117 ( .A1(n10957), .A2(n10956), .ZN(n10964) );
  INV_X1 U14118 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11172) );
  XNOR2_X1 U14119 ( .A(n10964), .B(n10958), .ZN(n14873) );
  NAND2_X1 U14120 ( .A1(n14873), .A2(n12496), .ZN(n10959) );
  INV_X1 U14121 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15229) );
  NAND2_X1 U14122 ( .A1(n10959), .A2(n15229), .ZN(n15109) );
  INV_X1 U14123 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15112) );
  NAND2_X1 U14124 ( .A1(n10960), .A2(n15112), .ZN(n14260) );
  NAND2_X1 U14125 ( .A1(n18910), .A2(n12496), .ZN(n10961) );
  NAND2_X1 U14126 ( .A1(n10961), .A2(n12422), .ZN(n12394) );
  AND2_X1 U14127 ( .A1(n14260), .A2(n12394), .ZN(n15106) );
  AND2_X1 U14128 ( .A1(n15109), .A2(n15106), .ZN(n12452) );
  AND2_X1 U14129 ( .A1(n12496), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10962) );
  NAND2_X1 U14130 ( .A1(n14873), .A2(n10962), .ZN(n15108) );
  INV_X1 U14131 ( .A(n15108), .ZN(n10963) );
  NAND2_X1 U14132 ( .A1(n10964), .A2(n11172), .ZN(n10966) );
  OR2_X2 U14133 ( .A1(n10966), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12445) );
  INV_X1 U14134 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11175) );
  NOR2_X1 U14135 ( .A1(n10803), .A2(n11175), .ZN(n10965) );
  AND2_X1 U14136 ( .A1(n10966), .A2(n10965), .ZN(n10967) );
  NOR2_X1 U14137 ( .A1(n12443), .A2(n10967), .ZN(n14858) );
  NAND2_X1 U14138 ( .A1(n14858), .A2(n12496), .ZN(n10968) );
  NAND2_X1 U14139 ( .A1(n10968), .A2(n15212), .ZN(n12454) );
  INV_X1 U14140 ( .A(n14858), .ZN(n10970) );
  NAND2_X1 U14141 ( .A1(n12496), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10969) );
  NAND2_X1 U14142 ( .A1(n12454), .A2(n12440), .ZN(n10971) );
  XNOR2_X1 U14143 ( .A(n10972), .B(n10971), .ZN(n15105) );
  INV_X1 U14144 ( .A(n10985), .ZN(n11005) );
  OAI21_X1 U14145 ( .B1(n10974), .B2(n11005), .A(n10973), .ZN(n10981) );
  AND2_X1 U14146 ( .A1(n16336), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10977) );
  AOI21_X1 U14147 ( .B1(n10981), .B2(n11011), .A(n11016), .ZN(n19954) );
  AND2_X1 U14148 ( .A1(n19283), .A2(n19968), .ZN(n13231) );
  INV_X1 U14149 ( .A(n13231), .ZN(n10983) );
  NOR2_X1 U14150 ( .A1(n10982), .A2(n10983), .ZN(n19957) );
  NAND2_X1 U14151 ( .A1(n19954), .A2(n19957), .ZN(n10998) );
  XNOR2_X1 U14152 ( .A(n10985), .B(n10984), .ZN(n11002) );
  AND2_X1 U14153 ( .A1(n10999), .A2(n11002), .ZN(n10986) );
  NAND2_X1 U14154 ( .A1(n11011), .A2(n10986), .ZN(n10988) );
  INV_X1 U14155 ( .A(n11016), .ZN(n10987) );
  INV_X1 U14156 ( .A(n11004), .ZN(n11003) );
  NAND3_X1 U14157 ( .A1(n11011), .A2(n10999), .A3(n11003), .ZN(n10989) );
  NAND3_X1 U14158 ( .A1(n16339), .A2(n15374), .A3(n10989), .ZN(n10994) );
  NAND2_X1 U14159 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12945) );
  INV_X1 U14160 ( .A(n12945), .ZN(n10990) );
  NAND2_X1 U14161 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n10990), .ZN(
        n10991) );
  NAND2_X1 U14162 ( .A1(n10991), .A2(n16358), .ZN(n16350) );
  INV_X1 U14163 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18876) );
  OAI21_X1 U14164 ( .B1(n10768), .B2(n16350), .A(n18876), .ZN(n10992) );
  AND2_X1 U14165 ( .A1(n10992), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19947) );
  INV_X1 U14166 ( .A(n19947), .ZN(n10993) );
  INV_X1 U14167 ( .A(n19956), .ZN(n10996) );
  INV_X1 U14168 ( .A(n10982), .ZN(n10995) );
  NAND3_X1 U14169 ( .A1(n10996), .A2(n10995), .A3(n11191), .ZN(n10997) );
  NAND2_X1 U14170 ( .A1(n10998), .A2(n10997), .ZN(n12398) );
  NAND2_X1 U14171 ( .A1(n19967), .A2(n11191), .ZN(n11000) );
  MUX2_X1 U14172 ( .A(n11000), .B(n11040), .S(n10999), .Z(n11010) );
  OAI211_X1 U14173 ( .C1(n11191), .C2(n11003), .A(n16351), .B(n11002), .ZN(
        n11007) );
  OAI21_X1 U14174 ( .B1(n11005), .B2(n11004), .A(n10568), .ZN(n11006) );
  OAI211_X1 U14175 ( .C1(n11001), .C2(n11008), .A(n11007), .B(n11006), .ZN(
        n11009) );
  NAND3_X1 U14176 ( .A1(n11010), .A2(n11011), .A3(n11009), .ZN(n11014) );
  INV_X1 U14177 ( .A(n11011), .ZN(n11012) );
  AOI21_X1 U14178 ( .B1(n10568), .B2(n11012), .A(n11016), .ZN(n11013) );
  NAND2_X1 U14179 ( .A1(n11014), .A2(n11013), .ZN(n11015) );
  MUX2_X1 U14180 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11015), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11020) );
  NAND2_X1 U14181 ( .A1(n16344), .A2(n11191), .ZN(n13396) );
  INV_X1 U14182 ( .A(n13396), .ZN(n11018) );
  NAND2_X1 U14183 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19822) );
  INV_X1 U14184 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18871) );
  NOR2_X1 U14185 ( .A1(n18871), .A2(n19852), .ZN(n19845) );
  NAND2_X1 U14186 ( .A1(n18871), .A2(n19852), .ZN(n19847) );
  INV_X1 U14187 ( .A(n19847), .ZN(n19837) );
  NOR3_X1 U14188 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19845), .A3(n19837), 
        .ZN(n19970) );
  NAND2_X1 U14189 ( .A1(n19822), .A2(n19970), .ZN(n13363) );
  INV_X1 U14190 ( .A(n13363), .ZN(n16345) );
  NAND3_X1 U14191 ( .A1(n11018), .A2(n11078), .A3(n16345), .ZN(n11036) );
  AOI21_X1 U14192 ( .B1(n11020), .B2(n16351), .A(n11019), .ZN(n11034) );
  NAND2_X1 U14193 ( .A1(n11201), .A2(n10499), .ZN(n11021) );
  NAND2_X1 U14194 ( .A1(n11021), .A2(n10544), .ZN(n11022) );
  NAND2_X1 U14195 ( .A1(n9710), .A2(n11022), .ZN(n11027) );
  AOI21_X1 U14196 ( .B1(n19968), .B2(n10547), .A(n11078), .ZN(n11024) );
  NAND2_X1 U14197 ( .A1(n11023), .A2(n19283), .ZN(n11091) );
  AOI21_X1 U14198 ( .B1(n11024), .B2(n11091), .A(n11077), .ZN(n11026) );
  NAND2_X1 U14199 ( .A1(n11029), .A2(n10547), .ZN(n11025) );
  NAND2_X1 U14200 ( .A1(n11025), .A2(n13231), .ZN(n11083) );
  NAND3_X1 U14201 ( .A1(n11027), .A2(n11026), .A3(n11083), .ZN(n11092) );
  NAND3_X1 U14202 ( .A1(n10553), .A2(n16339), .A3(n16345), .ZN(n11028) );
  OAI21_X1 U14203 ( .B1(n11029), .B2(n10499), .A(n11028), .ZN(n11030) );
  NOR2_X1 U14204 ( .A1(n11092), .A2(n11030), .ZN(n13365) );
  MUX2_X1 U14205 ( .A(n10553), .B(n11078), .S(n19283), .Z(n11031) );
  NAND3_X1 U14206 ( .A1(n11031), .A2(n16339), .A3(n19822), .ZN(n11032) );
  NAND2_X1 U14207 ( .A1(n13365), .A2(n11032), .ZN(n11033) );
  AOI21_X1 U14208 ( .B1(n11034), .B2(n13396), .A(n11033), .ZN(n11035) );
  NAND2_X1 U14209 ( .A1(n11036), .A2(n11035), .ZN(n11037) );
  NAND2_X1 U14210 ( .A1(n15374), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19828) );
  INV_X1 U14211 ( .A(n19828), .ZN(n11038) );
  NOR2_X1 U14212 ( .A1(n10982), .A2(n11040), .ZN(n19955) );
  XOR2_X1 U14213 ( .A(n11210), .B(n11042), .Z(n13422) );
  NAND2_X1 U14214 ( .A1(n11043), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13358) );
  XOR2_X1 U14215 ( .A(n11044), .B(n13356), .Z(n11045) );
  NOR2_X1 U14216 ( .A1(n13358), .A2(n11045), .ZN(n11046) );
  INV_X1 U14217 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14379) );
  XNOR2_X1 U14218 ( .A(n13358), .B(n11045), .ZN(n14378) );
  NOR2_X1 U14219 ( .A1(n14379), .A2(n14378), .ZN(n14377) );
  NOR2_X1 U14220 ( .A1(n11046), .A2(n14377), .ZN(n11047) );
  XNOR2_X1 U14221 ( .A(n13572), .B(n11047), .ZN(n13421) );
  NOR2_X1 U14222 ( .A1(n13422), .A2(n13421), .ZN(n13420) );
  NOR2_X1 U14223 ( .A1(n11047), .A2(n13572), .ZN(n11048) );
  OR2_X1 U14224 ( .A1(n13420), .A2(n11048), .ZN(n11049) );
  INV_X1 U14225 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16231) );
  XNOR2_X1 U14226 ( .A(n11049), .B(n16231), .ZN(n16229) );
  NAND2_X1 U14227 ( .A1(n11049), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11050) );
  NAND2_X1 U14228 ( .A1(n11054), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11053) );
  NAND2_X1 U14229 ( .A1(n11052), .A2(n11051), .ZN(n14037) );
  INV_X1 U14230 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14094) );
  INV_X1 U14231 ( .A(n11056), .ZN(n11058) );
  NAND2_X1 U14232 ( .A1(n15132), .A2(n16297), .ZN(n11066) );
  INV_X1 U14233 ( .A(n15132), .ZN(n11067) );
  NAND2_X1 U14234 ( .A1(n11067), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11068) );
  NAND2_X1 U14235 ( .A1(n11071), .A2(n12496), .ZN(n11070) );
  XNOR2_X1 U14236 ( .A(n11070), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16202) );
  NAND3_X1 U14237 ( .A1(n11071), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n12496), .ZN(n11072) );
  AND2_X1 U14238 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15336) );
  NAND2_X1 U14239 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15336), .ZN(
        n11367) );
  AND2_X1 U14240 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16261) );
  NAND2_X1 U14241 ( .A1(n16261), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16259) );
  NAND3_X1 U14242 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11073) );
  NOR2_X1 U14243 ( .A1(n16259), .A2(n11073), .ZN(n12423) );
  NAND2_X1 U14244 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n12423), .ZN(
        n14266) );
  NOR2_X1 U14245 ( .A1(n11367), .A2(n14266), .ZN(n12400) );
  NAND3_X1 U14246 ( .A1(n12400), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12577) );
  INV_X1 U14247 ( .A(n12577), .ZN(n11074) );
  NAND2_X1 U14248 ( .A1(n12591), .A2(n11074), .ZN(n15114) );
  AOI21_X1 U14249 ( .B1(n15212), .B2(n15114), .A(n15207), .ZN(n15103) );
  NAND2_X1 U14250 ( .A1(n11189), .A2(n19957), .ZN(n16307) );
  NOR2_X1 U14251 ( .A1(n10051), .A2(n11001), .ZN(n11075) );
  NAND2_X1 U14252 ( .A1(n11076), .A2(n11075), .ZN(n13144) );
  INV_X1 U14253 ( .A(n13142), .ZN(n13352) );
  OAI21_X1 U14254 ( .B1(n11077), .B2(n10499), .A(n13352), .ZN(n11080) );
  NAND2_X1 U14255 ( .A1(n11078), .A2(n19968), .ZN(n11079) );
  AND4_X1 U14256 ( .A1(n11081), .A2(n13144), .A3(n11080), .A4(n11079), .ZN(
        n11087) );
  NAND2_X1 U14257 ( .A1(n11082), .A2(n11191), .ZN(n13996) );
  NAND2_X1 U14258 ( .A1(n13996), .A2(n11083), .ZN(n11085) );
  NAND2_X1 U14259 ( .A1(n11085), .A2(n11084), .ZN(n11086) );
  NAND2_X1 U14260 ( .A1(n11087), .A2(n11086), .ZN(n11088) );
  AOI21_X1 U14261 ( .B1(n11089), .B2(n10579), .A(n11088), .ZN(n13720) );
  INV_X1 U14262 ( .A(n13728), .ZN(n13434) );
  NAND2_X1 U14263 ( .A1(n13720), .A2(n13434), .ZN(n11090) );
  NAND2_X1 U14264 ( .A1(n11189), .A2(n11090), .ZN(n15249) );
  NAND2_X1 U14265 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14385) );
  NOR2_X1 U14266 ( .A1(n13572), .A2(n14385), .ZN(n13574) );
  OR2_X1 U14267 ( .A1(n15249), .A2(n13574), .ZN(n13579) );
  NAND2_X1 U14268 ( .A1(n11189), .A2(n13143), .ZN(n15245) );
  NAND2_X1 U14269 ( .A1(n13572), .A2(n14385), .ZN(n13573) );
  NOR2_X1 U14270 ( .A1(n15245), .A2(n13573), .ZN(n13568) );
  INV_X1 U14271 ( .A(n13568), .ZN(n11094) );
  INV_X1 U14272 ( .A(n11189), .ZN(n11093) );
  NOR2_X2 U14273 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19934) );
  NAND2_X1 U14274 ( .A1(n19934), .A2(n15374), .ZN(n18868) );
  INV_X1 U14275 ( .A(n18868), .ZN(n13350) );
  AND2_X1 U14276 ( .A1(n13350), .A2(n19969), .ZN(n12404) );
  NAND2_X1 U14277 ( .A1(n11093), .A2(n9722), .ZN(n14380) );
  NAND2_X1 U14278 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11096), .ZN(
        n16311) );
  NAND2_X1 U14279 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14091) );
  NOR2_X1 U14280 ( .A1(n16311), .A2(n14091), .ZN(n11095) );
  NAND2_X1 U14281 ( .A1(n11095), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11097) );
  INV_X1 U14282 ( .A(n15247), .ZN(n15253) );
  NAND2_X1 U14283 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16288) );
  AND2_X1 U14284 ( .A1(n14099), .A2(n16288), .ZN(n11098) );
  INV_X1 U14285 ( .A(n15349), .ZN(n11100) );
  NAND2_X1 U14286 ( .A1(n15247), .A2(n12577), .ZN(n11099) );
  NAND2_X1 U14287 ( .A1(n11100), .A2(n11099), .ZN(n15213) );
  NAND2_X1 U14288 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11104) );
  AOI22_X1 U14289 ( .A1(n12543), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11103) );
  OAI211_X1 U14290 ( .C1(n12542), .C2(n10822), .A(n11104), .B(n11103), .ZN(
        n13743) );
  NAND2_X1 U14291 ( .A1(n13744), .A2(n13743), .ZN(n13745) );
  NAND2_X1 U14292 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11106) );
  AOI22_X1 U14293 ( .A1(n12543), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11105) );
  OAI211_X1 U14294 ( .C1(n13778), .C2(n12542), .A(n11106), .B(n11105), .ZN(
        n11107) );
  INV_X1 U14295 ( .A(n11107), .ZN(n13777) );
  NAND2_X1 U14296 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11112) );
  NAND2_X1 U14297 ( .A1(n12543), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11109) );
  NAND2_X1 U14298 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11108) );
  OAI211_X1 U14299 ( .C1(n12542), .C2(n19035), .A(n11109), .B(n11108), .ZN(
        n11110) );
  INV_X1 U14300 ( .A(n11110), .ZN(n11111) );
  NAND2_X1 U14301 ( .A1(n11112), .A2(n11111), .ZN(n13788) );
  NAND2_X1 U14302 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11114) );
  AOI22_X1 U14303 ( .A1(n12543), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11113) );
  OAI211_X1 U14304 ( .C1(n12542), .C2(n13819), .A(n11114), .B(n11113), .ZN(
        n13817) );
  NAND2_X1 U14305 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11116) );
  AOI22_X1 U14306 ( .A1(n12543), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11115) );
  OAI211_X1 U14307 ( .C1(n11117), .C2(n12542), .A(n11116), .B(n11115), .ZN(
        n13801) );
  INV_X1 U14308 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15350) );
  AOI22_X1 U14309 ( .A1(n12543), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11118) );
  OAI211_X1 U14310 ( .C1(n9892), .C2(n12542), .A(n11119), .B(n11118), .ZN(
        n11120) );
  INV_X1 U14311 ( .A(n11120), .ZN(n13797) );
  NAND2_X1 U14312 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11122) );
  AOI22_X1 U14313 ( .A1(n12543), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11121) );
  OAI211_X1 U14314 ( .C1(n12542), .C2(n18991), .A(n11122), .B(n11121), .ZN(
        n13881) );
  NAND2_X1 U14315 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11124) );
  AOI22_X1 U14316 ( .A1(n12543), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11123) );
  OAI211_X1 U14317 ( .C1(n13950), .C2(n12542), .A(n11124), .B(n11123), .ZN(
        n11125) );
  INV_X1 U14318 ( .A(n11125), .ZN(n13947) );
  INV_X1 U14319 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11128) );
  NAND2_X1 U14320 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11127) );
  AOI22_X1 U14321 ( .A1(n12543), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11126) );
  OAI211_X1 U14322 ( .C1(n11128), .C2(n12542), .A(n11127), .B(n11126), .ZN(
        n14341) );
  NAND2_X1 U14323 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14324 ( .A1(n12543), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11130) );
  NAND2_X1 U14325 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11129) );
  OAI211_X1 U14326 ( .C1(n12542), .C2(n11131), .A(n11130), .B(n11129), .ZN(
        n11132) );
  INV_X1 U14327 ( .A(n11132), .ZN(n11133) );
  NAND2_X1 U14328 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11140) );
  INV_X1 U14329 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11137) );
  NAND2_X1 U14330 ( .A1(n12543), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14331 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11135) );
  OAI211_X1 U14332 ( .C1(n12542), .C2(n11137), .A(n11136), .B(n11135), .ZN(
        n11138) );
  INV_X1 U14333 ( .A(n11138), .ZN(n11139) );
  NAND2_X1 U14334 ( .A1(n11140), .A2(n11139), .ZN(n14014) );
  NAND2_X1 U14335 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11146) );
  NAND2_X1 U14336 ( .A1(n12543), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11142) );
  NAND2_X1 U14337 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11141) );
  OAI211_X1 U14338 ( .C1(n12542), .C2(n11143), .A(n11142), .B(n11141), .ZN(
        n11144) );
  INV_X1 U14339 ( .A(n11144), .ZN(n11145) );
  INV_X1 U14340 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11149) );
  NAND2_X1 U14341 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11148) );
  AOI22_X1 U14342 ( .A1(n12543), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11147) );
  OAI211_X1 U14343 ( .C1(n12542), .C2(n11149), .A(n11148), .B(n11147), .ZN(
        n14122) );
  INV_X1 U14344 ( .A(n14122), .ZN(n11155) );
  NAND2_X1 U14345 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11154) );
  NAND2_X1 U14346 ( .A1(n12543), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U14347 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11150) );
  OAI211_X1 U14348 ( .C1(n12542), .C2(n14149), .A(n11151), .B(n11150), .ZN(
        n11152) );
  INV_X1 U14349 ( .A(n11152), .ZN(n11153) );
  NAND2_X1 U14350 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11162) );
  NAND2_X1 U14351 ( .A1(n12543), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11158) );
  NAND2_X1 U14352 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11157) );
  OAI211_X1 U14353 ( .C1(n12542), .C2(n11159), .A(n11158), .B(n11157), .ZN(
        n11160) );
  INV_X1 U14354 ( .A(n11160), .ZN(n11161) );
  AND2_X1 U14355 ( .A1(n11162), .A2(n11161), .ZN(n14235) );
  NAND2_X1 U14356 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11168) );
  NAND2_X1 U14357 ( .A1(n12543), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11164) );
  NAND2_X1 U14358 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11163) );
  OAI211_X1 U14359 ( .C1(n12542), .C2(n11165), .A(n11164), .B(n11163), .ZN(
        n11166) );
  INV_X1 U14360 ( .A(n11166), .ZN(n11167) );
  NAND2_X1 U14361 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11171) );
  AOI22_X1 U14362 ( .A1(n12543), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11170) );
  OAI211_X1 U14363 ( .C1(n12542), .C2(n11172), .A(n11171), .B(n11170), .ZN(
        n14151) );
  NAND2_X1 U14364 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11178) );
  NAND2_X1 U14365 ( .A1(n12543), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U14366 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11173) );
  OAI211_X1 U14367 ( .C1(n12542), .C2(n11175), .A(n11174), .B(n11173), .ZN(
        n11176) );
  INV_X1 U14368 ( .A(n11176), .ZN(n11177) );
  OR2_X1 U14369 ( .A1(n12510), .A2(n12508), .ZN(n14941) );
  NAND2_X1 U14370 ( .A1(n12510), .A2(n12508), .ZN(n11179) );
  NAND2_X1 U14371 ( .A1(n14941), .A2(n11179), .ZN(n15101) );
  NAND2_X1 U14372 ( .A1(n11180), .A2(n19283), .ZN(n11182) );
  INV_X1 U14373 ( .A(n13729), .ZN(n11181) );
  NAND2_X1 U14374 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  INV_X1 U14375 ( .A(n9722), .ZN(n15077) );
  NAND2_X1 U14376 ( .A1(n15077), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15096) );
  AND2_X1 U14377 ( .A1(n11184), .A2(n11185), .ZN(n16341) );
  INV_X1 U14378 ( .A(n16341), .ZN(n13721) );
  NAND2_X1 U14379 ( .A1(n11186), .A2(n11191), .ZN(n11187) );
  NAND2_X1 U14380 ( .A1(n13721), .A2(n11187), .ZN(n11188) );
  AND2_X2 U14381 ( .A1(n11189), .A2(n11188), .ZN(n16281) );
  INV_X1 U14382 ( .A(n11190), .ZN(n13147) );
  INV_X1 U14383 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18888) );
  OR2_X1 U14384 ( .A1(n11211), .A2(n18888), .ZN(n11195) );
  INV_X1 U14385 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13554) );
  NAND2_X1 U14386 ( .A1(n11191), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11192) );
  OAI211_X1 U14387 ( .C1(n10547), .C2(n13554), .A(n11192), .B(n19533), .ZN(
        n11193) );
  INV_X1 U14388 ( .A(n11193), .ZN(n11194) );
  NAND2_X1 U14389 ( .A1(n11195), .A2(n11194), .ZN(n13535) );
  MUX2_X1 U14390 ( .A(n10547), .B(n19950), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11197) );
  AND2_X1 U14391 ( .A1(n11196), .A2(n19533), .ZN(n11232) );
  NAND2_X1 U14392 ( .A1(n13146), .A2(n11232), .ZN(n11208) );
  AND2_X1 U14393 ( .A1(n11197), .A2(n11208), .ZN(n11198) );
  INV_X1 U14394 ( .A(n11232), .ZN(n11238) );
  INV_X1 U14395 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19210) );
  INV_X1 U14396 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19853) );
  OAI222_X1 U14397 ( .A1(n11238), .A2(n14379), .B1(n11350), .B2(n19210), .C1(
        n11211), .C2(n19853), .ZN(n11205) );
  NAND2_X1 U14398 ( .A1(n11201), .A2(n10547), .ZN(n11202) );
  MUX2_X1 U14399 ( .A(n11202), .B(n19943), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11203) );
  OAI21_X1 U14400 ( .B1(n11346), .B2(n11204), .A(n11203), .ZN(n13905) );
  NOR2_X1 U14401 ( .A1(n13906), .A2(n13905), .ZN(n11207) );
  NOR2_X1 U14402 ( .A1(n13534), .A2(n11205), .ZN(n11206) );
  NOR2_X2 U14403 ( .A1(n11207), .A2(n11206), .ZN(n11213) );
  NAND2_X1 U14404 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11209) );
  OAI211_X1 U14405 ( .C1(n11346), .C2(n11210), .A(n11209), .B(n11208), .ZN(
        n11212) );
  XNOR2_X1 U14406 ( .A(n11213), .B(n11212), .ZN(n13565) );
  INV_X1 U14407 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19208) );
  INV_X1 U14408 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19855) );
  OAI222_X1 U14409 ( .A1(n11238), .A2(n13572), .B1(n11350), .B2(n19208), .C1(
        n11211), .C2(n19855), .ZN(n13564) );
  NOR2_X1 U14410 ( .A1(n13565), .A2(n13564), .ZN(n13563) );
  INV_X1 U14411 ( .A(n13563), .ZN(n13707) );
  OR2_X1 U14412 ( .A1(n11213), .A2(n11212), .ZN(n13708) );
  INV_X1 U14413 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11214) );
  OR2_X1 U14414 ( .A1(n11211), .A2(n11214), .ZN(n11218) );
  AOI22_X1 U14415 ( .A1(n12564), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11216) );
  INV_X1 U14416 ( .A(n11350), .ZN(n12571) );
  NAND2_X1 U14417 ( .A1(n12571), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11215) );
  AND2_X1 U14418 ( .A1(n11216), .A2(n11215), .ZN(n11217) );
  OAI211_X1 U14419 ( .C1(n11346), .C2(n11219), .A(n11218), .B(n11217), .ZN(
        n13709) );
  AND2_X1 U14420 ( .A1(n13708), .A2(n13709), .ZN(n11220) );
  NAND2_X1 U14421 ( .A1(n13707), .A2(n11220), .ZN(n14040) );
  INV_X1 U14422 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11221) );
  OR2_X1 U14423 ( .A1(n11211), .A2(n11221), .ZN(n11225) );
  AOI22_X1 U14424 ( .A1(n12571), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12564), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11224) );
  OR2_X1 U14425 ( .A1(n11346), .A2(n11222), .ZN(n11223) );
  NOR2_X2 U14426 ( .A1(n14040), .A2(n14041), .ZN(n14098) );
  AOI22_X1 U14427 ( .A1(n12572), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11229) );
  INV_X1 U14428 ( .A(n11346), .ZN(n11227) );
  AOI22_X1 U14429 ( .A1(n11227), .A2(n11226), .B1(n12571), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U14430 ( .A1(n11229), .A2(n11228), .ZN(n14097) );
  NAND2_X1 U14431 ( .A1(n14098), .A2(n14097), .ZN(n14096) );
  OR2_X1 U14432 ( .A1(n11346), .A2(n11230), .ZN(n11231) );
  INV_X1 U14433 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19861) );
  OR2_X1 U14434 ( .A1(n11211), .A2(n19861), .ZN(n11234) );
  AOI22_X1 U14435 ( .A1(n12571), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12564), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11233) );
  NAND2_X1 U14436 ( .A1(n11234), .A2(n11233), .ZN(n15358) );
  AOI21_X1 U14437 ( .B1(n15359), .B2(n15358), .A(n11236), .ZN(n11237) );
  INV_X1 U14438 ( .A(n11237), .ZN(n16295) );
  INV_X1 U14439 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19196) );
  OAI222_X1 U14440 ( .A1(n16297), .A2(n11238), .B1(n11350), .B2(n19196), .C1(
        n11211), .C2(n19863), .ZN(n16294) );
  AOI22_X1 U14441 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11239), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14442 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14443 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14444 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12964), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11240) );
  NAND4_X1 U14445 ( .A1(n11243), .A2(n11242), .A3(n11241), .A4(n11240), .ZN(
        n11250) );
  AOI22_X1 U14446 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14447 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10775), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14448 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14449 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11245) );
  NAND4_X1 U14450 ( .A1(n11248), .A2(n11247), .A3(n11246), .A4(n11245), .ZN(
        n11249) );
  INV_X1 U14451 ( .A(n13808), .ZN(n11252) );
  AOI22_X1 U14452 ( .A1(n12571), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12564), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11251) );
  OAI21_X1 U14453 ( .B1(n11346), .B2(n11252), .A(n11251), .ZN(n11253) );
  AOI21_X1 U14454 ( .B1(n12572), .B2(P2_REIP_REG_8__SCAN_IN), .A(n11253), .ZN(
        n16280) );
  NOR2_X4 U14455 ( .A1(n16293), .A2(n16280), .ZN(n16279) );
  AOI22_X1 U14456 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12962), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14457 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n12963), .ZN(n11256) );
  AOI22_X1 U14458 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14459 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11254) );
  NAND4_X1 U14460 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11263) );
  AOI22_X1 U14461 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14462 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12970), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14463 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10775), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U14464 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11244), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11258) );
  NAND4_X1 U14465 ( .A1(n11261), .A2(n11260), .A3(n11259), .A4(n11258), .ZN(
        n11262) );
  NOR2_X1 U14466 ( .A1(n11263), .A2(n11262), .ZN(n12856) );
  INV_X1 U14467 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11264) );
  OR2_X1 U14468 ( .A1(n11211), .A2(n11264), .ZN(n11266) );
  AOI22_X1 U14469 ( .A1(n12571), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12564), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11265) );
  OAI211_X1 U14470 ( .C1(n11346), .C2(n12856), .A(n11266), .B(n11265), .ZN(
        n15352) );
  INV_X1 U14471 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11267) );
  OR2_X1 U14472 ( .A1(n11211), .A2(n11267), .ZN(n11280) );
  AOI22_X1 U14473 ( .A1(n12571), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U14474 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14475 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10775), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14476 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14477 ( .A1(n12971), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11268) );
  NAND4_X1 U14478 ( .A1(n11271), .A2(n11270), .A3(n11269), .A4(n11268), .ZN(
        n11277) );
  AOI22_X1 U14479 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U14480 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14481 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14482 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11272) );
  NAND4_X1 U14483 ( .A1(n11275), .A2(n11274), .A3(n11273), .A4(n11272), .ZN(
        n11276) );
  NOR2_X1 U14484 ( .A1(n11277), .A2(n11276), .ZN(n13879) );
  OR2_X1 U14485 ( .A1(n11346), .A2(n13879), .ZN(n11278) );
  AOI22_X1 U14486 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14487 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14488 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14489 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11281) );
  NAND4_X1 U14490 ( .A1(n11284), .A2(n11283), .A3(n11282), .A4(n11281), .ZN(
        n11290) );
  AOI22_X1 U14491 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11288) );
  AOI22_X1 U14492 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14493 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14494 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11285) );
  NAND4_X1 U14495 ( .A1(n11288), .A2(n11287), .A3(n11286), .A4(n11285), .ZN(
        n11289) );
  INV_X1 U14496 ( .A(n13943), .ZN(n11294) );
  INV_X1 U14497 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11291) );
  OR2_X1 U14498 ( .A1(n11211), .A2(n11291), .ZN(n11293) );
  AOI22_X1 U14499 ( .A1(n12571), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11292) );
  OAI211_X1 U14500 ( .C1(n11346), .C2(n11294), .A(n11293), .B(n11292), .ZN(
        n15335) );
  INV_X1 U14501 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11295) );
  OR2_X1 U14502 ( .A1(n11211), .A2(n11295), .ZN(n11309) );
  AOI22_X1 U14503 ( .A1(n12571), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14504 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12898), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14505 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10775), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11298) );
  AOI22_X1 U14506 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U14507 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11296) );
  NAND4_X1 U14508 ( .A1(n11299), .A2(n11298), .A3(n11297), .A4(n11296), .ZN(
        n11305) );
  AOI22_X1 U14509 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14510 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14511 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14512 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11300) );
  NAND4_X1 U14513 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n11304) );
  INV_X1 U14514 ( .A(n14345), .ZN(n11306) );
  OR2_X1 U14515 ( .A1(n11346), .A2(n11306), .ZN(n11307) );
  AOI22_X1 U14516 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14517 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14518 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14519 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11310) );
  NAND4_X1 U14520 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11319) );
  AOI22_X1 U14521 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14522 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14523 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14524 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11314) );
  NAND4_X1 U14525 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(
        n11318) );
  NOR2_X1 U14526 ( .A1(n11319), .A2(n11318), .ZN(n14006) );
  NAND2_X1 U14527 ( .A1(n12572), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14528 ( .A1(n12571), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11320) );
  OAI211_X1 U14529 ( .C1(n14006), .C2(n11346), .A(n11321), .B(n11320), .ZN(
        n14071) );
  AOI22_X1 U14530 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n12963), .ZN(n11325) );
  AOI22_X1 U14531 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14532 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n10723), .ZN(n11323) );
  AOI22_X1 U14533 ( .A1(n10768), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n12964), .ZN(n11322) );
  NAND4_X1 U14534 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11331) );
  AOI22_X1 U14535 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10722), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14536 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12970), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14537 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10775), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14538 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11244), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11326) );
  NAND4_X1 U14539 ( .A1(n11329), .A2(n11328), .A3(n11327), .A4(n11326), .ZN(
        n11330) );
  AOI22_X1 U14540 ( .A1(n12571), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11332) );
  OAI21_X1 U14541 ( .B1(n11346), .B2(n12862), .A(n11332), .ZN(n11333) );
  AOI21_X1 U14542 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n12572), .A(n11333), 
        .ZN(n16254) );
  AOI22_X1 U14543 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12962), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14544 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12963), .ZN(n11336) );
  AOI22_X1 U14545 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14546 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11334) );
  NAND4_X1 U14547 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11343) );
  AOI22_X1 U14548 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14549 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12970), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14550 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10775), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14551 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11244), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11338) );
  NAND4_X1 U14552 ( .A1(n11341), .A2(n11340), .A3(n11339), .A4(n11338), .ZN(
        n11342) );
  OR2_X1 U14553 ( .A1(n11343), .A2(n11342), .ZN(n14063) );
  INV_X1 U14554 ( .A(n14063), .ZN(n11347) );
  INV_X1 U14555 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n18940) );
  OR2_X1 U14556 ( .A1(n11211), .A2(n18940), .ZN(n11345) );
  AOI22_X1 U14557 ( .A1(n12571), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11344) );
  OAI211_X1 U14558 ( .C1(n11347), .C2(n11346), .A(n11345), .B(n11344), .ZN(
        n15279) );
  AND2_X2 U14559 ( .A1(n15280), .A2(n15279), .ZN(n15278) );
  INV_X1 U14560 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15264) );
  OR2_X1 U14561 ( .A1(n11211), .A2(n15264), .ZN(n11349) );
  AOI22_X1 U14562 ( .A1(n12571), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11348) );
  NAND2_X1 U14563 ( .A1(n11349), .A2(n11348), .ZN(n15262) );
  INV_X1 U14564 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n12405) );
  OR2_X1 U14565 ( .A1(n11211), .A2(n12405), .ZN(n11352) );
  AOI22_X1 U14566 ( .A1(n12571), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11351) );
  NAND2_X1 U14567 ( .A1(n11352), .A2(n11351), .ZN(n12424) );
  INV_X1 U14568 ( .A(n12424), .ZN(n11355) );
  INV_X1 U14569 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19877) );
  OR2_X1 U14570 ( .A1(n11211), .A2(n19877), .ZN(n11354) );
  AOI22_X1 U14571 ( .A1(n12571), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11353) );
  AND2_X1 U14572 ( .A1(n11354), .A2(n11353), .ZN(n15026) );
  OR2_X2 U14573 ( .A1(n15261), .A2(n11356), .ZN(n14264) );
  INV_X1 U14574 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15116) );
  OR2_X1 U14575 ( .A1(n11211), .A2(n15116), .ZN(n11358) );
  AOI22_X1 U14576 ( .A1(n12571), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11357) );
  AND2_X1 U14577 ( .A1(n11358), .A2(n11357), .ZN(n14861) );
  INV_X1 U14578 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19880) );
  OR2_X1 U14579 ( .A1(n11211), .A2(n19880), .ZN(n11360) );
  AOI22_X1 U14580 ( .A1(n12571), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11359) );
  AND2_X1 U14581 ( .A1(n11360), .A2(n11359), .ZN(n14263) );
  INV_X1 U14582 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19883) );
  OR2_X1 U14583 ( .A1(n11211), .A2(n19883), .ZN(n11363) );
  AOI22_X1 U14584 ( .A1(n12571), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11362) );
  NAND2_X1 U14585 ( .A1(n11363), .A2(n11362), .ZN(n11364) );
  OR2_X1 U14586 ( .A1(n14864), .A2(n11364), .ZN(n11365) );
  AND2_X1 U14587 ( .A1(n11365), .A2(n15217), .ZN(n15013) );
  NAND2_X1 U14588 ( .A1(n16281), .A2(n15013), .ZN(n11366) );
  OAI211_X1 U14589 ( .C1(n15101), .C2(n16283), .A(n15096), .B(n11366), .ZN(
        n11370) );
  INV_X1 U14590 ( .A(n11367), .ZN(n11369) );
  INV_X1 U14591 ( .A(n15245), .ZN(n13575) );
  OAI211_X1 U14592 ( .C1(n13575), .C2(n13574), .A(n13573), .B(n15247), .ZN(
        n11368) );
  INV_X1 U14593 ( .A(n11368), .ZN(n16312) );
  NAND2_X1 U14594 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16312), .ZN(
        n14092) );
  NOR2_X1 U14595 ( .A1(n14091), .A2(n14092), .ZN(n15362) );
  NAND2_X1 U14596 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15362), .ZN(
        n16287) );
  NAND2_X1 U14597 ( .A1(n11369), .A2(n15351), .ZN(n15319) );
  NOR2_X1 U14598 ( .A1(n15112), .A2(n14266), .ZN(n15230) );
  NAND3_X1 U14599 ( .A1(n16260), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15230), .ZN(n15211) );
  NOR2_X1 U14600 ( .A1(n15211), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15214) );
  AOI211_X1 U14601 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15213), .A(
        n11370), .B(n15214), .ZN(n11371) );
  OAI21_X1 U14602 ( .B1(n15105), .B2(n16315), .A(n11373), .ZN(P2_U3025) );
  INV_X1 U14603 ( .A(n11803), .ZN(n11374) );
  INV_X1 U14604 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14201) );
  INV_X1 U14605 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14514) );
  INV_X1 U14606 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12087) );
  INV_X1 U14607 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15713) );
  INV_X1 U14608 ( .A(n12161), .ZN(n11377) );
  INV_X1 U14609 ( .A(n12204), .ZN(n11380) );
  XNOR2_X1 U14610 ( .A(n13848), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14688) );
  INV_X1 U14611 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14612 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12103), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11386) );
  AOI22_X1 U14613 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11385) );
  AND2_X4 U14614 ( .A1(n11387), .A2(n13655), .ZN(n12004) );
  AND2_X4 U14615 ( .A1(n13673), .A2(n13655), .ZN(n12116) );
  AOI22_X1 U14616 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11384) );
  AND2_X2 U14617 ( .A1(n13655), .A2(n13647), .ZN(n11599) );
  AOI22_X1 U14618 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12097), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11383) );
  NAND4_X1 U14619 ( .A1(n11386), .A2(n11385), .A3(n11384), .A4(n11383), .ZN(
        n11397) );
  AOI22_X1 U14620 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11395) );
  AND2_X2 U14621 ( .A1(n11389), .A2(n13655), .ZN(n11537) );
  AOI22_X1 U14622 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11394) );
  AND3_X4 U14623 ( .A1(n13654), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n13473), .ZN(n11594) );
  AOI22_X1 U14624 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14625 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11392) );
  NAND4_X1 U14626 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(
        n11396) );
  NOR2_X1 U14627 ( .A1(n11397), .A2(n11396), .ZN(n12199) );
  AOI22_X1 U14628 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12103), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14629 ( .A1(n12102), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14630 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14631 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U14632 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11407) );
  AOI22_X1 U14633 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14634 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12125), .B1(
        n12097), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14635 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11594), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14636 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11402) );
  NAND4_X1 U14637 ( .A1(n11405), .A2(n11404), .A3(n11403), .A4(n11402), .ZN(
        n11406) );
  NOR2_X1 U14638 ( .A1(n11407), .A2(n11406), .ZN(n12178) );
  AOI22_X1 U14639 ( .A1(n12102), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14640 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14641 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14642 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11594), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11408) );
  NAND4_X1 U14643 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(
        n11417) );
  AOI22_X1 U14644 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14645 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12004), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14646 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14647 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11412) );
  NAND4_X1 U14648 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(
        n11416) );
  NOR2_X1 U14649 ( .A1(n11417), .A2(n11416), .ZN(n12157) );
  AOI22_X1 U14650 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14651 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U14652 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14653 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11418) );
  NAND4_X1 U14654 ( .A1(n11421), .A2(n11420), .A3(n11419), .A4(n11418), .ZN(
        n11427) );
  AOI22_X1 U14655 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14656 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14657 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14658 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11422) );
  NAND4_X1 U14659 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11426) );
  NOR2_X1 U14660 ( .A1(n11427), .A2(n11426), .ZN(n12140) );
  AOI22_X1 U14661 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14662 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14663 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14664 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11428) );
  NAND4_X1 U14665 ( .A1(n11431), .A2(n11430), .A3(n11429), .A4(n11428), .ZN(
        n11437) );
  AOI22_X1 U14666 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14667 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14668 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11594), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14669 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11432) );
  NAND4_X1 U14670 ( .A1(n11435), .A2(n11434), .A3(n11433), .A4(n11432), .ZN(
        n11436) );
  NOR2_X1 U14671 ( .A1(n11437), .A2(n11436), .ZN(n12139) );
  NOR2_X1 U14672 ( .A1(n12140), .A2(n12139), .ZN(n12151) );
  AOI22_X1 U14673 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14674 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14675 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14676 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11438) );
  NAND4_X1 U14677 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n11447) );
  AOI22_X1 U14678 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14679 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14680 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14681 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11442) );
  NAND4_X1 U14682 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11446) );
  OR2_X1 U14683 ( .A1(n11447), .A2(n11446), .ZN(n12150) );
  NAND2_X1 U14684 ( .A1(n12151), .A2(n12150), .ZN(n12158) );
  NOR2_X1 U14685 ( .A1(n12157), .A2(n12158), .ZN(n12168) );
  AOI22_X1 U14686 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14687 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14688 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14689 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11449) );
  NAND4_X1 U14690 ( .A1(n11452), .A2(n11451), .A3(n11450), .A4(n11449), .ZN(
        n11458) );
  AOI22_X1 U14691 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14692 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14693 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14694 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11453) );
  NAND4_X1 U14695 ( .A1(n11456), .A2(n11455), .A3(n11454), .A4(n11453), .ZN(
        n11457) );
  OR2_X1 U14696 ( .A1(n11458), .A2(n11457), .ZN(n12166) );
  NAND2_X1 U14697 ( .A1(n12168), .A2(n12166), .ZN(n12179) );
  NOR2_X1 U14698 ( .A1(n12178), .A2(n12179), .ZN(n12192) );
  AOI22_X1 U14699 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14700 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14701 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14702 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11459) );
  NAND4_X1 U14703 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n11469) );
  AOI22_X1 U14704 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11467) );
  AOI22_X1 U14705 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11466) );
  INV_X1 U14706 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14707 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14708 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11464) );
  NAND4_X1 U14709 ( .A1(n11467), .A2(n11466), .A3(n11465), .A4(n11464), .ZN(
        n11468) );
  OR2_X1 U14710 ( .A1(n11469), .A2(n11468), .ZN(n12191) );
  NAND2_X1 U14711 ( .A1(n12192), .A2(n12191), .ZN(n12200) );
  NOR2_X1 U14712 ( .A1(n12199), .A2(n12200), .ZN(n11481) );
  AOI22_X1 U14713 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14714 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14715 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14716 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11470) );
  NAND4_X1 U14717 ( .A1(n11473), .A2(n11472), .A3(n11471), .A4(n11470), .ZN(
        n11479) );
  AOI22_X1 U14718 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12023), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14719 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14720 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11474) );
  NAND4_X1 U14721 ( .A1(n11477), .A2(n11476), .A3(n11475), .A4(n11474), .ZN(
        n11478) );
  NOR2_X1 U14722 ( .A1(n11479), .A2(n11478), .ZN(n11480) );
  XOR2_X1 U14723 ( .A(n11481), .B(n11480), .Z(n11534) );
  AOI22_X1 U14724 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14725 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14726 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11646), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14727 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11482) );
  NAND4_X1 U14728 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11491) );
  AOI22_X1 U14729 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14730 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14731 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14732 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11567), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14733 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11490) );
  OR2_X2 U14734 ( .A1(n11491), .A2(n11490), .ZN(n11609) );
  NAND2_X1 U14735 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11495) );
  NAND2_X1 U14736 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11494) );
  NAND2_X1 U14737 ( .A1(n11567), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11493) );
  NAND2_X1 U14738 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11492) );
  NAND2_X1 U14739 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U14740 ( .A1(n11646), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11498) );
  NAND2_X1 U14741 ( .A1(n11542), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11497) );
  NAND2_X1 U14742 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11496) );
  NAND2_X1 U14743 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11503) );
  NAND2_X1 U14744 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11502) );
  NAND2_X1 U14745 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11501) );
  NAND2_X1 U14746 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14747 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11507) );
  NAND2_X1 U14748 ( .A1(n11647), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11506) );
  NAND2_X1 U14749 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11505) );
  NAND2_X1 U14750 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11504) );
  NAND4_X4 U14751 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n12209) );
  AOI22_X1 U14752 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14753 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11646), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14754 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14755 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11567), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11512) );
  NAND4_X1 U14756 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(
        n11521) );
  AOI22_X1 U14757 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14758 ( .A1(n11647), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14759 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14760 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11516) );
  NAND4_X1 U14761 ( .A1(n11519), .A2(n11518), .A3(n11517), .A4(n11516), .ZN(
        n11520) );
  AOI22_X1 U14762 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11599), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14763 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14764 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11567), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14765 ( .A1(n11646), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14766 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14767 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14768 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14769 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11528) );
  NAND2_X1 U14770 ( .A1(n11619), .A2(n11536), .ZN(n11611) );
  INV_X1 U14771 ( .A(n14829), .ZN(n11531) );
  NOR2_X1 U14772 ( .A1(n14425), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11532) );
  AOI211_X1 U14773 ( .C1(n12719), .C2(P1_EAX_REG_30__SCAN_IN), .A(n11532), .B(
        n12162), .ZN(n11533) );
  OAI21_X1 U14774 ( .B1(n11534), .B2(n12195), .A(n11533), .ZN(n11535) );
  OAI21_X1 U14775 ( .B1(n12198), .B2(n14688), .A(n11535), .ZN(n12208) );
  NAND2_X1 U14776 ( .A1(n11608), .A2(n11617), .ZN(n12212) );
  AOI22_X1 U14777 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14778 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14779 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11599), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14780 ( .A1(n11647), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14781 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14782 ( .A1(n11646), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14783 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14784 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11567), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11543) );
  NAND2_X1 U14785 ( .A1(n10090), .A2(n10091), .ZN(n11581) );
  INV_X2 U14786 ( .A(n11581), .ZN(n20213) );
  AOI21_X1 U14787 ( .B1(n11542), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n11547), .ZN(n11551) );
  AOI22_X1 U14788 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14789 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14790 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11567), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U14791 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11557) );
  AOI22_X1 U14792 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11646), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14793 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14794 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14795 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11552) );
  NAND4_X1 U14796 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11556) );
  NAND2_X1 U14797 ( .A1(n20213), .A2(n12600), .ZN(n12607) );
  INV_X1 U14798 ( .A(n12607), .ZN(n11558) );
  INV_X1 U14799 ( .A(n12764), .ZN(n11580) );
  NAND2_X1 U14800 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11562) );
  NAND2_X1 U14801 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11560) );
  NAND2_X1 U14802 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11559) );
  NAND2_X1 U14803 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11566) );
  NAND2_X1 U14804 ( .A1(n11646), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11565) );
  NAND2_X1 U14805 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11564) );
  NAND2_X1 U14806 ( .A1(n11647), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11563) );
  NAND2_X1 U14807 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11571) );
  NAND2_X1 U14808 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11570) );
  NAND2_X1 U14809 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11569) );
  NAND2_X1 U14810 ( .A1(n11567), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11568) );
  NAND2_X1 U14811 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11575) );
  NAND2_X1 U14812 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11574) );
  NAND2_X1 U14813 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11573) );
  NAND2_X1 U14814 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11572) );
  NAND4_X4 U14815 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n13854) );
  NAND2_X1 U14816 ( .A1(n11580), .A2(n13854), .ZN(n12785) );
  XNOR2_X1 U14817 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12761) );
  NOR2_X2 U14818 ( .A1(n11581), .A2(n12600), .ZN(n13662) );
  NAND2_X1 U14819 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11588) );
  NAND2_X1 U14820 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11586) );
  NAND2_X1 U14821 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11585) );
  NAND2_X1 U14822 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11593) );
  NAND2_X1 U14823 ( .A1(n11646), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11592) );
  NAND2_X1 U14824 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11591) );
  NAND2_X1 U14825 ( .A1(n11647), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11590) );
  NAND2_X1 U14826 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11598) );
  NAND2_X1 U14827 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11597) );
  NAND2_X1 U14828 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11596) );
  NAND2_X1 U14829 ( .A1(n11567), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11595) );
  NAND2_X1 U14830 ( .A1(n11537), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11603) );
  NAND2_X1 U14831 ( .A1(n11599), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11602) );
  NAND2_X1 U14832 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U14833 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11600) );
  NAND4_X4 U14835 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n13860) );
  NAND4_X1 U14836 ( .A1(n13662), .A2(n13852), .A3(n11608), .A4(n11790), .ZN(
        n12786) );
  OAI21_X1 U14837 ( .B1(n12785), .B2(n12761), .A(n12786), .ZN(n11616) );
  NAND2_X1 U14838 ( .A1(n11611), .A2(n11610), .ZN(n11612) );
  NAND2_X1 U14839 ( .A1(n12209), .A2(n11609), .ZN(n11613) );
  MUX2_X2 U14840 ( .A(n12778), .B(n11613), .S(n20213), .Z(n11614) );
  NAND2_X1 U14841 ( .A1(n11615), .A2(n11614), .ZN(n11618) );
  NOR2_X1 U14842 ( .A1(n11618), .A2(n15627), .ZN(n12722) );
  NAND2_X1 U14843 ( .A1(n12722), .A2(n13852), .ZN(n13677) );
  NAND2_X1 U14844 ( .A1(n13677), .A2(n12734), .ZN(n12777) );
  OAI21_X1 U14845 ( .B1(n11616), .B2(n12777), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11694) );
  NAND2_X1 U14846 ( .A1(n11581), .A2(n13854), .ZN(n12801) );
  NOR2_X1 U14847 ( .A1(n11636), .A2(n13662), .ZN(n11626) );
  NAND2_X1 U14848 ( .A1(n12792), .A2(n20196), .ZN(n11625) );
  NAND2_X1 U14849 ( .A1(n12336), .A2(n12607), .ZN(n12796) );
  NAND2_X1 U14850 ( .A1(n20196), .A2(n13860), .ZN(n13857) );
  INV_X1 U14851 ( .A(n11621), .ZN(n11622) );
  NAND2_X1 U14852 ( .A1(n11622), .A2(n20221), .ZN(n11623) );
  NAND2_X1 U14853 ( .A1(n11637), .A2(n14829), .ZN(n11624) );
  NAND2_X1 U14854 ( .A1(n16008), .A2(n20761), .ZN(n12714) );
  MUX2_X1 U14855 ( .A(n12714), .B(n12276), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11627) );
  OAI21_X1 U14856 ( .B1(n13852), .B2(n11628), .A(n12792), .ZN(n11640) );
  NAND2_X1 U14857 ( .A1(n13662), .A2(n20228), .ZN(n12800) );
  INV_X1 U14858 ( .A(n11630), .ZN(n11632) );
  INV_X1 U14859 ( .A(n11631), .ZN(n12677) );
  NAND2_X1 U14860 ( .A1(n11632), .A2(n12677), .ZN(n11634) );
  INV_X1 U14861 ( .A(n16008), .ZN(n14850) );
  NOR2_X1 U14862 ( .A1(n14850), .A2(n20761), .ZN(n11633) );
  NAND4_X1 U14863 ( .A1(n12800), .A2(n11634), .A3(n11633), .A4(n13857), .ZN(
        n11635) );
  NOR2_X1 U14864 ( .A1(n11636), .A2(n11635), .ZN(n11639) );
  NAND3_X1 U14865 ( .A1(n11637), .A2(n13860), .A3(n14829), .ZN(n11638) );
  NAND3_X1 U14866 ( .A1(n11640), .A2(n11639), .A3(n11638), .ZN(n11697) );
  INV_X1 U14867 ( .A(n11697), .ZN(n11641) );
  XNOR2_X1 U14868 ( .A(n11698), .B(n11641), .ZN(n11832) );
  NAND2_X1 U14869 ( .A1(n11832), .A2(n20761), .ZN(n11669) );
  AOI22_X1 U14870 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12103), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14871 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14872 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12097), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14873 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11642) );
  NAND4_X1 U14874 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11654) );
  AOI22_X1 U14875 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14876 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11650) );
  INV_X1 U14877 ( .A(n11647), .ZN(n11659) );
  INV_X1 U14878 ( .A(n11659), .ZN(n11648) );
  AOI22_X1 U14879 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11649) );
  NAND4_X1 U14880 ( .A1(n11652), .A2(n11651), .A3(n11650), .A4(n11649), .ZN(
        n11653) );
  AOI22_X1 U14881 ( .A1(n12004), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12103), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14882 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14883 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11655) );
  NAND4_X1 U14884 ( .A1(n11658), .A2(n11657), .A3(n11656), .A4(n11655), .ZN(
        n11666) );
  AOI22_X1 U14885 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12023), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14886 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14887 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12097), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14888 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11661) );
  NAND4_X1 U14889 ( .A1(n11664), .A2(n11663), .A3(n11662), .A4(n11661), .ZN(
        n11665) );
  XNOR2_X1 U14890 ( .A(n11671), .B(n12676), .ZN(n11667) );
  NAND2_X1 U14891 ( .A1(n11667), .A2(n11702), .ZN(n11668) );
  NAND2_X1 U14892 ( .A1(n11669), .A2(n11668), .ZN(n11830) );
  INV_X1 U14893 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11674) );
  NAND2_X1 U14894 ( .A1(n20221), .A2(n12676), .ZN(n11670) );
  OAI211_X1 U14895 ( .C1(n11671), .C2(n13854), .A(n11670), .B(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n11672) );
  INV_X1 U14896 ( .A(n11672), .ZN(n11673) );
  NAND2_X1 U14897 ( .A1(n11830), .A2(n11829), .ZN(n11676) );
  NAND2_X1 U14898 ( .A1(n11702), .A2(n12676), .ZN(n11675) );
  INV_X1 U14899 ( .A(n12676), .ZN(n11868) );
  NAND2_X1 U14900 ( .A1(n20196), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11736) );
  INV_X1 U14901 ( .A(n11736), .ZN(n11688) );
  AOI22_X1 U14902 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12125), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14903 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12023), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14904 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11678) );
  NAND4_X1 U14905 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11687) );
  AOI22_X1 U14906 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12103), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14907 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14908 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14909 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11682) );
  NAND4_X1 U14910 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11686) );
  AOI22_X1 U14911 ( .A1(n11702), .A2(n11868), .B1(n11688), .B2(n12606), .ZN(
        n11690) );
  NAND2_X1 U14912 ( .A1(n12270), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11689) );
  NAND2_X1 U14913 ( .A1(n11713), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11693) );
  NAND2_X1 U14914 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11716) );
  OAI21_X1 U14915 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11716), .ZN(n20519) );
  NAND2_X1 U14916 ( .A1(n15640), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11710) );
  OAI21_X1 U14917 ( .B1(n12714), .B2(n20519), .A(n11710), .ZN(n11691) );
  INV_X1 U14918 ( .A(n11691), .ZN(n11692) );
  NAND2_X1 U14919 ( .A1(n11693), .A2(n11692), .ZN(n11696) );
  XNOR2_X2 U14921 ( .A(n11696), .B(n11695), .ZN(n20297) );
  INV_X1 U14922 ( .A(n20297), .ZN(n11700) );
  INV_X1 U14923 ( .A(n11701), .ZN(n11699) );
  NAND2_X1 U14924 ( .A1(n11700), .A2(n11699), .ZN(n20243) );
  NAND2_X1 U14926 ( .A1(n20243), .A2(n11724), .ZN(n13934) );
  NAND2_X1 U14927 ( .A1(n11702), .A2(n12606), .ZN(n11703) );
  OAI21_X2 U14928 ( .B1(n13934), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11703), 
        .ZN(n11704) );
  INV_X1 U14929 ( .A(n11704), .ZN(n12605) );
  NAND2_X1 U14930 ( .A1(n11822), .A2(n12605), .ZN(n11709) );
  INV_X1 U14931 ( .A(n11705), .ZN(n11706) );
  NAND2_X1 U14932 ( .A1(n11709), .A2(n11708), .ZN(n11812) );
  INV_X1 U14933 ( .A(n11812), .ZN(n11741) );
  INV_X1 U14934 ( .A(n11695), .ZN(n11712) );
  NAND2_X1 U14935 ( .A1(n11710), .A2(n14831), .ZN(n11711) );
  NAND2_X1 U14936 ( .A1(n11712), .A2(n11711), .ZN(n11722) );
  NAND2_X1 U14937 ( .A1(n11724), .A2(n11722), .ZN(n11720) );
  INV_X1 U14939 ( .A(n12714), .ZN(n11743) );
  INV_X1 U14940 ( .A(n11716), .ZN(n11715) );
  NAND2_X1 U14941 ( .A1(n11715), .A2(n12247), .ZN(n20550) );
  NAND2_X1 U14942 ( .A1(n11716), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11717) );
  NAND2_X1 U14943 ( .A1(n20550), .A2(n11717), .ZN(n20205) );
  AND2_X1 U14944 ( .A1(n11743), .A2(n20205), .ZN(n11718) );
  NAND2_X1 U14945 ( .A1(n15640), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14946 ( .A1(n11723), .A2(n11721), .ZN(n11719) );
  NAND2_X1 U14947 ( .A1(n11720), .A2(n11719), .ZN(n11742) );
  NAND4_X1 U14948 ( .A1(n11724), .A2(n11723), .A3(n11722), .A4(n11721), .ZN(
        n11725) );
  NAND2_X1 U14949 ( .A1(n11742), .A2(n11725), .ZN(n13642) );
  AOI22_X1 U14950 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14951 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14952 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11726) );
  NAND4_X1 U14953 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11735) );
  AOI22_X1 U14954 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14955 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14956 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14957 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11730) );
  NAND4_X1 U14958 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n11734) );
  OAI22_X1 U14959 ( .A1(n13642), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12599), 
        .B2(n12671), .ZN(n11739) );
  OAI22_X1 U14960 ( .A1(n12259), .A2(n11737), .B1(n11736), .B2(n12599), .ZN(
        n11738) );
  XNOR2_X1 U14961 ( .A(n11739), .B(n11738), .ZN(n11813) );
  INV_X1 U14962 ( .A(n11813), .ZN(n11740) );
  NAND2_X2 U14963 ( .A1(n11741), .A2(n11740), .ZN(n11815) );
  NAND2_X1 U14964 ( .A1(n11714), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11745) );
  NOR3_X1 U14965 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12247), .A3(
        n20587), .ZN(n20425) );
  NAND2_X1 U14966 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20425), .ZN(
        n20420) );
  NAND3_X1 U14967 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20702) );
  NOR2_X1 U14968 ( .A1(n20628), .A2(n20702), .ZN(n20751) );
  AOI21_X1 U14969 ( .B1(n20420), .B2(n20549), .A(n20751), .ZN(n20455) );
  AOI22_X1 U14970 ( .A1(n20455), .A2(n11743), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15640), .ZN(n11744) );
  XNOR2_X2 U14971 ( .A(n13675), .B(n20336), .ZN(n13653) );
  INV_X1 U14972 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14973 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14974 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14975 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11749) );
  NAND4_X1 U14976 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n11758) );
  AOI22_X1 U14977 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14978 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14979 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14980 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11753) );
  NAND4_X1 U14981 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n11753), .ZN(
        n11757) );
  INV_X1 U14982 ( .A(n12632), .ZN(n11759) );
  OAI22_X1 U14983 ( .A1(n12259), .A2(n11760), .B1(n12268), .B2(n11759), .ZN(
        n11761) );
  OR2_X2 U14984 ( .A1(n11815), .A2(n11800), .ZN(n11802) );
  AOI22_X1 U14985 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12103), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14986 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12117), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14987 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11762) );
  NAND4_X1 U14988 ( .A1(n11765), .A2(n11764), .A3(n11763), .A4(n11762), .ZN(
        n11771) );
  AOI22_X1 U14989 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12024), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14990 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12023), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U14991 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14992 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11766) );
  NAND4_X1 U14993 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n11770) );
  AOI22_X1 U14994 ( .A1(n12270), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12232), .B2(n12642), .ZN(n11788) );
  NOR2_X2 U14995 ( .A1(n11802), .A2(n11788), .ZN(n11784) );
  AOI22_X1 U14996 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14997 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14998 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14999 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11772) );
  NAND4_X1 U15000 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11781) );
  AOI22_X1 U15001 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U15002 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U15003 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U15004 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11776) );
  NAND4_X1 U15005 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11780) );
  NAND2_X1 U15006 ( .A1(n12232), .A2(n12653), .ZN(n11782) );
  NAND2_X1 U15007 ( .A1(n11784), .A2(n11783), .ZN(n11864) );
  INV_X2 U15008 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20764) );
  INV_X1 U15009 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11786) );
  OAI21_X1 U15010 ( .B1(n11793), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n11858), .ZN(n20074) );
  AOI22_X1 U15011 ( .A1(n20074), .A2(n12162), .B1(n12718), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11785) );
  OAI21_X1 U15012 ( .B1(n12112), .B2(n11786), .A(n11785), .ZN(n11787) );
  AOI21_X1 U15013 ( .B1(n12641), .B2(n11994), .A(n11787), .ZN(n13814) );
  INV_X1 U15014 ( .A(n11788), .ZN(n11789) );
  XNOR2_X1 U15015 ( .A(n11802), .B(n11789), .ZN(n12631) );
  NAND2_X1 U15016 ( .A1(n11790), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11836) );
  INV_X1 U15017 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13674) );
  NAND2_X1 U15018 ( .A1(n20764), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11792) );
  NAND2_X1 U15019 ( .A1(n12719), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11791) );
  OAI211_X1 U15020 ( .C1(n11836), .C2(n13674), .A(n11792), .B(n11791), .ZN(
        n11798) );
  INV_X1 U15021 ( .A(n11793), .ZN(n11797) );
  INV_X1 U15022 ( .A(n11794), .ZN(n11806) );
  INV_X1 U15023 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11795) );
  NAND2_X1 U15024 ( .A1(n11806), .A2(n11795), .ZN(n11796) );
  NAND2_X1 U15025 ( .A1(n11797), .A2(n11796), .ZN(n20089) );
  MUX2_X1 U15026 ( .A(n11798), .B(n20089), .S(n12162), .Z(n11799) );
  AOI21_X1 U15027 ( .B1(n12631), .B2(n11994), .A(n11799), .ZN(n13813) );
  NAND2_X1 U15028 ( .A1(n11815), .A2(n11800), .ZN(n11801) );
  INV_X1 U15029 ( .A(n11994), .ZN(n11982) );
  NAND2_X1 U15030 ( .A1(n11804), .A2(n11803), .ZN(n11805) );
  NAND2_X1 U15031 ( .A1(n11806), .A2(n11805), .ZN(n20101) );
  AOI22_X1 U15032 ( .A1(n20101), .A2(n12162), .B1(n12718), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11808) );
  NAND2_X1 U15033 ( .A1(n12719), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11807) );
  OAI211_X1 U15034 ( .C1(n11836), .C2(n13669), .A(n11808), .B(n11807), .ZN(
        n11809) );
  INV_X1 U15035 ( .A(n11809), .ZN(n11810) );
  INV_X1 U15036 ( .A(n13752), .ZN(n11811) );
  NOR2_X1 U15037 ( .A1(n13813), .A2(n11811), .ZN(n11842) );
  NAND2_X1 U15038 ( .A1(n11813), .A2(n11812), .ZN(n11814) );
  NAND2_X1 U15039 ( .A1(n11815), .A2(n11814), .ZN(n12596) );
  XNOR2_X1 U15040 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13924) );
  AOI21_X1 U15041 ( .B1(n13843), .B2(n13924), .A(n12718), .ZN(n11818) );
  NAND2_X1 U15042 ( .A1(n12719), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11817) );
  OAI211_X1 U15043 ( .C1(n11836), .C2(n11816), .A(n11818), .B(n11817), .ZN(
        n11819) );
  INV_X1 U15044 ( .A(n11819), .ZN(n11820) );
  NAND2_X1 U15045 ( .A1(n12718), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11841) );
  INV_X1 U15046 ( .A(n11822), .ZN(n11823) );
  NAND2_X1 U15047 ( .A1(n9717), .A2(n11994), .ZN(n11828) );
  AOI22_X1 U15048 ( .A1(n12719), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20764), .ZN(n11826) );
  INV_X1 U15049 ( .A(n11836), .ZN(n11824) );
  NAND2_X1 U15050 ( .A1(n11824), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11825) );
  AND2_X1 U15051 ( .A1(n11826), .A2(n11825), .ZN(n11827) );
  NAND2_X1 U15052 ( .A1(n11828), .A2(n11827), .ZN(n13604) );
  NAND2_X1 U15053 ( .A1(n20579), .A2(n20228), .ZN(n11831) );
  NAND2_X1 U15054 ( .A1(n11831), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U15055 ( .A1(n20764), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11835) );
  NAND2_X1 U15056 ( .A1(n12719), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11834) );
  OAI211_X1 U15057 ( .C1(n11836), .C2(n13473), .A(n11835), .B(n11834), .ZN(
        n11837) );
  AOI21_X1 U15058 ( .B1(n11833), .B2(n11994), .A(n11837), .ZN(n11838) );
  OR2_X1 U15059 ( .A1(n13558), .A2(n11838), .ZN(n13559) );
  INV_X1 U15060 ( .A(n11838), .ZN(n13560) );
  OR2_X1 U15061 ( .A1(n13560), .A2(n12198), .ZN(n11839) );
  NAND2_X1 U15062 ( .A1(n13559), .A2(n11839), .ZN(n13603) );
  NAND2_X1 U15063 ( .A1(n13604), .A2(n13603), .ZN(n13608) );
  NAND3_X1 U15064 ( .A1(n11843), .A2(n11842), .A3(n13751), .ZN(n13812) );
  INV_X1 U15065 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U15066 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11542), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U15067 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U15068 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U15069 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11844) );
  NAND4_X1 U15070 ( .A1(n11847), .A2(n11846), .A3(n11845), .A4(n11844), .ZN(
        n11853) );
  AOI22_X1 U15071 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U15072 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U15073 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U15074 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11848) );
  NAND4_X1 U15075 ( .A1(n11851), .A2(n11850), .A3(n11849), .A4(n11848), .ZN(
        n11852) );
  NAND2_X1 U15076 ( .A1(n12232), .A2(n12662), .ZN(n11865) );
  OAI21_X1 U15077 ( .B1(n11854), .B2(n12259), .A(n11865), .ZN(n11855) );
  INV_X1 U15078 ( .A(n11855), .ZN(n11856) );
  NAND2_X1 U15079 ( .A1(n11864), .A2(n11856), .ZN(n12651) );
  INV_X1 U15080 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11862) );
  NAND2_X1 U15081 ( .A1(n11858), .A2(n11857), .ZN(n11860) );
  INV_X1 U15082 ( .A(n11871), .ZN(n11859) );
  NAND2_X1 U15083 ( .A1(n11860), .A2(n11859), .ZN(n20058) );
  AOI22_X1 U15084 ( .A1(n20058), .A2(n12162), .B1(n12718), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11861) );
  OAI21_X1 U15085 ( .B1(n12112), .B2(n11862), .A(n11861), .ZN(n11863) );
  INV_X1 U15086 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11869) );
  OAI22_X1 U15087 ( .A1(n12259), .A2(n11869), .B1(n12268), .B2(n11868), .ZN(
        n11870) );
  INV_X1 U15088 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11873) );
  OAI21_X1 U15089 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11871), .A(
        n11887), .ZN(n20047) );
  NAND2_X1 U15090 ( .A1(n20047), .A2(n12162), .ZN(n11872) );
  OAI21_X1 U15091 ( .B1(n11873), .B2(n12035), .A(n11872), .ZN(n11874) );
  AOI21_X1 U15092 ( .B1(n12719), .B2(P1_EAX_REG_7__SCAN_IN), .A(n11874), .ZN(
        n11875) );
  NAND2_X1 U15093 ( .A1(n13953), .A2(n13952), .ZN(n13951) );
  AOI22_X1 U15094 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U15095 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12097), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U15096 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11877) );
  NAND4_X1 U15097 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n11886) );
  AOI22_X1 U15098 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U15099 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U15100 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U15101 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11881) );
  NAND4_X1 U15102 ( .A1(n11884), .A2(n11883), .A3(n11882), .A4(n11881), .ZN(
        n11885) );
  OAI21_X1 U15103 ( .B1(n11886), .B2(n11885), .A(n11994), .ZN(n11891) );
  NAND2_X1 U15104 ( .A1(n12719), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11890) );
  XNOR2_X1 U15105 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11887), .ZN(
        n20032) );
  INV_X1 U15106 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20025) );
  OAI22_X1 U15107 ( .A1(n20032), .A2(n12198), .B1(n12035), .B2(n20025), .ZN(
        n11888) );
  INV_X1 U15108 ( .A(n11888), .ZN(n11889) );
  XNOR2_X1 U15109 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11893), .ZN(
        n20020) );
  INV_X1 U15110 ( .A(n20020), .ZN(n11908) );
  AOI22_X1 U15111 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12125), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U15112 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12103), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U15113 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U15114 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11894) );
  NAND4_X1 U15115 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n11903) );
  AOI22_X1 U15116 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U15117 ( .A1(n12102), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U15118 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12097), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11898) );
  NAND4_X1 U15119 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11902) );
  OAI21_X1 U15120 ( .B1(n11903), .B2(n11902), .A(n11994), .ZN(n11906) );
  NAND2_X1 U15121 ( .A1(n12719), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11905) );
  NAND2_X1 U15122 ( .A1(n12718), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11904) );
  NAND3_X1 U15123 ( .A1(n11906), .A2(n11905), .A3(n11904), .ZN(n11907) );
  AOI22_X1 U15124 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12125), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U15125 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12103), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U15126 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U15127 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11909) );
  NAND4_X1 U15128 ( .A1(n11912), .A2(n11911), .A3(n11910), .A4(n11909), .ZN(
        n11918) );
  AOI22_X1 U15129 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U15130 ( .A1(n12102), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15131 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15132 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12097), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11913) );
  NAND4_X1 U15133 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n11917) );
  NOR2_X1 U15134 ( .A1(n11918), .A2(n11917), .ZN(n11922) );
  XNOR2_X1 U15135 ( .A(n11919), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14190) );
  NAND2_X1 U15136 ( .A1(n14190), .A2(n12162), .ZN(n11921) );
  AOI22_X1 U15137 ( .A1(n12719), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12718), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11920) );
  OAI211_X1 U15138 ( .C1(n11922), .C2(n11982), .A(n11921), .B(n11920), .ZN(
        n14048) );
  AOI22_X1 U15139 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12023), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15140 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U15141 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15142 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U15143 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11932) );
  AOI22_X1 U15144 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12004), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15145 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15146 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U15147 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11927) );
  NAND4_X1 U15148 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11927), .ZN(
        n11931) );
  OR2_X1 U15149 ( .A1(n11932), .A2(n11931), .ZN(n11933) );
  NAND2_X1 U15150 ( .A1(n11994), .A2(n11933), .ZN(n14172) );
  INV_X1 U15151 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11936) );
  OAI21_X1 U15152 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11934), .A(
        n11964), .ZN(n15819) );
  NAND2_X1 U15153 ( .A1(n15819), .A2(n12162), .ZN(n11935) );
  OAI21_X1 U15154 ( .B1(n11936), .B2(n12035), .A(n11935), .ZN(n11937) );
  AOI21_X1 U15155 ( .B1(n12719), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11937), .ZN(
        n14141) );
  XNOR2_X1 U15156 ( .A(n11939), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15745) );
  AOI22_X1 U15157 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U15158 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U15159 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15160 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11940) );
  NAND4_X1 U15161 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11949) );
  AOI22_X1 U15162 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U15163 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12023), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U15164 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U15165 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11944) );
  NAND4_X1 U15166 ( .A1(n11947), .A2(n11946), .A3(n11945), .A4(n11944), .ZN(
        n11948) );
  OAI21_X1 U15167 ( .B1(n11949), .B2(n11948), .A(n11994), .ZN(n11952) );
  NAND2_X1 U15168 ( .A1(n12719), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U15169 ( .A1(n12718), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11950) );
  AND3_X1 U15170 ( .A1(n11952), .A2(n11951), .A3(n11950), .ZN(n11953) );
  OAI21_X1 U15171 ( .B1(n15745), .B2(n12198), .A(n11953), .ZN(n14159) );
  AOI22_X1 U15172 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12117), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15173 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12024), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U15174 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15175 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11954) );
  NAND4_X1 U15176 ( .A1(n11957), .A2(n11956), .A3(n11955), .A4(n11954), .ZN(
        n11963) );
  AOI22_X1 U15177 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12023), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15178 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12103), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11960) );
  AOI22_X1 U15179 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15180 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11958) );
  NAND4_X1 U15181 ( .A1(n11961), .A2(n11960), .A3(n11959), .A4(n11958), .ZN(
        n11962) );
  NOR2_X1 U15182 ( .A1(n11963), .A2(n11962), .ZN(n11969) );
  NAND2_X1 U15183 ( .A1(n12719), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11968) );
  XNOR2_X1 U15184 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11964), .ZN(
        n15808) );
  INV_X1 U15185 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11965) );
  OAI22_X1 U15186 ( .A1(n15808), .A2(n12198), .B1(n12035), .B2(n11965), .ZN(
        n11966) );
  INV_X1 U15187 ( .A(n11966), .ZN(n11967) );
  OAI211_X1 U15188 ( .C1(n11969), .C2(n11982), .A(n11968), .B(n11967), .ZN(
        n14160) );
  INV_X1 U15189 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14134) );
  XNOR2_X1 U15190 ( .A(n14134), .B(n11970), .ZN(n15798) );
  AOI22_X1 U15191 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15192 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U15193 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15194 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11971) );
  NAND4_X1 U15195 ( .A1(n11974), .A2(n11973), .A3(n11972), .A4(n11971), .ZN(
        n11980) );
  AOI22_X1 U15196 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15197 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15198 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15199 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U15200 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  NOR2_X1 U15201 ( .A1(n11980), .A2(n11979), .ZN(n11981) );
  OAI22_X1 U15202 ( .A1(n11982), .A2(n11981), .B1(n12035), .B2(n14134), .ZN(
        n11983) );
  AOI21_X1 U15203 ( .B1(n12719), .B2(P1_EAX_REG_14__SCAN_IN), .A(n11983), .ZN(
        n11984) );
  OAI21_X1 U15204 ( .B1(n15798), .B2(n12198), .A(n11984), .ZN(n14129) );
  XNOR2_X1 U15205 ( .A(n11985), .B(n14201), .ZN(n14230) );
  AOI22_X1 U15206 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15207 ( .A1(n12102), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15208 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U15209 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11986) );
  NAND4_X1 U15210 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n11996) );
  AOI22_X1 U15211 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12103), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15212 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12023), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15213 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15214 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11990) );
  NAND4_X1 U15215 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n11995) );
  OAI21_X1 U15216 ( .B1(n11996), .B2(n11995), .A(n11994), .ZN(n11999) );
  NAND2_X1 U15217 ( .A1(n12719), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11998) );
  NAND2_X1 U15218 ( .A1(n12718), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11997) );
  NAND3_X1 U15219 ( .A1(n11999), .A2(n11998), .A3(n11997), .ZN(n12000) );
  AOI21_X1 U15220 ( .B1(n14230), .B2(n13843), .A(n12000), .ZN(n14197) );
  INV_X1 U15221 ( .A(n14197), .ZN(n12001) );
  OR2_X1 U15222 ( .A1(n12002), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12003) );
  NAND2_X1 U15223 ( .A1(n12003), .A2(n12032), .ZN(n15789) );
  AOI22_X1 U15224 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12004), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15225 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U15226 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U15227 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12005) );
  NAND4_X1 U15228 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n12014) );
  AOI22_X1 U15229 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15230 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15231 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15232 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12009) );
  NAND4_X1 U15233 ( .A1(n12012), .A2(n12011), .A3(n12010), .A4(n12009), .ZN(
        n12013) );
  NOR2_X1 U15234 ( .A1(n12014), .A2(n12013), .ZN(n12017) );
  OAI21_X1 U15235 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20633), .A(
        n20764), .ZN(n12016) );
  NAND2_X1 U15236 ( .A1(n12719), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n12015) );
  OAI211_X1 U15237 ( .C1(n12195), .C2(n12017), .A(n12016), .B(n12015), .ZN(
        n12018) );
  OAI21_X1 U15238 ( .B1(n15789), .B2(n12198), .A(n12018), .ZN(n14531) );
  AOI22_X1 U15239 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9713), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15240 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15241 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15242 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12019) );
  NAND4_X1 U15243 ( .A1(n12022), .A2(n12021), .A3(n12020), .A4(n12019), .ZN(
        n12030) );
  AOI22_X1 U15244 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12023), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15245 ( .A1(n11647), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15246 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15247 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12025) );
  NAND4_X1 U15248 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12029) );
  OR2_X1 U15249 ( .A1(n12030), .A2(n12029), .ZN(n12031) );
  NAND2_X1 U15250 ( .A1(n12201), .A2(n12031), .ZN(n12038) );
  NAND2_X1 U15251 ( .A1(n14765), .A2(n12032), .ZN(n12034) );
  INV_X1 U15252 ( .A(n12033), .ZN(n12053) );
  OAI22_X1 U15253 ( .A1(n14769), .A2(n12198), .B1(n14765), .B2(n12035), .ZN(
        n12036) );
  AOI21_X1 U15254 ( .B1(n12719), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12036), .ZN(
        n12037) );
  NAND2_X1 U15255 ( .A1(n12038), .A2(n12037), .ZN(n14523) );
  AOI22_X1 U15256 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15257 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15258 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15259 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12039) );
  NAND4_X1 U15260 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12048) );
  AOI22_X1 U15261 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15262 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12097), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15263 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15264 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12043) );
  NAND4_X1 U15265 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12047) );
  NOR2_X1 U15266 ( .A1(n12048), .A2(n12047), .ZN(n12052) );
  OAI21_X1 U15267 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20633), .A(
        n20764), .ZN(n12049) );
  INV_X1 U15268 ( .A(n12049), .ZN(n12050) );
  AOI21_X1 U15269 ( .B1(n12719), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12050), .ZN(
        n12051) );
  OAI21_X1 U15270 ( .B1(n12195), .B2(n12052), .A(n12051), .ZN(n12057) );
  INV_X1 U15271 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12054) );
  NAND2_X1 U15272 ( .A1(n12054), .A2(n12053), .ZN(n12055) );
  AND2_X1 U15273 ( .A1(n12055), .A2(n12135), .ZN(n15731) );
  NAND2_X1 U15274 ( .A1(n15731), .A2(n12162), .ZN(n12056) );
  OR2_X1 U15275 ( .A1(n12058), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12059) );
  NAND2_X1 U15276 ( .A1(n12059), .A2(n12145), .ZN(n15773) );
  AOI22_X1 U15277 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12103), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15278 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12125), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15279 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15280 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12060) );
  NAND4_X1 U15281 ( .A1(n12063), .A2(n12062), .A3(n12061), .A4(n12060), .ZN(
        n12070) );
  AOI22_X1 U15282 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11647), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15283 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15284 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15285 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12065) );
  NAND4_X1 U15286 ( .A1(n12068), .A2(n12067), .A3(n12066), .A4(n12065), .ZN(
        n12069) );
  NOR2_X1 U15287 ( .A1(n12070), .A2(n12069), .ZN(n12071) );
  NOR2_X1 U15288 ( .A1(n12195), .A2(n12071), .ZN(n12074) );
  INV_X1 U15289 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14642) );
  NAND2_X1 U15290 ( .A1(n20764), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12072) );
  OAI211_X1 U15291 ( .C1(n12112), .C2(n14642), .A(n12198), .B(n12072), .ZN(
        n12073) );
  OAI22_X1 U15292 ( .A1(n15773), .A2(n12198), .B1(n12074), .B2(n12073), .ZN(
        n12075) );
  INV_X1 U15293 ( .A(n12075), .ZN(n14570) );
  AOI22_X1 U15294 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15295 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15296 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15297 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12076) );
  NAND4_X1 U15298 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12086) );
  AOI22_X1 U15299 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15300 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15301 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15302 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U15303 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12085) );
  NOR2_X1 U15304 ( .A1(n12086), .A2(n12085), .ZN(n12090) );
  AOI21_X1 U15305 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n12087), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12088) );
  AOI21_X1 U15306 ( .B1(n12719), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12088), .ZN(
        n12089) );
  OAI21_X1 U15307 ( .B1(n12195), .B2(n12090), .A(n12089), .ZN(n12092) );
  XNOR2_X1 U15308 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12094), .ZN(
        n14738) );
  NAND2_X1 U15309 ( .A1(n13843), .A2(n14738), .ZN(n12091) );
  NAND2_X1 U15310 ( .A1(n12092), .A2(n12091), .ZN(n14495) );
  OR2_X1 U15311 ( .A1(n12093), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12095) );
  NAND2_X1 U15312 ( .A1(n12095), .A2(n12094), .ZN(n15779) );
  AOI22_X1 U15313 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15314 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15315 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12023), .B1(
        n12097), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U15316 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12125), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12098) );
  NAND4_X1 U15317 ( .A1(n12101), .A2(n12100), .A3(n12099), .A4(n12098), .ZN(
        n12109) );
  AOI22_X1 U15318 ( .A1(n9713), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15319 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12103), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15320 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15321 ( .A1(n12123), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12104) );
  NAND4_X1 U15322 ( .A1(n12107), .A2(n12106), .A3(n12105), .A4(n12104), .ZN(
        n12108) );
  NOR2_X1 U15323 ( .A1(n12109), .A2(n12108), .ZN(n12110) );
  NOR2_X1 U15324 ( .A1(n12195), .A2(n12110), .ZN(n12114) );
  INV_X1 U15325 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14651) );
  NAND2_X1 U15326 ( .A1(n20764), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12111) );
  OAI211_X1 U15327 ( .C1(n12112), .C2(n14651), .A(n12198), .B(n12111), .ZN(
        n12113) );
  OAI22_X1 U15328 ( .A1(n15779), .A2(n12198), .B1(n12114), .B2(n12113), .ZN(
        n14583) );
  AOI22_X1 U15329 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12102), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15330 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15331 ( .A1(n11594), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12119) );
  NAND4_X1 U15332 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12119), .ZN(
        n12131) );
  AOI22_X1 U15333 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12123), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15334 ( .A1(n12023), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15335 ( .A1(n12125), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12124), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15336 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12126) );
  NAND4_X1 U15337 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12130) );
  NOR2_X1 U15338 ( .A1(n12131), .A2(n12130), .ZN(n12134) );
  AOI21_X1 U15339 ( .B1(n14514), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12132) );
  AOI21_X1 U15340 ( .B1(n12719), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12132), .ZN(
        n12133) );
  OAI21_X1 U15341 ( .B1(n12195), .B2(n12134), .A(n12133), .ZN(n12137) );
  XNOR2_X1 U15342 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12135), .ZN(
        n14747) );
  NAND2_X1 U15343 ( .A1(n14747), .A2(n13843), .ZN(n12136) );
  NAND2_X1 U15344 ( .A1(n12137), .A2(n12136), .ZN(n14507) );
  NOR2_X1 U15345 ( .A1(n14495), .A2(n14492), .ZN(n14493) );
  XOR2_X1 U15346 ( .A(n12140), .B(n12139), .Z(n12141) );
  NAND2_X1 U15347 ( .A1(n12141), .A2(n12201), .ZN(n12144) );
  AOI21_X1 U15348 ( .B1(n15713), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12142) );
  AOI21_X1 U15349 ( .B1(n12719), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12142), .ZN(
        n12143) );
  NAND2_X1 U15350 ( .A1(n12144), .A2(n12143), .ZN(n12147) );
  XNOR2_X1 U15351 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12145), .ZN(
        n15704) );
  NAND2_X1 U15352 ( .A1(n15704), .A2(n13843), .ZN(n12146) );
  OR2_X1 U15353 ( .A1(n12148), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12149) );
  NAND2_X1 U15354 ( .A1(n12149), .A2(n12161), .ZN(n15766) );
  XNOR2_X1 U15355 ( .A(n12151), .B(n12150), .ZN(n12155) );
  NAND2_X1 U15356 ( .A1(n20764), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12152) );
  NAND2_X1 U15357 ( .A1(n12198), .A2(n12152), .ZN(n12153) );
  AOI21_X1 U15358 ( .B1(n12719), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12153), .ZN(
        n12154) );
  OAI21_X1 U15359 ( .B1(n12155), .B2(n12195), .A(n12154), .ZN(n12156) );
  OAI21_X1 U15360 ( .B1(n15766), .B2(n12198), .A(n12156), .ZN(n14557) );
  XOR2_X1 U15361 ( .A(n12158), .B(n12157), .Z(n12159) );
  NAND2_X1 U15362 ( .A1(n12159), .A2(n12201), .ZN(n12165) );
  INV_X1 U15363 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14720) );
  OAI21_X1 U15364 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14720), .A(n12198), 
        .ZN(n12160) );
  AOI21_X1 U15365 ( .B1(n12719), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12160), .ZN(
        n12164) );
  XNOR2_X1 U15366 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n12161), .ZN(
        n14722) );
  AOI21_X1 U15367 ( .B1(n12165), .B2(n12164), .A(n12163), .ZN(n14480) );
  INV_X1 U15368 ( .A(n12166), .ZN(n12167) );
  XNOR2_X1 U15369 ( .A(n12168), .B(n12167), .ZN(n12169) );
  NAND2_X1 U15370 ( .A1(n12169), .A2(n12201), .ZN(n12177) );
  INV_X1 U15371 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12172) );
  AOI21_X1 U15372 ( .B1(n12172), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12170) );
  AOI21_X1 U15373 ( .B1(n12719), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12170), .ZN(
        n12176) );
  INV_X1 U15374 ( .A(n12171), .ZN(n12173) );
  NAND2_X1 U15375 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  NAND2_X1 U15376 ( .A1(n12184), .A2(n12174), .ZN(n14713) );
  NOR2_X1 U15377 ( .A1(n14713), .A2(n12198), .ZN(n12175) );
  AOI21_X1 U15378 ( .B1(n12177), .B2(n12176), .A(n12175), .ZN(n14468) );
  XOR2_X1 U15379 ( .A(n12179), .B(n12178), .Z(n12180) );
  NAND2_X1 U15380 ( .A1(n12180), .A2(n12201), .ZN(n12183) );
  AOI21_X1 U15381 ( .B1(n14295), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12181) );
  AOI21_X1 U15382 ( .B1(n12719), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12181), .ZN(
        n12182) );
  NAND2_X1 U15383 ( .A1(n12183), .A2(n12182), .ZN(n12187) );
  NAND2_X1 U15384 ( .A1(n12184), .A2(n14295), .ZN(n12185) );
  NAND2_X1 U15385 ( .A1(n14460), .A2(n13843), .ZN(n12186) );
  NAND2_X1 U15386 ( .A1(n12187), .A2(n12186), .ZN(n14292) );
  INV_X1 U15387 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12188) );
  NAND2_X1 U15388 ( .A1(n12189), .A2(n12188), .ZN(n12190) );
  NAND2_X1 U15389 ( .A1(n12204), .A2(n12190), .ZN(n14705) );
  XNOR2_X1 U15390 ( .A(n12192), .B(n12191), .ZN(n12196) );
  AOI21_X1 U15391 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20764), .A(
        n13843), .ZN(n12194) );
  NAND2_X1 U15392 ( .A1(n12719), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n12193) );
  OAI211_X1 U15393 ( .C1(n12196), .C2(n12195), .A(n12194), .B(n12193), .ZN(
        n12197) );
  OAI21_X1 U15394 ( .B1(n12198), .B2(n14705), .A(n12197), .ZN(n14444) );
  XOR2_X1 U15395 ( .A(n12200), .B(n12199), .Z(n12202) );
  NAND2_X1 U15396 ( .A1(n12202), .A2(n12201), .ZN(n12206) );
  INV_X1 U15397 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12715) );
  NOR2_X1 U15398 ( .A1(n12715), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12203) );
  AOI211_X1 U15399 ( .C1(n12719), .C2(P1_EAX_REG_29__SCAN_IN), .A(n13843), .B(
        n12203), .ZN(n12205) );
  XNOR2_X1 U15400 ( .A(n12204), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14435) );
  AOI22_X1 U15401 ( .A1(n12206), .A2(n12205), .B1(n13843), .B2(n14435), .ZN(
        n12709) );
  INV_X1 U15402 ( .A(n14690), .ZN(n14616) );
  NAND2_X1 U15403 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20628), .ZN(
        n12227) );
  OAI21_X1 U15404 ( .B1(n20628), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12227), .ZN(n12213) );
  INV_X1 U15405 ( .A(n12213), .ZN(n12210) );
  NAND2_X1 U15406 ( .A1(n12232), .A2(n12210), .ZN(n12211) );
  NAND2_X1 U15407 ( .A1(n12272), .A2(n12211), .ZN(n12218) );
  OAI211_X1 U15408 ( .C1(n20221), .C2(n12213), .A(n12212), .B(n13854), .ZN(
        n12216) );
  NAND2_X1 U15409 ( .A1(n11608), .A2(n13854), .ZN(n12215) );
  NAND2_X1 U15410 ( .A1(n12215), .A2(n12214), .ZN(n12239) );
  NAND2_X1 U15411 ( .A1(n12216), .A2(n12239), .ZN(n12217) );
  NAND2_X1 U15412 ( .A1(n12218), .A2(n12217), .ZN(n12226) );
  INV_X1 U15413 ( .A(n12226), .ZN(n12237) );
  NOR2_X1 U15414 ( .A1(n12209), .A2(n20761), .ZN(n12250) );
  AOI21_X1 U15415 ( .B1(n12232), .B2(n13860), .A(n12250), .ZN(n12223) );
  NAND2_X1 U15416 ( .A1(n20587), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12229) );
  NAND2_X1 U15417 ( .A1(n14831), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12219) );
  NAND2_X1 U15418 ( .A1(n12229), .A2(n12219), .ZN(n12228) );
  INV_X1 U15419 ( .A(n12227), .ZN(n12220) );
  XNOR2_X1 U15420 ( .A(n12228), .B(n12220), .ZN(n12725) );
  INV_X1 U15421 ( .A(n12725), .ZN(n12221) );
  NAND2_X1 U15422 ( .A1(n12270), .A2(n12221), .ZN(n12222) );
  INV_X1 U15423 ( .A(n12225), .ZN(n12236) );
  AOI21_X1 U15424 ( .B1(n12268), .B2(n12670), .A(n12725), .ZN(n12224) );
  OAI21_X1 U15425 ( .B1(n12226), .B2(n12225), .A(n12224), .ZN(n12235) );
  NAND2_X1 U15426 ( .A1(n12230), .A2(n12229), .ZN(n12246) );
  MUX2_X1 U15427 ( .A(n12247), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n11816), .Z(n12244) );
  XNOR2_X1 U15428 ( .A(n12246), .B(n12244), .ZN(n12726) );
  INV_X1 U15429 ( .A(n12726), .ZN(n12231) );
  NAND2_X1 U15430 ( .A1(n12270), .A2(n12231), .ZN(n12233) );
  NAND2_X1 U15431 ( .A1(n12232), .A2(n12726), .ZN(n12238) );
  NAND3_X1 U15432 ( .A1(n12233), .A2(n12239), .A3(n12238), .ZN(n12234) );
  OAI211_X1 U15433 ( .C1(n12237), .C2(n12236), .A(n12235), .B(n12234), .ZN(
        n12243) );
  INV_X1 U15434 ( .A(n12238), .ZN(n12241) );
  INV_X1 U15435 ( .A(n12239), .ZN(n12240) );
  NAND2_X1 U15436 ( .A1(n12241), .A2(n12240), .ZN(n12242) );
  NAND2_X1 U15437 ( .A1(n12243), .A2(n12242), .ZN(n12271) );
  INV_X1 U15438 ( .A(n12244), .ZN(n12245) );
  NAND2_X1 U15439 ( .A1(n12246), .A2(n12245), .ZN(n12249) );
  NAND2_X1 U15440 ( .A1(n12247), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12248) );
  NAND2_X1 U15441 ( .A1(n12249), .A2(n12248), .ZN(n12254) );
  XNOR2_X1 U15442 ( .A(n13669), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12251) );
  XNOR2_X1 U15443 ( .A(n12254), .B(n12251), .ZN(n12724) );
  NAND2_X1 U15444 ( .A1(n12271), .A2(n12724), .ZN(n12258) );
  INV_X1 U15445 ( .A(n12250), .ZN(n12256) );
  INV_X1 U15446 ( .A(n12251), .ZN(n12253) );
  NOR2_X1 U15447 ( .A1(n13669), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12252) );
  AOI21_X1 U15448 ( .B1(n12254), .B2(n12253), .A(n12252), .ZN(n12263) );
  NOR2_X1 U15449 ( .A1(n20188), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12255) );
  AND2_X1 U15450 ( .A1(n12263), .A2(n12255), .ZN(n12728) );
  NAND3_X1 U15451 ( .A1(n12256), .A2(n12728), .A3(n13860), .ZN(n12257) );
  NAND2_X1 U15452 ( .A1(n12258), .A2(n12257), .ZN(n12261) );
  NAND2_X1 U15453 ( .A1(n12259), .A2(n12728), .ZN(n12260) );
  NAND2_X1 U15454 ( .A1(n20188), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12262) );
  NAND2_X1 U15455 ( .A1(n12263), .A2(n12262), .ZN(n12265) );
  NAND2_X1 U15456 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13674), .ZN(
        n12264) );
  NAND2_X1 U15457 ( .A1(n12265), .A2(n12264), .ZN(n12729) );
  NOR2_X1 U15458 ( .A1(n12272), .A2(n12724), .ZN(n12266) );
  AOI21_X1 U15459 ( .B1(n20761), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n12266), .ZN(n12267) );
  OAI21_X1 U15460 ( .B1(n12268), .B2(n12729), .A(n12267), .ZN(n12269) );
  OR2_X1 U15461 ( .A1(n11621), .A2(n12214), .ZN(n12769) );
  NOR2_X1 U15462 ( .A1(n12277), .A2(n12769), .ZN(n13646) );
  NAND3_X1 U15463 ( .A1(n15646), .A2(n13460), .A3(n13646), .ZN(n12282) );
  INV_X1 U15464 ( .A(n12212), .ZN(n12280) );
  NOR2_X1 U15465 ( .A1(n11619), .A2(n19992), .ZN(n12279) );
  NAND4_X1 U15466 ( .A1(n13662), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12736) );
  INV_X2 U15467 ( .A(n12301), .ZN(n13380) );
  OR2_X1 U15468 ( .A1(n12736), .A2(n13380), .ZN(n12281) );
  NAND2_X1 U15469 ( .A1(n12356), .A2(n13935), .ZN(n12287) );
  INV_X1 U15470 ( .A(n12296), .ZN(n12300) );
  INV_X1 U15471 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13589) );
  NAND2_X1 U15472 ( .A1(n12373), .A2(n13589), .ZN(n12285) );
  OAI211_X1 U15473 ( .C1(n12284), .C2(P1_EBX_REG_1__SCAN_IN), .A(n12285), .B(
        n9907), .ZN(n12286) );
  NAND2_X1 U15474 ( .A1(n12287), .A2(n12286), .ZN(n12290) );
  NAND2_X1 U15475 ( .A1(n12373), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12289) );
  INV_X1 U15476 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13562) );
  NAND2_X1 U15477 ( .A1(n9907), .A2(n13562), .ZN(n12288) );
  NAND2_X1 U15478 ( .A1(n12289), .A2(n12288), .ZN(n13547) );
  INV_X1 U15479 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U15480 ( .A1(n12356), .A2(n13613), .ZN(n12293) );
  INV_X1 U15481 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12621) );
  NAND2_X1 U15482 ( .A1(n12373), .A2(n12621), .ZN(n12291) );
  OAI211_X1 U15483 ( .C1(n12284), .C2(P1_EBX_REG_2__SCAN_IN), .A(n12291), .B(
        n12329), .ZN(n12292) );
  AND2_X1 U15484 ( .A1(n12293), .A2(n12292), .ZN(n13610) );
  OR2_X1 U15485 ( .A1(n12371), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n12299) );
  NAND2_X1 U15486 ( .A1(n12329), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12297) );
  OAI211_X1 U15487 ( .C1(n13380), .C2(P1_EBX_REG_3__SCAN_IN), .A(n12373), .B(
        n12297), .ZN(n12298) );
  NAND2_X1 U15488 ( .A1(n12299), .A2(n12298), .ZN(n13754) );
  MUX2_X1 U15489 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12304) );
  INV_X2 U15490 ( .A(n12300), .ZN(n12373) );
  NAND2_X1 U15491 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13380), .ZN(
        n12302) );
  AND2_X1 U15492 ( .A1(n12351), .A2(n12302), .ZN(n12303) );
  NAND2_X1 U15493 ( .A1(n12304), .A2(n12303), .ZN(n13895) );
  OR2_X1 U15494 ( .A1(n12371), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U15495 ( .A1(n12329), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12305) );
  OAI211_X1 U15496 ( .C1(n13380), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12373), .B(
        n12305), .ZN(n12306) );
  AND2_X1 U15497 ( .A1(n12307), .A2(n12306), .ZN(n13894) );
  NAND2_X1 U15498 ( .A1(n13895), .A2(n13894), .ZN(n12308) );
  MUX2_X1 U15499 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12311) );
  NAND2_X1 U15500 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13380), .ZN(
        n12309) );
  AND2_X1 U15501 ( .A1(n12351), .A2(n12309), .ZN(n12310) );
  NAND2_X1 U15502 ( .A1(n12311), .A2(n12310), .ZN(n13956) );
  OR2_X1 U15503 ( .A1(n12371), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n12314) );
  NAND2_X1 U15504 ( .A1(n9907), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12312) );
  OAI211_X1 U15505 ( .C1(n13380), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12373), .B(
        n12312), .ZN(n12313) );
  AND2_X1 U15506 ( .A1(n12314), .A2(n12313), .ZN(n13955) );
  MUX2_X1 U15507 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12317) );
  NAND2_X1 U15508 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n13380), .ZN(
        n12316) );
  OR2_X1 U15509 ( .A1(n12371), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U15510 ( .A1(n12329), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12318) );
  OAI211_X1 U15511 ( .C1(n13380), .C2(P1_EBX_REG_9__SCAN_IN), .A(n12373), .B(
        n12318), .ZN(n12319) );
  NAND2_X1 U15512 ( .A1(n12320), .A2(n12319), .ZN(n14025) );
  MUX2_X1 U15513 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12323) );
  NAND2_X1 U15514 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n13380), .ZN(
        n12321) );
  AND2_X1 U15515 ( .A1(n12351), .A2(n12321), .ZN(n12322) );
  NAND2_X1 U15516 ( .A1(n12323), .A2(n12322), .ZN(n14053) );
  OR2_X1 U15517 ( .A1(n12371), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U15518 ( .A1(n9907), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12324) );
  OAI211_X1 U15519 ( .C1(n13380), .C2(P1_EBX_REG_11__SCAN_IN), .A(n12373), .B(
        n12324), .ZN(n12325) );
  MUX2_X1 U15520 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12328) );
  NAND2_X1 U15521 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n13380), .ZN(
        n12327) );
  OR2_X1 U15522 ( .A1(n12371), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n12332) );
  NAND2_X1 U15523 ( .A1(n12329), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12330) );
  OAI211_X1 U15524 ( .C1(n13380), .C2(P1_EBX_REG_13__SCAN_IN), .A(n12373), .B(
        n12330), .ZN(n12331) );
  NAND2_X1 U15525 ( .A1(n12332), .A2(n12331), .ZN(n14165) );
  MUX2_X1 U15526 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12335) );
  NAND2_X1 U15527 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n13380), .ZN(
        n12333) );
  AND2_X1 U15528 ( .A1(n12351), .A2(n12333), .ZN(n12334) );
  NAND2_X1 U15529 ( .A1(n12335), .A2(n12334), .ZN(n14132) );
  NAND2_X1 U15530 ( .A1(n14164), .A2(n14132), .ZN(n14198) );
  OR2_X1 U15531 ( .A1(n13546), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12338) );
  NAND2_X1 U15532 ( .A1(n13375), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n12337) );
  OAI211_X1 U15533 ( .C1(n12371), .C2(P1_EBX_REG_15__SCAN_IN), .A(n12338), .B(
        n12337), .ZN(n14199) );
  MUX2_X1 U15534 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12340) );
  NAND2_X1 U15535 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n13380), .ZN(
        n12339) );
  OR2_X1 U15536 ( .A1(n12371), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n12343) );
  OAI211_X1 U15537 ( .C1(n13380), .C2(P1_EBX_REG_17__SCAN_IN), .A(n12373), .B(
        n12341), .ZN(n12342) );
  NAND2_X1 U15538 ( .A1(n12343), .A2(n12342), .ZN(n14525) );
  INV_X1 U15539 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15728) );
  NAND2_X1 U15540 ( .A1(n12356), .A2(n15728), .ZN(n12346) );
  INV_X1 U15541 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15888) );
  NAND2_X1 U15542 ( .A1(n12373), .A2(n15888), .ZN(n12344) );
  OAI211_X1 U15543 ( .C1(n13380), .C2(P1_EBX_REG_18__SCAN_IN), .A(n12344), .B(
        n12329), .ZN(n12345) );
  NAND2_X1 U15544 ( .A1(n12346), .A2(n12345), .ZN(n14599) );
  OR2_X1 U15545 ( .A1(n12371), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n12349) );
  NAND2_X1 U15546 ( .A1(n9907), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12347) );
  OAI211_X1 U15547 ( .C1(n13380), .C2(P1_EBX_REG_19__SCAN_IN), .A(n12373), .B(
        n12347), .ZN(n12348) );
  NAND2_X1 U15548 ( .A1(n12349), .A2(n12348), .ZN(n14511) );
  MUX2_X1 U15549 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12352) );
  NAND2_X1 U15550 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13380), .ZN(
        n12350) );
  OR2_X1 U15551 ( .A1(n12371), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U15552 ( .A1(n12329), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12353) );
  OAI211_X1 U15553 ( .C1(n13380), .C2(P1_EBX_REG_21__SCAN_IN), .A(n12373), .B(
        n12353), .ZN(n12354) );
  AND2_X1 U15554 ( .A1(n12355), .A2(n12354), .ZN(n14496) );
  INV_X1 U15555 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14577) );
  NAND2_X1 U15556 ( .A1(n12356), .A2(n14577), .ZN(n12360) );
  INV_X1 U15557 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12357) );
  NAND2_X1 U15558 ( .A1(n12373), .A2(n12357), .ZN(n12358) );
  OAI211_X1 U15559 ( .C1(n13380), .C2(P1_EBX_REG_22__SCAN_IN), .A(n12358), .B(
        n12329), .ZN(n12359) );
  NAND2_X1 U15560 ( .A1(n12360), .A2(n12359), .ZN(n14573) );
  OR2_X1 U15561 ( .A1(n12371), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n12363) );
  NAND2_X1 U15562 ( .A1(n9907), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12361) );
  OAI211_X1 U15563 ( .C1(n13380), .C2(P1_EBX_REG_23__SCAN_IN), .A(n12373), .B(
        n12361), .ZN(n12362) );
  NAND2_X1 U15564 ( .A1(n12363), .A2(n12362), .ZN(n14567) );
  NAND2_X1 U15565 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n13380), .ZN(
        n12365) );
  MUX2_X1 U15566 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12364) );
  AND2_X1 U15567 ( .A1(n12365), .A2(n12364), .ZN(n14559) );
  OR2_X1 U15568 ( .A1(n12371), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n12368) );
  NAND2_X1 U15569 ( .A1(n9907), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12366) );
  OAI211_X1 U15570 ( .C1(n13380), .C2(P1_EBX_REG_25__SCAN_IN), .A(n12373), .B(
        n12366), .ZN(n12367) );
  NAND2_X1 U15571 ( .A1(n12368), .A2(n12367), .ZN(n14482) );
  MUX2_X1 U15572 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12370) );
  NAND2_X1 U15573 ( .A1(n13380), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12369) );
  NAND2_X1 U15574 ( .A1(n12370), .A2(n12369), .ZN(n14470) );
  OR2_X1 U15575 ( .A1(n12371), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n12375) );
  NAND2_X1 U15576 ( .A1(n12329), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12372) );
  OAI211_X1 U15577 ( .C1(n13380), .C2(P1_EBX_REG_27__SCAN_IN), .A(n12373), .B(
        n12372), .ZN(n12374) );
  NAND2_X1 U15578 ( .A1(n12375), .A2(n12374), .ZN(n14285) );
  MUX2_X1 U15579 ( .A(n12380), .B(n12373), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12377) );
  NAND2_X1 U15580 ( .A1(n12284), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12376) );
  AND2_X1 U15581 ( .A1(n12377), .A2(n12376), .ZN(n14454) );
  NOR2_X2 U15582 ( .A1(n14453), .A2(n14454), .ZN(n14452) );
  OR2_X1 U15583 ( .A1(n13546), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12379) );
  OR2_X1 U15584 ( .A1(n13380), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12378) );
  NAND2_X1 U15585 ( .A1(n12379), .A2(n12378), .ZN(n12381) );
  OAI22_X1 U15586 ( .A1(n12381), .A2(n13375), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12380), .ZN(n14404) );
  NAND2_X1 U15587 ( .A1(n14452), .A2(n14404), .ZN(n14406) );
  NAND2_X1 U15588 ( .A1(n14406), .A2(n13375), .ZN(n12384) );
  INV_X1 U15589 ( .A(n12381), .ZN(n12382) );
  NAND2_X1 U15590 ( .A1(n14452), .A2(n12382), .ZN(n12383) );
  NAND2_X1 U15591 ( .A1(n12384), .A2(n12383), .ZN(n12387) );
  NAND2_X1 U15592 ( .A1(n13546), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12386) );
  NAND2_X1 U15593 ( .A1(n13380), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12385) );
  NAND2_X1 U15594 ( .A1(n12386), .A2(n12385), .ZN(n12782) );
  INV_X1 U15595 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n12388) );
  OR2_X1 U15596 ( .A1(n14611), .A2(n12388), .ZN(n12389) );
  INV_X1 U15597 ( .A(n12392), .ZN(n12393) );
  NAND2_X1 U15598 ( .A1(n12393), .A2(n12394), .ZN(n14259) );
  INV_X1 U15599 ( .A(n14259), .ZN(n12396) );
  AOI21_X1 U15600 ( .B1(n12394), .B2(n14258), .A(n12393), .ZN(n12395) );
  AND2_X1 U15601 ( .A1(n19968), .A2(n16367), .ZN(n12397) );
  NAND2_X1 U15602 ( .A1(n12398), .A2(n12397), .ZN(n18875) );
  NAND2_X1 U15603 ( .A1(n12418), .A2(n19264), .ZN(n12417) );
  NAND2_X2 U15604 ( .A1(n16192), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15330) );
  INV_X1 U15605 ( .A(n12423), .ZN(n12399) );
  NOR2_X1 U15606 ( .A1(n15330), .A2(n12399), .ZN(n15127) );
  NAND2_X1 U15607 ( .A1(n12591), .A2(n12400), .ZN(n15113) );
  OAI21_X1 U15608 ( .B1(n15127), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15113), .ZN(n12431) );
  INV_X1 U15609 ( .A(n14236), .ZN(n12401) );
  AOI21_X1 U15610 ( .B1(n12402), .B2(n14121), .A(n12401), .ZN(n18914) );
  NOR2_X1 U15611 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14001) );
  OR2_X1 U15612 ( .A1(n19934), .A2(n14001), .ZN(n19935) );
  NAND2_X1 U15613 ( .A1(n19935), .A2(n19969), .ZN(n12403) );
  AND2_X1 U15614 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19936) );
  INV_X1 U15615 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12406) );
  OAI22_X1 U15616 ( .A1(n16239), .A2(n12406), .B1(n12405), .B2(n9722), .ZN(
        n12413) );
  INV_X1 U15617 ( .A(n12848), .ZN(n12408) );
  NAND2_X1 U15618 ( .A1(n19914), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12407) );
  NAND2_X1 U15619 ( .A1(n12408), .A2(n12407), .ZN(n13360) );
  AND2_X1 U15620 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12409) );
  AND2_X1 U15621 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12410) );
  AND2_X1 U15622 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12411) );
  INV_X1 U15623 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18921) );
  NOR2_X2 U15624 ( .A1(n13188), .A2(n18921), .ZN(n13189) );
  INV_X1 U15625 ( .A(n13172), .ZN(n13187) );
  OAI21_X1 U15626 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13189), .A(
        n13187), .ZN(n18908) );
  NOR2_X1 U15627 ( .A1(n19269), .A2(n18908), .ZN(n12412) );
  AOI211_X1 U15628 ( .C1(n18914), .C2(n19263), .A(n12413), .B(n12412), .ZN(
        n12414) );
  NAND2_X1 U15629 ( .A1(n12417), .A2(n12416), .ZN(P2_U2996) );
  NAND2_X1 U15630 ( .A1(n12418), .A2(n16301), .ZN(n12434) );
  AND2_X1 U15631 ( .A1(n14099), .A2(n15350), .ZN(n12419) );
  NOR2_X1 U15632 ( .A1(n15349), .A2(n12419), .ZN(n16269) );
  INV_X1 U15633 ( .A(n15336), .ZN(n12420) );
  NAND2_X1 U15634 ( .A1(n15247), .A2(n12420), .ZN(n12421) );
  NAND2_X1 U15635 ( .A1(n16269), .A2(n12421), .ZN(n16255) );
  AOI21_X1 U15636 ( .B1(n14266), .B2(n15247), .A(n16255), .ZN(n15228) );
  INV_X1 U15637 ( .A(n15228), .ZN(n12429) );
  INV_X1 U15638 ( .A(n18914), .ZN(n14213) );
  NAND3_X1 U15639 ( .A1(n16260), .A2(n12423), .A3(n12422), .ZN(n12427) );
  NOR2_X1 U15640 ( .A1(n15261), .A2(n15026), .ZN(n15028) );
  OR2_X1 U15641 ( .A1(n15028), .A2(n12424), .ZN(n12425) );
  AND2_X1 U15642 ( .A1(n14264), .A2(n12425), .ZN(n18913) );
  AOI22_X1 U15643 ( .A1(n16281), .A2(n18913), .B1(n15077), .B2(
        P2_REIP_REG_18__SCAN_IN), .ZN(n12426) );
  OAI211_X1 U15644 ( .C1(n14213), .C2(n16283), .A(n12427), .B(n12426), .ZN(
        n12428) );
  AOI21_X1 U15645 ( .B1(n12429), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12428), .ZN(n12430) );
  NAND2_X1 U15646 ( .A1(n12434), .A2(n12433), .ZN(P2_U3028) );
  AND4_X1 U15647 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n15296), .ZN(
        n12438) );
  AND4_X1 U15648 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n15108), .ZN(
        n15203) );
  INV_X1 U15649 ( .A(n15203), .ZN(n12459) );
  OR2_X1 U15650 ( .A1(n12441), .A2(n12459), .ZN(n12449) );
  NAND2_X1 U15651 ( .A1(n19300), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12442) );
  INV_X1 U15652 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n14945) );
  NAND2_X1 U15653 ( .A1(n12445), .A2(n12444), .ZN(n12446) );
  NAND2_X1 U15654 ( .A1(n12463), .A2(n12446), .ZN(n15601) );
  INV_X1 U15655 ( .A(n12450), .ZN(n12447) );
  NAND2_X1 U15656 ( .A1(n12447), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15201) );
  INV_X1 U15657 ( .A(n15201), .ZN(n12448) );
  NAND2_X1 U15658 ( .A1(n9719), .A2(n10077), .ZN(n15084) );
  INV_X1 U15659 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16242) );
  NAND2_X1 U15660 ( .A1(n12450), .A2(n16242), .ZN(n15200) );
  INV_X1 U15661 ( .A(n15200), .ZN(n12457) );
  AND4_X1 U15662 ( .A1(n12451), .A2(n16156), .A3(n15272), .A4(n15297), .ZN(
        n12453) );
  INV_X1 U15663 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12513) );
  XNOR2_X1 U15664 ( .A(n12463), .B(n9815), .ZN(n16109) );
  NAND2_X1 U15665 ( .A1(n16109), .A2(n12496), .ZN(n12461) );
  XNOR2_X1 U15666 ( .A(n12461), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15086) );
  AND2_X1 U15667 ( .A1(n15083), .A2(n15086), .ZN(n12460) );
  NAND2_X1 U15668 ( .A1(n15084), .A2(n12460), .ZN(n15085) );
  INV_X1 U15669 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16244) );
  OR2_X1 U15670 ( .A1(n12461), .A2(n16244), .ZN(n12462) );
  INV_X1 U15671 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14923) );
  NAND2_X1 U15672 ( .A1(n19300), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12464) );
  OAI21_X1 U15673 ( .B1(n12465), .B2(n12464), .A(n12473), .ZN(n12466) );
  OR2_X1 U15674 ( .A1(n12468), .A2(n12466), .ZN(n16101) );
  INV_X1 U15675 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15190) );
  NOR2_X1 U15676 ( .A1(n12467), .A2(n15190), .ZN(n15074) );
  NAND2_X1 U15677 ( .A1(n12467), .A2(n15190), .ZN(n15072) );
  OAI21_X2 U15678 ( .B1(n15076), .B2(n15074), .A(n15072), .ZN(n14318) );
  INV_X1 U15679 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14912) );
  NOR2_X1 U15680 ( .A1(n12468), .A2(n14912), .ZN(n12469) );
  NAND2_X1 U15681 ( .A1(n19300), .A2(n12469), .ZN(n12470) );
  AND2_X1 U15682 ( .A1(n12473), .A2(n12470), .ZN(n12471) );
  NAND2_X1 U15683 ( .A1(n12474), .A2(n12471), .ZN(n16086) );
  OR2_X1 U15684 ( .A1(n16086), .A2(n12494), .ZN(n12472) );
  INV_X1 U15685 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14329) );
  NAND2_X1 U15686 ( .A1(n12472), .A2(n14329), .ZN(n15061) );
  NOR2_X1 U15687 ( .A1(n12479), .A2(n10937), .ZN(n12477) );
  NAND3_X1 U15688 ( .A1(n19300), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n12474), 
        .ZN(n12475) );
  NAND2_X1 U15689 ( .A1(n12477), .A2(n12475), .ZN(n16073) );
  XNOR2_X1 U15690 ( .A(n12487), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15064) );
  NAND2_X1 U15691 ( .A1(n15061), .A2(n15064), .ZN(n12476) );
  NAND2_X1 U15692 ( .A1(n19300), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12478) );
  INV_X1 U15693 ( .A(n12478), .ZN(n12481) );
  NAND2_X1 U15694 ( .A1(n12481), .A2(n12480), .ZN(n12482) );
  INV_X1 U15695 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12534) );
  NOR2_X1 U15696 ( .A1(n10803), .A2(n12534), .ZN(n12483) );
  NOR2_X2 U15697 ( .A1(n12484), .A2(n12483), .ZN(n12491) );
  NAND2_X1 U15698 ( .A1(n12484), .A2(n12483), .ZN(n12485) );
  NAND2_X1 U15699 ( .A1(n12486), .A2(n12485), .ZN(n13220) );
  INV_X1 U15700 ( .A(n12487), .ZN(n12488) );
  NAND2_X1 U15701 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12489) );
  NAND2_X1 U15702 ( .A1(n19300), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12490) );
  XNOR2_X1 U15703 ( .A(n12491), .B(n12490), .ZN(n12495) );
  INV_X1 U15704 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15046) );
  OAI21_X1 U15705 ( .B1(n12495), .B2(n12494), .A(n15046), .ZN(n15041) );
  NAND2_X1 U15706 ( .A1(n15042), .A2(n15041), .ZN(n14299) );
  NAND2_X1 U15707 ( .A1(n19300), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12492) );
  XNOR2_X1 U15708 ( .A(n16023), .B(n12492), .ZN(n12493) );
  AOI21_X1 U15709 ( .B1(n12493), .B2(n12496), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14300) );
  INV_X1 U15710 ( .A(n12493), .ZN(n16039) );
  INV_X1 U15711 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12576) );
  INV_X1 U15712 ( .A(n12495), .ZN(n16048) );
  NAND3_X1 U15713 ( .A1(n16048), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12496), .ZN(n15040) );
  INV_X1 U15714 ( .A(n15040), .ZN(n12497) );
  NOR2_X1 U15715 ( .A1(n9769), .A2(n12497), .ZN(n12498) );
  NOR2_X1 U15716 ( .A1(n12499), .A2(n9949), .ZN(n12500) );
  XOR2_X1 U15717 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12500), .Z(
        n12501) );
  XNOR2_X1 U15718 ( .A(n12502), .B(n12501), .ZN(n14317) );
  NAND2_X1 U15719 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12507) );
  NAND2_X1 U15720 ( .A1(n12543), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12504) );
  NAND2_X1 U15721 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12503) );
  OAI211_X1 U15722 ( .C1(n12542), .C2(n14945), .A(n12504), .B(n12503), .ZN(
        n12505) );
  INV_X1 U15723 ( .A(n12505), .ZN(n12506) );
  AND2_X1 U15724 ( .A1(n12507), .A2(n12506), .ZN(n14940) );
  NAND2_X1 U15725 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12512) );
  AOI22_X1 U15726 ( .A1(n12543), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12511) );
  OAI211_X1 U15727 ( .C1(n12542), .C2(n12513), .A(n12512), .B(n12511), .ZN(
        n14931) );
  NAND2_X1 U15728 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12518) );
  NAND2_X1 U15729 ( .A1(n12543), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12515) );
  NAND2_X1 U15730 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12514) );
  OAI211_X1 U15731 ( .C1(n12542), .C2(n14923), .A(n12515), .B(n12514), .ZN(
        n12516) );
  INV_X1 U15732 ( .A(n12516), .ZN(n12517) );
  NAND2_X1 U15733 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12523) );
  NAND2_X1 U15734 ( .A1(n12543), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12520) );
  NAND2_X1 U15735 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12519) );
  OAI211_X1 U15736 ( .C1(n12542), .C2(n14912), .A(n12520), .B(n12519), .ZN(
        n12521) );
  INV_X1 U15737 ( .A(n12521), .ZN(n12522) );
  AND2_X1 U15738 ( .A1(n12523), .A2(n12522), .ZN(n14321) );
  NAND2_X1 U15739 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12529) );
  INV_X1 U15740 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12526) );
  NAND2_X1 U15741 ( .A1(n12543), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12525) );
  NAND2_X1 U15742 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12524) );
  OAI211_X1 U15743 ( .C1(n12542), .C2(n12526), .A(n12525), .B(n12524), .ZN(
        n12527) );
  INV_X1 U15744 ( .A(n12527), .ZN(n12528) );
  NAND2_X1 U15745 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12531) );
  AOI22_X1 U15746 ( .A1(n12543), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12530) );
  OAI211_X1 U15747 ( .C1(n12542), .C2(n10231), .A(n12531), .B(n12530), .ZN(
        n14896) );
  NAND2_X1 U15748 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12533) );
  AOI22_X1 U15749 ( .A1(n12543), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12532) );
  OAI211_X1 U15750 ( .C1(n12542), .C2(n12534), .A(n12533), .B(n12532), .ZN(
        n13223) );
  INV_X1 U15751 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12537) );
  NAND2_X1 U15752 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12536) );
  AOI22_X1 U15753 ( .A1(n12543), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12535) );
  OAI211_X1 U15754 ( .C1(n12542), .C2(n12537), .A(n12536), .B(n12535), .ZN(
        n14877) );
  INV_X1 U15755 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12541) );
  NAND2_X1 U15756 ( .A1(n12538), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12540) );
  AOI22_X1 U15757 ( .A1(n12543), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12539) );
  OAI211_X1 U15758 ( .C1(n12542), .C2(n12541), .A(n12540), .B(n12539), .ZN(
        n14304) );
  INV_X1 U15759 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U15760 ( .A1(n12543), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12546) );
  NAND2_X1 U15761 ( .A1(n12544), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12545) );
  OAI211_X1 U15762 ( .C1(n11102), .C2(n13180), .A(n12546), .B(n12545), .ZN(
        n12547) );
  INV_X1 U15763 ( .A(n12547), .ZN(n12548) );
  INV_X1 U15764 ( .A(n16283), .ZN(n12589) );
  INV_X1 U15765 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12550) );
  OR2_X1 U15766 ( .A1(n11211), .A2(n12550), .ZN(n12552) );
  AOI22_X1 U15767 ( .A1(n12571), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12551) );
  NAND2_X1 U15768 ( .A1(n12552), .A2(n12551), .ZN(n15216) );
  INV_X1 U15769 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19886) );
  OR2_X1 U15770 ( .A1(n11211), .A2(n19886), .ZN(n12554) );
  AOI22_X1 U15771 ( .A1(n12571), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12553) );
  AND2_X1 U15772 ( .A1(n12554), .A2(n12553), .ZN(n15004) );
  INV_X1 U15773 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n12555) );
  OR2_X1 U15774 ( .A1(n11211), .A2(n12555), .ZN(n12557) );
  AOI22_X1 U15775 ( .A1(n12571), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12556) );
  NAND2_X1 U15776 ( .A1(n12557), .A2(n12556), .ZN(n14996) );
  INV_X1 U15777 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19889) );
  OR2_X1 U15778 ( .A1(n11211), .A2(n19889), .ZN(n12559) );
  AOI22_X1 U15779 ( .A1(n12571), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12558) );
  AND2_X1 U15780 ( .A1(n12559), .A2(n12558), .ZN(n14323) );
  INV_X1 U15781 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15066) );
  OR2_X1 U15782 ( .A1(n11211), .A2(n15066), .ZN(n12561) );
  AOI22_X1 U15783 ( .A1(n12571), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11232), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12560) );
  AND2_X1 U15784 ( .A1(n12561), .A2(n12560), .ZN(n14977) );
  INV_X1 U15785 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19893) );
  OR2_X1 U15786 ( .A1(n11211), .A2(n19893), .ZN(n12563) );
  AOI22_X1 U15787 ( .A1(n11200), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11232), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12562) );
  NAND2_X1 U15788 ( .A1(n12563), .A2(n12562), .ZN(n14967) );
  AND2_X2 U15789 ( .A1(n14966), .A2(n14967), .ZN(n13227) );
  INV_X1 U15790 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19894) );
  OR2_X1 U15791 ( .A1(n11211), .A2(n19894), .ZN(n12566) );
  AOI22_X1 U15792 ( .A1(n11200), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12565) );
  NAND2_X1 U15793 ( .A1(n12566), .A2(n12565), .ZN(n13228) );
  INV_X1 U15794 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19896) );
  OR2_X1 U15795 ( .A1(n11211), .A2(n19896), .ZN(n12568) );
  AOI22_X1 U15796 ( .A1(n11200), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11232), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12567) );
  AND2_X1 U15797 ( .A1(n12568), .A2(n12567), .ZN(n14950) );
  INV_X1 U15798 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n14308) );
  OR2_X1 U15799 ( .A1(n11211), .A2(n14308), .ZN(n12570) );
  AOI22_X1 U15800 ( .A1(n11200), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12564), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12569) );
  AND2_X1 U15801 ( .A1(n12570), .A2(n12569), .ZN(n13159) );
  AOI222_X1 U15802 ( .A1(n12572), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11232), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n12571), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n12573) );
  NAND2_X1 U15803 ( .A1(n15077), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14311) );
  INV_X1 U15804 ( .A(n14311), .ZN(n12574) );
  AOI21_X1 U15805 ( .B1(n19101), .B2(n16281), .A(n12574), .ZN(n12587) );
  NAND3_X1 U15806 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15191) );
  NOR3_X1 U15807 ( .A1(n15211), .A2(n15191), .A3(n15190), .ZN(n15179) );
  AND2_X1 U15808 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12581) );
  NAND2_X1 U15809 ( .A1(n15179), .A2(n12581), .ZN(n15157) );
  INV_X1 U15810 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15173) );
  NOR2_X1 U15811 ( .A1(n12575), .A2(n15173), .ZN(n14361) );
  NAND2_X1 U15812 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n14361), .ZN(
        n14305) );
  NOR4_X1 U15813 ( .A1(n15157), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14305), .A4(n12576), .ZN(n12586) );
  INV_X1 U15814 ( .A(n14099), .ZN(n12585) );
  INV_X1 U15815 ( .A(n14305), .ZN(n12584) );
  NOR2_X1 U15816 ( .A1(n12577), .A2(n15191), .ZN(n12590) );
  INV_X1 U15817 ( .A(n12590), .ZN(n12578) );
  NAND2_X1 U15818 ( .A1(n14099), .A2(n12578), .ZN(n12579) );
  NAND2_X1 U15819 ( .A1(n12579), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12580) );
  NOR2_X1 U15820 ( .A1(n15349), .A2(n12580), .ZN(n15189) );
  OR2_X1 U15821 ( .A1(n15189), .A2(n12585), .ZN(n15184) );
  INV_X1 U15822 ( .A(n12581), .ZN(n12582) );
  NAND2_X1 U15823 ( .A1(n14099), .A2(n12582), .ZN(n12583) );
  OAI211_X1 U15824 ( .C1(n12585), .C2(n12584), .A(n15167), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14306) );
  NAND2_X1 U15825 ( .A1(n12587), .A2(n10079), .ZN(n12588) );
  NAND2_X1 U15826 ( .A1(n15044), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12593) );
  OAI211_X1 U15827 ( .C1(n14317), .C2(n16315), .A(n12595), .B(n12594), .ZN(
        P2_U3015) );
  INV_X1 U15828 ( .A(n12596), .ZN(n12597) );
  NAND2_X1 U15829 ( .A1(n12597), .A2(n12670), .ZN(n12604) );
  NAND2_X1 U15830 ( .A1(n12606), .A2(n12613), .ZN(n12598) );
  NAND2_X1 U15831 ( .A1(n12598), .A2(n12599), .ZN(n12633) );
  OAI21_X1 U15832 ( .B1(n12599), .B2(n12598), .A(n12633), .ZN(n12602) );
  NAND2_X1 U15833 ( .A1(n20196), .A2(n12600), .ZN(n12612) );
  INV_X1 U15834 ( .A(n12612), .ZN(n12601) );
  AOI21_X1 U15835 ( .B1(n12602), .B2(n12677), .A(n12601), .ZN(n12603) );
  NAND2_X1 U15836 ( .A1(n12604), .A2(n12603), .ZN(n13691) );
  NAND2_X1 U15837 ( .A1(n12605), .A2(n13860), .ZN(n12611) );
  XNOR2_X1 U15838 ( .A(n12606), .B(n12613), .ZN(n12608) );
  OAI211_X1 U15839 ( .C1(n11631), .C2(n12608), .A(n11558), .B(n12209), .ZN(
        n12609) );
  INV_X1 U15840 ( .A(n12609), .ZN(n12610) );
  NAND2_X1 U15841 ( .A1(n12611), .A2(n12610), .ZN(n12617) );
  INV_X1 U15842 ( .A(n12670), .ZN(n12627) );
  OAI21_X1 U15843 ( .B1(n11631), .B2(n12613), .A(n12612), .ZN(n12614) );
  INV_X1 U15844 ( .A(n12614), .ZN(n12615) );
  NAND2_X1 U15845 ( .A1(n13587), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12620) );
  INV_X1 U15846 ( .A(n13544), .ZN(n12618) );
  NAND2_X1 U15847 ( .A1(n12618), .A2(n12617), .ZN(n12619) );
  NAND2_X1 U15848 ( .A1(n13691), .A2(n13690), .ZN(n12624) );
  NAND2_X1 U15849 ( .A1(n12622), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12623) );
  INV_X1 U15850 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12625) );
  XNOR2_X1 U15851 ( .A(n12628), .B(n12625), .ZN(n13764) );
  XNOR2_X1 U15852 ( .A(n12633), .B(n12632), .ZN(n12626) );
  OAI22_X1 U15853 ( .A1(n20193), .A2(n12627), .B1(n11631), .B2(n12626), .ZN(
        n13766) );
  NAND2_X1 U15854 ( .A1(n13764), .A2(n13766), .ZN(n12630) );
  NAND2_X1 U15855 ( .A1(n12628), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12629) );
  NAND2_X1 U15856 ( .A1(n12630), .A2(n12629), .ZN(n13822) );
  NAND2_X1 U15857 ( .A1(n12631), .A2(n12670), .ZN(n12636) );
  NAND2_X1 U15858 ( .A1(n12633), .A2(n12632), .ZN(n12644) );
  XNOR2_X1 U15859 ( .A(n12644), .B(n12642), .ZN(n12634) );
  NAND2_X1 U15860 ( .A1(n12634), .A2(n12677), .ZN(n12635) );
  NAND2_X1 U15861 ( .A1(n12636), .A2(n12635), .ZN(n12638) );
  INV_X1 U15862 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12637) );
  XNOR2_X1 U15863 ( .A(n12638), .B(n12637), .ZN(n13824) );
  NAND2_X1 U15864 ( .A1(n13822), .A2(n13824), .ZN(n12640) );
  NAND2_X1 U15865 ( .A1(n12638), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12639) );
  NAND2_X1 U15866 ( .A1(n12640), .A2(n12639), .ZN(n13886) );
  NAND2_X1 U15867 ( .A1(n12641), .A2(n12670), .ZN(n12647) );
  INV_X1 U15868 ( .A(n12642), .ZN(n12643) );
  OR2_X1 U15869 ( .A1(n12644), .A2(n12643), .ZN(n12652) );
  XNOR2_X1 U15870 ( .A(n12652), .B(n12653), .ZN(n12645) );
  NAND2_X1 U15871 ( .A1(n12645), .A2(n12677), .ZN(n12646) );
  NAND2_X1 U15872 ( .A1(n12647), .A2(n12646), .ZN(n12648) );
  INV_X1 U15873 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13898) );
  XNOR2_X1 U15874 ( .A(n12648), .B(n13898), .ZN(n13888) );
  NAND2_X1 U15875 ( .A1(n13886), .A2(n13888), .ZN(n12650) );
  NAND2_X1 U15876 ( .A1(n12648), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12649) );
  NAND2_X1 U15877 ( .A1(n12650), .A2(n12649), .ZN(n15826) );
  NAND3_X1 U15878 ( .A1(n12674), .A2(n12651), .A3(n12670), .ZN(n12657) );
  INV_X1 U15879 ( .A(n12652), .ZN(n12654) );
  NAND2_X1 U15880 ( .A1(n12654), .A2(n12653), .ZN(n12661) );
  XNOR2_X1 U15881 ( .A(n12661), .B(n12662), .ZN(n12655) );
  NAND2_X1 U15882 ( .A1(n12655), .A2(n12677), .ZN(n12656) );
  NAND2_X1 U15883 ( .A1(n12658), .A2(n15986), .ZN(n15829) );
  NAND2_X1 U15884 ( .A1(n15826), .A2(n15829), .ZN(n12660) );
  INV_X1 U15885 ( .A(n12658), .ZN(n12659) );
  NAND2_X1 U15886 ( .A1(n12659), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15828) );
  NAND2_X1 U15887 ( .A1(n12660), .A2(n15828), .ZN(n15820) );
  INV_X1 U15888 ( .A(n12661), .ZN(n12663) );
  NAND2_X1 U15889 ( .A1(n12663), .A2(n12662), .ZN(n12675) );
  XNOR2_X1 U15890 ( .A(n12675), .B(n12676), .ZN(n12664) );
  AND2_X1 U15891 ( .A1(n12664), .A2(n12677), .ZN(n12665) );
  NAND2_X1 U15892 ( .A1(n15821), .A2(n15997), .ZN(n12666) );
  NAND2_X1 U15893 ( .A1(n15820), .A2(n12666), .ZN(n12669) );
  INV_X1 U15894 ( .A(n15821), .ZN(n12667) );
  NAND2_X1 U15895 ( .A1(n12667), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12668) );
  NAND2_X1 U15896 ( .A1(n12670), .A2(n12676), .ZN(n12672) );
  NOR2_X1 U15897 ( .A1(n12672), .A2(n12671), .ZN(n12673) );
  INV_X1 U15898 ( .A(n12675), .ZN(n12678) );
  NAND3_X1 U15899 ( .A1(n12678), .A2(n12677), .A3(n12676), .ZN(n12679) );
  NAND2_X1 U15900 ( .A1(n9712), .A2(n12679), .ZN(n13989) );
  INV_X1 U15901 ( .A(n13989), .ZN(n12681) );
  INV_X1 U15902 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15992) );
  NAND2_X1 U15903 ( .A1(n12681), .A2(n15992), .ZN(n12682) );
  NAND2_X1 U15904 ( .A1(n10011), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12684) );
  INV_X1 U15905 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15983) );
  NAND2_X1 U15906 ( .A1(n9711), .A2(n15983), .ZN(n12685) );
  NAND2_X1 U15907 ( .A1(n9757), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15793) );
  INV_X1 U15908 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15937) );
  NAND2_X1 U15909 ( .A1(n9712), .A2(n15937), .ZN(n12686) );
  NAND2_X1 U15910 ( .A1(n15790), .A2(n14775), .ZN(n15803) );
  NAND2_X1 U15911 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12687) );
  NAND2_X1 U15912 ( .A1(n9711), .A2(n12687), .ZN(n14773) );
  AND2_X1 U15913 ( .A1(n15803), .A2(n14773), .ZN(n12688) );
  NAND2_X1 U15914 ( .A1(n14776), .A2(n12688), .ZN(n15791) );
  INV_X1 U15915 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12689) );
  AND2_X1 U15916 ( .A1(n9711), .A2(n12689), .ZN(n12690) );
  INV_X1 U15917 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15889) );
  XNOR2_X1 U15918 ( .A(n9712), .B(n15889), .ZN(n15784) );
  INV_X1 U15919 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15976) );
  INV_X1 U15920 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15940) );
  NAND2_X1 U15921 ( .A1(n15976), .A2(n15940), .ZN(n12693) );
  NAND2_X1 U15922 ( .A1(n10011), .A2(n12693), .ZN(n14771) );
  NAND2_X1 U15923 ( .A1(n10011), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15804) );
  NAND2_X1 U15924 ( .A1(n10011), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12694) );
  AND2_X1 U15925 ( .A1(n15793), .A2(n12694), .ZN(n12695) );
  NAND2_X1 U15926 ( .A1(n10011), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14225) );
  NAND2_X1 U15927 ( .A1(n14224), .A2(n14225), .ZN(n15780) );
  NOR2_X1 U15928 ( .A1(n15780), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12696) );
  NAND2_X1 U15929 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  NAND2_X1 U15930 ( .A1(n10011), .A2(n15888), .ZN(n15675) );
  NAND2_X1 U15931 ( .A1(n9711), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12699) );
  INV_X1 U15932 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15679) );
  AND3_X1 U15933 ( .A1(n15874), .A2(n15888), .A3(n15679), .ZN(n12700) );
  INV_X1 U15934 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12701) );
  INV_X1 U15935 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15762) );
  INV_X1 U15936 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12813) );
  NAND2_X1 U15937 ( .A1(n15762), .A2(n12813), .ZN(n14695) );
  NAND2_X1 U15938 ( .A1(n14718), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14282) );
  NOR2_X1 U15939 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14800) );
  NAND2_X1 U15940 ( .A1(n14681), .A2(n10011), .ZN(n12705) );
  NAND3_X1 U15941 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14693) );
  NAND2_X1 U15942 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14794) );
  OR2_X1 U15943 ( .A1(n14693), .A2(n14794), .ZN(n12704) );
  XNOR2_X1 U15944 ( .A(n9711), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12706) );
  XNOR2_X1 U15945 ( .A(n12757), .B(n12706), .ZN(n14799) );
  INV_X1 U15946 ( .A(n12791), .ZN(n12708) );
  NAND2_X1 U15947 ( .A1(n14829), .A2(n20196), .ZN(n12707) );
  NAND3_X1 U15948 ( .A1(n12708), .A2(n11558), .A3(n12707), .ZN(n15628) );
  OR2_X1 U15949 ( .A1(n15646), .A2(n15628), .ZN(n12732) );
  NAND3_X1 U15950 ( .A1(n20761), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16013) );
  INV_X1 U15951 ( .A(n16013), .ZN(n12711) );
  NOR2_X2 U15952 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20636) );
  NAND2_X1 U15953 ( .A1(n20698), .A2(n12714), .ZN(n20863) );
  NAND2_X1 U15954 ( .A1(n20863), .A2(n20761), .ZN(n12712) );
  NAND2_X1 U15955 ( .A1(n20761), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15641) );
  NAND2_X1 U15956 ( .A1(n20633), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12713) );
  NAND2_X1 U15957 ( .A1(n15641), .A2(n12713), .ZN(n20164) );
  OR2_X2 U15958 ( .A1(n12714), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20177) );
  INV_X2 U15959 ( .A(n20177), .ZN(n16000) );
  NAND2_X1 U15960 ( .A1(n16000), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14792) );
  OAI21_X1 U15961 ( .B1(n15837), .B2(n12715), .A(n14792), .ZN(n12716) );
  AOI21_X1 U15962 ( .B1(n14435), .B2(n15809), .A(n12716), .ZN(n12717) );
  AOI22_X1 U15963 ( .A1(n12719), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12718), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12720) );
  NAND3_X1 U15964 ( .A1(n12726), .A2(n12725), .A3(n12724), .ZN(n12727) );
  OR2_X1 U15965 ( .A1(n12728), .A2(n12727), .ZN(n12730) );
  NAND2_X1 U15966 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20864) );
  NAND3_X1 U15967 ( .A1(n12723), .A2(n13386), .A3(n20864), .ZN(n12731) );
  NAND2_X1 U15968 ( .A1(n12732), .A2(n12731), .ZN(n12733) );
  NAND2_X1 U15969 ( .A1(n12733), .A2(n13852), .ZN(n13451) );
  INV_X1 U15970 ( .A(n20864), .ZN(n15671) );
  OR2_X1 U15971 ( .A1(n15646), .A2(n15671), .ZN(n15644) );
  OR2_X1 U15972 ( .A1(n15644), .A2(n12734), .ZN(n12735) );
  INV_X1 U15973 ( .A(n13852), .ZN(n13644) );
  NAND3_X1 U15974 ( .A1(n14411), .A2(n20234), .A3(n14670), .ZN(n12755) );
  NOR4_X1 U15975 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12742) );
  NOR4_X1 U15976 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12741) );
  NOR4_X1 U15977 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12740) );
  NOR4_X1 U15978 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12739) );
  AND4_X1 U15979 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n12739), .ZN(
        n12747) );
  NOR4_X1 U15980 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12745) );
  NOR4_X1 U15981 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12744) );
  NOR4_X1 U15982 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12743) );
  INV_X1 U15983 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20785) );
  AND4_X1 U15984 ( .A1(n12745), .A2(n12744), .A3(n12743), .A4(n20785), .ZN(
        n12746) );
  NAND2_X1 U15985 ( .A1(n12747), .A2(n12746), .ZN(n12748) );
  NOR3_X1 U15986 ( .A1(n14666), .A2(n20189), .A3(n11610), .ZN(n12749) );
  AOI22_X1 U15987 ( .A1(n14675), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14666), .ZN(n12750) );
  INV_X1 U15988 ( .A(n12750), .ZN(n12753) );
  NOR2_X1 U15989 ( .A1(n11610), .A2(n20190), .ZN(n12751) );
  NAND2_X1 U15990 ( .A1(n14670), .A2(n12751), .ZN(n14673) );
  INV_X1 U15991 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16462) );
  NOR2_X1 U15992 ( .A1(n14673), .A2(n16462), .ZN(n12752) );
  NOR2_X1 U15993 ( .A1(n12753), .A2(n12752), .ZN(n12754) );
  NAND2_X1 U15994 ( .A1(n12755), .A2(n12754), .ZN(P1_U2873) );
  INV_X1 U15995 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12821) );
  MUX2_X1 U15996 ( .A(n12756), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .S(
        n9712), .Z(n12758) );
  INV_X1 U15997 ( .A(n12761), .ZN(n12762) );
  NAND2_X1 U15998 ( .A1(n12762), .A2(n20772), .ZN(n15674) );
  AOI21_X1 U15999 ( .B1(n13860), .B2(n15674), .A(n15671), .ZN(n12763) );
  NAND2_X1 U16000 ( .A1(n13386), .A2(n12763), .ZN(n12768) );
  INV_X1 U16001 ( .A(n15674), .ZN(n15638) );
  OAI21_X1 U16002 ( .B1(n13860), .B2(n15638), .A(n20864), .ZN(n13856) );
  OAI211_X1 U16003 ( .C1(n13464), .C2(n13856), .A(n13854), .B(n11610), .ZN(
        n12765) );
  INV_X1 U16004 ( .A(n12765), .ZN(n12766) );
  OR2_X1 U16005 ( .A1(n15646), .A2(n12766), .ZN(n12767) );
  MUX2_X1 U16006 ( .A(n12768), .B(n12767), .S(n20213), .Z(n12775) );
  INV_X1 U16007 ( .A(n12769), .ZN(n12773) );
  NAND2_X1 U16008 ( .A1(n12723), .A2(n20196), .ZN(n13387) );
  INV_X1 U16009 ( .A(n15628), .ZN(n12771) );
  AND2_X1 U16010 ( .A1(n12769), .A2(n13854), .ZN(n12770) );
  NAND2_X1 U16011 ( .A1(n11637), .A2(n12770), .ZN(n12795) );
  NAND2_X1 U16012 ( .A1(n12771), .A2(n12795), .ZN(n12772) );
  AOI21_X1 U16013 ( .B1(n15646), .B2(n12773), .A(n13456), .ZN(n12774) );
  NAND2_X1 U16014 ( .A1(n12775), .A2(n12774), .ZN(n12776) );
  INV_X1 U16015 ( .A(n12777), .ZN(n12780) );
  BUF_X1 U16016 ( .A(n12778), .Z(n12797) );
  NOR2_X1 U16017 ( .A1(n12797), .A2(n13852), .ZN(n12779) );
  OR2_X1 U16018 ( .A1(n15628), .A2(n12779), .ZN(n13384) );
  OAI211_X1 U16019 ( .C1(n20221), .C2(n12786), .A(n12780), .B(n13384), .ZN(
        n12781) );
  AOI22_X1 U16020 ( .A1(n13546), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13380), .ZN(n12783) );
  OAI22_X1 U16021 ( .A1(n12785), .A2(n13860), .B1(n11536), .B2(n12786), .ZN(
        n12787) );
  NAND2_X1 U16022 ( .A1(n20228), .A2(n11581), .ZN(n12788) );
  NAND2_X1 U16023 ( .A1(n12788), .A2(n11619), .ZN(n12789) );
  OR2_X1 U16024 ( .A1(n12789), .A2(n13662), .ZN(n12790) );
  AOI22_X1 U16025 ( .A1(n12791), .A2(n13375), .B1(n13860), .B2(n12790), .ZN(
        n12794) );
  NAND2_X1 U16026 ( .A1(n12792), .A2(n13852), .ZN(n12793) );
  NAND3_X1 U16027 ( .A1(n12795), .A2(n12794), .A3(n12793), .ZN(n13467) );
  INV_X1 U16028 ( .A(n13467), .ZN(n12802) );
  OAI211_X1 U16029 ( .C1(n12797), .C2(n13857), .A(n9743), .B(n12796), .ZN(
        n13465) );
  NAND2_X1 U16030 ( .A1(n13465), .A2(n12798), .ZN(n12799) );
  NAND4_X1 U16031 ( .A1(n12802), .A2(n12801), .A3(n12800), .A4(n12799), .ZN(
        n12803) );
  NAND2_X1 U16032 ( .A1(n12807), .A2(n12803), .ZN(n15914) );
  INV_X1 U16033 ( .A(n13857), .ZN(n12804) );
  NAND2_X1 U16034 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15863) );
  NAND3_X1 U16035 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13889) );
  NOR3_X1 U16036 ( .A1(n12621), .A2(n13589), .A3(n13889), .ZN(n15964) );
  NAND3_X1 U16037 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15968) );
  NOR3_X1 U16038 ( .A1(n15976), .A2(n15983), .A3(n15968), .ZN(n15941) );
  NAND2_X1 U16039 ( .A1(n15964), .A2(n15941), .ZN(n15942) );
  NOR3_X1 U16040 ( .A1(n14775), .A2(n15940), .A3(n15942), .ZN(n15878) );
  NAND3_X1 U16041 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15881) );
  NOR4_X1 U16042 ( .A1(n15888), .A2(n15937), .A3(n12689), .A4(n15881), .ZN(
        n12805) );
  NAND2_X1 U16043 ( .A1(n15878), .A2(n12805), .ZN(n15681) );
  INV_X1 U16044 ( .A(n15966), .ZN(n15943) );
  AOI21_X1 U16045 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13768) );
  NOR2_X1 U16046 ( .A1(n13768), .A2(n13889), .ZN(n15965) );
  NAND3_X1 U16047 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15941), .A3(
        n15965), .ZN(n15944) );
  NOR2_X1 U16048 ( .A1(n14775), .A2(n15944), .ZN(n15917) );
  NAND2_X1 U16049 ( .A1(n12805), .A2(n15917), .ZN(n15682) );
  NAND2_X1 U16050 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12806) );
  AOI211_X1 U16051 ( .C1(n15681), .C2(n15943), .A(n15682), .B(n12806), .ZN(
        n12808) );
  INV_X1 U16052 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20172) );
  NOR2_X1 U16053 ( .A1(n16000), .A2(n12807), .ZN(n15919) );
  AOI21_X1 U16054 ( .B1(n15685), .B2(n20172), .A(n15919), .ZN(n15946) );
  OAI21_X1 U16055 ( .B1(n13892), .B2(n12808), .A(n15946), .ZN(n15861) );
  AOI21_X1 U16056 ( .B1(n15985), .B2(n15863), .A(n15861), .ZN(n15860) );
  OAI21_X1 U16057 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15916), .A(
        n15860), .ZN(n15851) );
  NAND2_X1 U16058 ( .A1(n15928), .A2(n14693), .ZN(n12811) );
  AOI22_X1 U16059 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(n15916), .B2(n15914), .ZN(
        n12809) );
  INV_X1 U16060 ( .A(n12809), .ZN(n12810) );
  NAND2_X1 U16061 ( .A1(n12811), .A2(n12810), .ZN(n12812) );
  NOR2_X1 U16062 ( .A1(n15851), .A2(n12812), .ZN(n15838) );
  NAND2_X1 U16063 ( .A1(n15838), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14811) );
  OR2_X1 U16064 ( .A1(n14811), .A2(n12813), .ZN(n12814) );
  NAND2_X1 U16065 ( .A1(n15838), .A2(n13892), .ZN(n12817) );
  NAND2_X1 U16066 ( .A1(n12814), .A2(n12817), .ZN(n14284) );
  NAND2_X1 U16067 ( .A1(n12817), .A2(n14794), .ZN(n12815) );
  NAND2_X1 U16068 ( .A1(n14284), .A2(n12815), .ZN(n14797) );
  OAI21_X1 U16069 ( .B1(n13892), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12816) );
  OR2_X1 U16070 ( .A1(n14797), .A2(n12816), .ZN(n14787) );
  AND3_X1 U16071 ( .A1(n14787), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12817), .ZN(n12818) );
  NOR2_X1 U16072 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15928), .ZN(
        n13594) );
  NOR2_X1 U16073 ( .A1(n15966), .A2(n13594), .ZN(n15850) );
  NAND2_X1 U16074 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15850), .ZN(
        n20186) );
  NAND3_X1 U16075 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n15875), .ZN(n15862) );
  INV_X1 U16076 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14697) );
  NOR2_X1 U16077 ( .A1(n14693), .A2(n14697), .ZN(n12819) );
  NAND2_X1 U16078 ( .A1(n15846), .A2(n12819), .ZN(n14802) );
  INV_X1 U16079 ( .A(n14794), .ZN(n14801) );
  NAND2_X1 U16080 ( .A1(n14801), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12820) );
  NOR2_X1 U16081 ( .A1(n14802), .A2(n12820), .ZN(n14788) );
  NOR2_X1 U16082 ( .A1(n12821), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12822) );
  INV_X1 U16083 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14421) );
  NOR2_X1 U16084 ( .A1(n20177), .A2(n14421), .ZN(n14349) );
  AOI21_X1 U16085 ( .B1(n14788), .B2(n12822), .A(n14349), .ZN(n12823) );
  NAND2_X1 U16086 ( .A1(n12824), .A2(n12848), .ZN(n12828) );
  NAND2_X1 U16087 ( .A1(n10549), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12825) );
  INV_X1 U16088 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19533) );
  AND2_X1 U16089 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19380) );
  NAND2_X1 U16090 ( .A1(n19380), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19273) );
  INV_X1 U16091 ( .A(n19380), .ZN(n19625) );
  NAND2_X1 U16092 ( .A1(n19625), .A2(n19933), .ZN(n12826) );
  AND2_X1 U16093 ( .A1(n19273), .A2(n12826), .ZN(n19418) );
  AND2_X1 U16094 ( .A1(n19418), .A2(n19934), .ZN(n19412) );
  AOI21_X1 U16095 ( .B1(n12845), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n19412), .ZN(n12827) );
  NAND2_X1 U16096 ( .A1(n12828), .A2(n12827), .ZN(n12830) );
  NAND2_X1 U16097 ( .A1(n12830), .A2(n12829), .ZN(n12841) );
  OAI21_X1 U16098 ( .B1(n12830), .B2(n12829), .A(n12841), .ZN(n13699) );
  INV_X1 U16099 ( .A(n13699), .ZN(n12840) );
  NAND2_X1 U16100 ( .A1(n12845), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12831) );
  NAND2_X1 U16101 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19943), .ZN(
        n19679) );
  NAND2_X1 U16102 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19950), .ZN(
        n19593) );
  NAND2_X1 U16103 ( .A1(n19679), .A2(n19593), .ZN(n19718) );
  NAND2_X1 U16104 ( .A1(n19934), .A2(n19718), .ZN(n19599) );
  NAND2_X1 U16105 ( .A1(n12831), .A2(n19599), .ZN(n12832) );
  AOI22_X1 U16106 ( .A1(n12845), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19934), .B2(n19950), .ZN(n12833) );
  INV_X1 U16107 ( .A(n13023), .ZN(n13071) );
  INV_X1 U16108 ( .A(n15375), .ZN(n12836) );
  NAND2_X1 U16109 ( .A1(n12836), .A2(n12835), .ZN(n12837) );
  INV_X1 U16110 ( .A(n13700), .ZN(n12839) );
  NAND2_X1 U16111 ( .A1(n12840), .A2(n12839), .ZN(n12842) );
  NAND2_X1 U16112 ( .A1(n12842), .A2(n12841), .ZN(n13599) );
  NAND2_X1 U16113 ( .A1(n19273), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12843) );
  NOR2_X1 U16114 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19933), .ZN(
        n19413) );
  NAND2_X1 U16115 ( .A1(n19380), .A2(n19413), .ZN(n19535) );
  NAND2_X1 U16116 ( .A1(n12843), .A2(n19535), .ZN(n12844) );
  AOI22_X1 U16117 ( .A1(n12845), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19934), .B2(n12844), .ZN(n12847) );
  INV_X1 U16118 ( .A(n12847), .ZN(n12849) );
  AND2_X1 U16119 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12850) );
  INV_X1 U16120 ( .A(n13740), .ZN(n12852) );
  NOR2_X1 U16121 ( .A1(n12854), .A2(n12850), .ZN(n12851) );
  NOR2_X2 U16122 ( .A1(n12852), .A2(n12851), .ZN(n13598) );
  NAND2_X1 U16123 ( .A1(n13599), .A2(n13598), .ZN(n13600) );
  NAND2_X1 U16124 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10549), .ZN(
        n12853) );
  NAND2_X1 U16125 ( .A1(n12854), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12855) );
  INV_X1 U16126 ( .A(n13879), .ZN(n12858) );
  INV_X1 U16127 ( .A(n12856), .ZN(n13794) );
  NAND2_X1 U16128 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13783) );
  NOR2_X1 U16129 ( .A1(n19319), .A2(n13783), .ZN(n13805) );
  AND2_X1 U16130 ( .A1(n13808), .A2(n13805), .ZN(n12857) );
  AND2_X1 U16131 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13804) );
  AOI22_X1 U16132 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U16133 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12865) );
  AOI22_X1 U16134 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U16135 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12863) );
  NAND4_X1 U16136 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n12872) );
  AOI22_X1 U16137 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U16138 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12869) );
  AOI22_X1 U16139 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12868) );
  AOI22_X1 U16140 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12867) );
  NAND4_X1 U16141 ( .A1(n12870), .A2(n12869), .A3(n12868), .A4(n12867), .ZN(
        n12871) );
  NOR2_X1 U16142 ( .A1(n12872), .A2(n12871), .ZN(n14210) );
  AOI22_X1 U16143 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10768), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U16144 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n12963), .ZN(n12875) );
  AOI22_X1 U16145 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12874) );
  AOI22_X1 U16146 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12873) );
  NAND4_X1 U16147 ( .A1(n12876), .A2(n12875), .A3(n12874), .A4(n12873), .ZN(
        n12882) );
  AOI22_X1 U16148 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U16149 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12970), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U16150 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10775), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U16151 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11244), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12877) );
  NAND4_X1 U16152 ( .A1(n12880), .A2(n12879), .A3(n12878), .A4(n12877), .ZN(
        n12881) );
  NOR2_X1 U16153 ( .A1(n12882), .A2(n12881), .ZN(n14124) );
  NOR2_X1 U16154 ( .A1(n14210), .A2(n14124), .ZN(n12893) );
  AOI22_X1 U16155 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U16156 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12885) );
  AOI22_X1 U16157 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12884) );
  AOI22_X1 U16158 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12883) );
  NAND4_X1 U16159 ( .A1(n12886), .A2(n12885), .A3(n12884), .A4(n12883), .ZN(
        n12892) );
  AOI22_X1 U16160 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16161 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16162 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U16163 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12887) );
  NAND4_X1 U16164 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n12887), .ZN(
        n12891) );
  OR2_X1 U16165 ( .A1(n12892), .A2(n12891), .ZN(n14144) );
  AND2_X1 U16166 ( .A1(n12893), .A2(n14144), .ZN(n14206) );
  AOI22_X1 U16167 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12897) );
  AOI22_X1 U16168 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U16169 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U16170 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12894) );
  NAND4_X1 U16171 ( .A1(n12897), .A2(n12896), .A3(n12895), .A4(n12894), .ZN(
        n12910) );
  INV_X1 U16172 ( .A(n12898), .ZN(n12903) );
  INV_X1 U16173 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12902) );
  INV_X1 U16174 ( .A(n12899), .ZN(n12901) );
  INV_X1 U16175 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12900) );
  OAI22_X1 U16176 ( .A1(n12903), .A2(n12902), .B1(n12901), .B2(n12900), .ZN(
        n12904) );
  INV_X1 U16177 ( .A(n12904), .ZN(n12908) );
  AOI22_X1 U16178 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U16179 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U16180 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12905) );
  NAND4_X1 U16181 ( .A1(n12908), .A2(n12907), .A3(n12906), .A4(n12905), .ZN(
        n12909) );
  NOR2_X1 U16182 ( .A1(n12910), .A2(n12909), .ZN(n14240) );
  INV_X1 U16183 ( .A(n14240), .ZN(n12911) );
  AND2_X1 U16184 ( .A1(n14206), .A2(n12911), .ZN(n12912) );
  AND2_X1 U16185 ( .A1(n12912), .A2(n14063), .ZN(n12913) );
  AND2_X2 U16186 ( .A1(n14015), .A2(n12913), .ZN(n14153) );
  AOI22_X1 U16187 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16188 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U16189 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U16190 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12914) );
  NAND4_X1 U16191 ( .A1(n12917), .A2(n12916), .A3(n12915), .A4(n12914), .ZN(
        n12923) );
  AOI22_X1 U16192 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U16193 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U16194 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U16195 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12918) );
  NAND4_X1 U16196 ( .A1(n12921), .A2(n12920), .A3(n12919), .A4(n12918), .ZN(
        n12922) );
  OR2_X1 U16197 ( .A1(n12923), .A2(n12922), .ZN(n14154) );
  AOI22_X1 U16198 ( .A1(n12962), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10768), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U16199 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U16200 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U16201 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12924) );
  NAND4_X1 U16202 ( .A1(n12927), .A2(n12926), .A3(n12925), .A4(n12924), .ZN(
        n12933) );
  AOI22_X1 U16203 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16204 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U16205 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U16206 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12928) );
  NAND4_X1 U16207 ( .A1(n12931), .A2(n12930), .A3(n12929), .A4(n12928), .ZN(
        n12932) );
  NOR2_X1 U16208 ( .A1(n12933), .A2(n12932), .ZN(n14221) );
  INV_X1 U16209 ( .A(n14221), .ZN(n12934) );
  AOI22_X1 U16210 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10768), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U16211 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12963), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U16212 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U16213 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12935) );
  NAND4_X1 U16214 ( .A1(n12938), .A2(n12937), .A3(n12936), .A4(n12935), .ZN(
        n12944) );
  AOI22_X1 U16215 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U16216 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12970), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U16217 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10775), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16218 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11244), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12939) );
  NAND4_X1 U16219 ( .A1(n12942), .A2(n12941), .A3(n12940), .A4(n12939), .ZN(
        n12943) );
  NOR2_X1 U16220 ( .A1(n12944), .A2(n12943), .ZN(n14938) );
  AOI22_X1 U16221 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13130), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12952) );
  INV_X1 U16222 ( .A(n13125), .ZN(n13101) );
  INV_X1 U16223 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12947) );
  OAI21_X1 U16224 ( .B1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n12945), .ZN(n13124) );
  NAND2_X1 U16225 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12946) );
  OAI211_X1 U16226 ( .C1(n13101), .C2(n12947), .A(n13124), .B(n12946), .ZN(
        n12948) );
  INV_X1 U16227 ( .A(n12948), .ZN(n12951) );
  AOI22_X1 U16228 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U16229 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13118), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12949) );
  NAND4_X1 U16230 ( .A1(n12952), .A2(n12951), .A3(n12950), .A4(n12949), .ZN(
        n12961) );
  AOI22_X1 U16231 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13082), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12959) );
  INV_X1 U16232 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12954) );
  INV_X1 U16233 ( .A(n13124), .ZN(n13119) );
  NAND2_X1 U16234 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12953) );
  OAI211_X1 U16235 ( .C1(n13101), .C2(n12954), .A(n13119), .B(n12953), .ZN(
        n12955) );
  INV_X1 U16236 ( .A(n12955), .ZN(n12958) );
  AOI22_X1 U16237 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U16238 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13118), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12956) );
  NAND4_X1 U16239 ( .A1(n12959), .A2(n12958), .A3(n12957), .A4(n12956), .ZN(
        n12960) );
  NAND2_X1 U16240 ( .A1(n12961), .A2(n12960), .ZN(n13004) );
  NOR2_X1 U16241 ( .A1(n19283), .A2(n13004), .ZN(n12979) );
  AOI22_X1 U16242 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10768), .B1(
        n12962), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U16243 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n12963), .ZN(n12968) );
  AOI22_X1 U16244 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16245 ( .A1(n10722), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12966) );
  NAND4_X1 U16246 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        n12978) );
  AOI22_X1 U16247 ( .A1(n12898), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12899), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12976) );
  AOI22_X1 U16248 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12970), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U16249 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10775), .B1(
        n12971), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U16250 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11244), .B1(
        n12972), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12973) );
  NAND4_X1 U16251 ( .A1(n12976), .A2(n12975), .A3(n12974), .A4(n12973), .ZN(
        n12977) );
  NOR2_X1 U16252 ( .A1(n12978), .A2(n12977), .ZN(n12997) );
  XNOR2_X1 U16253 ( .A(n12979), .B(n12997), .ZN(n13002) );
  XNOR2_X1 U16254 ( .A(n12980), .B(n13002), .ZN(n14930) );
  INV_X1 U16255 ( .A(n13004), .ZN(n12998) );
  NAND2_X1 U16256 ( .A1(n19283), .A2(n12998), .ZN(n14929) );
  OR2_X2 U16257 ( .A1(n14930), .A2(n14929), .ZN(n14927) );
  AOI22_X1 U16258 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13132), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12987) );
  INV_X1 U16259 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12982) );
  NAND2_X1 U16260 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12981) );
  OAI211_X1 U16261 ( .C1(n13101), .C2(n12982), .A(n13124), .B(n12981), .ZN(
        n12983) );
  INV_X1 U16262 ( .A(n12983), .ZN(n12986) );
  AOI22_X1 U16263 ( .A1(n13130), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16264 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12984) );
  NAND4_X1 U16265 ( .A1(n12987), .A2(n12986), .A3(n12985), .A4(n12984), .ZN(
        n12996) );
  AOI22_X1 U16266 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13082), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12994) );
  NAND2_X1 U16267 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12988) );
  OAI211_X1 U16268 ( .C1(n13101), .C2(n12989), .A(n13119), .B(n12988), .ZN(
        n12990) );
  INV_X1 U16269 ( .A(n12990), .ZN(n12993) );
  AOI22_X1 U16270 ( .A1(n13130), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16271 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12991) );
  NAND4_X1 U16272 ( .A1(n12994), .A2(n12993), .A3(n12992), .A4(n12991), .ZN(
        n12995) );
  AND2_X1 U16273 ( .A1(n12996), .A2(n12995), .ZN(n13003) );
  INV_X1 U16274 ( .A(n12997), .ZN(n12999) );
  AND2_X1 U16275 ( .A1(n12999), .A2(n12998), .ZN(n13000) );
  NAND2_X1 U16276 ( .A1(n13000), .A2(n13003), .ZN(n13006) );
  OAI211_X1 U16277 ( .C1(n13003), .C2(n13000), .A(n13006), .B(n13023), .ZN(
        n14916) );
  INV_X1 U16278 ( .A(n13002), .ZN(n13005) );
  NAND2_X1 U16279 ( .A1(n19283), .A2(n13003), .ZN(n14919) );
  INV_X1 U16280 ( .A(n13006), .ZN(n13024) );
  AOI22_X1 U16281 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13132), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13013) );
  INV_X1 U16282 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13008) );
  NAND2_X1 U16283 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13007) );
  OAI211_X1 U16284 ( .C1(n13101), .C2(n13008), .A(n13124), .B(n13007), .ZN(
        n13009) );
  INV_X1 U16285 ( .A(n13009), .ZN(n13012) );
  AOI22_X1 U16286 ( .A1(n13130), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U16287 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13010) );
  NAND4_X1 U16288 ( .A1(n13013), .A2(n13012), .A3(n13011), .A4(n13010), .ZN(
        n13022) );
  AOI22_X1 U16289 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13132), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13020) );
  INV_X1 U16290 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13015) );
  NAND2_X1 U16291 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13014) );
  OAI211_X1 U16292 ( .C1(n13101), .C2(n13015), .A(n13119), .B(n13014), .ZN(
        n13016) );
  INV_X1 U16293 ( .A(n13016), .ZN(n13019) );
  AOI22_X1 U16294 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U16295 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9737), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13017) );
  NAND4_X1 U16296 ( .A1(n13020), .A2(n13019), .A3(n13018), .A4(n13017), .ZN(
        n13021) );
  AND2_X1 U16297 ( .A1(n13022), .A2(n13021), .ZN(n13025) );
  NAND2_X1 U16298 ( .A1(n13024), .A2(n13025), .ZN(n13048) );
  OAI211_X1 U16299 ( .C1(n13024), .C2(n13025), .A(n13048), .B(n13023), .ZN(
        n13028) );
  INV_X1 U16300 ( .A(n13025), .ZN(n13026) );
  NOR2_X1 U16301 ( .A1(n11191), .A2(n13026), .ZN(n14910) );
  INV_X1 U16302 ( .A(n13027), .ZN(n13030) );
  AOI22_X1 U16303 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13082), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U16304 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13032) );
  OAI211_X1 U16305 ( .C1(n13101), .C2(n13033), .A(n13124), .B(n13032), .ZN(
        n13034) );
  INV_X1 U16306 ( .A(n13034), .ZN(n13037) );
  AOI22_X1 U16307 ( .A1(n13130), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U16308 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13035) );
  NAND4_X1 U16309 ( .A1(n13038), .A2(n13037), .A3(n13036), .A4(n13035), .ZN(
        n13047) );
  AOI22_X1 U16310 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13132), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13045) );
  INV_X1 U16311 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13040) );
  NAND2_X1 U16312 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13039) );
  OAI211_X1 U16313 ( .C1(n13101), .C2(n13040), .A(n13119), .B(n13039), .ZN(
        n13041) );
  INV_X1 U16314 ( .A(n13041), .ZN(n13044) );
  AOI22_X1 U16315 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U16316 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13042) );
  NAND4_X1 U16317 ( .A1(n13045), .A2(n13044), .A3(n13043), .A4(n13042), .ZN(
        n13046) );
  NAND2_X1 U16318 ( .A1(n13047), .A2(n13046), .ZN(n13050) );
  AOI21_X1 U16319 ( .B1(n13048), .B2(n13050), .A(n13071), .ZN(n13049) );
  OR2_X1 U16320 ( .A1(n13048), .A2(n13050), .ZN(n13072) );
  NAND2_X1 U16321 ( .A1(n13049), .A2(n13072), .ZN(n13052) );
  NOR2_X1 U16322 ( .A1(n11191), .A2(n13050), .ZN(n14900) );
  AOI22_X1 U16323 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13082), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13061) );
  INV_X1 U16324 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13056) );
  NAND2_X1 U16325 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13055) );
  OAI211_X1 U16326 ( .C1(n13101), .C2(n13056), .A(n13124), .B(n13055), .ZN(
        n13057) );
  INV_X1 U16327 ( .A(n13057), .ZN(n13060) );
  AOI22_X1 U16328 ( .A1(n13130), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U16329 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13058) );
  NAND4_X1 U16330 ( .A1(n13061), .A2(n13060), .A3(n13059), .A4(n13058), .ZN(
        n13070) );
  AOI22_X1 U16331 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13082), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13068) );
  INV_X1 U16332 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13063) );
  NAND2_X1 U16333 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13062) );
  OAI211_X1 U16334 ( .C1(n13101), .C2(n13063), .A(n13119), .B(n13062), .ZN(
        n13064) );
  INV_X1 U16335 ( .A(n13064), .ZN(n13067) );
  AOI22_X1 U16336 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16337 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9737), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13065) );
  NAND4_X1 U16338 ( .A1(n13068), .A2(n13067), .A3(n13066), .A4(n13065), .ZN(
        n13069) );
  NAND2_X1 U16339 ( .A1(n13070), .A2(n13069), .ZN(n13074) );
  NOR2_X1 U16340 ( .A1(n13072), .A2(n13074), .ZN(n14885) );
  AOI211_X1 U16341 ( .C1(n13072), .C2(n13074), .A(n13071), .B(n14885), .ZN(
        n13073) );
  NOR2_X1 U16342 ( .A1(n11196), .A2(n13074), .ZN(n14894) );
  AOI22_X1 U16343 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13082), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U16344 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13075) );
  OAI211_X1 U16345 ( .C1(n13101), .C2(n13076), .A(n13124), .B(n13075), .ZN(
        n13077) );
  INV_X1 U16346 ( .A(n13077), .ZN(n13080) );
  AOI22_X1 U16347 ( .A1(n13130), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13079) );
  AOI22_X1 U16348 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13078) );
  NAND4_X1 U16349 ( .A1(n13081), .A2(n13080), .A3(n13079), .A4(n13078), .ZN(
        n13091) );
  AOI22_X1 U16350 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13082), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13089) );
  INV_X1 U16351 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13084) );
  NAND2_X1 U16352 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13083) );
  OAI211_X1 U16353 ( .C1(n13101), .C2(n13084), .A(n13119), .B(n13083), .ZN(
        n13085) );
  INV_X1 U16354 ( .A(n13085), .ZN(n13088) );
  AOI22_X1 U16355 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16356 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13086) );
  NAND4_X1 U16357 ( .A1(n13089), .A2(n13088), .A3(n13087), .A4(n13086), .ZN(
        n13090) );
  NAND2_X1 U16358 ( .A1(n13091), .A2(n13090), .ZN(n13109) );
  AOI21_X1 U16359 ( .B1(n14893), .B2(n14887), .A(n13109), .ZN(n14880) );
  AOI22_X1 U16360 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13130), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13098) );
  NAND2_X1 U16361 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13092) );
  OAI211_X1 U16362 ( .C1(n13101), .C2(n13093), .A(n13124), .B(n13092), .ZN(
        n13094) );
  INV_X1 U16363 ( .A(n13094), .ZN(n13097) );
  AOI22_X1 U16364 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U16365 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13095) );
  NAND4_X1 U16366 ( .A1(n13098), .A2(n13097), .A3(n13096), .A4(n13095), .ZN(
        n13108) );
  AOI22_X1 U16367 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9708), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13106) );
  INV_X1 U16368 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13100) );
  NAND2_X1 U16369 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13099) );
  OAI211_X1 U16370 ( .C1(n13101), .C2(n13100), .A(n13119), .B(n13099), .ZN(
        n13102) );
  INV_X1 U16371 ( .A(n13102), .ZN(n13105) );
  AOI22_X1 U16372 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U16373 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13103) );
  NAND4_X1 U16374 ( .A1(n13106), .A2(n13105), .A3(n13104), .A4(n13103), .ZN(
        n13107) );
  NAND2_X1 U16375 ( .A1(n13108), .A2(n13107), .ZN(n13112) );
  INV_X1 U16376 ( .A(n13109), .ZN(n14888) );
  AND2_X1 U16377 ( .A1(n11196), .A2(n14888), .ZN(n13110) );
  NAND2_X1 U16378 ( .A1(n14885), .A2(n13110), .ZN(n13111) );
  NOR2_X1 U16379 ( .A1(n13111), .A2(n13112), .ZN(n13113) );
  AOI21_X1 U16380 ( .B1(n13112), .B2(n13111), .A(n13113), .ZN(n14879) );
  NAND2_X1 U16381 ( .A1(n14880), .A2(n14879), .ZN(n14881) );
  INV_X1 U16382 ( .A(n13113), .ZN(n13114) );
  NAND2_X1 U16383 ( .A1(n14881), .A2(n13114), .ZN(n13141) );
  AOI22_X1 U16384 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13130), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13116) );
  NAND2_X1 U16385 ( .A1(n13131), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13115) );
  OAI211_X1 U16386 ( .C1(n13117), .C2(n19319), .A(n13116), .B(n13115), .ZN(
        n13138) );
  INV_X1 U16387 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16388 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13118), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13121) );
  AOI21_X1 U16389 ( .B1(n13125), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n13119), .ZN(n13120) );
  OAI211_X1 U16390 ( .C1(n13122), .C2(n13129), .A(n13121), .B(n13120), .ZN(
        n13137) );
  INV_X1 U16391 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16392 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13123), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13127) );
  AOI21_X1 U16393 ( .B1(n13125), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n13124), .ZN(n13126) );
  OAI211_X1 U16394 ( .C1(n13129), .C2(n13128), .A(n13127), .B(n13126), .ZN(
        n13136) );
  AOI22_X1 U16395 ( .A1(n9723), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9708), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U16396 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13131), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13133) );
  NAND2_X1 U16397 ( .A1(n13134), .A2(n13133), .ZN(n13135) );
  OAI22_X1 U16398 ( .A1(n13138), .A2(n13137), .B1(n13136), .B2(n13135), .ZN(
        n13139) );
  INV_X1 U16399 ( .A(n13139), .ZN(n13140) );
  XNOR2_X1 U16400 ( .A(n13141), .B(n13140), .ZN(n14410) );
  AND2_X1 U16401 ( .A1(n11186), .A2(n16339), .ZN(n16348) );
  AND2_X1 U16402 ( .A1(n13142), .A2(n19822), .ZN(n16346) );
  AOI22_X1 U16403 ( .A1(n13143), .A2(n16344), .B1(n16348), .B2(n16346), .ZN(
        n13366) );
  NAND2_X1 U16404 ( .A1(n13366), .A2(n13144), .ZN(n13145) );
  NOR4_X1 U16405 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n13151) );
  NOR4_X1 U16406 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n13150) );
  NOR4_X1 U16407 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13149) );
  NOR4_X1 U16408 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13148) );
  NAND4_X1 U16409 ( .A1(n13151), .A2(n13150), .A3(n13149), .A4(n13148), .ZN(
        n13156) );
  NOR4_X1 U16410 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13154) );
  NOR4_X1 U16411 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n13153) );
  NOR4_X1 U16412 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n13152) );
  INV_X1 U16413 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19857) );
  NAND4_X1 U16414 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n19857), .ZN(
        n13155) );
  OAI21_X1 U16415 ( .B1(n13156), .B2(n13155), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13157) );
  MUX2_X1 U16416 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n16122), .Z(n19230) );
  AOI21_X1 U16417 ( .B1(n13159), .B2(n14952), .A(n13158), .ZN(n16041) );
  INV_X1 U16418 ( .A(n16041), .ZN(n13162) );
  NAND2_X1 U16419 ( .A1(n19132), .A2(n13160), .ZN(n16124) );
  INV_X1 U16420 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13161) );
  OAI22_X1 U16421 ( .A1(n13162), .A2(n16124), .B1(n19132), .B2(n13161), .ZN(
        n13163) );
  AOI21_X1 U16422 ( .B1(n19105), .B2(n19230), .A(n13163), .ZN(n13165) );
  NAND2_X1 U16423 ( .A1(n19132), .A2(n9848), .ZN(n13553) );
  NOR2_X2 U16424 ( .A1(n13553), .A2(n16122), .ZN(n19106) );
  NOR2_X2 U16425 ( .A1(n13553), .A2(n16121), .ZN(n19107) );
  AOI22_X1 U16426 ( .A1(n19106), .A2(BUF1_REG_30__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n13164) );
  OAI21_X1 U16427 ( .B1(n14410), .B2(n19162), .A(n13166), .ZN(P2_U2889) );
  NOR3_X1 U16428 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20861), .ZN(n13168) );
  NOR4_X1 U16429 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13167) );
  NAND4_X1 U16430 ( .A1(n20189), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13168), .A4(
        n13167), .ZN(U214) );
  INV_X1 U16431 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19952) );
  NOR2_X1 U16432 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n19952), .ZN(n13170) );
  NOR4_X1 U16433 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13169) );
  NAND4_X1 U16434 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13170), .A3(n13169), .A4(
        n19902), .ZN(n13171) );
  NOR2_X1 U16435 ( .A1(n16122), .A2(n13171), .ZN(n16461) );
  NAND2_X1 U16436 ( .A1(n16461), .A2(U214), .ZN(U212) );
  NOR2_X1 U16437 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13171), .ZN(n16534)
         );
  AND2_X1 U16438 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13173) );
  INV_X1 U16439 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16085) );
  NAND2_X1 U16440 ( .A1(n13182), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13177) );
  INV_X1 U16441 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15056) );
  INV_X1 U16442 ( .A(n13175), .ZN(n13207) );
  NAND2_X1 U16443 ( .A1(n13207), .A2(n9862), .ZN(n13176) );
  NAND2_X1 U16444 ( .A1(n15047), .A2(n13176), .ZN(n14370) );
  INV_X1 U16445 ( .A(n14370), .ZN(n13210) );
  OR2_X1 U16446 ( .A1(n13182), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13178) );
  NAND2_X1 U16447 ( .A1(n13177), .A2(n13178), .ZN(n15067) );
  INV_X1 U16448 ( .A(n15067), .ZN(n16071) );
  INV_X1 U16449 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15048) );
  INV_X1 U16450 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13179) );
  AOI21_X1 U16451 ( .B1(n16085), .B2(n13181), .A(n13182), .ZN(n16084) );
  OAI21_X1 U16452 ( .B1(n13183), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n13181), .ZN(n15080) );
  INV_X1 U16453 ( .A(n15080), .ZN(n16099) );
  AOI21_X1 U16454 ( .B1(n13174), .B2(n13184), .A(n13183), .ZN(n16108) );
  OAI21_X1 U16455 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13186), .A(
        n13184), .ZN(n16141) );
  INV_X1 U16456 ( .A(n16141), .ZN(n15605) );
  INV_X1 U16457 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15097) );
  NAND2_X1 U16458 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n13185), .ZN(
        n13205) );
  AOI21_X1 U16459 ( .B1(n15097), .B2(n13205), .A(n13186), .ZN(n15099) );
  INV_X1 U16460 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14272) );
  AOI21_X1 U16461 ( .B1(n14272), .B2(n13187), .A(n13185), .ZN(n18897) );
  AOI21_X1 U16462 ( .B1(n18921), .B2(n13188), .A(n13189), .ZN(n18920) );
  AOI21_X1 U16463 ( .B1(n18941), .B2(n13203), .A(n13190), .ZN(n18949) );
  INV_X1 U16464 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16170) );
  AND2_X1 U16465 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n13191), .ZN(
        n13204) );
  AOI21_X1 U16466 ( .B1(n16170), .B2(n13202), .A(n13204), .ZN(n16163) );
  AOI21_X1 U16467 ( .B1(n18978), .B2(n13200), .A(n13192), .ZN(n18984) );
  INV_X1 U16468 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19001) );
  NAND2_X1 U16469 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n13193), .ZN(
        n13199) );
  AOI21_X1 U16470 ( .B1(n19001), .B2(n13199), .A(n13201), .ZN(n19007) );
  INV_X1 U16471 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15139) );
  NAND2_X1 U16472 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n13198), .ZN(
        n13197) );
  AOI21_X1 U16473 ( .B1(n15139), .B2(n13197), .A(n13193), .ZN(n19025) );
  AOI21_X1 U16474 ( .B1(n16225), .B2(n13196), .A(n13198), .ZN(n19052) );
  AOI21_X1 U16475 ( .B1(n16240), .B2(n13195), .A(n13194), .ZN(n16226) );
  AOI22_X1 U16476 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n10835), .B1(n19077), 
        .B2(n19969), .ZN(n19076) );
  AOI22_X1 U16477 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14379), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19969), .ZN(n13904) );
  NOR2_X1 U16478 ( .A1(n19076), .A2(n13904), .ZN(n13903) );
  OAI21_X1 U16479 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13195), .ZN(n13831) );
  NAND2_X1 U16480 ( .A1(n13903), .A2(n13831), .ZN(n13704) );
  NOR2_X1 U16481 ( .A1(n16226), .A2(n13704), .ZN(n19068) );
  OAI21_X1 U16482 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13194), .A(
        n13196), .ZN(n19268) );
  NAND2_X1 U16483 ( .A1(n19068), .A2(n19268), .ZN(n19050) );
  OAI21_X1 U16484 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13198), .A(
        n13197), .ZN(n19040) );
  OAI21_X1 U16485 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13193), .A(
        n13199), .ZN(n19017) );
  NOR2_X1 U16486 ( .A1(n19007), .A2(n19005), .ZN(n18993) );
  OAI21_X1 U16487 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13201), .A(
        n13200), .ZN(n18994) );
  NAND2_X1 U16488 ( .A1(n18993), .A2(n18994), .ZN(n18982) );
  OAI21_X1 U16489 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13192), .A(
        n13202), .ZN(n18972) );
  OAI21_X1 U16490 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13204), .A(
        n13203), .ZN(n18962) );
  NOR2_X1 U16491 ( .A1(n18949), .A2(n18948), .ZN(n18934) );
  OAI21_X1 U16492 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13190), .A(
        n13188), .ZN(n18935) );
  NAND2_X1 U16493 ( .A1(n18934), .A2(n18935), .ZN(n18918) );
  OR2_X1 U16494 ( .A1(n13185), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13206) );
  AND2_X1 U16495 ( .A1(n13206), .A2(n13205), .ZN(n14868) );
  INV_X1 U16496 ( .A(n14868), .ZN(n15117) );
  NOR2_X1 U16497 ( .A1(n19069), .A2(n15603), .ZN(n16107) );
  NOR2_X1 U16498 ( .A1(n16084), .A2(n16082), .ZN(n16083) );
  NOR2_X1 U16499 ( .A1(n19069), .A2(n16083), .ZN(n16070) );
  NOR2_X1 U16500 ( .A1(n16071), .A2(n16070), .ZN(n16069) );
  NOR2_X1 U16501 ( .A1(n16069), .A2(n19069), .ZN(n16063) );
  AOI21_X1 U16502 ( .B1(n15056), .B2(n13177), .A(n13175), .ZN(n16064) );
  NOR4_X4 U16503 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n15374), .ZN(n19055) );
  AOI211_X1 U16504 ( .C1(n13210), .C2(n13209), .A(n19825), .B(n16029), .ZN(
        n13235) );
  NAND2_X1 U16505 ( .A1(n16339), .A2(n16367), .ZN(n13348) );
  OR2_X1 U16506 ( .A1(n13211), .A2(n13348), .ZN(n13349) );
  NOR2_X1 U16507 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13363), .ZN(n13230) );
  INV_X1 U16508 ( .A(n13230), .ZN(n13212) );
  NAND2_X1 U16509 ( .A1(n19245), .A2(n13212), .ZN(n16026) );
  INV_X1 U16510 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19914) );
  AND2_X1 U16511 ( .A1(n19822), .A2(n19914), .ZN(n13213) );
  NOR2_X1 U16512 ( .A1(n13349), .A2(n13213), .ZN(n13219) );
  INV_X1 U16513 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14876) );
  NAND2_X1 U16514 ( .A1(n13219), .A2(n14876), .ZN(n13214) );
  NAND2_X2 U16515 ( .A1(n16026), .A2(n13214), .ZN(n19058) );
  NAND2_X1 U16516 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19973), .ZN(n19820) );
  NOR2_X1 U16517 ( .A1(n19828), .A2(n19820), .ZN(n16366) );
  NAND2_X1 U16518 ( .A1(n9722), .A2(n19825), .ZN(n13215) );
  OR2_X1 U16519 ( .A1(n16366), .A2(n13215), .ZN(n13216) );
  AOI22_X1 U16520 ( .A1(n19058), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19081), .ZN(n13217) );
  INV_X1 U16521 ( .A(n13217), .ZN(n13234) );
  AND2_X1 U16522 ( .A1(n11191), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13218) );
  OAI22_X1 U16523 ( .A1(n13220), .A2(n19063), .B1(n9862), .B2(n19079), .ZN(
        n13233) );
  NOR2_X1 U16524 ( .A1(n13222), .A2(n13223), .ZN(n13224) );
  NAND2_X1 U16525 ( .A1(n11191), .A2(n19822), .ZN(n13225) );
  OR2_X1 U16526 ( .A1(n13227), .A2(n13228), .ZN(n13229) );
  NAND2_X1 U16527 ( .A1(n13226), .A2(n13229), .ZN(n14362) );
  AND2_X1 U16528 ( .A1(n13231), .A2(n13230), .ZN(n16369) );
  OAI22_X1 U16529 ( .A1(n14890), .A2(n19075), .B1(n14362), .B2(n19083), .ZN(
        n13232) );
  OR4_X1 U16530 ( .A1(n13235), .A2(n13234), .A3(n13233), .A4(n13232), .ZN(
        P2_U2827) );
  NOR2_X1 U16531 ( .A1(n18162), .A2(n18735), .ZN(n17844) );
  NOR2_X1 U16532 ( .A1(n16398), .A2(n18191), .ZN(n13242) );
  NOR2_X1 U16533 ( .A1(n13236), .A2(n13242), .ZN(n18858) );
  AOI21_X1 U16534 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18150) );
  INV_X1 U16535 ( .A(n18150), .ZN(n13251) );
  NAND2_X1 U16536 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15485) );
  INV_X1 U16537 ( .A(n15485), .ZN(n13252) );
  INV_X1 U16538 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18828) );
  INV_X1 U16539 ( .A(n13239), .ZN(n18645) );
  NOR3_X1 U16540 ( .A1(n18850), .A2(n13240), .A3(n18631), .ZN(n13249) );
  INV_X1 U16541 ( .A(n13241), .ZN(n18667) );
  OAI21_X1 U16542 ( .B1(n18226), .B2(n18667), .A(n13242), .ZN(n13265) );
  AOI21_X1 U16543 ( .B1(n13243), .B2(n13265), .A(n18204), .ZN(n13244) );
  AOI21_X1 U16544 ( .B1(n13245), .B2(n18204), .A(n13244), .ZN(n13246) );
  INV_X1 U16545 ( .A(n13246), .ZN(n13248) );
  NOR3_X2 U16546 ( .A1(n13249), .A2(n13248), .A3(n13247), .ZN(n18644) );
  AOI21_X1 U16547 ( .B1(n18668), .B2(n18828), .A(n18145), .ZN(n16452) );
  AOI22_X1 U16548 ( .A1(n18664), .A2(n13251), .B1(n13252), .B2(n16452), .ZN(
        n18128) );
  INV_X1 U16549 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18127) );
  NAND2_X1 U16550 ( .A1(n18666), .A2(n18828), .ZN(n17974) );
  INV_X1 U16551 ( .A(n17974), .ZN(n18149) );
  OAI22_X1 U16552 ( .A1(n18145), .A2(n13252), .B1(n18144), .B2(n13251), .ZN(
        n13253) );
  NOR3_X1 U16553 ( .A1(n18149), .A2(n18127), .A3(n13253), .ZN(n18135) );
  INV_X1 U16554 ( .A(n13254), .ZN(n13257) );
  AOI211_X1 U16555 ( .C1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(n18831), .A(
        n13256), .B(n13255), .ZN(n13259) );
  AOI21_X1 U16556 ( .B1(n13257), .B2(n13259), .A(n16554), .ZN(n18638) );
  NOR2_X1 U16557 ( .A1(n18850), .A2(n18217), .ZN(n13262) );
  AOI22_X1 U16558 ( .A1(n18638), .A2(n13262), .B1(n13261), .B2(n18635), .ZN(
        n13271) );
  INV_X1 U16559 ( .A(n16554), .ZN(n18637) );
  NOR2_X1 U16560 ( .A1(n13269), .A2(n18850), .ZN(n13272) );
  AOI21_X1 U16561 ( .B1(n13269), .B2(n18850), .A(n13272), .ZN(n13263) );
  AOI21_X1 U16562 ( .B1(n18848), .B2(n13263), .A(n18722), .ZN(n16553) );
  OAI211_X1 U16563 ( .C1(n13269), .C2(n18213), .A(n18637), .B(n16553), .ZN(
        n13264) );
  INV_X1 U16564 ( .A(n13264), .ZN(n13268) );
  OAI211_X1 U16565 ( .C1(n16546), .C2(n13267), .A(n13266), .B(n13265), .ZN(
        n14246) );
  AOI211_X1 U16566 ( .C1(n18635), .C2(n15394), .A(n13268), .B(n14246), .ZN(
        n13270) );
  AOI221_X4 U16567 ( .B1(n13271), .B2(n13270), .C1(n13269), .C2(n13270), .A(
        n18697), .ZN(n18169) );
  AOI211_X1 U16568 ( .C1(n18128), .C2(n18127), .A(n18135), .B(n18159), .ZN(
        n13339) );
  NAND2_X1 U16569 ( .A1(n16380), .A2(n18169), .ZN(n18173) );
  AOI22_X1 U16570 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U16571 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15508), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13286) );
  INV_X1 U16572 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17220) );
  AOI22_X1 U16573 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13275) );
  OAI21_X1 U16574 ( .B1(n9761), .B2(n17220), .A(n13275), .ZN(n13284) );
  AOI22_X1 U16575 ( .A1(n13288), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13276), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U16576 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16577 ( .A1(n13278), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U16578 ( .A1(n13289), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13279) );
  NAND4_X1 U16579 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n13283) );
  AOI211_X1 U16580 ( .C1(n17175), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n13284), .B(n13283), .ZN(n13285) );
  NAND3_X1 U16581 ( .A1(n13287), .A2(n13286), .A3(n13285), .ZN(n17370) );
  AOI22_X1 U16582 ( .A1(n13288), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n10188), .ZN(n13301) );
  AOI22_X1 U16583 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17177), .B1(
        n13274), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U16584 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n13290), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13289), .ZN(n13291) );
  OAI21_X1 U16585 ( .B1(n15511), .B2(n15438), .A(n13291), .ZN(n13292) );
  INV_X1 U16586 ( .A(n13292), .ZN(n13298) );
  AOI22_X1 U16587 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17174), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U16588 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n13293), .ZN(n13296) );
  AOI22_X1 U16589 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17116), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U16590 ( .A1(n13278), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17080), .ZN(n13294) );
  XNOR2_X1 U16591 ( .A(n17370), .B(n13329), .ZN(n13303) );
  NAND2_X1 U16592 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13303), .ZN(
        n13315) );
  NAND2_X1 U16593 ( .A1(n13329), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13314) );
  AOI22_X1 U16594 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13307) );
  AOI22_X1 U16595 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15508), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U16596 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U16597 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13304) );
  NAND4_X1 U16598 ( .A1(n13307), .A2(n13306), .A3(n13305), .A4(n13304), .ZN(
        n13313) );
  AOI22_X1 U16599 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13311) );
  AOI22_X1 U16600 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U16601 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17116), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U16602 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13308) );
  NAND4_X1 U16603 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n13308), .ZN(
        n13312) );
  NOR2_X1 U16604 ( .A1(n17871), .A2(n18828), .ZN(n17870) );
  NAND2_X1 U16605 ( .A1(n17865), .A2(n17870), .ZN(n17864) );
  NAND2_X1 U16606 ( .A1(n13314), .A2(n17864), .ZN(n17851) );
  NAND2_X1 U16607 ( .A1(n17852), .A2(n17851), .ZN(n17850) );
  NAND2_X1 U16608 ( .A1(n13315), .A2(n17850), .ZN(n15559) );
  AOI22_X1 U16609 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13319) );
  AOI22_X1 U16610 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U16611 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U16612 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13316) );
  NAND4_X1 U16613 ( .A1(n13319), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n13325) );
  AOI22_X1 U16614 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15508), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U16615 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13322) );
  AOI22_X1 U16616 ( .A1(n15523), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U16617 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13320) );
  NAND4_X1 U16618 ( .A1(n13323), .A2(n13322), .A3(n13321), .A4(n13320), .ZN(
        n13324) );
  NAND2_X1 U16619 ( .A1(n17376), .A2(n17370), .ZN(n15552) );
  XOR2_X1 U16620 ( .A(n17364), .B(n15552), .Z(n15560) );
  OAI21_X1 U16621 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13327), .A(
        n15561), .ZN(n17841) );
  NOR2_X1 U16622 ( .A1(n18173), .A2(n17841), .ZN(n13338) );
  NOR2_X1 U16623 ( .A1(n18153), .A2(n18159), .ZN(n18126) );
  XOR2_X1 U16624 ( .A(n17364), .B(n15507), .Z(n15535) );
  XNOR2_X1 U16625 ( .A(n18127), .B(n15535), .ZN(n13336) );
  XNOR2_X1 U16626 ( .A(n13330), .B(n17370), .ZN(n13333) );
  NAND2_X1 U16627 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13333), .ZN(
        n13334) );
  INV_X1 U16628 ( .A(n17871), .ZN(n17862) );
  AOI21_X1 U16629 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17376), .A(
        n17862), .ZN(n13332) );
  NOR2_X1 U16630 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17376), .ZN(
        n13331) );
  AOI221_X1 U16631 ( .B1(n17862), .B2(n17376), .C1(n13332), .C2(n18828), .A(
        n13331), .ZN(n17855) );
  XOR2_X1 U16632 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13333), .Z(
        n17854) );
  NAND2_X1 U16633 ( .A1(n17855), .A2(n17854), .ZN(n17853) );
  NAND2_X1 U16634 ( .A1(n13334), .A2(n17853), .ZN(n13335) );
  NAND2_X1 U16635 ( .A1(n13336), .A2(n13335), .ZN(n15536) );
  OAI21_X1 U16636 ( .B1(n13336), .B2(n13335), .A(n15536), .ZN(n17842) );
  OAI22_X1 U16637 ( .A1(n18127), .A2(n18133), .B1(n18175), .B2(n17842), .ZN(
        n13337) );
  OR4_X1 U16638 ( .A1(n17844), .A2(n13339), .A3(n13338), .A4(n13337), .ZN(
        P3_U2859) );
  AOI211_X1 U16639 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16643), .A(n16634), .B(
        n16911), .ZN(n13347) );
  OAI21_X1 U16640 ( .B1(n16894), .B2(n16631), .A(n16912), .ZN(n16638) );
  AOI221_X1 U16641 ( .B1(n13340), .B2(n18774), .C1(n16902), .C2(n18774), .A(
        n16638), .ZN(n13346) );
  AOI211_X1 U16642 ( .C1(n13343), .C2(n13342), .A(n13341), .B(n18704), .ZN(
        n13345) );
  INV_X1 U16643 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16975) );
  OAI22_X1 U16644 ( .A1(n9872), .A2(n16891), .B1(n16975), .B2(n16910), .ZN(
        n13344) );
  OR4_X1 U16645 ( .A1(n13347), .A2(n13346), .A3(n13345), .A4(n13344), .ZN(
        P3_U2648) );
  NOR2_X1 U16646 ( .A1(n9710), .A2(n13348), .ZN(n19066) );
  INV_X1 U16647 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19984) );
  OAI211_X1 U16648 ( .C1(n19066), .C2(n19984), .A(n13349), .B(n18868), .ZN(
        P2_U2814) );
  INV_X1 U16649 ( .A(n18870), .ZN(n19965) );
  OAI21_X1 U16650 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n13350), .A(n19965), 
        .ZN(n13351) );
  OAI21_X1 U16651 ( .B1(n13352), .B2(n19965), .A(n13351), .ZN(P2_U3612) );
  INV_X1 U16652 ( .A(n13353), .ZN(n19087) );
  NOR2_X1 U16653 ( .A1(n19087), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13354) );
  NOR2_X1 U16654 ( .A1(n13355), .A2(n13354), .ZN(n13541) );
  OR2_X1 U16655 ( .A1(n13356), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13357) );
  NAND2_X1 U16656 ( .A1(n13358), .A2(n13357), .ZN(n13530) );
  NAND2_X1 U16657 ( .A1(n15077), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13531) );
  OAI21_X1 U16658 ( .B1(n16219), .B2(n13530), .A(n13531), .ZN(n13359) );
  AOI21_X1 U16659 ( .B1(n19264), .B2(n13541), .A(n13359), .ZN(n13362) );
  OAI21_X1 U16660 ( .B1(n19258), .B2(n13360), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13361) );
  OAI211_X1 U16661 ( .C1(n16214), .C2(n10622), .A(n13362), .B(n13361), .ZN(
        P2_U3014) );
  OR2_X1 U16662 ( .A1(n9710), .A2(n13363), .ZN(n13368) );
  INV_X1 U16663 ( .A(n16344), .ZN(n13364) );
  NAND2_X1 U16664 ( .A1(n13364), .A2(n16341), .ZN(n13435) );
  AND2_X1 U16665 ( .A1(n13435), .A2(n13365), .ZN(n13367) );
  OAI211_X1 U16666 ( .C1(n13368), .C2(n13396), .A(n13367), .B(n13366), .ZN(
        n16359) );
  NAND2_X1 U16667 ( .A1(n16359), .A2(n16367), .ZN(n13370) );
  NOR2_X1 U16668 ( .A1(n15374), .A2(n19973), .ZN(n13977) );
  NAND2_X1 U16669 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13977), .ZN(n16378) );
  INV_X1 U16670 ( .A(n16378), .ZN(n15691) );
  AOI22_X1 U16671 ( .A1(n15691), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n19969), .ZN(n13369) );
  NAND2_X1 U16672 ( .A1(n13370), .A2(n13369), .ZN(n15391) );
  INV_X1 U16673 ( .A(n16350), .ZN(n13371) );
  INV_X1 U16674 ( .A(n14001), .ZN(n19916) );
  NOR4_X1 U16675 ( .A1(n9710), .A2(n13371), .A3(n11196), .A4(n19916), .ZN(
        n13372) );
  NAND2_X1 U16676 ( .A1(n15391), .A2(n13372), .ZN(n13373) );
  OAI21_X1 U16677 ( .B1(n15391), .B2(n16358), .A(n13373), .ZN(P2_U3595) );
  NOR2_X1 U16678 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20698), .ZN(n19987) );
  INV_X1 U16679 ( .A(n13386), .ZN(n13374) );
  NOR2_X1 U16680 ( .A1(n13387), .A2(n13374), .ZN(n13378) );
  NAND2_X1 U16681 ( .A1(n13460), .A2(n13378), .ZN(n19986) );
  OAI21_X1 U16682 ( .B1(n19987), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13847), 
        .ZN(n13377) );
  INV_X1 U16683 ( .A(n13847), .ZN(n20862) );
  OAI21_X1 U16684 ( .B1(n13852), .B2(n13375), .A(n20862), .ZN(n13376) );
  NAND2_X1 U16685 ( .A1(n13377), .A2(n13376), .ZN(P1_U3487) );
  INV_X1 U16686 ( .A(n12785), .ZN(n15639) );
  NOR2_X1 U16687 ( .A1(n13378), .A2(n15639), .ZN(n13379) );
  AOI21_X1 U16688 ( .B1(n15646), .B2(n13644), .A(n13379), .ZN(n19991) );
  NAND3_X1 U16689 ( .A1(n13644), .A2(n12284), .A3(n15674), .ZN(n13381) );
  NAND2_X1 U16690 ( .A1(n13381), .A2(n20864), .ZN(n20865) );
  AND2_X1 U16691 ( .A1(n19991), .A2(n20865), .ZN(n15633) );
  NOR2_X1 U16692 ( .A1(n15633), .A2(n19992), .ZN(n19999) );
  INV_X1 U16693 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13394) );
  INV_X1 U16694 ( .A(n13646), .ZN(n13390) );
  NAND3_X1 U16695 ( .A1(n13382), .A2(n11558), .A3(n13854), .ZN(n13383) );
  NAND2_X1 U16696 ( .A1(n13384), .A2(n13383), .ZN(n13385) );
  NAND2_X1 U16697 ( .A1(n15646), .A2(n13385), .ZN(n13389) );
  OR2_X1 U16698 ( .A1(n13387), .A2(n13386), .ZN(n13388) );
  OAI211_X1 U16699 ( .C1(n15646), .C2(n13390), .A(n13389), .B(n13388), .ZN(
        n13391) );
  NAND2_X1 U16700 ( .A1(n13391), .A2(n11619), .ZN(n15626) );
  INV_X1 U16701 ( .A(n15626), .ZN(n13392) );
  NAND2_X1 U16702 ( .A1(n19999), .A2(n13392), .ZN(n13393) );
  OAI21_X1 U16703 ( .B1(n19999), .B2(n13394), .A(n13393), .ZN(P1_U3484) );
  INV_X1 U16704 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19177) );
  INV_X1 U16705 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n19176) );
  AOI22_X1 U16706 ( .A1(n16121), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16122), .ZN(n19114) );
  OAI222_X1 U16707 ( .A1(n13449), .A2(n19177), .B1(n13444), .B2(n19176), .C1(
        n19254), .C2(n19114), .ZN(P2_U2982) );
  INV_X1 U16708 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13401) );
  INV_X1 U16709 ( .A(n16367), .ZN(n18873) );
  OR2_X1 U16710 ( .A1(n9710), .A2(n18873), .ZN(n13395) );
  OAI21_X1 U16711 ( .B1(n13396), .B2(n13395), .A(n13449), .ZN(n13397) );
  NAND2_X1 U16712 ( .A1(n19203), .A2(n13398), .ZN(n19168) );
  NAND2_X1 U16713 ( .A1(n13977), .A2(n19969), .ZN(n19966) );
  INV_X1 U16714 ( .A(n19966), .ZN(n13399) );
  CLKBUF_X1 U16715 ( .A(n13399), .Z(n19212) );
  AOI22_X1 U16716 ( .A1(n19212), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13400) );
  OAI21_X1 U16717 ( .B1(n13401), .B2(n19168), .A(n13400), .ZN(P2_U2932) );
  INV_X1 U16718 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U16719 ( .A1(n19212), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13402) );
  OAI21_X1 U16720 ( .B1(n13403), .B2(n19168), .A(n13402), .ZN(P2_U2934) );
  INV_X1 U16721 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13405) );
  AOI22_X1 U16722 ( .A1(n19212), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13404) );
  OAI21_X1 U16723 ( .B1(n13405), .B2(n19168), .A(n13404), .ZN(P2_U2929) );
  INV_X1 U16724 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U16725 ( .A1(n19212), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13406) );
  OAI21_X1 U16726 ( .B1(n13407), .B2(n19168), .A(n13406), .ZN(P2_U2935) );
  INV_X1 U16727 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U16728 ( .A1(n19212), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13408) );
  OAI21_X1 U16729 ( .B1(n14972), .B2(n19168), .A(n13408), .ZN(P2_U2924) );
  AOI22_X1 U16730 ( .A1(n19212), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13409) );
  OAI21_X1 U16731 ( .B1(n13446), .B2(n19168), .A(n13409), .ZN(P2_U2927) );
  INV_X1 U16732 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U16733 ( .A1(n19212), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13410) );
  OAI21_X1 U16734 ( .B1(n13411), .B2(n19168), .A(n13410), .ZN(P2_U2922) );
  INV_X1 U16735 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14989) );
  AOI22_X1 U16736 ( .A1(n19212), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13412) );
  OAI21_X1 U16737 ( .B1(n14989), .B2(n19168), .A(n13412), .ZN(P2_U2926) );
  INV_X1 U16738 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13414) );
  AOI22_X1 U16739 ( .A1(n19212), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13413) );
  OAI21_X1 U16740 ( .B1(n13414), .B2(n19168), .A(n13413), .ZN(P2_U2931) );
  INV_X1 U16741 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13416) );
  INV_X1 U16742 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13415) );
  OAI222_X1 U16743 ( .A1(n19168), .A2(n13416), .B1(n19205), .B2(n16530), .C1(
        n13415), .C2(n19966), .ZN(P2_U2930) );
  INV_X1 U16744 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13418) );
  INV_X1 U16745 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13417) );
  OAI222_X1 U16746 ( .A1(n19168), .A2(n13418), .B1(n19205), .B2(n16532), .C1(
        n13417), .C2(n19966), .ZN(P2_U2928) );
  INV_X1 U16747 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14960) );
  INV_X1 U16748 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n13419) );
  OAI222_X1 U16749 ( .A1(n19168), .A2(n14960), .B1(n19966), .B2(n13419), .C1(
        n19205), .C2(n16537), .ZN(P2_U2923) );
  AOI21_X1 U16750 ( .B1(n13422), .B2(n13421), .A(n13420), .ZN(n13576) );
  NAND2_X1 U16751 ( .A1(n13424), .A2(n13423), .ZN(n13567) );
  AND3_X1 U16752 ( .A1(n13566), .A2(n19264), .A3(n13567), .ZN(n13427) );
  AND2_X1 U16753 ( .A1(n15077), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13569) );
  AOI21_X1 U16754 ( .B1(n19258), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13569), .ZN(n13425) );
  OAI21_X1 U16755 ( .B1(n19269), .B2(n13831), .A(n13425), .ZN(n13426) );
  AOI211_X1 U16756 ( .C1(n13576), .C2(n19260), .A(n13427), .B(n13426), .ZN(
        n13428) );
  OAI21_X1 U16757 ( .B1(n9853), .B2(n16214), .A(n13428), .ZN(P2_U3012) );
  NOR2_X1 U16758 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13430) );
  OAI21_X1 U16759 ( .B1(n13431), .B2(n13430), .A(n13429), .ZN(n13432) );
  INV_X1 U16760 ( .A(n13432), .ZN(n13433) );
  NAND2_X1 U16761 ( .A1(n13435), .A2(n13434), .ZN(n13436) );
  NAND2_X1 U16762 ( .A1(n14936), .A2(n10547), .ZN(n14926) );
  MUX2_X1 U16763 ( .A(n10622), .B(n19090), .S(n14907), .Z(n13437) );
  OAI21_X1 U16764 ( .B1(n19945), .B2(n14926), .A(n13437), .ZN(P2_U2887) );
  OR2_X2 U16765 ( .A1(n19988), .A2(n13860), .ZN(n13617) );
  INV_X1 U16766 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14216) );
  AND2_X1 U16767 ( .A1(n11631), .A2(n15671), .ZN(n13438) );
  NAND2_X1 U16768 ( .A1(n20151), .A2(n13860), .ZN(n13475) );
  INV_X1 U16769 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13439) );
  NOR2_X1 U16770 ( .A1(n20190), .A2(n13439), .ZN(n13440) );
  AOI21_X1 U16771 ( .B1(DATAI_15_), .B2(n20190), .A(n13440), .ZN(n14217) );
  OAI222_X1 U16772 ( .A1(n13617), .A2(n14216), .B1(n13475), .B2(n14217), .C1(
        n20151), .C2(n20113), .ZN(P1_U2967) );
  INV_X1 U16773 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20117) );
  MUX2_X1 U16774 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20189), .Z(
        n14401) );
  INV_X1 U16775 ( .A(n14401), .ZN(n13441) );
  NOR2_X1 U16776 ( .A1(n13475), .A2(n13441), .ZN(n20148) );
  INV_X1 U16777 ( .A(n20148), .ZN(n13443) );
  NAND2_X1 U16778 ( .A1(n20152), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n13442) );
  OAI211_X1 U16779 ( .C1(n20117), .C2(n13617), .A(n13443), .B(n13442), .ZN(
        P1_U2965) );
  INV_X2 U16780 ( .A(n13444), .ZN(n19246) );
  NAND2_X1 U16781 ( .A1(n19246), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13445) );
  MUX2_X1 U16782 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n16122), .Z(n19128) );
  NAND2_X1 U16783 ( .A1(n19231), .A2(n19128), .ZN(n13447) );
  OAI211_X1 U16784 ( .C1(n13446), .C2(n13449), .A(n13445), .B(n13447), .ZN(
        P2_U2960) );
  INV_X1 U16785 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19194) );
  NAND2_X1 U16786 ( .A1(n19246), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13448) );
  OAI211_X1 U16787 ( .C1(n19194), .C2(n13449), .A(n13448), .B(n13447), .ZN(
        P2_U2975) );
  INV_X1 U16788 ( .A(n15644), .ZN(n13450) );
  AND2_X1 U16789 ( .A1(n15638), .A2(n13450), .ZN(n13453) );
  NAND3_X1 U16790 ( .A1(n13451), .A2(n13464), .A3(n13666), .ZN(n13452) );
  OAI21_X1 U16791 ( .B1(n13454), .B2(n13453), .A(n13452), .ZN(n13459) );
  NOR2_X1 U16792 ( .A1(n13857), .A2(n11581), .ZN(n13455) );
  OR2_X1 U16793 ( .A1(n13456), .A2(n13455), .ZN(n13457) );
  AOI21_X1 U16794 ( .B1(n15646), .B2(n13646), .A(n13457), .ZN(n13458) );
  NAND2_X1 U16795 ( .A1(n13459), .A2(n13458), .ZN(n15614) );
  NAND2_X1 U16796 ( .A1(n15614), .A2(n13460), .ZN(n13462) );
  NAND2_X1 U16797 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16021) );
  NOR2_X1 U16798 ( .A1(n20761), .A2(n16021), .ZN(n13681) );
  NAND2_X1 U16799 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13681), .ZN(n13461) );
  NAND2_X1 U16800 ( .A1(n13462), .A2(n13461), .ZN(n16007) );
  AND2_X1 U16801 ( .A1(n20761), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13463) );
  OR2_X1 U16802 ( .A1(n16007), .A2(n13463), .ZN(n16011) );
  INV_X1 U16803 ( .A(n16011), .ZN(n13472) );
  AOI21_X1 U16804 ( .B1(n15612), .B2(n16008), .A(n13472), .ZN(n13474) );
  INV_X1 U16805 ( .A(n11833), .ZN(n13871) );
  OR2_X1 U16806 ( .A1(n13465), .A2(n11580), .ZN(n13466) );
  NOR2_X1 U16807 ( .A1(n13467), .A2(n13466), .ZN(n13469) );
  OAI21_X1 U16808 ( .B1(n12723), .B2(n11608), .A(n13852), .ZN(n13468) );
  AND2_X1 U16809 ( .A1(n13469), .A2(n13468), .ZN(n14833) );
  OAI22_X1 U16810 ( .A1(n13871), .A2(n14833), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14829), .ZN(n15611) );
  INV_X1 U16811 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20593) );
  OAI22_X1 U16812 ( .A1(n20760), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14848), .ZN(n13470) );
  AOI21_X1 U16813 ( .B1(n15611), .B2(n16008), .A(n13470), .ZN(n13471) );
  OAI22_X1 U16814 ( .A1(n13474), .A2(n13473), .B1(n13472), .B2(n13471), .ZN(
        P1_U3474) );
  INV_X1 U16815 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13625) );
  MUX2_X1 U16816 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20189), .Z(
        n14623) );
  NAND2_X1 U16817 ( .A1(n13524), .A2(n14623), .ZN(n20154) );
  NAND2_X1 U16818 ( .A1(n20152), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13476) );
  OAI211_X1 U16819 ( .C1(n13625), .C2(n13617), .A(n20154), .B(n13476), .ZN(
        P1_U2948) );
  NAND2_X1 U16820 ( .A1(n20190), .A2(DATAI_2_), .ZN(n13478) );
  NAND2_X1 U16821 ( .A1(n20189), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13477) );
  AND2_X1 U16822 ( .A1(n13478), .A2(n13477), .ZN(n20214) );
  INV_X1 U16823 ( .A(n20214), .ZN(n13479) );
  NAND2_X1 U16824 ( .A1(n13524), .A2(n13479), .ZN(n13484) );
  INV_X1 U16825 ( .A(n13617), .ZN(n20153) );
  AOI22_X1 U16826 ( .A1(n20153), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20152), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13480) );
  NAND2_X1 U16827 ( .A1(n13484), .A2(n13480), .ZN(P1_U2939) );
  MUX2_X1 U16828 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20189), .Z(
        n14629) );
  NAND2_X1 U16829 ( .A1(n13524), .A2(n14629), .ZN(n13486) );
  AOI22_X1 U16830 ( .A1(n20153), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20152), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13481) );
  NAND2_X1 U16831 ( .A1(n13486), .A2(n13481), .ZN(P1_U2947) );
  MUX2_X1 U16832 ( .A(DATAI_0_), .B(BUF1_REG_0__SCAN_IN), .S(n20189), .Z(
        n20203) );
  NAND2_X1 U16833 ( .A1(n13524), .A2(n20203), .ZN(n13488) );
  AOI22_X1 U16834 ( .A1(n20153), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20152), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13482) );
  NAND2_X1 U16835 ( .A1(n13488), .A2(n13482), .ZN(P1_U2937) );
  INV_X1 U16836 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20141) );
  NAND2_X1 U16837 ( .A1(n20152), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n13483) );
  OAI211_X1 U16838 ( .C1(n20141), .C2(n13617), .A(n13484), .B(n13483), .ZN(
        P1_U2954) );
  INV_X1 U16839 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20124) );
  NAND2_X1 U16840 ( .A1(n20152), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n13485) );
  OAI211_X1 U16841 ( .C1(n20124), .C2(n13617), .A(n13486), .B(n13485), .ZN(
        P1_U2962) );
  INV_X1 U16842 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20147) );
  NAND2_X1 U16843 ( .A1(n20152), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n13487) );
  OAI211_X1 U16844 ( .C1(n20147), .C2(n13617), .A(n13488), .B(n13487), .ZN(
        P1_U2952) );
  INV_X1 U16845 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20137) );
  NAND2_X1 U16846 ( .A1(n20190), .A2(DATAI_4_), .ZN(n13490) );
  NAND2_X1 U16847 ( .A1(n20189), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13489) );
  AND2_X1 U16848 ( .A1(n13490), .A2(n13489), .ZN(n20222) );
  INV_X1 U16849 ( .A(n20222), .ZN(n13491) );
  NAND2_X1 U16850 ( .A1(n13524), .A2(n13491), .ZN(n13501) );
  NAND2_X1 U16851 ( .A1(n20152), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n13492) );
  OAI211_X1 U16852 ( .C1(n20137), .C2(n13617), .A(n13501), .B(n13492), .ZN(
        P1_U2956) );
  NAND2_X1 U16853 ( .A1(n20190), .A2(DATAI_5_), .ZN(n13494) );
  NAND2_X1 U16854 ( .A1(n20189), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13493) );
  AND2_X1 U16855 ( .A1(n13494), .A2(n13493), .ZN(n20225) );
  INV_X1 U16856 ( .A(n20225), .ZN(n14647) );
  NAND2_X1 U16857 ( .A1(n13524), .A2(n14647), .ZN(n13503) );
  NAND2_X1 U16858 ( .A1(n20152), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n13495) );
  OAI211_X1 U16859 ( .C1(n11786), .C2(n13617), .A(n13503), .B(n13495), .ZN(
        P1_U2957) );
  NAND2_X1 U16860 ( .A1(n20190), .A2(DATAI_6_), .ZN(n13497) );
  NAND2_X1 U16861 ( .A1(n20189), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13496) );
  AND2_X1 U16862 ( .A1(n13497), .A2(n13496), .ZN(n20229) );
  INV_X1 U16863 ( .A(n20229), .ZN(n13498) );
  NAND2_X1 U16864 ( .A1(n13524), .A2(n13498), .ZN(n13505) );
  NAND2_X1 U16865 ( .A1(n20152), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13499) );
  OAI211_X1 U16866 ( .C1(n14642), .C2(n13617), .A(n13505), .B(n13499), .ZN(
        P1_U2943) );
  NAND2_X1 U16867 ( .A1(n20152), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13500) );
  OAI211_X1 U16868 ( .C1(n14651), .C2(n13617), .A(n13501), .B(n13500), .ZN(
        P1_U2941) );
  INV_X1 U16869 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13633) );
  NAND2_X1 U16870 ( .A1(n20152), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13502) );
  OAI211_X1 U16871 ( .C1(n13633), .C2(n13617), .A(n13503), .B(n13502), .ZN(
        P1_U2942) );
  NAND2_X1 U16872 ( .A1(n20152), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n13504) );
  OAI211_X1 U16873 ( .C1(n11862), .C2(n13617), .A(n13505), .B(n13504), .ZN(
        P1_U2958) );
  INV_X1 U16874 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13629) );
  INV_X1 U16875 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n14957) );
  NOR2_X1 U16876 ( .A1(n20190), .A2(n14957), .ZN(n13506) );
  AOI21_X1 U16877 ( .B1(DATAI_12_), .B2(n20190), .A(n13506), .ZN(n14618) );
  INV_X1 U16878 ( .A(n14618), .ZN(n13507) );
  NAND2_X1 U16879 ( .A1(n13524), .A2(n13507), .ZN(n13512) );
  NAND2_X1 U16880 ( .A1(n20152), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13508) );
  OAI211_X1 U16881 ( .C1(n13629), .C2(n13617), .A(n13512), .B(n13508), .ZN(
        P1_U2949) );
  INV_X1 U16882 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20126) );
  MUX2_X1 U16883 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20189), .Z(
        n14632) );
  NAND2_X1 U16884 ( .A1(n13524), .A2(n14632), .ZN(n13519) );
  NAND2_X1 U16885 ( .A1(n20152), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n13509) );
  OAI211_X1 U16886 ( .C1(n20126), .C2(n13617), .A(n13519), .B(n13509), .ZN(
        P1_U2961) );
  INV_X1 U16887 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13636) );
  MUX2_X1 U16888 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20189), .Z(
        n14636) );
  NAND2_X1 U16889 ( .A1(n13524), .A2(n14636), .ZN(n13514) );
  NAND2_X1 U16890 ( .A1(n20152), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13510) );
  OAI211_X1 U16891 ( .C1(n13636), .C2(n13617), .A(n13514), .B(n13510), .ZN(
        P1_U2945) );
  INV_X1 U16892 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20119) );
  NAND2_X1 U16893 ( .A1(n20152), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n13511) );
  OAI211_X1 U16894 ( .C1(n20119), .C2(n13617), .A(n13512), .B(n13511), .ZN(
        P1_U2964) );
  INV_X1 U16895 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20128) );
  NAND2_X1 U16896 ( .A1(n20152), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13513) );
  OAI211_X1 U16897 ( .C1(n20128), .C2(n13617), .A(n13514), .B(n13513), .ZN(
        P1_U2960) );
  INV_X1 U16898 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13620) );
  MUX2_X1 U16899 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20189), .Z(
        n14613) );
  NAND2_X1 U16900 ( .A1(n13524), .A2(n14613), .ZN(n13517) );
  NAND2_X1 U16901 ( .A1(n20152), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13515) );
  OAI211_X1 U16902 ( .C1(n13620), .C2(n13617), .A(n13517), .B(n13515), .ZN(
        P1_U2951) );
  INV_X1 U16903 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20115) );
  NAND2_X1 U16904 ( .A1(n20152), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n13516) );
  OAI211_X1 U16905 ( .C1(n20115), .C2(n13617), .A(n13517), .B(n13516), .ZN(
        P1_U2966) );
  INV_X1 U16906 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13627) );
  NAND2_X1 U16907 ( .A1(n20152), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13518) );
  OAI211_X1 U16908 ( .C1(n13627), .C2(n13617), .A(n13519), .B(n13518), .ZN(
        P1_U2946) );
  INV_X1 U16909 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20143) );
  MUX2_X1 U16910 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n20189), .Z(
        n20210) );
  NAND2_X1 U16911 ( .A1(n13524), .A2(n20210), .ZN(n13523) );
  NAND2_X1 U16912 ( .A1(n20152), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n13520) );
  OAI211_X1 U16913 ( .C1(n20143), .C2(n13617), .A(n13523), .B(n13520), .ZN(
        P1_U2953) );
  INV_X1 U16914 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20139) );
  MUX2_X1 U16915 ( .A(DATAI_3_), .B(BUF1_REG_3__SCAN_IN), .S(n20189), .Z(
        n20218) );
  NAND2_X1 U16916 ( .A1(n13524), .A2(n20218), .ZN(n13527) );
  NAND2_X1 U16917 ( .A1(n20152), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n13521) );
  OAI211_X1 U16918 ( .C1(n20139), .C2(n13617), .A(n13527), .B(n13521), .ZN(
        P1_U2955) );
  INV_X1 U16919 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U16920 ( .A1(n20152), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13522) );
  OAI211_X1 U16921 ( .C1(n13623), .C2(n13617), .A(n13523), .B(n13522), .ZN(
        P1_U2938) );
  INV_X1 U16922 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13638) );
  MUX2_X1 U16923 ( .A(DATAI_7_), .B(BUF1_REG_7__SCAN_IN), .S(n20189), .Z(
        n20237) );
  NAND2_X1 U16924 ( .A1(n13524), .A2(n20237), .ZN(n13529) );
  NAND2_X1 U16925 ( .A1(n20152), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13525) );
  OAI211_X1 U16926 ( .C1(n13638), .C2(n13617), .A(n13529), .B(n13525), .ZN(
        P1_U2944) );
  INV_X1 U16927 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13631) );
  NAND2_X1 U16928 ( .A1(n20152), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13526) );
  OAI211_X1 U16929 ( .C1(n13631), .C2(n13617), .A(n13527), .B(n13526), .ZN(
        P1_U2940) );
  INV_X1 U16930 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20130) );
  NAND2_X1 U16931 ( .A1(n20152), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n13528) );
  OAI211_X1 U16932 ( .C1(n20130), .C2(n13617), .A(n13529), .B(n13528), .ZN(
        P1_U2959) );
  NOR2_X1 U16933 ( .A1(n16307), .A2(n13530), .ZN(n13533) );
  OAI21_X1 U16934 ( .B1(n14380), .B2(n10835), .A(n13531), .ZN(n13532) );
  AOI211_X1 U16935 ( .C1(n12589), .C2(n19094), .A(n13533), .B(n13532), .ZN(
        n13543) );
  INV_X1 U16936 ( .A(n13534), .ZN(n13539) );
  INV_X1 U16937 ( .A(n13535), .ZN(n13536) );
  NAND2_X1 U16938 ( .A1(n13537), .A2(n13536), .ZN(n13538) );
  NAND2_X1 U16939 ( .A1(n13539), .A2(n13538), .ZN(n19084) );
  INV_X1 U16940 ( .A(n19084), .ZN(n13540) );
  AOI22_X1 U16941 ( .A1(n16301), .A2(n13541), .B1(n16281), .B2(n13540), .ZN(
        n13542) );
  OAI211_X1 U16942 ( .C1(n15253), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13543), .B(n13542), .ZN(P2_U3046) );
  AOI21_X1 U16943 ( .B1(n9817), .B2(n20172), .A(n12618), .ZN(n20168) );
  NAND2_X1 U16944 ( .A1(n15916), .A2(n15914), .ZN(n13545) );
  AND2_X1 U16945 ( .A1(n13545), .A2(n20172), .ZN(n13591) );
  OR2_X1 U16946 ( .A1(n13546), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13548) );
  NAND2_X1 U16947 ( .A1(n13548), .A2(n13547), .ZN(n13866) );
  OAI21_X1 U16948 ( .B1(n15928), .B2(n15919), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13550) );
  INV_X1 U16949 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13549) );
  OR2_X1 U16950 ( .A1(n20177), .A2(n13549), .ZN(n20169) );
  OAI211_X1 U16951 ( .C1(n20179), .C2(n13866), .A(n13550), .B(n20169), .ZN(
        n13551) );
  AOI211_X1 U16952 ( .C1(n20168), .C2(n20182), .A(n13591), .B(n13551), .ZN(
        n13552) );
  INV_X1 U16953 ( .A(n13552), .ZN(P1_U3031) );
  INV_X1 U16954 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16512) );
  INV_X1 U16955 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18186) );
  AOI22_X1 U16956 ( .A1(n16121), .A2(n16512), .B1(n18186), .B2(n16122), .ZN(
        n19104) );
  NAND2_X1 U16957 ( .A1(n14999), .A2(n13553), .ZN(n19134) );
  OAI22_X1 U16958 ( .A1(n16124), .A2(n19084), .B1(n19132), .B2(n13554), .ZN(
        n13556) );
  NOR2_X1 U16959 ( .A1(n19945), .A2(n19084), .ZN(n19161) );
  AOI211_X1 U16960 ( .C1(n19945), .C2(n19084), .A(n19162), .B(n19161), .ZN(
        n13555) );
  AOI211_X1 U16961 ( .C1(n19104), .C2(n19134), .A(n13556), .B(n13555), .ZN(
        n13557) );
  INV_X1 U16962 ( .A(n13557), .ZN(P2_U2919) );
  INV_X1 U16963 ( .A(n13558), .ZN(n13561) );
  OAI21_X1 U16964 ( .B1(n13561), .B2(n13560), .A(n13559), .ZN(n20171) );
  OAI222_X1 U16965 ( .A1(n13866), .A2(n14612), .B1(n14611), .B2(n13562), .C1(
        n20171), .C2(n14595), .ZN(P1_U2872) );
  AOI21_X1 U16966 ( .B1(n13565), .B2(n13564), .A(n13563), .ZN(n19137) );
  INV_X1 U16967 ( .A(n19137), .ZN(n19931) );
  NAND3_X1 U16968 ( .A1(n16301), .A2(n13567), .A3(n13566), .ZN(n13571) );
  NOR2_X1 U16969 ( .A1(n13569), .A2(n13568), .ZN(n13570) );
  OAI211_X1 U16970 ( .C1(n14380), .C2(n13572), .A(n13571), .B(n13570), .ZN(
        n13581) );
  INV_X1 U16971 ( .A(n13573), .ZN(n13578) );
  AOI22_X1 U16972 ( .A1(n13576), .A2(n16274), .B1(n13575), .B2(n13574), .ZN(
        n13577) );
  OAI21_X1 U16973 ( .B1(n13579), .B2(n13578), .A(n13577), .ZN(n13580) );
  AOI211_X1 U16974 ( .C1(n19931), .C2(n16281), .A(n13581), .B(n13580), .ZN(
        n13582) );
  OAI21_X1 U16975 ( .B1(n9853), .B2(n16283), .A(n13582), .ZN(P2_U3044) );
  MUX2_X1 U16976 ( .A(n14399), .B(n13585), .S(n14907), .Z(n13586) );
  OAI21_X1 U16977 ( .B1(n19937), .B2(n14926), .A(n13586), .ZN(P2_U2886) );
  XNOR2_X1 U16978 ( .A(n13588), .B(n13589), .ZN(n20156) );
  XNOR2_X1 U16979 ( .A(n13590), .B(n13380), .ZN(n13605) );
  OAI21_X1 U16980 ( .B1(n15919), .B2(n13591), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13593) );
  INV_X1 U16981 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20852) );
  NOR2_X1 U16982 ( .A1(n20177), .A2(n20852), .ZN(n20161) );
  INV_X1 U16983 ( .A(n20161), .ZN(n13592) );
  OAI211_X1 U16984 ( .C1(n20179), .C2(n13605), .A(n13593), .B(n13592), .ZN(
        n13596) );
  NOR3_X1 U16985 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13892), .A3(
        n13594), .ZN(n13595) );
  AOI211_X1 U16986 ( .C1(n20182), .C2(n20156), .A(n13596), .B(n13595), .ZN(
        n13597) );
  INV_X1 U16987 ( .A(n13597), .ZN(P1_U3030) );
  NAND2_X1 U16988 ( .A1(n10640), .A2(n14936), .ZN(n13602) );
  NAND2_X1 U16989 ( .A1(n14884), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13601) );
  OAI211_X1 U16990 ( .C1(n19323), .C2(n14926), .A(n13602), .B(n13601), .ZN(
        P2_U2884) );
  OAI21_X1 U16991 ( .B1(n13604), .B2(n13603), .A(n13608), .ZN(n20163) );
  OAI22_X1 U16992 ( .A1(n14612), .A2(n13605), .B1(n13935), .B2(n14611), .ZN(
        n13606) );
  INV_X1 U16993 ( .A(n13606), .ZN(n13607) );
  OAI21_X1 U16994 ( .B1(n20163), .B2(n14595), .A(n13607), .ZN(P1_U2871) );
  OAI21_X1 U16995 ( .B1(n10075), .B2(n11840), .A(n13609), .ZN(n13933) );
  INV_X1 U16996 ( .A(n13933), .ZN(n13694) );
  NAND2_X1 U16997 ( .A1(n13611), .A2(n13610), .ZN(n13612) );
  NAND2_X1 U16998 ( .A1(n13755), .A2(n13612), .ZN(n20178) );
  OAI22_X1 U16999 ( .A1(n14612), .A2(n20178), .B1(n13613), .B2(n14611), .ZN(
        n13614) );
  AOI21_X1 U17000 ( .B1(n13694), .B2(n13760), .A(n13614), .ZN(n13615) );
  INV_X1 U17001 ( .A(n13615), .ZN(P1_U2870) );
  OR3_X1 U17002 ( .A1(n15646), .A2(n19992), .A3(n13666), .ZN(n13616) );
  NAND2_X1 U17003 ( .A1(n13617), .A2(n13616), .ZN(n13618) );
  NAND2_X1 U17004 ( .A1(n20120), .A2(n13854), .ZN(n20109) );
  OR2_X1 U17005 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16021), .ZN(n20133) );
  NOR2_X4 U17006 ( .A1(n20120), .A2(n9726), .ZN(n20144) );
  AOI22_X1 U17007 ( .A1(n9726), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13619) );
  OAI21_X1 U17008 ( .B1(n13620), .B2(n20109), .A(n13619), .ZN(P1_U2906) );
  INV_X1 U17009 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14659) );
  AOI22_X1 U17010 ( .A1(n9726), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13621) );
  OAI21_X1 U17011 ( .B1(n14659), .B2(n20109), .A(n13621), .ZN(P1_U2918) );
  AOI22_X1 U17012 ( .A1(n9726), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13622) );
  OAI21_X1 U17013 ( .B1(n13623), .B2(n20109), .A(n13622), .ZN(P1_U2919) );
  AOI22_X1 U17014 ( .A1(n9726), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13624) );
  OAI21_X1 U17015 ( .B1(n13625), .B2(n20109), .A(n13624), .ZN(P1_U2909) );
  AOI22_X1 U17016 ( .A1(n9726), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13626) );
  OAI21_X1 U17017 ( .B1(n13627), .B2(n20109), .A(n13626), .ZN(P1_U2911) );
  AOI22_X1 U17018 ( .A1(n9726), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13628) );
  OAI21_X1 U17019 ( .B1(n13629), .B2(n20109), .A(n13628), .ZN(P1_U2908) );
  AOI22_X1 U17020 ( .A1(n9726), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13630) );
  OAI21_X1 U17021 ( .B1(n13631), .B2(n20109), .A(n13630), .ZN(P1_U2917) );
  AOI22_X1 U17022 ( .A1(n9726), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13632) );
  OAI21_X1 U17023 ( .B1(n13633), .B2(n20109), .A(n13632), .ZN(P1_U2915) );
  AOI22_X1 U17024 ( .A1(n9726), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13634) );
  OAI21_X1 U17025 ( .B1(n14642), .B2(n20109), .A(n13634), .ZN(P1_U2914) );
  AOI22_X1 U17026 ( .A1(n9726), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13635) );
  OAI21_X1 U17027 ( .B1(n13636), .B2(n20109), .A(n13635), .ZN(P1_U2912) );
  AOI22_X1 U17028 ( .A1(n9726), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13637) );
  OAI21_X1 U17029 ( .B1(n13638), .B2(n20109), .A(n13637), .ZN(P1_U2913) );
  AOI22_X1 U17030 ( .A1(n9726), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13639) );
  OAI21_X1 U17031 ( .B1(n14651), .B2(n20109), .A(n13639), .ZN(P1_U2916) );
  INV_X1 U17032 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14671) );
  AOI22_X1 U17033 ( .A1(n9726), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13640) );
  OAI21_X1 U17034 ( .B1(n14671), .B2(n20109), .A(n13640), .ZN(P1_U2920) );
  INV_X1 U17035 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14627) );
  AOI22_X1 U17036 ( .A1(n9726), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13641) );
  OAI21_X1 U17037 ( .B1(n14627), .B2(n20109), .A(n13641), .ZN(P1_U2910) );
  INV_X1 U17038 ( .A(n13643), .ZN(n20199) );
  INV_X1 U17039 ( .A(n14833), .ZN(n13668) );
  XNOR2_X1 U17040 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13651) );
  NOR2_X1 U17041 ( .A1(n15628), .A2(n13644), .ZN(n13645) );
  OR2_X1 U17042 ( .A1(n13646), .A2(n13645), .ZN(n13659) );
  XNOR2_X1 U17043 ( .A(n14834), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13648) );
  NAND2_X1 U17044 ( .A1(n13659), .A2(n13648), .ZN(n13650) );
  INV_X1 U17045 ( .A(n13648), .ZN(n14841) );
  NAND3_X1 U17046 ( .A1(n14833), .A2(n13662), .A3(n14841), .ZN(n13649) );
  OAI211_X1 U17047 ( .C1(n13666), .C2(n13651), .A(n13650), .B(n13649), .ZN(
        n13652) );
  AOI21_X1 U17048 ( .B1(n20199), .B2(n13668), .A(n13652), .ZN(n14845) );
  MUX2_X1 U17049 ( .A(n11816), .B(n14845), .S(n15614), .Z(n15621) );
  NAND2_X1 U17050 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n19998), .ZN(n13670) );
  OAI22_X1 U17051 ( .A1(n15621), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n13670), 
        .B2(n11816), .ZN(n13672) );
  XNOR2_X1 U17052 ( .A(n13654), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13665) );
  MUX2_X1 U17053 ( .A(n13655), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14834), .Z(n13657) );
  NOR2_X1 U17054 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  NAND2_X1 U17055 ( .A1(n13659), .A2(n13658), .ZN(n13664) );
  NAND2_X1 U17056 ( .A1(n14834), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13660) );
  NAND2_X1 U17057 ( .A1(n13660), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13661) );
  NAND2_X1 U17058 ( .A1(n11659), .A2(n13661), .ZN(n14847) );
  NAND3_X1 U17059 ( .A1(n14833), .A2(n13662), .A3(n14847), .ZN(n13663) );
  OAI211_X1 U17060 ( .C1(n13666), .C2(n13665), .A(n13664), .B(n13663), .ZN(
        n13667) );
  AOI21_X1 U17061 ( .B1(n13653), .B2(n13668), .A(n13667), .ZN(n14851) );
  MUX2_X1 U17062 ( .A(n13669), .B(n14851), .S(n15614), .Z(n15625) );
  NAND2_X1 U17063 ( .A1(n15625), .A2(n13670), .ZN(n13671) );
  OAI211_X1 U17064 ( .C1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n20760), .A(
        n13672), .B(n13671), .ZN(n15634) );
  NOR2_X1 U17065 ( .A1(n13674), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13679) );
  INV_X1 U17066 ( .A(n20336), .ZN(n20584) );
  NOR2_X1 U17067 ( .A1(n13675), .A2(n20584), .ZN(n13676) );
  XNOR2_X1 U17068 ( .A(n13676), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20076) );
  OR2_X1 U17069 ( .A1(n20076), .A2(n13677), .ZN(n16006) );
  NAND2_X1 U17070 ( .A1(n16006), .A2(n15614), .ZN(n13678) );
  MUX2_X1 U17071 ( .A(n13679), .B(n13678), .S(n20760), .Z(n13680) );
  OAI21_X1 U17072 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15614), .A(
        n13680), .ZN(n15629) );
  OAI21_X1 U17073 ( .B1(n15634), .B2(n13673), .A(n15629), .ZN(n13696) );
  OAI21_X1 U17074 ( .B1(n13696), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13681), .ZN(
        n13682) );
  NOR2_X1 U17075 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20867) );
  INV_X1 U17076 ( .A(n16021), .ZN(n16019) );
  NAND2_X1 U17077 ( .A1(n13682), .A2(n20342), .ZN(n20187) );
  NOR2_X1 U17078 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20760), .ZN(n14823) );
  OR2_X1 U17079 ( .A1(n9717), .A2(n20698), .ZN(n13684) );
  NAND2_X1 U17080 ( .A1(n20636), .A2(n20633), .ZN(n20582) );
  NAND2_X1 U17081 ( .A1(n13684), .A2(n20582), .ZN(n20556) );
  INV_X1 U17082 ( .A(n20556), .ZN(n13686) );
  AND2_X1 U17083 ( .A1(n20636), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13685) );
  NAND2_X1 U17084 ( .A1(n9717), .A2(n13685), .ZN(n20703) );
  MUX2_X1 U17085 ( .A(n13686), .B(n20703), .S(n20192), .Z(n13687) );
  OAI21_X1 U17086 ( .B1(n14823), .B2(n13643), .A(n13687), .ZN(n13688) );
  NAND2_X1 U17087 ( .A1(n20187), .A2(n13688), .ZN(n13689) );
  OAI21_X1 U17088 ( .B1(n20187), .B2(n12247), .A(n13689), .ZN(P1_U3476) );
  XNOR2_X1 U17089 ( .A(n13691), .B(n13690), .ZN(n20176) );
  AOI22_X1 U17090 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13692) );
  OAI21_X1 U17091 ( .B1(n20157), .B2(n13924), .A(n13692), .ZN(n13693) );
  AOI21_X1 U17092 ( .B1(n13694), .B2(n15799), .A(n13693), .ZN(n13695) );
  OAI21_X1 U17093 ( .B1(n20158), .B2(n20176), .A(n13695), .ZN(P1_U2997) );
  NOR2_X1 U17094 ( .A1(n13696), .A2(n16021), .ZN(n15649) );
  OAI22_X1 U17095 ( .A1(n20579), .A2(n20698), .B1(n13871), .B2(n14823), .ZN(
        n13697) );
  OAI21_X1 U17096 ( .B1(n15649), .B2(n13697), .A(n20187), .ZN(n13698) );
  OAI21_X1 U17097 ( .B1(n20187), .B2(n20628), .A(n13698), .ZN(P1_U3478) );
  MUX2_X1 U17098 ( .A(n9853), .B(n13701), .S(n14907), .Z(n13702) );
  OAI21_X1 U17099 ( .B1(n19929), .B2(n14926), .A(n13702), .ZN(P2_U2885) );
  INV_X1 U17100 ( .A(n19066), .ZN(n19096) );
  NAND2_X1 U17101 ( .A1(n9716), .A2(n13704), .ZN(n13705) );
  XNOR2_X1 U17102 ( .A(n16226), .B(n13705), .ZN(n13706) );
  NAND2_X1 U17103 ( .A1(n13706), .A2(n19055), .ZN(n13719) );
  AND2_X1 U17104 ( .A1(n13708), .A2(n13707), .ZN(n13710) );
  OR2_X1 U17105 ( .A1(n13710), .A2(n13709), .ZN(n13711) );
  NAND2_X1 U17106 ( .A1(n13711), .A2(n14040), .ZN(n19923) );
  INV_X1 U17107 ( .A(n19058), .ZN(n19091) );
  OAI22_X1 U17108 ( .A1(n19091), .A2(n13712), .B1(n16240), .B2(n19079), .ZN(
        n13715) );
  OAI22_X1 U17109 ( .A1(n13713), .A2(n19063), .B1(n19034), .B2(n11214), .ZN(
        n13714) );
  NOR2_X1 U17110 ( .A1(n13715), .A2(n13714), .ZN(n13716) );
  OAI21_X1 U17111 ( .B1(n19923), .B2(n19083), .A(n13716), .ZN(n13717) );
  AOI21_X1 U17112 ( .B1(n19093), .B2(n10640), .A(n13717), .ZN(n13718) );
  OAI211_X1 U17113 ( .C1(n19096), .C2(n19323), .A(n13719), .B(n13718), .ZN(
        P2_U2852) );
  INV_X1 U17114 ( .A(n19323), .ZN(n19920) );
  INV_X1 U17115 ( .A(n15390), .ZN(n16370) );
  INV_X1 U17116 ( .A(n13720), .ZN(n15386) );
  NAND2_X1 U17117 ( .A1(n10640), .A2(n15386), .ZN(n13735) );
  NAND2_X1 U17118 ( .A1(n13721), .A2(n16343), .ZN(n15380) );
  INV_X1 U17119 ( .A(n15381), .ZN(n13722) );
  NAND2_X1 U17120 ( .A1(n15380), .A2(n13722), .ZN(n13724) );
  AOI21_X1 U17121 ( .B1(n11180), .B2(n13725), .A(n10665), .ZN(n13723) );
  NAND2_X1 U17122 ( .A1(n13724), .A2(n13723), .ZN(n13732) );
  NAND2_X1 U17123 ( .A1(n15380), .A2(n15381), .ZN(n13730) );
  INV_X1 U17124 ( .A(n13725), .ZN(n13726) );
  NAND2_X1 U17125 ( .A1(n11180), .A2(n13726), .ZN(n15384) );
  OAI21_X1 U17126 ( .B1(n13729), .B2(n13728), .A(n13727), .ZN(n15379) );
  NAND3_X1 U17127 ( .A1(n13730), .A2(n15384), .A3(n15379), .ZN(n13731) );
  MUX2_X1 U17128 ( .A(n13732), .B(n13731), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13733) );
  INV_X1 U17129 ( .A(n13733), .ZN(n13734) );
  NAND2_X1 U17130 ( .A1(n13735), .A2(n13734), .ZN(n16321) );
  AOI22_X1 U17131 ( .A1(n19920), .A2(n16370), .B1(n14001), .B2(n16321), .ZN(
        n13737) );
  INV_X1 U17132 ( .A(n15391), .ZN(n14004) );
  NAND2_X1 U17133 ( .A1(n14004), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13736) );
  OAI21_X1 U17134 ( .B1(n13737), .B2(n14004), .A(n13736), .ZN(P2_U3596) );
  NAND2_X1 U17135 ( .A1(n13738), .A2(n13804), .ZN(n13784) );
  INV_X1 U17136 ( .A(n13804), .ZN(n13739) );
  NAND3_X1 U17137 ( .A1(n13741), .A2(n13740), .A3(n13739), .ZN(n13742) );
  NAND2_X1 U17138 ( .A1(n13784), .A2(n13742), .ZN(n19145) );
  OR2_X1 U17139 ( .A1(n13744), .A2(n13743), .ZN(n13746) );
  NAND2_X1 U17140 ( .A1(n13746), .A2(n13745), .ZN(n19259) );
  MUX2_X1 U17141 ( .A(n19259), .B(n10822), .S(n14907), .Z(n13747) );
  OAI21_X1 U17142 ( .B1(n19145), .B2(n14926), .A(n13747), .ZN(P2_U2883) );
  NAND2_X1 U17143 ( .A1(n11621), .A2(n11619), .ZN(n13748) );
  OAI222_X1 U17144 ( .A1(n13933), .A2(n14679), .B1(n14218), .B2(n20214), .C1(
        n14670), .C2(n20141), .ZN(P1_U2902) );
  INV_X1 U17145 ( .A(n20210), .ZN(n13749) );
  OAI222_X1 U17146 ( .A1(n20163), .A2(n14679), .B1(n14218), .B2(n13749), .C1(
        n14670), .C2(n20143), .ZN(P1_U2903) );
  INV_X1 U17147 ( .A(n20203), .ZN(n13750) );
  OAI222_X1 U17148 ( .A1(n20171), .A2(n14679), .B1(n14218), .B2(n13750), .C1(
        n14670), .C2(n20147), .ZN(P1_U2904) );
  NAND2_X1 U17149 ( .A1(n13751), .A2(n13752), .ZN(n13916) );
  OR2_X1 U17150 ( .A1(n13751), .A2(n13752), .ZN(n13753) );
  AND2_X1 U17151 ( .A1(n13916), .A2(n13753), .ZN(n20105) );
  NAND2_X1 U17152 ( .A1(n13755), .A2(n13754), .ZN(n13756) );
  AND2_X1 U17153 ( .A1(n13893), .A2(n13756), .ZN(n20100) );
  INV_X1 U17154 ( .A(n20100), .ZN(n13758) );
  INV_X1 U17155 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13757) );
  OAI22_X1 U17156 ( .A1(n14612), .A2(n13758), .B1(n13757), .B2(n14611), .ZN(
        n13759) );
  AOI21_X1 U17157 ( .B1(n20105), .B2(n13760), .A(n13759), .ZN(n13761) );
  INV_X1 U17158 ( .A(n13761), .ZN(P1_U2869) );
  INV_X1 U17159 ( .A(n20105), .ZN(n13763) );
  AOI22_X1 U17160 ( .A1(n14173), .A2(n20218), .B1(P1_EAX_REG_3__SCAN_IN), .B2(
        n14666), .ZN(n13762) );
  OAI21_X1 U17161 ( .B1(n13763), .B2(n14679), .A(n13762), .ZN(P1_U2901) );
  XNOR2_X1 U17162 ( .A(n13765), .B(n13766), .ZN(n13776) );
  INV_X1 U17163 ( .A(n13768), .ZN(n13767) );
  NOR2_X1 U17164 ( .A1(n15916), .A2(n13767), .ZN(n20181) );
  OAI21_X1 U17165 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n15966), .A(
        n15946), .ZN(n20173) );
  AOI211_X1 U17166 ( .C1(n12621), .C2(n15943), .A(n20181), .B(n20173), .ZN(
        n13890) );
  INV_X1 U17167 ( .A(n13890), .ZN(n13828) );
  NOR2_X1 U17168 ( .A1(n13768), .A2(n15939), .ZN(n13899) );
  AOI22_X1 U17169 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13828), .B1(
        n13899), .B2(n12625), .ZN(n13771) );
  INV_X1 U17170 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13769) );
  NOR2_X1 U17171 ( .A1(n20177), .A2(n13769), .ZN(n13772) );
  AOI21_X1 U17172 ( .B1(n15999), .B2(n20100), .A(n13772), .ZN(n13770) );
  OAI211_X1 U17173 ( .C1(n15988), .C2(n13776), .A(n13771), .B(n13770), .ZN(
        P1_U3028) );
  AOI21_X1 U17174 ( .B1(n20165), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13772), .ZN(n13773) );
  OAI21_X1 U17175 ( .B1(n20157), .B2(n20101), .A(n13773), .ZN(n13774) );
  AOI21_X1 U17176 ( .B1(n20105), .B2(n15799), .A(n13774), .ZN(n13775) );
  OAI21_X1 U17177 ( .B1(n13776), .B2(n20158), .A(n13775), .ZN(P1_U2996) );
  XOR2_X1 U17178 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13784), .Z(n13781)
         );
  AOI21_X1 U17179 ( .B1(n13777), .B2(n13745), .A(n13787), .ZN(n19053) );
  NOR2_X1 U17180 ( .A1(n14936), .A2(n13778), .ZN(n13779) );
  AOI21_X1 U17181 ( .B1(n19053), .B2(n14936), .A(n13779), .ZN(n13780) );
  OAI21_X1 U17182 ( .B1(n13781), .B2(n14926), .A(n13780), .ZN(P2_U2882) );
  INV_X1 U17183 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13782) );
  NOR2_X1 U17184 ( .A1(n13784), .A2(n13782), .ZN(n13785) );
  OR2_X1 U17185 ( .A1(n13784), .A2(n13783), .ZN(n13816) );
  OAI211_X1 U17186 ( .C1(n13785), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14939), .B(n13816), .ZN(n13791) );
  NOR2_X1 U17187 ( .A1(n13788), .A2(n13787), .ZN(n13789) );
  OR2_X1 U17188 ( .A1(n13786), .A2(n13789), .ZN(n15149) );
  INV_X1 U17189 ( .A(n15149), .ZN(n19042) );
  NAND2_X1 U17190 ( .A1(n19042), .A2(n14936), .ZN(n13790) );
  OAI211_X1 U17191 ( .C1(n14936), .C2(n19035), .A(n13791), .B(n13790), .ZN(
        P2_U2881) );
  NAND2_X1 U17192 ( .A1(n13738), .A2(n13792), .ZN(n13807) );
  INV_X1 U17193 ( .A(n13807), .ZN(n13795) );
  NAND2_X1 U17194 ( .A1(n13738), .A2(n13793), .ZN(n13878) );
  OAI211_X1 U17195 ( .C1(n13795), .C2(n13794), .A(n14939), .B(n13878), .ZN(
        n13799) );
  AOI21_X1 U17196 ( .B1(n13797), .B2(n13802), .A(n13796), .ZN(n19009) );
  NAND2_X1 U17197 ( .A1(n19009), .A2(n14936), .ZN(n13798) );
  OAI211_X1 U17198 ( .C1(n14936), .C2(n9892), .A(n13799), .B(n13798), .ZN(
        P2_U2878) );
  OR2_X1 U17199 ( .A1(n13800), .A2(n13801), .ZN(n13803) );
  NAND2_X1 U17200 ( .A1(n13803), .A2(n13802), .ZN(n19023) );
  AND2_X1 U17201 ( .A1(n13738), .A2(n13804), .ZN(n13806) );
  AND2_X1 U17202 ( .A1(n13806), .A2(n13805), .ZN(n13809) );
  OAI211_X1 U17203 ( .C1(n13809), .C2(n13808), .A(n13807), .B(n14939), .ZN(
        n13811) );
  NAND2_X1 U17204 ( .A1(n14884), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13810) );
  OAI211_X1 U17205 ( .C1(n19023), .C2(n14907), .A(n13811), .B(n13810), .ZN(
        P2_U2879) );
  OR2_X1 U17206 ( .A1(n13916), .A2(n13813), .ZN(n13914) );
  NAND2_X1 U17207 ( .A1(n13814), .A2(n13914), .ZN(n13815) );
  NAND2_X1 U17208 ( .A1(n13812), .A2(n13815), .ZN(n20068) );
  OAI222_X1 U17209 ( .A1(n20068), .A2(n14679), .B1(n14218), .B2(n20225), .C1(
        n14670), .C2(n11786), .ZN(P1_U2899) );
  XOR2_X1 U17210 ( .A(n13816), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13821)
         );
  NOR2_X1 U17211 ( .A1(n13786), .A2(n13817), .ZN(n13818) );
  OR2_X1 U17212 ( .A1(n13800), .A2(n13818), .ZN(n19029) );
  MUX2_X1 U17213 ( .A(n19029), .B(n13819), .S(n14907), .Z(n13820) );
  OAI21_X1 U17214 ( .B1(n13821), .B2(n14926), .A(n13820), .ZN(P2_U2880) );
  XNOR2_X1 U17215 ( .A(n13823), .B(n13824), .ZN(n13921) );
  NAND2_X1 U17216 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13825) );
  OAI211_X1 U17217 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13899), .B(n13825), .ZN(n13830) );
  INV_X1 U17218 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20786) );
  NOR2_X1 U17219 ( .A1(n20177), .A2(n20786), .ZN(n13917) );
  INV_X1 U17220 ( .A(n13895), .ZN(n13826) );
  XNOR2_X1 U17221 ( .A(n13893), .B(n13826), .ZN(n20080) );
  NOR2_X1 U17222 ( .A1(n20179), .A2(n20080), .ZN(n13827) );
  AOI211_X1 U17223 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n13828), .A(
        n13917), .B(n13827), .ZN(n13829) );
  OAI211_X1 U17224 ( .C1(n15988), .C2(n13921), .A(n13830), .B(n13829), .ZN(
        P1_U3027) );
  NOR2_X1 U17225 ( .A1(n19069), .A2(n13903), .ZN(n13832) );
  XNOR2_X1 U17226 ( .A(n13832), .B(n13831), .ZN(n13833) );
  NAND2_X1 U17227 ( .A1(n13833), .A2(n19055), .ZN(n13841) );
  INV_X1 U17228 ( .A(n13834), .ZN(n13836) );
  AOI22_X1 U17229 ( .A1(n19081), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n19058), .ZN(n13835) );
  OAI21_X1 U17230 ( .B1(n13836), .B2(n19063), .A(n13835), .ZN(n13839) );
  INV_X1 U17231 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13837) );
  OAI22_X1 U17232 ( .A1(n19137), .A2(n19083), .B1(n13837), .B2(n19079), .ZN(
        n13838) );
  AOI211_X1 U17233 ( .C1(n19093), .C2(n15387), .A(n13839), .B(n13838), .ZN(
        n13840) );
  OAI211_X1 U17234 ( .C1(n19096), .C2(n19929), .A(n13841), .B(n13840), .ZN(
        P2_U2853) );
  NAND2_X1 U17235 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20867), .ZN(n16015) );
  AND2_X1 U17236 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20761), .ZN(n13842) );
  NAND2_X1 U17237 ( .A1(n13843), .A2(n13842), .ZN(n13844) );
  OAI211_X1 U17238 ( .C1(n16015), .C2(n20761), .A(n20177), .B(n13844), .ZN(
        n13845) );
  INV_X1 U17239 ( .A(n13845), .ZN(n13846) );
  NAND2_X1 U17240 ( .A1(n13848), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13850) );
  INV_X1 U17241 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13849) );
  NOR2_X1 U17242 ( .A1(n14351), .A2(n20760), .ZN(n13851) );
  AND3_X1 U17243 ( .A1(n14458), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n13852), 
        .ZN(n13853) );
  INV_X1 U17244 ( .A(n20104), .ZN(n13941) );
  AND2_X1 U17245 ( .A1(n13854), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13855) );
  NAND2_X1 U17246 ( .A1(n14458), .A2(n13855), .ZN(n13865) );
  OR2_X1 U17247 ( .A1(n13856), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13859) );
  NOR2_X1 U17248 ( .A1(n13857), .A2(n20764), .ZN(n13858) );
  AND2_X1 U17249 ( .A1(n14458), .A2(n13858), .ZN(n20077) );
  INV_X1 U17250 ( .A(n20077), .ZN(n20095) );
  INV_X1 U17251 ( .A(n13859), .ZN(n13862) );
  AND2_X1 U17252 ( .A1(n13860), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13861) );
  NAND2_X1 U17253 ( .A1(n20864), .A2(n20633), .ZN(n13863) );
  NAND2_X1 U17254 ( .A1(n13863), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13864) );
  INV_X1 U17255 ( .A(n13866), .ZN(n13867) );
  AOI22_X1 U17256 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(n20093), .B1(n20099), .B2(
        n13867), .ZN(n13870) );
  OAI21_X1 U17257 ( .B1(n20092), .B2(n20102), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13869) );
  OAI211_X1 U17258 ( .C1(n20095), .C2(n13871), .A(n13870), .B(n13869), .ZN(
        n13872) );
  AOI21_X1 U17259 ( .B1(n15737), .B2(P1_REIP_REG_0__SCAN_IN), .A(n13872), .ZN(
        n13873) );
  OAI21_X1 U17260 ( .B1(n13941), .B2(n20171), .A(n13873), .ZN(P1_U2840) );
  INV_X1 U17261 ( .A(n13874), .ZN(n13875) );
  XNOR2_X1 U17262 ( .A(n13812), .B(n13875), .ZN(n20052) );
  INV_X1 U17263 ( .A(n20052), .ZN(n13885) );
  XOR2_X1 U17264 ( .A(n13956), .B(n13957), .Z(n20049) );
  AOI22_X1 U17265 ( .A1(n20049), .A2(n14607), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14568), .ZN(n13876) );
  OAI21_X1 U17266 ( .B1(n13885), .B2(n14595), .A(n13876), .ZN(P1_U2866) );
  AND2_X1 U17267 ( .A1(n13738), .A2(n13877), .ZN(n13944) );
  AOI211_X1 U17268 ( .C1(n13879), .C2(n13878), .A(n14926), .B(n13944), .ZN(
        n13880) );
  INV_X1 U17269 ( .A(n13880), .ZN(n13884) );
  OR2_X1 U17270 ( .A1(n13881), .A2(n13796), .ZN(n13882) );
  NAND2_X1 U17271 ( .A1(n13882), .A2(n13946), .ZN(n18999) );
  INV_X1 U17272 ( .A(n18999), .ZN(n16193) );
  NAND2_X1 U17273 ( .A1(n16193), .A2(n14936), .ZN(n13883) );
  OAI211_X1 U17274 ( .C1(n14936), .C2(n18991), .A(n13884), .B(n13883), .ZN(
        P2_U2877) );
  OAI222_X1 U17275 ( .A1(n14679), .A2(n13885), .B1(n14218), .B2(n20229), .C1(
        n14670), .C2(n11862), .ZN(P1_U2898) );
  XNOR2_X1 U17276 ( .A(n13888), .B(n13887), .ZN(n15833) );
  INV_X1 U17277 ( .A(n13889), .ZN(n13891) );
  OAI21_X1 U17278 ( .B1(n13892), .B2(n13891), .A(n13890), .ZN(n16001) );
  INV_X1 U17279 ( .A(n13893), .ZN(n13896) );
  AOI21_X1 U17280 ( .B1(n13896), .B2(n13895), .A(n13894), .ZN(n13897) );
  OR2_X1 U17281 ( .A1(n13897), .A2(n13957), .ZN(n20061) );
  NAND4_X1 U17282 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n13899), .A4(n13898), .ZN(
        n13900) );
  NAND2_X1 U17283 ( .A1(n16000), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n15835) );
  OAI211_X1 U17284 ( .C1(n20179), .C2(n20061), .A(n13900), .B(n15835), .ZN(
        n13901) );
  AOI21_X1 U17285 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16001), .A(
        n13901), .ZN(n13902) );
  OAI21_X1 U17286 ( .B1(n15988), .B2(n15833), .A(n13902), .ZN(P1_U3026) );
  NOR2_X1 U17287 ( .A1(n9715), .A2(n19825), .ZN(n18947) );
  INV_X1 U17288 ( .A(n18947), .ZN(n19078) );
  AOI211_X1 U17289 ( .C1(n19076), .C2(n13904), .A(n19069), .B(n13903), .ZN(
        n14000) );
  NAND2_X1 U17290 ( .A1(n14000), .A2(n19055), .ZN(n13913) );
  XNOR2_X1 U17291 ( .A(n13906), .B(n13905), .ZN(n19941) );
  NOR2_X1 U17292 ( .A1(n19063), .A2(n14383), .ZN(n13909) );
  AOI22_X1 U17293 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9707), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n19058), .ZN(n13907) );
  OAI21_X1 U17294 ( .B1(n19034), .B2(n19853), .A(n13907), .ZN(n13908) );
  AOI211_X1 U17295 ( .C1(n19941), .C2(n19019), .A(n13909), .B(n13908), .ZN(
        n13910) );
  OAI21_X1 U17296 ( .B1(n14399), .B2(n19075), .A(n13910), .ZN(n13911) );
  AOI21_X1 U17297 ( .B1(n19917), .B2(n19066), .A(n13911), .ZN(n13912) );
  OAI211_X1 U17298 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19078), .A(
        n13913), .B(n13912), .ZN(P2_U2854) );
  INV_X1 U17299 ( .A(n13914), .ZN(n13915) );
  AOI21_X1 U17300 ( .B1(n13813), .B2(n13916), .A(n13915), .ZN(n20085) );
  AOI21_X1 U17301 ( .B1(n20165), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13917), .ZN(n13918) );
  OAI21_X1 U17302 ( .B1(n20157), .B2(n20089), .A(n13918), .ZN(n13919) );
  AOI21_X1 U17303 ( .B1(n20085), .B2(n15799), .A(n13919), .ZN(n13920) );
  OAI21_X1 U17304 ( .B1(n13921), .B2(n20158), .A(n13920), .ZN(P1_U2995) );
  INV_X1 U17305 ( .A(n20085), .ZN(n13923) );
  OAI222_X1 U17306 ( .A1(n13923), .A2(n14679), .B1(n14218), .B2(n20222), .C1(
        n14670), .C2(n20137), .ZN(P1_U2900) );
  INV_X1 U17307 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13922) );
  OAI222_X1 U17308 ( .A1(n13923), .A2(n14595), .B1(n14612), .B2(n20080), .C1(
        n14611), .C2(n13922), .ZN(P1_U2868) );
  NAND2_X1 U17309 ( .A1(n20784), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13928) );
  INV_X1 U17310 ( .A(n13924), .ZN(n13925) );
  AOI22_X1 U17311 ( .A1(n13925), .A2(n20102), .B1(n20092), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13927) );
  NAND2_X1 U17312 ( .A1(n20093), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13926) );
  OAI211_X1 U17313 ( .C1(n13928), .C2(n20091), .A(n13927), .B(n13926), .ZN(
        n13931) );
  INV_X1 U17314 ( .A(n14458), .ZN(n14500) );
  AOI21_X1 U17315 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .A(n20091), .ZN(n13929) );
  NOR2_X1 U17316 ( .A1(n14500), .A2(n13929), .ZN(n20108) );
  OAI22_X1 U17317 ( .A1(n20108), .A2(n20784), .B1(n20081), .B2(n20178), .ZN(
        n13930) );
  AOI211_X1 U17318 ( .C1(n20199), .C2(n20077), .A(n13931), .B(n13930), .ZN(
        n13932) );
  OAI21_X1 U17319 ( .B1(n13941), .B2(n13933), .A(n13932), .ZN(P1_U2838) );
  INV_X1 U17320 ( .A(n20392), .ZN(n20659) );
  OAI22_X1 U17321 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n20091), .B1(n20024), 
        .B2(n13935), .ZN(n13939) );
  NAND2_X1 U17322 ( .A1(n20099), .A2(n13590), .ZN(n13937) );
  AOI22_X1 U17323 ( .A1(n20092), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14500), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13936) );
  OAI211_X1 U17324 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20088), .A(
        n13937), .B(n13936), .ZN(n13938) );
  AOI211_X1 U17325 ( .C1(n20659), .C2(n20077), .A(n13939), .B(n13938), .ZN(
        n13940) );
  OAI21_X1 U17326 ( .B1(n20163), .B2(n13941), .A(n13940), .ZN(P1_U2839) );
  INV_X1 U17327 ( .A(n14346), .ZN(n13942) );
  OAI211_X1 U17328 ( .C1(n13944), .C2(n13943), .A(n13942), .B(n14939), .ZN(
        n13949) );
  AOI21_X1 U17329 ( .B1(n13947), .B2(n13946), .A(n13945), .ZN(n18986) );
  NAND2_X1 U17330 ( .A1(n18986), .A2(n14936), .ZN(n13948) );
  OAI211_X1 U17331 ( .C1(n14936), .C2(n13950), .A(n13949), .B(n13948), .ZN(
        P2_U2876) );
  OR2_X1 U17332 ( .A1(n13953), .A2(n13952), .ZN(n13954) );
  AND2_X1 U17333 ( .A1(n13951), .A2(n13954), .ZN(n20044) );
  INV_X1 U17334 ( .A(n20044), .ZN(n13962) );
  INV_X1 U17335 ( .A(n14031), .ZN(n13959) );
  AOI21_X1 U17336 ( .B1(n13957), .B2(n13956), .A(n13955), .ZN(n13958) );
  NOR2_X1 U17337 ( .A1(n13959), .A2(n13958), .ZN(n20038) );
  AOI22_X1 U17338 ( .A1(n20038), .A2(n14607), .B1(n14568), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n13960) );
  OAI21_X1 U17339 ( .B1(n13962), .B2(n14595), .A(n13960), .ZN(P1_U2865) );
  AOI22_X1 U17340 ( .A1(n14173), .A2(n20237), .B1(P1_EAX_REG_7__SCAN_IN), .B2(
        n14666), .ZN(n13961) );
  OAI21_X1 U17341 ( .B1(n13962), .B2(n14679), .A(n13961), .ZN(P1_U2897) );
  XNOR2_X1 U17342 ( .A(n19929), .B(n19137), .ZN(n13967) );
  INV_X1 U17343 ( .A(n19941), .ZN(n13963) );
  NAND2_X1 U17344 ( .A1(n19937), .A2(n13963), .ZN(n13964) );
  OAI21_X1 U17345 ( .B1(n19937), .B2(n13963), .A(n13964), .ZN(n19160) );
  NOR2_X1 U17346 ( .A1(n19160), .A2(n19161), .ZN(n19159) );
  INV_X1 U17347 ( .A(n13964), .ZN(n13965) );
  NOR2_X1 U17348 ( .A1(n19159), .A2(n13965), .ZN(n13966) );
  NOR2_X1 U17349 ( .A1(n13966), .A2(n13967), .ZN(n19136) );
  AOI21_X1 U17350 ( .B1(n13967), .B2(n13966), .A(n19136), .ZN(n13970) );
  INV_X1 U17351 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16505) );
  INV_X1 U17352 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18198) );
  AOI22_X1 U17353 ( .A1(n16121), .A2(n16505), .B1(n18198), .B2(n16122), .ZN(
        n16131) );
  AOI22_X1 U17354 ( .A1(n19134), .A2(n16131), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19157), .ZN(n13969) );
  NAND2_X1 U17355 ( .A1(n19931), .A2(n19158), .ZN(n13968) );
  OAI211_X1 U17356 ( .C1(n13970), .C2(n19162), .A(n13969), .B(n13968), .ZN(
        P2_U2917) );
  INV_X1 U17357 ( .A(n13971), .ZN(n13972) );
  AOI21_X1 U17358 ( .B1(n13973), .B2(n13951), .A(n13972), .ZN(n13993) );
  INV_X1 U17359 ( .A(n13993), .ZN(n20030) );
  AOI22_X1 U17360 ( .A1(n14173), .A2(n14636), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14666), .ZN(n13974) );
  OAI21_X1 U17361 ( .B1(n20030), .B2(n14679), .A(n13974), .ZN(P1_U2896) );
  NAND2_X1 U17362 ( .A1(n19323), .A2(n14106), .ZN(n19506) );
  OAI21_X1 U17363 ( .B1(n19486), .B2(n19521), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13982) );
  NAND2_X1 U17364 ( .A1(n19718), .A2(n19413), .ZN(n13985) );
  INV_X1 U17365 ( .A(n19413), .ZN(n19496) );
  NOR2_X1 U17366 ( .A1(n19496), .A2(n19593), .ZN(n19489) );
  INV_X1 U17367 ( .A(n19489), .ZN(n13975) );
  NAND2_X1 U17368 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13975), .ZN(n13976) );
  NOR2_X1 U17369 ( .A1(n10757), .A2(n13976), .ZN(n13984) );
  NOR2_X1 U17370 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19975) );
  INV_X1 U17371 ( .A(n19975), .ZN(n13979) );
  INV_X1 U17372 ( .A(n13977), .ZN(n13978) );
  NAND2_X1 U17373 ( .A1(n13979), .A2(n13978), .ZN(n13980) );
  OAI21_X1 U17374 ( .B1(n19489), .B2(n19533), .A(n19768), .ZN(n13981) );
  AOI211_X1 U17375 ( .C1(n13982), .C2(n13985), .A(n13984), .B(n13981), .ZN(
        n19475) );
  INV_X1 U17376 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13988) );
  AOI22_X1 U17377 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19314), .ZN(n19729) );
  AOI22_X1 U17378 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19314), .ZN(n19773) );
  AOI22_X1 U17379 ( .A1(n19521), .A2(n19770), .B1(n19486), .B2(n19715), .ZN(
        n13987) );
  INV_X1 U17380 ( .A(n19820), .ZN(n19681) );
  AOI211_X2 U17381 ( .C1(n19973), .C2(n13985), .A(n19681), .B(n13984), .ZN(
        n19490) );
  INV_X1 U17382 ( .A(n19104), .ZN(n19234) );
  NOR2_X2 U17383 ( .A1(n19234), .A2(n19357), .ZN(n19762) );
  NOR2_X2 U17384 ( .A1(n16351), .A2(n19310), .ZN(n19761) );
  AOI22_X1 U17385 ( .A1(n19490), .A2(n19762), .B1(n19761), .B2(n19489), .ZN(
        n13986) );
  OAI211_X1 U17386 ( .C1(n19475), .C2(n13988), .A(n13987), .B(n13986), .ZN(
        P2_U3096) );
  INV_X1 U17387 ( .A(n20032), .ZN(n13991) );
  AOI22_X1 U17388 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13990) );
  OAI21_X1 U17389 ( .B1(n20157), .B2(n13991), .A(n13990), .ZN(n13992) );
  AOI21_X1 U17390 ( .B1(n13993), .B2(n15799), .A(n13992), .ZN(n13994) );
  OAI21_X1 U17391 ( .B1(n15987), .B2(n20158), .A(n13994), .ZN(P1_U2991) );
  NAND2_X1 U17392 ( .A1(n13995), .A2(n15386), .ZN(n13999) );
  NAND2_X1 U17393 ( .A1(n10563), .A2(n13996), .ZN(n15370) );
  XNOR2_X1 U17394 ( .A(n15369), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13997) );
  AOI22_X1 U17395 ( .A1(n9855), .A2(n11180), .B1(n15370), .B2(n13997), .ZN(
        n13998) );
  AND2_X1 U17396 ( .A1(n13999), .A2(n13998), .ZN(n16326) );
  INV_X1 U17397 ( .A(n16326), .ZN(n14002) );
  OAI22_X1 U17398 ( .A1(n9716), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19076), .B2(n19069), .ZN(n15372) );
  NOR2_X1 U17399 ( .A1(n15374), .A2(n15372), .ZN(n15377) );
  AOI21_X1 U17400 ( .B1(n19069), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n14000), .ZN(n15388) );
  AOI222_X1 U17401 ( .A1(n14002), .A2(n14001), .B1(n15377), .B2(n15388), .C1(
        n16370), .C2(n19917), .ZN(n14005) );
  NAND2_X1 U17402 ( .A1(n14004), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14003) );
  OAI21_X1 U17403 ( .B1(n14005), .B2(n14004), .A(n14003), .ZN(P2_U3600) );
  OAI211_X1 U17404 ( .C1(n12861), .C2(n12860), .A(n14939), .B(n14007), .ZN(
        n14013) );
  NAND2_X1 U17405 ( .A1(n14008), .A2(n14342), .ZN(n14011) );
  INV_X1 U17406 ( .A(n14009), .ZN(n14010) );
  NAND2_X1 U17407 ( .A1(n16167), .A2(n14936), .ZN(n14012) );
  OAI211_X1 U17408 ( .C1(n14936), .C2(n11131), .A(n14013), .B(n14012), .ZN(
        P2_U2874) );
  OAI21_X1 U17409 ( .B1(n14014), .B2(n14009), .A(n14065), .ZN(n18966) );
  INV_X1 U17410 ( .A(n14007), .ZN(n14018) );
  INV_X1 U17411 ( .A(n14015), .ZN(n14016) );
  OAI211_X1 U17412 ( .C1(n14018), .C2(n14017), .A(n14016), .B(n14939), .ZN(
        n14020) );
  NAND2_X1 U17413 ( .A1(n14884), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14019) );
  OAI211_X1 U17414 ( .C1(n18966), .C2(n14907), .A(n14020), .B(n14019), .ZN(
        P2_U2873) );
  AND2_X1 U17415 ( .A1(n13971), .A2(n14021), .ZN(n14023) );
  OR2_X1 U17416 ( .A1(n14023), .A2(n14022), .ZN(n20019) );
  AOI22_X1 U17417 ( .A1(n14173), .A2(n14632), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14666), .ZN(n14024) );
  OAI21_X1 U17418 ( .B1(n20019), .B2(n14679), .A(n14024), .ZN(P1_U2895) );
  AND2_X1 U17419 ( .A1(n14033), .A2(n14025), .ZN(n14026) );
  OR2_X1 U17420 ( .A1(n14026), .A2(n9804), .ZN(n15977) );
  INV_X1 U17421 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14027) );
  OAI22_X1 U17422 ( .A1(n15977), .A2(n14612), .B1(n14027), .B2(n14611), .ZN(
        n14028) );
  INV_X1 U17423 ( .A(n14028), .ZN(n14029) );
  OAI21_X1 U17424 ( .B1(n20019), .B2(n14609), .A(n14029), .ZN(P1_U2863) );
  NAND2_X1 U17425 ( .A1(n14031), .A2(n14030), .ZN(n14032) );
  NAND2_X1 U17426 ( .A1(n14033), .A2(n14032), .ZN(n20036) );
  INV_X1 U17427 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14034) );
  OAI222_X1 U17428 ( .A1(n20036), .A2(n14612), .B1(n14611), .B2(n14034), .C1(
        n14609), .C2(n20030), .ZN(P1_U2864) );
  XOR2_X1 U17429 ( .A(n14036), .B(n14035), .Z(n19265) );
  INV_X1 U17430 ( .A(n19265), .ZN(n14047) );
  XNOR2_X1 U17431 ( .A(n14037), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14038) );
  XNOR2_X1 U17432 ( .A(n14039), .B(n14038), .ZN(n19261) );
  AOI21_X1 U17433 ( .B1(n14041), .B2(n14040), .A(n14098), .ZN(n19143) );
  AOI22_X1 U17434 ( .A1(n16281), .A2(n19143), .B1(n15077), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n14042) );
  OAI21_X1 U17435 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14092), .A(
        n14042), .ZN(n14045) );
  NAND3_X1 U17436 ( .A1(n14099), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        n16311), .ZN(n14043) );
  OAI21_X1 U17437 ( .B1(n19259), .B2(n16283), .A(n14043), .ZN(n14044) );
  AOI211_X1 U17438 ( .C1(n19261), .C2(n16274), .A(n14045), .B(n14044), .ZN(
        n14046) );
  OAI21_X1 U17439 ( .B1(n14047), .B2(n16315), .A(n14046), .ZN(P2_U3042) );
  INV_X1 U17440 ( .A(n14022), .ZN(n14050) );
  AOI21_X1 U17441 ( .B1(n10019), .B2(n14050), .A(n9720), .ZN(n14192) );
  INV_X1 U17442 ( .A(n14192), .ZN(n14061) );
  AOI22_X1 U17443 ( .A1(n14173), .A2(n14629), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14666), .ZN(n14051) );
  OAI21_X1 U17444 ( .B1(n14061), .B2(n14679), .A(n14051), .ZN(P1_U2894) );
  NAND2_X1 U17445 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14131) );
  NAND4_X1 U17446 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14413)
         );
  INV_X1 U17447 ( .A(n14413), .ZN(n14055) );
  NAND4_X1 U17448 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n14414)
         );
  NOR2_X1 U17449 ( .A1(n14500), .A2(n14414), .ZN(n20059) );
  AOI21_X1 U17450 ( .B1(n14055), .B2(n20059), .A(n20060), .ZN(n20027) );
  AOI21_X1 U17451 ( .B1(n14131), .B2(n15737), .A(n20027), .ZN(n15759) );
  INV_X1 U17452 ( .A(n15759), .ZN(n15736) );
  INV_X1 U17453 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14052) );
  OAI22_X1 U17454 ( .A1(n20088), .A2(n14190), .B1(n20024), .B2(n14052), .ZN(
        n14059) );
  NOR2_X1 U17455 ( .A1(n9804), .A2(n14053), .ZN(n14054) );
  OR2_X1 U17456 ( .A1(n9742), .A2(n14054), .ZN(n15972) );
  INV_X1 U17457 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20796) );
  NAND2_X1 U17458 ( .A1(n14055), .A2(n20067), .ZN(n20013) );
  NOR3_X1 U17459 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20796), .A3(n20013), 
        .ZN(n14056) );
  AOI211_X1 U17460 ( .C1(n20092), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16000), .B(n14056), .ZN(n14057) );
  OAI21_X1 U17461 ( .B1(n20081), .B2(n15972), .A(n14057), .ZN(n14058) );
  AOI211_X1 U17462 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n15736), .A(n14059), 
        .B(n14058), .ZN(n14060) );
  OAI21_X1 U17463 ( .B1(n14061), .B2(n20029), .A(n14060), .ZN(P1_U2830) );
  OAI222_X1 U17464 ( .A1(n15972), .A2(n14612), .B1(n14611), .B2(n14052), .C1(
        n14609), .C2(n14061), .ZN(P1_U2862) );
  INV_X1 U17465 ( .A(n14207), .ZN(n14062) );
  OAI211_X1 U17466 ( .C1(n14015), .C2(n14063), .A(n14062), .B(n14939), .ZN(
        n14068) );
  NAND2_X1 U17467 ( .A1(n14065), .A2(n14064), .ZN(n14066) );
  AND2_X1 U17468 ( .A1(n14146), .A2(n14066), .ZN(n18952) );
  NAND2_X1 U17469 ( .A1(n18952), .A2(n14936), .ZN(n14067) );
  OAI211_X1 U17470 ( .C1(n14936), .C2(n11143), .A(n14068), .B(n14067), .ZN(
        P2_U2872) );
  NOR2_X1 U17471 ( .A1(n19069), .A2(n19825), .ZN(n16030) );
  INV_X1 U17472 ( .A(n16030), .ZN(n19099) );
  NOR2_X1 U17473 ( .A1(n18957), .A2(n19099), .ZN(n18963) );
  NAND2_X1 U17474 ( .A1(n16163), .A2(n14069), .ZN(n14073) );
  INV_X1 U17475 ( .A(n16167), .ZN(n15304) );
  OAI21_X1 U17476 ( .B1(n14071), .B2(n15314), .A(n16253), .ZN(n19119) );
  OAI22_X1 U17477 ( .A1(n15304), .A2(n19075), .B1(n19119), .B2(n19083), .ZN(
        n14072) );
  AOI21_X1 U17478 ( .B1(n18963), .B2(n14073), .A(n14072), .ZN(n14077) );
  INV_X1 U17479 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19871) );
  AOI22_X1 U17480 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n9707), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19058), .ZN(n14074) );
  OAI211_X1 U17481 ( .C1(n19871), .C2(n19034), .A(n14074), .B(n9722), .ZN(
        n14075) );
  AOI21_X1 U17482 ( .B1(n16163), .B2(n18947), .A(n14075), .ZN(n14076) );
  OAI211_X1 U17483 ( .C1(n14078), .C2(n19063), .A(n14077), .B(n14076), .ZN(
        P2_U2842) );
  XNOR2_X1 U17484 ( .A(n9711), .B(n15983), .ZN(n14079) );
  XNOR2_X1 U17485 ( .A(n14080), .B(n14079), .ZN(n15979) );
  OAI22_X1 U17486 ( .A1(n15837), .A2(n20016), .B1(n20177), .B2(n20796), .ZN(
        n14082) );
  NOR2_X1 U17487 ( .A1(n20019), .A2(n20191), .ZN(n14081) );
  AOI211_X1 U17488 ( .C1(n15809), .C2(n20020), .A(n14082), .B(n14081), .ZN(
        n14083) );
  OAI21_X1 U17489 ( .B1(n15979), .B2(n20158), .A(n14083), .ZN(P1_U2990) );
  XNOR2_X1 U17490 ( .A(n14085), .B(n14084), .ZN(n16221) );
  OAI21_X1 U17491 ( .B1(n14089), .B2(n14087), .A(n14086), .ZN(n14088) );
  OAI21_X1 U17492 ( .B1(n14090), .B2(n14089), .A(n14088), .ZN(n16218) );
  INV_X1 U17493 ( .A(n16218), .ZN(n14104) );
  INV_X1 U17494 ( .A(n14091), .ZN(n14093) );
  AOI211_X1 U17495 ( .C1(n14095), .C2(n14094), .A(n14093), .B(n14092), .ZN(
        n14103) );
  OAI21_X1 U17496 ( .B1(n14098), .B2(n14097), .A(n14096), .ZN(n19141) );
  INV_X1 U17497 ( .A(n16281), .ZN(n16306) );
  AOI22_X1 U17498 ( .A1(n12589), .A2(n19053), .B1(n15077), .B2(
        P2_REIP_REG_5__SCAN_IN), .ZN(n14101) );
  NAND3_X1 U17499 ( .A1(n14099), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n16311), .ZN(n14100) );
  OAI211_X1 U17500 ( .C1(n19141), .C2(n16306), .A(n14101), .B(n14100), .ZN(
        n14102) );
  AOI211_X1 U17501 ( .C1(n14104), .C2(n16274), .A(n14103), .B(n14102), .ZN(
        n14105) );
  OAI21_X1 U17502 ( .B1(n16315), .B2(n16221), .A(n14105), .ZN(P2_U3041) );
  NOR2_X2 U17503 ( .A1(n19713), .A2(n19676), .ZN(n19709) );
  NOR2_X2 U17504 ( .A1(n19675), .A2(n19915), .ZN(n19670) );
  OAI21_X1 U17505 ( .B1(n19709), .B2(n19670), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14112) );
  INV_X1 U17506 ( .A(n19718), .ZN(n19411) );
  NAND3_X1 U17507 ( .A1(n19418), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n19411), .ZN(n14111) );
  NOR2_X1 U17508 ( .A1(n19926), .A2(n19933), .ZN(n19717) );
  NAND2_X1 U17509 ( .A1(n19717), .A2(n19943), .ZN(n19684) );
  NOR2_X1 U17510 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19684), .ZN(
        n19668) );
  INV_X1 U17511 ( .A(n19668), .ZN(n14107) );
  NAND2_X1 U17512 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n14107), .ZN(n14108) );
  NOR2_X1 U17513 ( .A1(n14109), .A2(n14108), .ZN(n14113) );
  OAI21_X1 U17514 ( .B1(n19668), .B2(n19533), .A(n19768), .ZN(n14110) );
  INV_X1 U17515 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U17516 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19314), .ZN(n19735) );
  AOI22_X1 U17517 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19314), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19315), .ZN(n19785) );
  AOI22_X1 U17518 ( .A1(n19709), .A2(n19782), .B1(n19670), .B2(n19732), .ZN(
        n14116) );
  NAND4_X1 U17519 ( .A1(n19418), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n19411), .A4(n19533), .ZN(n14114) );
  AOI21_X1 U17520 ( .B1(n19973), .B2(n14114), .A(n14113), .ZN(n19669) );
  INV_X1 U17521 ( .A(n16131), .ZN(n19237) );
  NOR2_X2 U17522 ( .A1(n19237), .A2(n19357), .ZN(n19781) );
  NOR2_X2 U17523 ( .A1(n10544), .A2(n19310), .ZN(n19780) );
  AOI22_X1 U17524 ( .A1(n19669), .A2(n19781), .B1(n19668), .B2(n19780), .ZN(
        n14115) );
  OAI211_X1 U17525 ( .C1(n19674), .C2(n14117), .A(n14116), .B(n14115), .ZN(
        P2_U3146) );
  INV_X1 U17526 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14120) );
  AOI22_X1 U17527 ( .A1(n19709), .A2(n19770), .B1(n19670), .B2(n19715), .ZN(
        n14119) );
  AOI22_X1 U17528 ( .A1(n19669), .A2(n19762), .B1(n19761), .B2(n19668), .ZN(
        n14118) );
  OAI211_X1 U17529 ( .C1(n19674), .C2(n14120), .A(n14119), .B(n14118), .ZN(
        P2_U3144) );
  OAI21_X1 U17530 ( .B1(n14147), .B2(n14122), .A(n14121), .ZN(n15241) );
  NAND2_X1 U17531 ( .A1(n14207), .A2(n14144), .ZN(n14143) );
  OR2_X1 U17532 ( .A1(n14143), .A2(n14124), .ZN(n14209) );
  INV_X1 U17533 ( .A(n14209), .ZN(n14123) );
  AOI21_X1 U17534 ( .B1(n14124), .B2(n14143), .A(n14123), .ZN(n15024) );
  NAND2_X1 U17535 ( .A1(n15024), .A2(n14939), .ZN(n14126) );
  NAND2_X1 U17536 ( .A1(n14884), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14125) );
  OAI211_X1 U17537 ( .C1(n15241), .C2(n14907), .A(n14126), .B(n14125), .ZN(
        P2_U2870) );
  OR2_X1 U17538 ( .A1(n14128), .A2(n14129), .ZN(n14130) );
  AND2_X1 U17539 ( .A1(n14127), .A2(n14130), .ZN(n15800) );
  INV_X1 U17540 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20805) );
  INV_X1 U17541 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20804) );
  INV_X1 U17542 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20802) );
  INV_X1 U17543 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20800) );
  NOR4_X1 U17544 ( .A1(n20805), .A2(n20804), .A3(n20802), .A4(n20800), .ZN(
        n14412) );
  OAI21_X1 U17545 ( .B1(n14412), .B2(n20060), .A(n15759), .ZN(n14533) );
  NOR2_X1 U17546 ( .A1(n14131), .A2(n20013), .ZN(n15756) );
  NAND3_X1 U17547 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n15756), .ZN(n15741) );
  OAI21_X1 U17548 ( .B1(n20804), .B2(n15741), .A(n20805), .ZN(n14138) );
  OR2_X1 U17549 ( .A1(n14164), .A2(n14132), .ZN(n14133) );
  NAND2_X1 U17550 ( .A1(n14198), .A2(n14133), .ZN(n15921) );
  OAI22_X1 U17551 ( .A1(n14134), .A2(n20064), .B1(n20081), .B2(n15921), .ZN(
        n14137) );
  AOI22_X1 U17552 ( .A1(n20093), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n20102), 
        .B2(n15798), .ZN(n14135) );
  NAND2_X1 U17553 ( .A1(n20177), .A2(n14135), .ZN(n14136) );
  AOI211_X1 U17554 ( .C1(n14533), .C2(n14138), .A(n14137), .B(n14136), .ZN(
        n14139) );
  OAI21_X1 U17555 ( .B1(n14180), .B2(n20029), .A(n14139), .ZN(P1_U2826) );
  AOI22_X1 U17556 ( .A1(n14173), .A2(n14613), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14666), .ZN(n14140) );
  OAI21_X1 U17557 ( .B1(n14180), .B2(n14679), .A(n14140), .ZN(P1_U2890) );
  OAI21_X1 U17558 ( .B1(n9720), .B2(n11938), .A(n14142), .ZN(n14171) );
  OAI21_X1 U17559 ( .B1(n14171), .B2(n14172), .A(n14142), .ZN(n14161) );
  XNOR2_X1 U17560 ( .A(n14161), .B(n14160), .ZN(n15812) );
  OAI222_X1 U17561 ( .A1(n15812), .A2(n14679), .B1(n14218), .B2(n14618), .C1(
        n20119), .C2(n14670), .ZN(P1_U2892) );
  OAI21_X1 U17562 ( .B1(n14207), .B2(n14144), .A(n14143), .ZN(n19108) );
  AND2_X1 U17563 ( .A1(n14146), .A2(n14145), .ZN(n14148) );
  MUX2_X1 U17564 ( .A(n18939), .B(n14149), .S(n14907), .Z(n14150) );
  OAI21_X1 U17565 ( .B1(n19108), .B2(n14926), .A(n14150), .ZN(P2_U2871) );
  OR2_X1 U17566 ( .A1(n14237), .A2(n14151), .ZN(n14152) );
  NAND2_X1 U17567 ( .A1(n12510), .A2(n14152), .ZN(n15235) );
  OR2_X1 U17568 ( .A1(n14153), .A2(n14154), .ZN(n14156) );
  AND2_X1 U17569 ( .A1(n14156), .A2(n14155), .ZN(n16127) );
  NAND2_X1 U17570 ( .A1(n16127), .A2(n14939), .ZN(n14158) );
  NAND2_X1 U17571 ( .A1(n14884), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14157) );
  OAI211_X1 U17572 ( .C1(n15235), .C2(n14907), .A(n14158), .B(n14157), .ZN(
        P2_U2867) );
  AOI21_X1 U17573 ( .B1(n14161), .B2(n14160), .A(n14159), .ZN(n14162) );
  NOR2_X1 U17574 ( .A1(n14162), .A2(n14128), .ZN(n14781) );
  INV_X1 U17575 ( .A(n14781), .ZN(n15742) );
  AOI22_X1 U17576 ( .A1(n14173), .A2(n14401), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14666), .ZN(n14163) );
  OAI21_X1 U17577 ( .B1(n15742), .B2(n14679), .A(n14163), .ZN(P1_U2891) );
  AOI21_X1 U17578 ( .B1(n14165), .B2(n14169), .A(n14164), .ZN(n15933) );
  AOI22_X1 U17579 ( .A1(n15933), .A2(n14607), .B1(n14568), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14166) );
  OAI21_X1 U17580 ( .B1(n15742), .B2(n14595), .A(n14166), .ZN(P1_U2859) );
  NAND2_X1 U17581 ( .A1(n14175), .A2(n14167), .ZN(n14168) );
  NAND2_X1 U17582 ( .A1(n14169), .A2(n14168), .ZN(n15956) );
  INV_X1 U17583 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14170) );
  OAI222_X1 U17584 ( .A1(n15956), .A2(n14612), .B1(n14611), .B2(n14170), .C1(
        n14609), .C2(n15812), .ZN(P1_U2860) );
  XOR2_X1 U17585 ( .A(n14172), .B(n14171), .Z(n15816) );
  INV_X1 U17586 ( .A(n15816), .ZN(n14179) );
  AOI22_X1 U17587 ( .A1(n14173), .A2(n14623), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14666), .ZN(n14174) );
  OAI21_X1 U17588 ( .B1(n14179), .B2(n14679), .A(n14174), .ZN(P1_U2893) );
  OAI21_X1 U17589 ( .B1(n9742), .B2(n14176), .A(n14175), .ZN(n14177) );
  INV_X1 U17590 ( .A(n14177), .ZN(n15958) );
  AOI22_X1 U17591 ( .A1(n15958), .A2(n14607), .B1(n14568), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n14178) );
  OAI21_X1 U17592 ( .B1(n14179), .B2(n14609), .A(n14178), .ZN(P1_U2861) );
  INV_X1 U17593 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14181) );
  OAI222_X1 U17594 ( .A1(n15921), .A2(n14612), .B1(n14611), .B2(n14181), .C1(
        n14609), .C2(n14180), .ZN(P1_U2858) );
  NAND2_X1 U17595 ( .A1(n14186), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14185) );
  XNOR2_X1 U17596 ( .A(n14183), .B(n15976), .ZN(n14184) );
  MUX2_X1 U17597 ( .A(n14185), .B(n14184), .S(n9712), .Z(n14188) );
  NOR3_X1 U17598 ( .A1(n14186), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9712), .ZN(n15813) );
  INV_X1 U17599 ( .A(n15813), .ZN(n14187) );
  NAND2_X1 U17600 ( .A1(n14188), .A2(n14187), .ZN(n15974) );
  INV_X1 U17601 ( .A(n15974), .ZN(n14194) );
  AOI22_X1 U17602 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14189) );
  OAI21_X1 U17603 ( .B1(n20157), .B2(n14190), .A(n14189), .ZN(n14191) );
  AOI21_X1 U17604 ( .B1(n14192), .B2(n15799), .A(n14191), .ZN(n14193) );
  OAI21_X1 U17605 ( .B1(n14194), .B2(n20158), .A(n14193), .ZN(P1_U2989) );
  INV_X1 U17606 ( .A(n14195), .ZN(n14196) );
  AOI21_X1 U17607 ( .B1(n14197), .B2(n14127), .A(n14196), .ZN(n14232) );
  INV_X1 U17608 ( .A(n14232), .ZN(n14219) );
  NAND2_X1 U17609 ( .A1(n14412), .A2(n15756), .ZN(n14524) );
  NOR2_X1 U17610 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14524), .ZN(n14534) );
  AOI21_X1 U17611 ( .B1(n14199), .B2(n14198), .A(n9967), .ZN(n15909) );
  AOI22_X1 U17612 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(n20093), .B1(n20099), 
        .B2(n15909), .ZN(n14200) );
  OAI211_X1 U17613 ( .C1(n20064), .C2(n14201), .A(n14200), .B(n20177), .ZN(
        n14204) );
  NAND2_X1 U17614 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14533), .ZN(n14202) );
  OAI21_X1 U17615 ( .B1(n20088), .B2(n14230), .A(n14202), .ZN(n14203) );
  NOR3_X1 U17616 ( .A1(n14534), .A2(n14204), .A3(n14203), .ZN(n14205) );
  OAI21_X1 U17617 ( .B1(n14219), .B2(n20029), .A(n14205), .ZN(P1_U2825) );
  NAND2_X1 U17618 ( .A1(n14207), .A2(n14206), .ZN(n14239) );
  INV_X1 U17619 ( .A(n14239), .ZN(n14208) );
  AOI21_X1 U17620 ( .B1(n14210), .B2(n14209), .A(n14208), .ZN(n16132) );
  NAND2_X1 U17621 ( .A1(n16132), .A2(n14939), .ZN(n14212) );
  NAND2_X1 U17622 ( .A1(n14884), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14211) );
  OAI211_X1 U17623 ( .C1(n14213), .C2(n14884), .A(n14212), .B(n14211), .ZN(
        P2_U2869) );
  INV_X1 U17624 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14215) );
  INV_X1 U17625 ( .A(n15909), .ZN(n14214) );
  OAI222_X1 U17626 ( .A1(n14219), .A2(n14595), .B1(n14611), .B2(n14215), .C1(
        n14214), .C2(n14612), .ZN(P1_U2857) );
  OAI222_X1 U17627 ( .A1(n14219), .A2(n14679), .B1(n14218), .B2(n14217), .C1(
        n14670), .C2(n14216), .ZN(P1_U2889) );
  INV_X1 U17628 ( .A(n14937), .ZN(n14220) );
  AOI21_X1 U17629 ( .B1(n14221), .B2(n14155), .A(n14220), .ZN(n15012) );
  NAND2_X1 U17630 ( .A1(n15012), .A2(n14939), .ZN(n14223) );
  NAND2_X1 U17631 ( .A1(n14884), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14222) );
  OAI211_X1 U17632 ( .C1(n15101), .C2(n14907), .A(n14223), .B(n14222), .ZN(
        P2_U2866) );
  NAND2_X1 U17633 ( .A1(n15783), .A2(n14224), .ZN(n14228) );
  INV_X1 U17634 ( .A(n15781), .ZN(n14226) );
  NAND2_X1 U17635 ( .A1(n14226), .A2(n14225), .ZN(n14227) );
  XNOR2_X1 U17636 ( .A(n14228), .B(n14227), .ZN(n15910) );
  INV_X1 U17637 ( .A(n15910), .ZN(n14234) );
  AOI22_X1 U17638 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14229) );
  OAI21_X1 U17639 ( .B1(n20157), .B2(n14230), .A(n14229), .ZN(n14231) );
  AOI21_X1 U17640 ( .B1(n14232), .B2(n15799), .A(n14231), .ZN(n14233) );
  OAI21_X1 U17641 ( .B1(n14234), .B2(n20158), .A(n14233), .ZN(P1_U2984) );
  AND2_X1 U17642 ( .A1(n14236), .A2(n14235), .ZN(n14238) );
  OR2_X1 U17643 ( .A1(n14238), .A2(n14237), .ZN(n18901) );
  AOI21_X1 U17644 ( .B1(n14240), .B2(n14239), .A(n14153), .ZN(n15018) );
  NAND2_X1 U17645 ( .A1(n15018), .A2(n14939), .ZN(n14242) );
  NAND2_X1 U17646 ( .A1(n14884), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14241) );
  OAI211_X1 U17647 ( .C1(n18901), .C2(n14884), .A(n14242), .B(n14241), .ZN(
        P2_U2868) );
  INV_X1 U17648 ( .A(n18863), .ZN(n18813) );
  NAND2_X1 U17649 ( .A1(n14252), .A2(n18643), .ZN(n14243) );
  NAND2_X1 U17650 ( .A1(n18632), .A2(n14243), .ZN(n18641) );
  NOR2_X1 U17651 ( .A1(n18813), .A2(n18641), .ZN(n14251) );
  NOR2_X1 U17652 ( .A1(n16554), .A2(n18722), .ZN(n14247) );
  NAND2_X1 U17653 ( .A1(n18850), .A2(n17454), .ZN(n18691) );
  AOI21_X1 U17654 ( .B1(n14245), .B2(n18691), .A(n18848), .ZN(n17385) );
  AOI21_X1 U17655 ( .B1(n14247), .B2(n17385), .A(n14246), .ZN(n14249) );
  NAND2_X1 U17656 ( .A1(n15396), .A2(n18635), .ZN(n14248) );
  OAI221_X1 U17657 ( .B1(n18632), .B2(n17454), .C1(n18632), .C2(n16398), .A(
        n14247), .ZN(n15694) );
  NAND3_X1 U17658 ( .A1(n14249), .A2(n14248), .A3(n15694), .ZN(n18665) );
  NOR2_X1 U17659 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18803), .ZN(n18190) );
  NAND3_X1 U17660 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18801)
         );
  NOR2_X1 U17661 ( .A1(n18180), .A2(n18801), .ZN(n14250) );
  AOI211_X1 U17662 ( .C1(n18846), .C2(n18665), .A(n18190), .B(n14250), .ZN(
        n18832) );
  MUX2_X1 U17663 ( .A(n14251), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18832), .Z(P3_U3284) );
  NAND3_X1 U17664 ( .A1(n17180), .A2(n14252), .A3(n18643), .ZN(n18179) );
  NOR2_X1 U17665 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18179), .ZN(n14254) );
  NOR2_X1 U17666 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18853) );
  NOR2_X1 U17667 ( .A1(n18810), .A2(n18862), .ZN(n18177) );
  NOR2_X1 U17668 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18803), .ZN(
        n18826) );
  INV_X1 U17669 ( .A(n18826), .ZN(n18812) );
  OAI21_X1 U17670 ( .B1(n18853), .B2(n18177), .A(n18812), .ZN(n18189) );
  OAI21_X1 U17671 ( .B1(n14254), .B2(n18801), .A(n18231), .ZN(n18185) );
  INV_X1 U17672 ( .A(n18185), .ZN(n14255) );
  NAND2_X1 U17673 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17846) );
  INV_X1 U17674 ( .A(n17846), .ZN(n17667) );
  NAND2_X1 U17675 ( .A1(n18862), .A2(n18803), .ZN(n16549) );
  AND2_X1 U17676 ( .A1(n18813), .A2(n16549), .ZN(n18845) );
  NOR2_X1 U17677 ( .A1(n17667), .A2(n18845), .ZN(n15482) );
  AOI21_X1 U17678 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15482), .ZN(n15483) );
  NOR2_X1 U17679 ( .A1(n14255), .A2(n15483), .ZN(n14257) );
  NOR3_X1 U17680 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18849), .ZN(n18543) );
  NOR2_X1 U17681 ( .A1(n18803), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18230) );
  OR2_X1 U17682 ( .A1(n18230), .A2(n14255), .ZN(n15481) );
  OR2_X1 U17683 ( .A1(n18543), .A2(n15481), .ZN(n14256) );
  MUX2_X1 U17684 ( .A(n14257), .B(n14256), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  XNOR2_X1 U17685 ( .A(n15113), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14276) );
  OR2_X1 U17686 ( .A1(n14264), .A2(n14263), .ZN(n14862) );
  NAND2_X1 U17687 ( .A1(n14264), .A2(n14263), .ZN(n14265) );
  NAND2_X1 U17688 ( .A1(n15077), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n14271) );
  OAI21_X1 U17689 ( .B1(n18901), .B2(n16283), .A(n14271), .ZN(n14267) );
  NOR3_X1 U17690 ( .A1(n15319), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14266), .ZN(n15226) );
  AOI211_X1 U17691 ( .C1(n16281), .C2(n18902), .A(n14267), .B(n15226), .ZN(
        n14268) );
  OAI21_X1 U17692 ( .B1(n15228), .B2(n15112), .A(n14268), .ZN(n14269) );
  AOI21_X1 U17693 ( .B1(n14276), .B2(n16274), .A(n14269), .ZN(n14270) );
  OAI21_X1 U17694 ( .B1(n14278), .B2(n16315), .A(n14270), .ZN(P2_U3027) );
  OAI21_X1 U17695 ( .B1(n16239), .B2(n14272), .A(n14271), .ZN(n14273) );
  AOI21_X1 U17696 ( .B1(n18897), .B2(n16227), .A(n14273), .ZN(n14274) );
  OAI21_X1 U17697 ( .B1(n16214), .B2(n18901), .A(n14274), .ZN(n14275) );
  AOI21_X1 U17698 ( .B1(n14276), .B2(n19260), .A(n14275), .ZN(n14277) );
  OAI21_X1 U17699 ( .B1(n14278), .B2(n16220), .A(n14277), .ZN(P2_U2995) );
  INV_X1 U17700 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14279) );
  OAI22_X1 U17701 ( .A1(n14612), .A2(n20061), .B1(n14279), .B2(n14611), .ZN(
        n14280) );
  INV_X1 U17702 ( .A(n14280), .ZN(n14281) );
  OAI21_X1 U17703 ( .B1(n20068), .B2(n14595), .A(n14281), .ZN(P1_U2867) );
  MUX2_X1 U17704 ( .A(n9744), .B(n9779), .S(n9711), .Z(n14283) );
  XNOR2_X1 U17705 ( .A(n14283), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14298) );
  INV_X1 U17706 ( .A(n14284), .ZN(n14807) );
  NAND2_X1 U17707 ( .A1(n14469), .A2(n14285), .ZN(n14286) );
  NAND2_X1 U17708 ( .A1(n14453), .A2(n14286), .ZN(n14551) );
  NAND2_X1 U17709 ( .A1(n16000), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14293) );
  OAI21_X1 U17710 ( .B1(n14551), .B2(n20179), .A(n14293), .ZN(n14288) );
  NOR2_X1 U17711 ( .A1(n14802), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14287) );
  AOI211_X1 U17712 ( .C1(n14807), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14288), .B(n14287), .ZN(n14289) );
  OAI21_X1 U17713 ( .B1(n14298), .B2(n15988), .A(n14289), .ZN(P1_U3004) );
  INV_X1 U17714 ( .A(n14443), .ZN(n14291) );
  AOI21_X1 U17715 ( .B1(n14292), .B2(n14290), .A(n14291), .ZN(n14457) );
  NAND2_X1 U17716 ( .A1(n15809), .A2(n14460), .ZN(n14294) );
  OAI211_X1 U17717 ( .C1(n15837), .C2(n14295), .A(n14294), .B(n14293), .ZN(
        n14296) );
  AOI21_X1 U17718 ( .B1(n14457), .B2(n15799), .A(n14296), .ZN(n14297) );
  OAI21_X1 U17719 ( .B1(n20158), .B2(n14298), .A(n14297), .ZN(P1_U2972) );
  NAND2_X1 U17720 ( .A1(n14299), .A2(n15040), .ZN(n14302) );
  NOR2_X1 U17721 ( .A1(n14300), .A2(n9769), .ZN(n14301) );
  XNOR2_X1 U17722 ( .A(n14302), .B(n14301), .ZN(n15039) );
  NOR2_X1 U17723 ( .A1(n15157), .A2(n14305), .ZN(n14307) );
  OAI21_X1 U17724 ( .B1(n14307), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14306), .ZN(n14309) );
  NOR2_X1 U17725 ( .A1(n9722), .A2(n14308), .ZN(n15034) );
  NAND2_X1 U17726 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14310) );
  OAI211_X1 U17727 ( .C1(n19269), .C2(n14312), .A(n14311), .B(n14310), .ZN(
        n14313) );
  INV_X1 U17728 ( .A(n14313), .ZN(n14314) );
  OAI21_X1 U17729 ( .B1(n14317), .B2(n16220), .A(n14316), .ZN(P2_U2983) );
  NAND2_X1 U17730 ( .A1(n15061), .A2(n15063), .ZN(n14319) );
  XNOR2_X1 U17731 ( .A(n14318), .B(n14319), .ZN(n14340) );
  NOR2_X1 U17732 ( .A1(n15184), .A2(n14329), .ZN(n14327) );
  INV_X1 U17733 ( .A(n14903), .ZN(n14320) );
  AOI21_X1 U17734 ( .B1(n14321), .B2(n14920), .A(n14320), .ZN(n16093) );
  INV_X1 U17735 ( .A(n16093), .ZN(n14334) );
  NAND2_X1 U17736 ( .A1(n14322), .A2(n14323), .ZN(n14324) );
  NAND2_X1 U17737 ( .A1(n14978), .A2(n14324), .ZN(n16090) );
  INV_X1 U17738 ( .A(n16090), .ZN(n14991) );
  AOI22_X1 U17739 ( .A1(n16281), .A2(n14991), .B1(P2_REIP_REG_25__SCAN_IN), 
        .B2(n15077), .ZN(n14325) );
  OAI21_X1 U17740 ( .B1(n14334), .B2(n16283), .A(n14325), .ZN(n14326) );
  AOI211_X1 U17741 ( .C1(n15179), .C2(n14329), .A(n14327), .B(n14326), .ZN(
        n14333) );
  INV_X1 U17742 ( .A(n14328), .ZN(n14330) );
  NAND2_X1 U17743 ( .A1(n14330), .A2(n14329), .ZN(n14337) );
  NAND3_X1 U17744 ( .A1(n14337), .A2(n16274), .A3(n14331), .ZN(n14332) );
  OAI211_X1 U17745 ( .C1(n14340), .C2(n16315), .A(n14333), .B(n14332), .ZN(
        P2_U3021) );
  OAI22_X1 U17746 ( .A1(n16239), .A2(n16085), .B1(n19889), .B2(n9722), .ZN(
        n14336) );
  NOR2_X1 U17747 ( .A1(n14334), .A2(n16214), .ZN(n14335) );
  AOI211_X1 U17748 ( .C1(n16227), .C2(n16084), .A(n14336), .B(n14335), .ZN(
        n14339) );
  NAND3_X1 U17749 ( .A1(n14337), .A2(n19260), .A3(n14331), .ZN(n14338) );
  OAI211_X1 U17750 ( .C1(n14340), .C2(n16220), .A(n14339), .B(n14338), .ZN(
        P2_U2989) );
  OR2_X1 U17751 ( .A1(n14341), .A2(n13945), .ZN(n14343) );
  NAND2_X1 U17752 ( .A1(n14343), .A2(n14342), .ZN(n18977) );
  OAI211_X1 U17753 ( .C1(n14346), .C2(n14345), .A(n14344), .B(n14939), .ZN(
        n14348) );
  NAND2_X1 U17754 ( .A1(n14884), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14347) );
  OAI211_X1 U17755 ( .C1(n18977), .C2(n14907), .A(n14348), .B(n14347), .ZN(
        P2_U2875) );
  AOI21_X1 U17756 ( .B1(n20165), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14349), .ZN(n14350) );
  OAI21_X1 U17757 ( .B1(n20157), .B2(n14351), .A(n14350), .ZN(n14352) );
  AOI21_X1 U17758 ( .B1(n14411), .B2(n15799), .A(n14352), .ZN(n14353) );
  OAI21_X1 U17759 ( .B1(n14354), .B2(n20158), .A(n14353), .ZN(P1_U2968) );
  NAND2_X1 U17760 ( .A1(n9778), .A2(n14355), .ZN(n14356) );
  XNOR2_X1 U17761 ( .A(n14358), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14359) );
  XNOR2_X1 U17762 ( .A(n14360), .B(n14359), .ZN(n14376) );
  OAI21_X1 U17763 ( .B1(n15157), .B2(n14361), .A(n15167), .ZN(n15160) );
  INV_X1 U17764 ( .A(n15157), .ZN(n15174) );
  INV_X1 U17765 ( .A(n14361), .ZN(n15156) );
  NAND3_X1 U17766 ( .A1(n15174), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15156), .ZN(n14364) );
  INV_X1 U17767 ( .A(n14362), .ZN(n14962) );
  NOR2_X1 U17768 ( .A1(n9722), .A2(n19894), .ZN(n14368) );
  AOI21_X1 U17769 ( .B1(n16281), .B2(n14962), .A(n14368), .ZN(n14363) );
  OAI211_X1 U17770 ( .C1(n14890), .C2(n16283), .A(n14364), .B(n14363), .ZN(
        n14366) );
  NOR2_X1 U17771 ( .A1(n14371), .A2(n16307), .ZN(n14365) );
  OAI21_X1 U17772 ( .B1(n14376), .B2(n16315), .A(n14367), .ZN(P2_U3018) );
  INV_X1 U17773 ( .A(n14890), .ZN(n14374) );
  AOI21_X1 U17774 ( .B1(n19258), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14368), .ZN(n14369) );
  OAI21_X1 U17775 ( .B1(n19269), .B2(n14370), .A(n14369), .ZN(n14373) );
  NOR2_X1 U17776 ( .A1(n14371), .A2(n16219), .ZN(n14372) );
  OAI21_X1 U17777 ( .B1(n14376), .B2(n16220), .A(n14375), .ZN(P2_U2986) );
  AOI21_X1 U17778 ( .B1(n14379), .B2(n14378), .A(n14377), .ZN(n14391) );
  NAND2_X1 U17779 ( .A1(n15077), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n14393) );
  OAI21_X1 U17780 ( .B1(n14380), .B2(n14379), .A(n14393), .ZN(n14389) );
  OAI21_X1 U17781 ( .B1(n14383), .B2(n14382), .A(n14381), .ZN(n14384) );
  XNOR2_X1 U17782 ( .A(n14384), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14392) );
  AOI22_X1 U17783 ( .A1(n16301), .A2(n14392), .B1(n16281), .B2(n19941), .ZN(
        n14387) );
  OAI211_X1 U17784 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15247), .B(n14385), .ZN(n14386) );
  NAND2_X1 U17785 ( .A1(n14387), .A2(n14386), .ZN(n14388) );
  AOI211_X1 U17786 ( .C1(n16274), .C2(n14391), .A(n14389), .B(n14388), .ZN(
        n14390) );
  OAI21_X1 U17787 ( .B1(n14399), .B2(n16283), .A(n14390), .ZN(P2_U3045) );
  INV_X1 U17788 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14397) );
  INV_X1 U17789 ( .A(n14391), .ZN(n14395) );
  AOI22_X1 U17790 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19258), .B1(
        n19264), .B2(n14392), .ZN(n14394) );
  OAI211_X1 U17791 ( .C1(n16219), .C2(n14395), .A(n14394), .B(n14393), .ZN(
        n14396) );
  AOI21_X1 U17792 ( .B1(n16227), .B2(n14397), .A(n14396), .ZN(n14398) );
  OAI21_X1 U17793 ( .B1(n14399), .B2(n16214), .A(n14398), .ZN(P2_U3013) );
  INV_X1 U17794 ( .A(n14400), .ZN(n14433) );
  AOI22_X1 U17795 ( .A1(n14667), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14666), .ZN(n14403) );
  NOR3_X2 U17796 ( .A1(n14666), .A2(n20234), .A3(n12209), .ZN(n14676) );
  AOI22_X1 U17797 ( .A1(n14676), .A2(n14401), .B1(n14675), .B2(DATAI_29_), 
        .ZN(n14402) );
  OAI211_X1 U17798 ( .C1(n14400), .C2(n14679), .A(n14403), .B(n14402), .ZN(
        P1_U2875) );
  INV_X1 U17799 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14407) );
  OR2_X1 U17800 ( .A1(n14452), .A2(n14404), .ZN(n14405) );
  NAND2_X1 U17801 ( .A1(n14406), .A2(n14405), .ZN(n14793) );
  OAI222_X1 U17802 ( .A1(n14407), .A2(n14611), .B1(n14612), .B2(n14793), .C1(
        n14400), .C2(n14595), .ZN(P1_U2843) );
  NOR2_X1 U17803 ( .A1(n16047), .A2(n14907), .ZN(n14408) );
  AOI21_X1 U17804 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14907), .A(n14408), .ZN(
        n14409) );
  OAI21_X1 U17805 ( .B1(n14410), .B2(n14926), .A(n14409), .ZN(P2_U2857) );
  INV_X1 U17806 ( .A(n14411), .ZN(n14424) );
  INV_X1 U17807 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20824) );
  INV_X1 U17808 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20814) );
  NAND4_X1 U17809 ( .A1(n14412), .A2(P1_REIP_REG_17__SCAN_IN), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_15__SCAN_IN), .ZN(n14509) );
  NOR3_X1 U17810 ( .A1(n14414), .A2(n14413), .A3(n14509), .ZN(n14415) );
  NAND4_X1 U17811 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .A4(n14415), .ZN(n15705) );
  NOR2_X1 U17812 ( .A1(n20814), .A2(n15705), .ZN(n14499) );
  INV_X1 U17813 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20818) );
  INV_X1 U17814 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20817) );
  NOR2_X1 U17815 ( .A1(n20818), .A2(n20817), .ZN(n15706) );
  NAND4_X1 U17816 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n14499), .A4(n15706), .ZN(n15698) );
  NOR2_X1 U17817 ( .A1(n20824), .A2(n15698), .ZN(n14484) );
  NAND3_X1 U17818 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .A3(n14484), .ZN(n14461) );
  INV_X1 U17819 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14416) );
  NOR2_X1 U17820 ( .A1(n14461), .A2(n14416), .ZN(n14445) );
  NAND2_X1 U17821 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n14445), .ZN(n14446) );
  INV_X1 U17822 ( .A(n14446), .ZN(n14434) );
  AND2_X1 U17823 ( .A1(n14458), .A2(n14434), .ZN(n14417) );
  NOR2_X1 U17824 ( .A1(n20060), .A2(n14417), .ZN(n14451) );
  AOI21_X1 U17825 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(P1_REIP_REG_29__SCAN_IN), 
        .A(n20091), .ZN(n14418) );
  NOR2_X1 U17826 ( .A1(n14451), .A2(n14418), .ZN(n14427) );
  AOI22_X1 U17827 ( .A1(n20093), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20092), .ZN(n14420) );
  INV_X1 U17828 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20831) );
  NOR3_X1 U17829 ( .A1(n20091), .A2(n14446), .A3(n20831), .ZN(n14426) );
  NAND3_X1 U17830 ( .A1(n14426), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n14421), 
        .ZN(n14419) );
  OAI211_X1 U17831 ( .C1(n14427), .C2(n14421), .A(n14420), .B(n14419), .ZN(
        n14422) );
  AOI21_X1 U17832 ( .B1(n14546), .B2(n20099), .A(n14422), .ZN(n14423) );
  OAI21_X1 U17833 ( .B1(n14424), .B2(n20029), .A(n14423), .ZN(P1_U2809) );
  NAND2_X1 U17834 ( .A1(n14690), .A2(n20051), .ZN(n14432) );
  OAI22_X1 U17835 ( .A1(n14425), .A2(n20064), .B1(n20088), .B2(n14688), .ZN(
        n14430) );
  INV_X1 U17836 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14686) );
  INV_X1 U17837 ( .A(n14426), .ZN(n14428) );
  AOI21_X1 U17838 ( .B1(n14686), .B2(n14428), .A(n14427), .ZN(n14429) );
  AOI211_X1 U17839 ( .C1(n20093), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14430), .B(
        n14429), .ZN(n14431) );
  OAI211_X1 U17840 ( .C1(n20081), .C2(n14784), .A(n14432), .B(n14431), .ZN(
        P1_U2810) );
  NAND2_X1 U17841 ( .A1(n14433), .A2(n20051), .ZN(n14441) );
  NAND2_X1 U17842 ( .A1(n20831), .A2(n14434), .ZN(n14438) );
  AOI22_X1 U17843 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20092), .B1(
        n20102), .B2(n14435), .ZN(n14437) );
  NAND2_X1 U17844 ( .A1(n20093), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14436) );
  OAI211_X1 U17845 ( .C1(n20091), .C2(n14438), .A(n14437), .B(n14436), .ZN(
        n14439) );
  AOI21_X1 U17846 ( .B1(n14451), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14439), 
        .ZN(n14440) );
  OAI211_X1 U17847 ( .C1(n20081), .C2(n14793), .A(n14441), .B(n14440), .ZN(
        P1_U2811) );
  AOI21_X1 U17848 ( .B1(n14444), .B2(n14443), .A(n14442), .ZN(n14707) );
  INV_X1 U17849 ( .A(n14707), .ZN(n14622) );
  INV_X1 U17850 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14550) );
  INV_X1 U17851 ( .A(n20091), .ZN(n15696) );
  NAND3_X1 U17852 ( .A1(n15696), .A2(n14446), .A3(n14445), .ZN(n14449) );
  INV_X1 U17853 ( .A(n14705), .ZN(n14447) );
  AOI22_X1 U17854 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20092), .B1(
        n20102), .B2(n14447), .ZN(n14448) );
  OAI211_X1 U17855 ( .C1(n14550), .C2(n20024), .A(n14449), .B(n14448), .ZN(
        n14450) );
  AOI21_X1 U17856 ( .B1(n14451), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14450), 
        .ZN(n14456) );
  AOI21_X1 U17857 ( .B1(n14454), .B2(n14453), .A(n14452), .ZN(n14549) );
  NAND2_X1 U17858 ( .A1(n14549), .A2(n20099), .ZN(n14455) );
  OAI211_X1 U17859 ( .C1(n14622), .C2(n20029), .A(n14456), .B(n14455), .ZN(
        P1_U2812) );
  INV_X1 U17860 ( .A(n14457), .ZN(n14626) );
  INV_X1 U17861 ( .A(n14461), .ZN(n14459) );
  OAI21_X1 U17862 ( .B1(n20091), .B2(n14459), .A(n14458), .ZN(n14471) );
  INV_X1 U17863 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14552) );
  AOI22_X1 U17864 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20092), .B1(
        n20102), .B2(n14460), .ZN(n14463) );
  OR3_X1 U17865 ( .A1(n20091), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14461), .ZN(
        n14462) );
  OAI211_X1 U17866 ( .C1(n14552), .C2(n20024), .A(n14463), .B(n14462), .ZN(
        n14465) );
  NOR2_X1 U17867 ( .A1(n14551), .A2(n20081), .ZN(n14464) );
  AOI211_X1 U17868 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14471), .A(n14465), 
        .B(n14464), .ZN(n14466) );
  OAI21_X1 U17869 ( .B1(n14626), .B2(n20029), .A(n14466), .ZN(P1_U2813) );
  OAI21_X1 U17870 ( .B1(n14467), .B2(n14468), .A(n14290), .ZN(n14717) );
  OAI21_X1 U17871 ( .B1(n14481), .B2(n14470), .A(n14469), .ZN(n14553) );
  INV_X1 U17872 ( .A(n14553), .ZN(n14817) );
  INV_X1 U17873 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14554) );
  AND3_X1 U17874 ( .A1(n15696), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14484), 
        .ZN(n14472) );
  OAI21_X1 U17875 ( .B1(n14472), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14471), 
        .ZN(n14475) );
  INV_X1 U17876 ( .A(n14713), .ZN(n14473) );
  AOI22_X1 U17877 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20092), .B1(
        n20102), .B2(n14473), .ZN(n14474) );
  OAI211_X1 U17878 ( .C1(n14554), .C2(n20024), .A(n14475), .B(n14474), .ZN(
        n14476) );
  AOI21_X1 U17879 ( .B1(n14817), .B2(n20099), .A(n14476), .ZN(n14477) );
  OAI21_X1 U17880 ( .B1(n14717), .B2(n20029), .A(n14477), .ZN(P1_U2814) );
  INV_X1 U17881 ( .A(n14467), .ZN(n14479) );
  OAI21_X1 U17882 ( .B1(n14480), .B2(n14478), .A(n14479), .ZN(n14725) );
  OAI21_X1 U17883 ( .B1(n14500), .B2(n15698), .A(n15737), .ZN(n15707) );
  OAI21_X1 U17884 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n20091), .A(n15707), 
        .ZN(n14490) );
  AOI21_X1 U17885 ( .B1(n14482), .B2(n14561), .A(n14481), .ZN(n15841) );
  INV_X1 U17886 ( .A(n15841), .ZN(n14488) );
  INV_X1 U17887 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14483) );
  OAI22_X1 U17888 ( .A1(n14720), .A2(n20064), .B1(n14483), .B2(n20024), .ZN(
        n14486) );
  AND3_X1 U17889 ( .A1(n20826), .A2(n15696), .A3(n14484), .ZN(n14485) );
  AOI211_X1 U17890 ( .C1(n20102), .C2(n14722), .A(n14486), .B(n14485), .ZN(
        n14487) );
  OAI21_X1 U17891 ( .B1(n14488), .B2(n20081), .A(n14487), .ZN(n14489) );
  AOI21_X1 U17892 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n14490), .A(n14489), 
        .ZN(n14491) );
  OAI21_X1 U17893 ( .B1(n14725), .B2(n20029), .A(n14491), .ZN(P1_U2815) );
  INV_X1 U17894 ( .A(n14494), .ZN(n14598) );
  AND2_X1 U17895 ( .A1(n14494), .A2(n14493), .ZN(n14571) );
  AOI21_X1 U17896 ( .B1(n14495), .B2(n14586), .A(n14571), .ZN(n14742) );
  INV_X1 U17897 ( .A(n14742), .ZN(n14650) );
  NOR2_X1 U17898 ( .A1(n14589), .A2(n14496), .ZN(n14497) );
  OR2_X1 U17899 ( .A1(n14574), .A2(n14497), .ZN(n15656) );
  AOI22_X1 U17900 ( .A1(n20092), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20102), .B2(n14738), .ZN(n14498) );
  OAI21_X1 U17901 ( .B1(n15656), .B2(n20081), .A(n14498), .ZN(n14504) );
  NAND2_X1 U17902 ( .A1(n14499), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14501) );
  AOI21_X1 U17903 ( .B1(n15696), .B2(n14501), .A(n14500), .ZN(n15722) );
  INV_X1 U17904 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14580) );
  OAI22_X1 U17905 ( .A1(n15722), .A2(n20818), .B1(n14580), .B2(n20024), .ZN(
        n14503) );
  NOR3_X1 U17906 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n20091), .A3(n14501), 
        .ZN(n14502) );
  NOR3_X1 U17907 ( .A1(n14504), .A2(n14503), .A3(n14502), .ZN(n14505) );
  OAI21_X1 U17908 ( .B1(n14650), .B2(n20029), .A(n14505), .ZN(P1_U2819) );
  INV_X1 U17909 ( .A(n14584), .ZN(n14506) );
  AOI21_X1 U17910 ( .B1(n14507), .B2(n14598), .A(n14506), .ZN(n14748) );
  INV_X1 U17911 ( .A(n14748), .ZN(n14658) );
  NAND3_X1 U17912 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14508) );
  NOR3_X1 U17913 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14508), .A3(n14524), 
        .ZN(n15730) );
  INV_X1 U17914 ( .A(n14509), .ZN(n14510) );
  OAI21_X1 U17915 ( .B1(n14510), .B2(n20060), .A(n15759), .ZN(n15732) );
  OAI21_X1 U17916 ( .B1(n15730), .B2(n15732), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14518) );
  NAND2_X1 U17917 ( .A1(n14602), .A2(n14511), .ZN(n14512) );
  AND2_X1 U17918 ( .A1(n14588), .A2(n14512), .ZN(n15870) );
  NOR3_X1 U17919 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n20091), .A3(n15705), 
        .ZN(n14516) );
  AOI22_X1 U17920 ( .A1(n14747), .A2(n20102), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n20093), .ZN(n14513) );
  OAI211_X1 U17921 ( .C1(n20064), .C2(n14514), .A(n14513), .B(n20177), .ZN(
        n14515) );
  AOI211_X1 U17922 ( .C1(n20099), .C2(n15870), .A(n14516), .B(n14515), .ZN(
        n14517) );
  OAI211_X1 U17923 ( .C1(n14658), .C2(n20029), .A(n14518), .B(n14517), .ZN(
        P1_U2821) );
  INV_X1 U17924 ( .A(n14521), .ZN(n14522) );
  OAI21_X1 U17925 ( .B1(n14520), .B2(n14523), .A(n14522), .ZN(n14766) );
  INV_X1 U17926 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20808) );
  NOR2_X1 U17927 ( .A1(n20808), .A2(n14524), .ZN(n14532) );
  OAI221_X1 U17928 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), .C1(P1_REIP_REG_17__SCAN_IN), .C2(n14532), .A(n15732), .ZN(n14530) );
  AND2_X1 U17929 ( .A1(n14540), .A2(n14525), .ZN(n14526) );
  NOR2_X1 U17930 ( .A1(n14600), .A2(n14526), .ZN(n15892) );
  AOI22_X1 U17931 ( .A1(n14769), .A2(n20102), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n20093), .ZN(n14527) );
  OAI211_X1 U17932 ( .C1(n20064), .C2(n14765), .A(n14527), .B(n20177), .ZN(
        n14528) );
  AOI21_X1 U17933 ( .B1(n15892), .B2(n20099), .A(n14528), .ZN(n14529) );
  OAI211_X1 U17934 ( .C1(n14766), .C2(n20029), .A(n14530), .B(n14529), .ZN(
        P1_U2823) );
  AOI21_X1 U17935 ( .B1(n14531), .B2(n14195), .A(n14520), .ZN(n15786) );
  INV_X1 U17936 ( .A(n15786), .ZN(n14680) );
  INV_X1 U17937 ( .A(n14532), .ZN(n14536) );
  NOR2_X1 U17938 ( .A1(n14534), .A2(n14533), .ZN(n14535) );
  MUX2_X1 U17939 ( .A(n14536), .B(n14535), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n14545) );
  NAND2_X1 U17940 ( .A1(n14538), .A2(n14537), .ZN(n14539) );
  NAND2_X1 U17941 ( .A1(n14540), .A2(n14539), .ZN(n15907) );
  OAI22_X1 U17942 ( .A1(n15789), .A2(n20088), .B1(n20081), .B2(n15907), .ZN(
        n14543) );
  INV_X1 U17943 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14541) );
  OAI21_X1 U17944 ( .B1(n20064), .B2(n14541), .A(n20177), .ZN(n14542) );
  AOI211_X1 U17945 ( .C1(n20093), .C2(P1_EBX_REG_16__SCAN_IN), .A(n14543), .B(
        n14542), .ZN(n14544) );
  OAI211_X1 U17946 ( .C1(n14680), .C2(n20029), .A(n14545), .B(n14544), .ZN(
        P1_U2824) );
  INV_X1 U17947 ( .A(n14546), .ZN(n14548) );
  INV_X1 U17948 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14547) );
  OAI22_X1 U17949 ( .A1(n14548), .A2(n14612), .B1(n14547), .B2(n14611), .ZN(
        P1_U2841) );
  INV_X1 U17950 ( .A(n14549), .ZN(n14804) );
  OAI222_X1 U17951 ( .A1(n14550), .A2(n14611), .B1(n14612), .B2(n14804), .C1(
        n14622), .C2(n14609), .ZN(P1_U2844) );
  OAI222_X1 U17952 ( .A1(n14552), .A2(n14611), .B1(n14612), .B2(n14551), .C1(
        n14626), .C2(n14609), .ZN(P1_U2845) );
  OAI222_X1 U17953 ( .A1(n14554), .A2(n14611), .B1(n14612), .B2(n14553), .C1(
        n14717), .C2(n14609), .ZN(P1_U2846) );
  AOI22_X1 U17954 ( .A1(n15841), .A2(n14607), .B1(n14568), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14555) );
  OAI21_X1 U17955 ( .B1(n14725), .B2(n14609), .A(n14555), .ZN(P1_U2847) );
  AND2_X1 U17956 ( .A1(n14556), .A2(n14557), .ZN(n14558) );
  NOR2_X1 U17957 ( .A1(n14478), .A2(n14558), .ZN(n15763) );
  INV_X1 U17958 ( .A(n15763), .ZN(n14639) );
  INV_X1 U17959 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14562) );
  NAND2_X1 U17960 ( .A1(n14565), .A2(n14559), .ZN(n14560) );
  NAND2_X1 U17961 ( .A1(n14561), .A2(n14560), .ZN(n15853) );
  OAI222_X1 U17962 ( .A1(n14609), .A2(n14639), .B1(n14611), .B2(n14562), .C1(
        n14612), .C2(n15853), .ZN(P1_U2848) );
  INV_X1 U17963 ( .A(n14563), .ZN(n14564) );
  OAI21_X1 U17964 ( .B1(n14564), .B2(n10074), .A(n14556), .ZN(n15709) );
  INV_X1 U17965 ( .A(n14565), .ZN(n14566) );
  AOI21_X1 U17966 ( .B1(n14567), .B2(n14576), .A(n14566), .ZN(n15856) );
  AOI22_X1 U17967 ( .A1(n15856), .A2(n14607), .B1(n14568), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n14569) );
  OAI21_X1 U17968 ( .B1(n15709), .B2(n14609), .A(n14569), .ZN(P1_U2849) );
  OR2_X1 U17969 ( .A1(n14571), .A2(n14570), .ZN(n14572) );
  AND2_X1 U17970 ( .A1(n14572), .A2(n14563), .ZN(n15770) );
  OR2_X1 U17971 ( .A1(n14574), .A2(n14573), .ZN(n14575) );
  NAND2_X1 U17972 ( .A1(n14576), .A2(n14575), .ZN(n15868) );
  OAI22_X1 U17973 ( .A1(n15868), .A2(n14612), .B1(n14577), .B2(n14611), .ZN(
        n14578) );
  INV_X1 U17974 ( .A(n14578), .ZN(n14579) );
  OAI21_X1 U17975 ( .B1(n15714), .B2(n14595), .A(n14579), .ZN(P1_U2850) );
  OAI22_X1 U17976 ( .A1(n15656), .A2(n14612), .B1(n14580), .B2(n14611), .ZN(
        n14581) );
  INV_X1 U17977 ( .A(n14581), .ZN(n14582) );
  OAI21_X1 U17978 ( .B1(n14650), .B2(n14609), .A(n14582), .ZN(P1_U2851) );
  NAND2_X1 U17979 ( .A1(n14584), .A2(n14583), .ZN(n14585) );
  INV_X1 U17980 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14591) );
  AND2_X1 U17981 ( .A1(n14588), .A2(n14587), .ZN(n14590) );
  OR2_X1 U17982 ( .A1(n14590), .A2(n14589), .ZN(n15721) );
  OAI222_X1 U17983 ( .A1(n14609), .A2(n14655), .B1(n14611), .B2(n14591), .C1(
        n14612), .C2(n15721), .ZN(P1_U2852) );
  INV_X1 U17984 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14592) );
  NOR2_X1 U17985 ( .A1(n14611), .A2(n14592), .ZN(n14593) );
  AOI21_X1 U17986 ( .B1(n15870), .B2(n14607), .A(n14593), .ZN(n14594) );
  OAI21_X1 U17987 ( .B1(n14658), .B2(n14595), .A(n14594), .ZN(P1_U2853) );
  OR2_X1 U17988 ( .A1(n14521), .A2(n14596), .ZN(n14597) );
  OR2_X1 U17989 ( .A1(n14600), .A2(n14599), .ZN(n14601) );
  NAND2_X1 U17990 ( .A1(n14602), .A2(n14601), .ZN(n15882) );
  OAI22_X1 U17991 ( .A1(n15882), .A2(n14612), .B1(n15728), .B2(n14611), .ZN(
        n14603) );
  INV_X1 U17992 ( .A(n14603), .ZN(n14604) );
  OAI21_X1 U17993 ( .B1(n14665), .B2(n14609), .A(n14604), .ZN(P1_U2854) );
  INV_X1 U17994 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14605) );
  NOR2_X1 U17995 ( .A1(n14611), .A2(n14605), .ZN(n14606) );
  AOI21_X1 U17996 ( .B1(n15892), .B2(n14607), .A(n14606), .ZN(n14608) );
  OAI21_X1 U17997 ( .B1(n14766), .B2(n14609), .A(n14608), .ZN(P1_U2855) );
  INV_X1 U17998 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14610) );
  OAI222_X1 U17999 ( .A1(n15907), .A2(n14612), .B1(n14611), .B2(n14610), .C1(
        n14609), .C2(n14680), .ZN(P1_U2856) );
  AOI22_X1 U18000 ( .A1(n14667), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14666), .ZN(n14615) );
  AOI22_X1 U18001 ( .A1(n14676), .A2(n14613), .B1(n14675), .B2(DATAI_30_), 
        .ZN(n14614) );
  OAI211_X1 U18002 ( .C1(n14616), .C2(n14679), .A(n14615), .B(n14614), .ZN(
        P1_U2874) );
  INV_X1 U18003 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16466) );
  NOR2_X1 U18004 ( .A1(n14673), .A2(n16466), .ZN(n14620) );
  INV_X1 U18005 ( .A(n14676), .ZN(n14661) );
  INV_X1 U18006 ( .A(n14675), .ZN(n14617) );
  OAI22_X1 U18007 ( .A1(n14661), .A2(n14618), .B1(n14617), .B2(n10337), .ZN(
        n14619) );
  AOI211_X1 U18008 ( .C1(n14666), .C2(P1_EAX_REG_28__SCAN_IN), .A(n14620), .B(
        n14619), .ZN(n14621) );
  OAI21_X1 U18009 ( .B1(n14622), .B2(n14679), .A(n14621), .ZN(P1_U2876) );
  AOI22_X1 U18010 ( .A1(n14667), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14666), .ZN(n14625) );
  AOI22_X1 U18011 ( .A1(n14676), .A2(n14623), .B1(n14675), .B2(DATAI_27_), 
        .ZN(n14624) );
  OAI211_X1 U18012 ( .C1(n14626), .C2(n14679), .A(n14625), .B(n14624), .ZN(
        P1_U2877) );
  INV_X1 U18013 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16470) );
  OAI22_X1 U18014 ( .A1(n14673), .A2(n16470), .B1(n14627), .B2(n14670), .ZN(
        n14628) );
  INV_X1 U18015 ( .A(n14628), .ZN(n14631) );
  AOI22_X1 U18016 ( .A1(n14676), .A2(n14629), .B1(n14675), .B2(DATAI_26_), 
        .ZN(n14630) );
  OAI211_X1 U18017 ( .C1(n14717), .C2(n14679), .A(n14631), .B(n14630), .ZN(
        P1_U2878) );
  AOI22_X1 U18018 ( .A1(n14667), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14666), .ZN(n14634) );
  AOI22_X1 U18019 ( .A1(n14676), .A2(n14632), .B1(n14675), .B2(DATAI_25_), 
        .ZN(n14633) );
  OAI211_X1 U18020 ( .C1(n14725), .C2(n14679), .A(n14634), .B(n14633), .ZN(
        P1_U2879) );
  INV_X1 U18021 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16475) );
  OAI22_X1 U18022 ( .A1(n14673), .A2(n16475), .B1(n13636), .B2(n14670), .ZN(
        n14635) );
  INV_X1 U18023 ( .A(n14635), .ZN(n14638) );
  AOI22_X1 U18024 ( .A1(n14676), .A2(n14636), .B1(n14675), .B2(DATAI_24_), 
        .ZN(n14637) );
  OAI211_X1 U18025 ( .C1(n14639), .C2(n14679), .A(n14638), .B(n14637), .ZN(
        P1_U2880) );
  AOI22_X1 U18026 ( .A1(n14667), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14666), .ZN(n14641) );
  AOI22_X1 U18027 ( .A1(n14676), .A2(n20237), .B1(n14675), .B2(DATAI_23_), 
        .ZN(n14640) );
  OAI211_X1 U18028 ( .C1(n15709), .C2(n14679), .A(n14641), .B(n14640), .ZN(
        P1_U2881) );
  INV_X1 U18029 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14643) );
  OAI22_X1 U18030 ( .A1(n14673), .A2(n14643), .B1(n14642), .B2(n14670), .ZN(
        n14645) );
  NOR2_X1 U18031 ( .A1(n14661), .A2(n20229), .ZN(n14644) );
  AOI211_X1 U18032 ( .C1(n14675), .C2(DATAI_22_), .A(n14645), .B(n14644), .ZN(
        n14646) );
  OAI21_X1 U18033 ( .B1(n15714), .B2(n14679), .A(n14646), .ZN(P1_U2882) );
  AOI22_X1 U18034 ( .A1(n14667), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14666), .ZN(n14649) );
  AOI22_X1 U18035 ( .A1(n14676), .A2(n14647), .B1(n14675), .B2(DATAI_21_), 
        .ZN(n14648) );
  OAI211_X1 U18036 ( .C1(n14650), .C2(n14679), .A(n14649), .B(n14648), .ZN(
        P1_U2883) );
  INV_X1 U18037 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16480) );
  OAI22_X1 U18038 ( .A1(n14673), .A2(n16480), .B1(n14651), .B2(n14670), .ZN(
        n14653) );
  NOR2_X1 U18039 ( .A1(n14661), .A2(n20222), .ZN(n14652) );
  AOI211_X1 U18040 ( .C1(n14675), .C2(DATAI_20_), .A(n14653), .B(n14652), .ZN(
        n14654) );
  OAI21_X1 U18041 ( .B1(n14655), .B2(n14679), .A(n14654), .ZN(P1_U2884) );
  AOI22_X1 U18042 ( .A1(n14667), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14666), .ZN(n14657) );
  AOI22_X1 U18043 ( .A1(n14676), .A2(n20218), .B1(n14675), .B2(DATAI_19_), 
        .ZN(n14656) );
  OAI211_X1 U18044 ( .C1(n14658), .C2(n14679), .A(n14657), .B(n14656), .ZN(
        P1_U2885) );
  INV_X1 U18045 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14660) );
  OAI22_X1 U18046 ( .A1(n14673), .A2(n14660), .B1(n14659), .B2(n14670), .ZN(
        n14663) );
  NOR2_X1 U18047 ( .A1(n14661), .A2(n20214), .ZN(n14662) );
  AOI211_X1 U18048 ( .C1(n14675), .C2(DATAI_18_), .A(n14663), .B(n14662), .ZN(
        n14664) );
  OAI21_X1 U18049 ( .B1(n14665), .B2(n14679), .A(n14664), .ZN(P1_U2886) );
  AOI22_X1 U18050 ( .A1(n14667), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14666), .ZN(n14669) );
  AOI22_X1 U18051 ( .A1(n14676), .A2(n20210), .B1(n14675), .B2(DATAI_17_), 
        .ZN(n14668) );
  OAI211_X1 U18052 ( .C1(n14766), .C2(n14679), .A(n14669), .B(n14668), .ZN(
        P1_U2887) );
  INV_X1 U18053 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14672) );
  OAI22_X1 U18054 ( .A1(n14673), .A2(n14672), .B1(n14671), .B2(n14670), .ZN(
        n14674) );
  INV_X1 U18055 ( .A(n14674), .ZN(n14678) );
  AOI22_X1 U18056 ( .A1(n14676), .A2(n20203), .B1(n14675), .B2(DATAI_16_), 
        .ZN(n14677) );
  OAI211_X1 U18057 ( .C1(n14680), .C2(n14679), .A(n14678), .B(n14677), .ZN(
        P1_U2888) );
  NOR2_X1 U18058 ( .A1(n14681), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14684) );
  NOR2_X1 U18059 ( .A1(n14682), .A2(n12756), .ZN(n14683) );
  MUX2_X1 U18060 ( .A(n14684), .B(n14683), .S(n9712), .Z(n14685) );
  XNOR2_X1 U18061 ( .A(n14685), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14791) );
  NOR2_X1 U18062 ( .A1(n20177), .A2(n14686), .ZN(n14785) );
  AOI21_X1 U18063 ( .B1(n20165), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14785), .ZN(n14687) );
  OAI21_X1 U18064 ( .B1(n20157), .B2(n14688), .A(n14687), .ZN(n14689) );
  AOI21_X1 U18065 ( .B1(n14690), .B2(n15799), .A(n14689), .ZN(n14691) );
  OAI21_X1 U18066 ( .B1(n20158), .B2(n14791), .A(n14691), .ZN(P1_U2969) );
  INV_X1 U18067 ( .A(n14727), .ZN(n14694) );
  INV_X1 U18068 ( .A(n14693), .ZN(n14812) );
  NOR2_X1 U18069 ( .A1(n10011), .A2(n14812), .ZN(n14710) );
  NOR3_X1 U18070 ( .A1(n14695), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14696) );
  MUX2_X1 U18071 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14697), .S(
        n9711), .Z(n14698) );
  NAND2_X1 U18072 ( .A1(n16000), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14803) );
  NAND2_X1 U18073 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14704) );
  OAI211_X1 U18074 ( .C1(n20157), .C2(n14705), .A(n14803), .B(n14704), .ZN(
        n14706) );
  AOI21_X1 U18075 ( .B1(n14707), .B2(n15799), .A(n14706), .ZN(n14708) );
  OAI21_X1 U18076 ( .B1(n20158), .B2(n14809), .A(n14708), .ZN(P1_U2971) );
  AOI21_X1 U18077 ( .B1(n9711), .B2(n14727), .A(n14709), .ZN(n14711) );
  NOR2_X1 U18078 ( .A1(n14711), .A2(n14710), .ZN(n14712) );
  XOR2_X1 U18079 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14712), .Z(
        n14810) );
  NAND2_X1 U18080 ( .A1(n14810), .A2(n20167), .ZN(n14716) );
  INV_X1 U18081 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20828) );
  NOR2_X1 U18082 ( .A1(n20177), .A2(n20828), .ZN(n14816) );
  NOR2_X1 U18083 ( .A1(n20157), .A2(n14713), .ZN(n14714) );
  AOI211_X1 U18084 ( .C1(n20165), .C2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14816), .B(n14714), .ZN(n14715) );
  OAI211_X1 U18085 ( .C1(n20191), .C2(n14717), .A(n14716), .B(n14715), .ZN(
        P1_U2973) );
  NOR2_X1 U18086 ( .A1(n14727), .A2(n9712), .ZN(n15761) );
  INV_X1 U18087 ( .A(n15761), .ZN(n14731) );
  NAND2_X1 U18088 ( .A1(n14718), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15760) );
  NAND2_X1 U18089 ( .A1(n15840), .A2(n20167), .ZN(n14724) );
  OAI22_X1 U18090 ( .A1(n15837), .A2(n14720), .B1(n20177), .B2(n20826), .ZN(
        n14721) );
  AOI21_X1 U18091 ( .B1(n15809), .B2(n14722), .A(n14721), .ZN(n14723) );
  OAI211_X1 U18092 ( .C1(n20191), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        P1_U2974) );
  NAND2_X1 U18093 ( .A1(n9711), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14729) );
  INV_X1 U18094 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14726) );
  MUX2_X1 U18095 ( .A(n14726), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .S(
        n9711), .Z(n14728) );
  MUX2_X1 U18096 ( .A(n14729), .B(n14728), .S(n14727), .Z(n14730) );
  OAI21_X1 U18097 ( .B1(n14731), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14730), .ZN(n15857) );
  NAND2_X1 U18098 ( .A1(n15857), .A2(n20167), .ZN(n14735) );
  INV_X1 U18099 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14732) );
  OAI22_X1 U18100 ( .A1(n15837), .A2(n15713), .B1(n20177), .B2(n14732), .ZN(
        n14733) );
  AOI21_X1 U18101 ( .B1(n15809), .B2(n15704), .A(n14733), .ZN(n14734) );
  OAI211_X1 U18102 ( .C1(n20191), .C2(n15709), .A(n14735), .B(n14734), .ZN(
        P1_U2976) );
  NAND2_X1 U18103 ( .A1(n9775), .A2(n9711), .ZN(n15678) );
  AOI22_X1 U18104 ( .A1(n15678), .A2(n14736), .B1(n9712), .B2(n15679), .ZN(
        n14737) );
  XNOR2_X1 U18105 ( .A(n14737), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15655) );
  INV_X1 U18106 ( .A(n14738), .ZN(n14740) );
  AOI22_X1 U18107 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n14739) );
  OAI21_X1 U18108 ( .B1(n20157), .B2(n14740), .A(n14739), .ZN(n14741) );
  AOI21_X1 U18109 ( .B1(n14742), .B2(n15799), .A(n14741), .ZN(n14743) );
  OAI21_X1 U18110 ( .B1(n20158), .B2(n15655), .A(n14743), .ZN(P1_U2978) );
  OR2_X1 U18111 ( .A1(n14744), .A2(n14751), .ZN(n14752) );
  MUX2_X1 U18112 ( .A(n9757), .B(n15675), .S(n14752), .Z(n14745) );
  XNOR2_X1 U18113 ( .A(n14745), .B(n15874), .ZN(n15869) );
  OAI22_X1 U18114 ( .A1(n15837), .A2(n14514), .B1(n20177), .B2(n20814), .ZN(
        n14746) );
  AOI21_X1 U18115 ( .B1(n15809), .B2(n14747), .A(n14746), .ZN(n14750) );
  NAND2_X1 U18116 ( .A1(n14748), .A2(n15799), .ZN(n14749) );
  OAI211_X1 U18117 ( .C1(n15869), .C2(n20158), .A(n14750), .B(n14749), .ZN(
        P1_U2980) );
  INV_X1 U18118 ( .A(n14744), .ZN(n14754) );
  INV_X1 U18119 ( .A(n14751), .ZN(n14753) );
  OAI21_X1 U18120 ( .B1(n14754), .B2(n14753), .A(n14752), .ZN(n15883) );
  INV_X1 U18121 ( .A(n15731), .ZN(n14756) );
  AOI22_X1 U18122 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14755) );
  OAI21_X1 U18123 ( .B1(n20157), .B2(n14756), .A(n14755), .ZN(n14757) );
  AOI21_X1 U18124 ( .B1(n15733), .B2(n15799), .A(n14757), .ZN(n14758) );
  OAI21_X1 U18125 ( .B1(n15883), .B2(n20158), .A(n14758), .ZN(P1_U2981) );
  INV_X1 U18126 ( .A(n14759), .ZN(n14760) );
  NOR3_X1 U18127 ( .A1(n14760), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15780), .ZN(n14762) );
  OAI21_X1 U18128 ( .B1(n14762), .B2(n9712), .A(n14761), .ZN(n14763) );
  XOR2_X1 U18129 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n14763), .Z(
        n15891) );
  INV_X1 U18130 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14764) );
  OAI22_X1 U18131 ( .A1(n15837), .A2(n14765), .B1(n20177), .B2(n14764), .ZN(
        n14768) );
  NOR2_X1 U18132 ( .A1(n14766), .A2(n20191), .ZN(n14767) );
  AOI211_X1 U18133 ( .C1(n15809), .C2(n14769), .A(n14768), .B(n14767), .ZN(
        n14770) );
  OAI21_X1 U18134 ( .B1(n20158), .B2(n15891), .A(n14770), .ZN(P1_U2982) );
  INV_X1 U18135 ( .A(n14183), .ZN(n14774) );
  INV_X1 U18136 ( .A(n14771), .ZN(n14772) );
  AOI21_X1 U18137 ( .B1(n14774), .B2(n14773), .A(n14772), .ZN(n15807) );
  OAI211_X1 U18138 ( .C1(n14775), .C2(n9712), .A(n15807), .B(n15803), .ZN(
        n15805) );
  NAND2_X1 U18139 ( .A1(n15805), .A2(n15803), .ZN(n14777) );
  XNOR2_X1 U18140 ( .A(n14777), .B(n14776), .ZN(n15934) );
  INV_X1 U18141 ( .A(n15934), .ZN(n14783) );
  INV_X1 U18142 ( .A(n15745), .ZN(n14779) );
  AOI22_X1 U18143 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14778) );
  OAI21_X1 U18144 ( .B1(n20157), .B2(n14779), .A(n14778), .ZN(n14780) );
  AOI21_X1 U18145 ( .B1(n14781), .B2(n15799), .A(n14780), .ZN(n14782) );
  OAI21_X1 U18146 ( .B1(n14783), .B2(n20158), .A(n14782), .ZN(P1_U2986) );
  INV_X1 U18147 ( .A(n14784), .ZN(n14786) );
  AOI21_X1 U18148 ( .B1(n14786), .B2(n15999), .A(n14785), .ZN(n14790) );
  OAI21_X1 U18149 ( .B1(n14788), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14787), .ZN(n14789) );
  OAI211_X1 U18150 ( .C1(n14791), .C2(n15988), .A(n14790), .B(n14789), .ZN(
        P1_U3001) );
  OAI21_X1 U18151 ( .B1(n14793), .B2(n20179), .A(n14792), .ZN(n14796) );
  NOR3_X1 U18152 ( .A1(n14802), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14794), .ZN(n14795) );
  AOI211_X1 U18153 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14797), .A(
        n14796), .B(n14795), .ZN(n14798) );
  OAI21_X1 U18154 ( .B1(n14799), .B2(n15988), .A(n14798), .ZN(P1_U3002) );
  NOR3_X1 U18155 ( .A1(n14802), .A2(n14801), .A3(n14800), .ZN(n14806) );
  OAI21_X1 U18156 ( .B1(n14804), .B2(n20179), .A(n14803), .ZN(n14805) );
  AOI211_X1 U18157 ( .C1(n14807), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14806), .B(n14805), .ZN(n14808) );
  OAI21_X1 U18158 ( .B1(n14809), .B2(n15988), .A(n14808), .ZN(P1_U3003) );
  INV_X1 U18159 ( .A(n14810), .ZN(n14819) );
  NAND4_X1 U18160 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n15846), .A4(n12813), .ZN(
        n15843) );
  INV_X1 U18161 ( .A(n14811), .ZN(n14814) );
  AOI21_X1 U18162 ( .B1(n15846), .B2(n14812), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14813) );
  AOI21_X1 U18163 ( .B1(n15843), .B2(n14814), .A(n14813), .ZN(n14815) );
  AOI211_X1 U18164 ( .C1(n15999), .C2(n14817), .A(n14816), .B(n14815), .ZN(
        n14818) );
  OAI21_X1 U18165 ( .B1(n14819), .B2(n15988), .A(n14818), .ZN(P1_U3005) );
  OAI21_X1 U18166 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9717), .A(n20556), 
        .ZN(n14820) );
  OAI21_X1 U18167 ( .B1(n14823), .B2(n20392), .A(n14820), .ZN(n14821) );
  MUX2_X1 U18168 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14821), .S(
        n20187), .Z(P1_U3477) );
  INV_X1 U18169 ( .A(n20193), .ZN(n14822) );
  OR2_X1 U18170 ( .A1(n20192), .A2(n11800), .ZN(n20704) );
  NOR2_X1 U18171 ( .A1(n20704), .A2(n9717), .ZN(n20580) );
  AOI211_X1 U18172 ( .C1(n14822), .C2(n20633), .A(n20580), .B(n20553), .ZN(
        n14827) );
  INV_X1 U18173 ( .A(n14823), .ZN(n14825) );
  INV_X1 U18174 ( .A(n11800), .ZN(n14824) );
  NOR2_X1 U18175 ( .A1(n20427), .A2(n20703), .ZN(n20424) );
  AOI21_X1 U18176 ( .B1(n13653), .B2(n14825), .A(n20424), .ZN(n14826) );
  OAI21_X1 U18177 ( .B1(n14827), .B2(n20698), .A(n14826), .ZN(n14828) );
  MUX2_X1 U18178 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n14828), .S(
        n20187), .Z(P1_U3475) );
  NOR3_X1 U18179 ( .A1(n14829), .A2(n14834), .A3(n13673), .ZN(n14830) );
  AOI21_X1 U18180 ( .B1(n15612), .B2(n14831), .A(n14830), .ZN(n14832) );
  OAI21_X1 U18181 ( .B1(n20392), .B2(n14833), .A(n14832), .ZN(n15613) );
  INV_X1 U18182 ( .A(n15613), .ZN(n14838) );
  AOI22_X1 U18183 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13589), .B2(n12760), .ZN(
        n14843) );
  INV_X1 U18184 ( .A(n14843), .ZN(n14836) );
  NOR2_X1 U18185 ( .A1(n20760), .A2(n20172), .ZN(n14842) );
  NOR3_X1 U18186 ( .A1(n13673), .A2(n14834), .A3(n14848), .ZN(n14835) );
  AOI21_X1 U18187 ( .B1(n14836), .B2(n14842), .A(n14835), .ZN(n14837) );
  OAI21_X1 U18188 ( .B1(n14838), .B2(n14850), .A(n14837), .ZN(n14839) );
  MUX2_X1 U18189 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14839), .S(
        n16011), .Z(P1_U3473) );
  AOI22_X1 U18190 ( .A1(n14843), .A2(n14842), .B1(n14841), .B2(n14840), .ZN(
        n14844) );
  OAI21_X1 U18191 ( .B1(n14845), .B2(n14850), .A(n14844), .ZN(n14846) );
  MUX2_X1 U18192 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14846), .S(
        n16011), .Z(P1_U3472) );
  INV_X1 U18193 ( .A(n14847), .ZN(n14849) );
  OAI22_X1 U18194 ( .A1(n14851), .A2(n14850), .B1(n14849), .B2(n14848), .ZN(
        n14852) );
  MUX2_X1 U18195 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14852), .S(
        n16011), .Z(P1_U3469) );
  AOI211_X1 U18196 ( .C1(n15099), .C2(n14865), .A(n14853), .B(n19825), .ZN(
        n14855) );
  OAI22_X1 U18197 ( .A1(n19883), .A2(n19034), .B1(n15097), .B2(n19079), .ZN(
        n14854) );
  AOI211_X1 U18198 ( .C1(P2_EBX_REG_21__SCAN_IN), .C2(n19058), .A(n14855), .B(
        n14854), .ZN(n14860) );
  INV_X1 U18199 ( .A(n15013), .ZN(n14856) );
  OAI22_X1 U18200 ( .A1(n15101), .A2(n19075), .B1(n14856), .B2(n19083), .ZN(
        n14857) );
  AOI21_X1 U18201 ( .B1(n14858), .B2(n19086), .A(n14857), .ZN(n14859) );
  NAND2_X1 U18202 ( .A1(n14860), .A2(n14859), .ZN(P2_U2834) );
  AND2_X1 U18203 ( .A1(n14862), .A2(n14861), .ZN(n14863) );
  OR2_X1 U18204 ( .A1(n14864), .A2(n14863), .ZN(n16125) );
  OAI211_X1 U18205 ( .C1(n15117), .C2(n14866), .A(n14865), .B(n19055), .ZN(
        n14867) );
  OAI21_X1 U18206 ( .B1(n19083), .B2(n16125), .A(n14867), .ZN(n14872) );
  AOI22_X1 U18207 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19081), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9707), .ZN(n14870) );
  AOI22_X1 U18208 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19058), .B1(n14868), 
        .B2(n18947), .ZN(n14869) );
  OAI211_X1 U18209 ( .C1(n15235), .C2(n19075), .A(n14870), .B(n14869), .ZN(
        n14871) );
  AOI211_X1 U18210 ( .C1(n19086), .C2(n14873), .A(n14872), .B(n14871), .ZN(
        n14874) );
  INV_X1 U18211 ( .A(n14874), .ZN(P2_U2835) );
  NAND2_X1 U18212 ( .A1(n9974), .A2(n14936), .ZN(n14875) );
  OAI21_X1 U18213 ( .B1(n14936), .B2(n14876), .A(n14875), .ZN(P2_U2856) );
  OR2_X1 U18214 ( .A1(n13221), .A2(n14877), .ZN(n14878) );
  OR2_X1 U18215 ( .A1(n14880), .A2(n14879), .ZN(n14946) );
  NAND3_X1 U18216 ( .A1(n14946), .A2(n14881), .A3(n14939), .ZN(n14883) );
  NAND2_X1 U18217 ( .A1(n14884), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14882) );
  OAI211_X1 U18218 ( .C1(n14884), .C2(n16058), .A(n14883), .B(n14882), .ZN(
        P2_U2858) );
  INV_X1 U18219 ( .A(n14885), .ZN(n14886) );
  NAND2_X1 U18220 ( .A1(n14887), .A2(n14886), .ZN(n14889) );
  XNOR2_X1 U18221 ( .A(n14889), .B(n14888), .ZN(n14965) );
  NOR2_X1 U18222 ( .A1(n14890), .A2(n14907), .ZN(n14891) );
  AOI21_X1 U18223 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14907), .A(n14891), .ZN(
        n14892) );
  OAI21_X1 U18224 ( .B1(n14965), .B2(n14926), .A(n14892), .ZN(P2_U2859) );
  OAI21_X1 U18225 ( .B1(n14895), .B2(n14894), .A(n14893), .ZN(n14976) );
  NOR2_X1 U18226 ( .A1(n14904), .A2(n14896), .ZN(n14897) );
  MUX2_X1 U18227 ( .A(n16068), .B(n10231), .S(n14907), .Z(n14898) );
  OAI21_X1 U18228 ( .B1(n14976), .B2(n14926), .A(n14898), .ZN(P2_U2860) );
  OAI21_X1 U18229 ( .B1(n14901), .B2(n14900), .A(n14899), .ZN(n14985) );
  AND2_X1 U18230 ( .A1(n14903), .A2(n14902), .ZN(n14905) );
  OR2_X1 U18231 ( .A1(n14905), .A2(n14904), .ZN(n16077) );
  NOR2_X1 U18232 ( .A1(n16077), .A2(n14907), .ZN(n14906) );
  AOI21_X1 U18233 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n14907), .A(n14906), .ZN(
        n14908) );
  OAI21_X1 U18234 ( .B1(n14985), .B2(n14926), .A(n14908), .ZN(P2_U2861) );
  OAI21_X1 U18235 ( .B1(n14911), .B2(n14910), .A(n14909), .ZN(n14994) );
  NOR2_X1 U18236 ( .A1(n14936), .A2(n14912), .ZN(n14913) );
  AOI21_X1 U18237 ( .B1(n16093), .B2(n14936), .A(n14913), .ZN(n14914) );
  OAI21_X1 U18238 ( .B1(n14994), .B2(n14926), .A(n14914), .ZN(P2_U2862) );
  INV_X1 U18239 ( .A(n14915), .ZN(n14917) );
  AOI21_X1 U18240 ( .B1(n14917), .B2(n14916), .A(n9776), .ZN(n14918) );
  XOR2_X1 U18241 ( .A(n14919), .B(n14918), .Z(n15003) );
  INV_X1 U18242 ( .A(n14920), .ZN(n14921) );
  AOI21_X1 U18243 ( .B1(n14922), .B2(n14933), .A(n14921), .ZN(n16096) );
  NOR2_X1 U18244 ( .A1(n14936), .A2(n14923), .ZN(n14924) );
  AOI21_X1 U18245 ( .B1(n16096), .B2(n14936), .A(n14924), .ZN(n14925) );
  OAI21_X1 U18246 ( .B1(n15003), .B2(n14926), .A(n14925), .ZN(P2_U2863) );
  INV_X1 U18247 ( .A(n14927), .ZN(n14928) );
  AOI21_X1 U18248 ( .B1(n14930), .B2(n14929), .A(n14928), .ZN(n15010) );
  NAND2_X1 U18249 ( .A1(n15010), .A2(n14939), .ZN(n14935) );
  OR2_X1 U18250 ( .A1(n9783), .A2(n14931), .ZN(n14932) );
  AND2_X1 U18251 ( .A1(n14933), .A2(n14932), .ZN(n16248) );
  NAND2_X1 U18252 ( .A1(n16248), .A2(n14936), .ZN(n14934) );
  OAI211_X1 U18253 ( .C1(n14936), .C2(n12513), .A(n14935), .B(n14934), .ZN(
        P2_U2864) );
  AOI21_X1 U18254 ( .B1(n14938), .B2(n14937), .A(n12980), .ZN(n16117) );
  NAND2_X1 U18255 ( .A1(n16117), .A2(n14939), .ZN(n14944) );
  AND2_X1 U18256 ( .A1(n14941), .A2(n14940), .ZN(n14942) );
  OR2_X1 U18257 ( .A1(n14942), .A2(n9783), .ZN(n15222) );
  NAND2_X1 U18258 ( .A1(n16137), .A2(n14936), .ZN(n14943) );
  OAI211_X1 U18259 ( .C1(n14936), .C2(n14945), .A(n14944), .B(n14943), .ZN(
        P2_U2865) );
  NAND3_X1 U18260 ( .A1(n14946), .A2(n14881), .A3(n19146), .ZN(n14956) );
  INV_X1 U18261 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16490) );
  OR2_X1 U18262 ( .A1(n16122), .A2(n16490), .ZN(n14948) );
  NAND2_X1 U18263 ( .A1(n16122), .A2(BUF2_REG_13__SCAN_IN), .ZN(n14947) );
  AND2_X1 U18264 ( .A1(n14948), .A2(n14947), .ZN(n19255) );
  INV_X1 U18265 ( .A(n19255), .ZN(n14949) );
  AOI22_X1 U18266 ( .A1(n19105), .A2(n14949), .B1(n19157), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n14955) );
  AOI22_X1 U18267 ( .A1(n19106), .A2(BUF1_REG_29__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14954) );
  NAND2_X1 U18268 ( .A1(n13226), .A2(n14950), .ZN(n14951) );
  NAND2_X1 U18269 ( .A1(n14952), .A2(n14951), .ZN(n16051) );
  INV_X1 U18270 ( .A(n16051), .ZN(n15153) );
  NAND2_X1 U18271 ( .A1(n15153), .A2(n19158), .ZN(n14953) );
  NAND4_X1 U18272 ( .A1(n14956), .A2(n14955), .A3(n14954), .A4(n14953), .ZN(
        P2_U2890) );
  OR2_X1 U18273 ( .A1(n16122), .A2(n14957), .ZN(n14959) );
  NAND2_X1 U18274 ( .A1(n16122), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14958) );
  AND2_X1 U18275 ( .A1(n14959), .A2(n14958), .ZN(n19252) );
  OAI22_X1 U18276 ( .A1(n14999), .A2(n19252), .B1(n19132), .B2(n14960), .ZN(
        n14961) );
  AOI21_X1 U18277 ( .B1(n19158), .B2(n14962), .A(n14961), .ZN(n14964) );
  AOI22_X1 U18278 ( .A1(n19106), .A2(BUF1_REG_28__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n14963) );
  OAI211_X1 U18279 ( .C1(n14965), .C2(n19162), .A(n14964), .B(n14963), .ZN(
        P2_U2891) );
  NOR2_X1 U18280 ( .A1(n14966), .A2(n14967), .ZN(n14968) );
  OR2_X1 U18281 ( .A1(n13227), .A2(n14968), .ZN(n16062) );
  INV_X1 U18282 ( .A(n16062), .ZN(n15168) );
  INV_X1 U18283 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14969) );
  OR2_X1 U18284 ( .A1(n16122), .A2(n14969), .ZN(n14971) );
  NAND2_X1 U18285 ( .A1(n16122), .A2(BUF2_REG_11__SCAN_IN), .ZN(n14970) );
  AND2_X1 U18286 ( .A1(n14971), .A2(n14970), .ZN(n19250) );
  OAI22_X1 U18287 ( .A1(n14999), .A2(n19250), .B1(n19132), .B2(n14972), .ZN(
        n14973) );
  AOI21_X1 U18288 ( .B1(n19158), .B2(n15168), .A(n14973), .ZN(n14975) );
  AOI22_X1 U18289 ( .A1(n19106), .A2(BUF1_REG_27__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n14974) );
  OAI211_X1 U18290 ( .C1(n14976), .C2(n19162), .A(n14975), .B(n14974), .ZN(
        P2_U2892) );
  AND2_X1 U18291 ( .A1(n14978), .A2(n14977), .ZN(n14979) );
  NOR2_X1 U18292 ( .A1(n14966), .A2(n14979), .ZN(n16080) );
  MUX2_X1 U18293 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n16122), .Z(n19224) );
  INV_X1 U18294 ( .A(n19224), .ZN(n14981) );
  INV_X1 U18295 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14980) );
  OAI22_X1 U18296 ( .A1(n14999), .A2(n14981), .B1(n19132), .B2(n14980), .ZN(
        n14982) );
  AOI21_X1 U18297 ( .B1(n19158), .B2(n16080), .A(n14982), .ZN(n14984) );
  AOI22_X1 U18298 ( .A1(n19106), .A2(BUF1_REG_26__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n14983) );
  OAI211_X1 U18299 ( .C1(n14985), .C2(n19162), .A(n14984), .B(n14983), .ZN(
        P2_U2893) );
  INV_X1 U18300 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14986) );
  OR2_X1 U18301 ( .A1(n16122), .A2(n14986), .ZN(n14988) );
  NAND2_X1 U18302 ( .A1(n16122), .A2(BUF2_REG_9__SCAN_IN), .ZN(n14987) );
  AND2_X1 U18303 ( .A1(n14988), .A2(n14987), .ZN(n19244) );
  OAI22_X1 U18304 ( .A1(n14999), .A2(n19244), .B1(n19132), .B2(n14989), .ZN(
        n14990) );
  AOI21_X1 U18305 ( .B1(n19158), .B2(n14991), .A(n14990), .ZN(n14993) );
  AOI22_X1 U18306 ( .A1(n19106), .A2(BUF1_REG_25__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n14992) );
  OAI211_X1 U18307 ( .C1(n14994), .C2(n19162), .A(n14993), .B(n14992), .ZN(
        P2_U2894) );
  OR2_X1 U18308 ( .A1(n14995), .A2(n14996), .ZN(n14997) );
  AND2_X1 U18309 ( .A1(n14322), .A2(n14997), .ZN(n16095) );
  INV_X1 U18310 ( .A(n19128), .ZN(n14998) );
  OAI22_X1 U18311 ( .A1(n14999), .A2(n14998), .B1(n19132), .B2(n13446), .ZN(
        n15000) );
  AOI21_X1 U18312 ( .B1(n19158), .B2(n16095), .A(n15000), .ZN(n15002) );
  AOI22_X1 U18313 ( .A1(n19106), .A2(BUF1_REG_24__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15001) );
  OAI211_X1 U18314 ( .C1(n15003), .C2(n19162), .A(n15002), .B(n15001), .ZN(
        P2_U2895) );
  AND2_X1 U18315 ( .A1(n15219), .A2(n15004), .ZN(n15005) );
  OR2_X1 U18316 ( .A1(n15005), .A2(n14995), .ZN(n16243) );
  AOI22_X1 U18317 ( .A1(n19106), .A2(BUF1_REG_23__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U18318 ( .A1(n16121), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16122), .ZN(n19313) );
  INV_X1 U18319 ( .A(n19313), .ZN(n15006) );
  AOI22_X1 U18320 ( .A1(n19105), .A2(n15006), .B1(n19157), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15007) );
  OAI211_X1 U18321 ( .C1(n16124), .C2(n16243), .A(n15008), .B(n15007), .ZN(
        n15009) );
  AOI21_X1 U18322 ( .B1(n15010), .B2(n19146), .A(n15009), .ZN(n15011) );
  INV_X1 U18323 ( .A(n15011), .ZN(P2_U2896) );
  NAND2_X1 U18324 ( .A1(n15012), .A2(n19146), .ZN(n15017) );
  AOI22_X1 U18325 ( .A1(n16121), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16122), .ZN(n19302) );
  INV_X1 U18326 ( .A(n19302), .ZN(n19135) );
  AOI22_X1 U18327 ( .A1(n19105), .A2(n19135), .B1(n19157), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15016) );
  AOI22_X1 U18328 ( .A1(n19106), .A2(BUF1_REG_21__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15015) );
  NAND2_X1 U18329 ( .A1(n15013), .A2(n19158), .ZN(n15014) );
  NAND4_X1 U18330 ( .A1(n15017), .A2(n15016), .A3(n15015), .A4(n15014), .ZN(
        P2_U2898) );
  NAND2_X1 U18331 ( .A1(n15018), .A2(n19146), .ZN(n15023) );
  AOI22_X1 U18332 ( .A1(n16121), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16122), .ZN(n19292) );
  INV_X1 U18333 ( .A(n19292), .ZN(n15019) );
  AOI22_X1 U18334 ( .A1(n19105), .A2(n15019), .B1(n19157), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15022) );
  AOI22_X1 U18335 ( .A1(n19106), .A2(BUF1_REG_19__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15021) );
  NAND2_X1 U18336 ( .A1(n19158), .A2(n18902), .ZN(n15020) );
  NAND4_X1 U18337 ( .A1(n15023), .A2(n15022), .A3(n15021), .A4(n15020), .ZN(
        P2_U2900) );
  NAND2_X1 U18338 ( .A1(n15024), .A2(n19146), .ZN(n15032) );
  AOI22_X1 U18339 ( .A1(n16121), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16122), .ZN(n19284) );
  INV_X1 U18340 ( .A(n19284), .ZN(n15025) );
  AOI22_X1 U18341 ( .A1(n19105), .A2(n15025), .B1(n19157), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15031) );
  AOI22_X1 U18342 ( .A1(n19106), .A2(BUF1_REG_17__SCAN_IN), .B1(n19107), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n15030) );
  AND2_X1 U18343 ( .A1(n15261), .A2(n15026), .ZN(n15027) );
  NOR2_X1 U18344 ( .A1(n15028), .A2(n15027), .ZN(n18926) );
  NAND2_X1 U18345 ( .A1(n19158), .A2(n18926), .ZN(n15029) );
  NAND4_X1 U18346 ( .A1(n15032), .A2(n15031), .A3(n15030), .A4(n15029), .ZN(
        P2_U2902) );
  XNOR2_X1 U18347 ( .A(n9812), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16028) );
  NOR2_X1 U18348 ( .A1(n19269), .A2(n16028), .ZN(n15033) );
  AOI211_X1 U18349 ( .C1(n19258), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15034), .B(n15033), .ZN(n15035) );
  OAI21_X1 U18350 ( .B1(n16047), .B2(n16214), .A(n15035), .ZN(n15036) );
  AOI21_X1 U18351 ( .B1(n15037), .B2(n19260), .A(n15036), .ZN(n15038) );
  OAI21_X1 U18352 ( .B1(n15039), .B2(n16220), .A(n15038), .ZN(P2_U2984) );
  NAND2_X1 U18353 ( .A1(n15041), .A2(n15040), .ZN(n15043) );
  XOR2_X1 U18354 ( .A(n15043), .B(n15042), .Z(n15164) );
  AOI21_X1 U18355 ( .B1(n15046), .B2(n15045), .A(n15044), .ZN(n15161) );
  AOI21_X1 U18356 ( .B1(n15048), .B2(n15047), .A(n9812), .ZN(n16054) );
  NAND2_X1 U18357 ( .A1(n15077), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15155) );
  OAI21_X1 U18358 ( .B1(n16239), .B2(n15048), .A(n15155), .ZN(n15049) );
  AOI21_X1 U18359 ( .B1(n16227), .B2(n16054), .A(n15049), .ZN(n15050) );
  OAI21_X1 U18360 ( .B1(n16058), .B2(n16214), .A(n15050), .ZN(n15051) );
  AOI21_X1 U18361 ( .B1(n15161), .B2(n19260), .A(n15051), .ZN(n15052) );
  OAI21_X1 U18362 ( .B1(n15164), .B2(n16220), .A(n15052), .ZN(P2_U2985) );
  OAI21_X1 U18363 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n9759), .A(
        n10036), .ZN(n15177) );
  INV_X1 U18364 ( .A(n15054), .ZN(n15166) );
  NAND2_X1 U18365 ( .A1(n15055), .A2(n15173), .ZN(n15165) );
  NAND3_X1 U18366 ( .A1(n15166), .A2(n19264), .A3(n15165), .ZN(n15060) );
  NAND2_X1 U18367 ( .A1(n15077), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15170) );
  OAI21_X1 U18368 ( .B1(n16239), .B2(n15056), .A(n15170), .ZN(n15058) );
  NOR2_X1 U18369 ( .A1(n16068), .A2(n16214), .ZN(n15057) );
  AOI211_X1 U18370 ( .C1(n16227), .C2(n16064), .A(n15058), .B(n15057), .ZN(
        n15059) );
  OAI211_X1 U18371 ( .C1(n16219), .C2(n15177), .A(n15060), .B(n15059), .ZN(
        P2_U2987) );
  INV_X1 U18372 ( .A(n15061), .ZN(n15062) );
  AOI21_X1 U18373 ( .B1(n14318), .B2(n15063), .A(n15062), .ZN(n15065) );
  XNOR2_X1 U18374 ( .A(n15065), .B(n15064), .ZN(n15188) );
  AOI21_X1 U18375 ( .B1(n10038), .B2(n14331), .A(n9759), .ZN(n15186) );
  NOR2_X1 U18376 ( .A1(n9722), .A2(n15066), .ZN(n15181) );
  NOR2_X1 U18377 ( .A1(n19269), .A2(n15067), .ZN(n15068) );
  AOI211_X1 U18378 ( .C1(n19258), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15181), .B(n15068), .ZN(n15069) );
  OAI21_X1 U18379 ( .B1(n16077), .B2(n16214), .A(n15069), .ZN(n15070) );
  AOI21_X1 U18380 ( .B1(n15186), .B2(n19260), .A(n15070), .ZN(n15071) );
  OAI21_X1 U18381 ( .B1(n15188), .B2(n16220), .A(n15071), .ZN(P2_U2988) );
  INV_X1 U18382 ( .A(n15072), .ZN(n15073) );
  NOR2_X1 U18383 ( .A1(n15074), .A2(n15073), .ZN(n15075) );
  XNOR2_X1 U18384 ( .A(n15076), .B(n15075), .ZN(n15199) );
  AOI21_X1 U18385 ( .B1(n15190), .B2(n15089), .A(n14328), .ZN(n15197) );
  NAND2_X1 U18386 ( .A1(n16096), .A2(n19263), .ZN(n15079) );
  AOI22_X1 U18387 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n15077), .ZN(n15078) );
  OAI211_X1 U18388 ( .C1(n19269), .C2(n15080), .A(n15079), .B(n15078), .ZN(
        n15081) );
  AOI21_X1 U18389 ( .B1(n15197), .B2(n19260), .A(n15081), .ZN(n15082) );
  OAI21_X1 U18390 ( .B1(n15199), .B2(n16220), .A(n15082), .ZN(P2_U2990) );
  AND2_X1 U18391 ( .A1(n15084), .A2(n15083), .ZN(n15087) );
  OAI21_X1 U18392 ( .B1(n15087), .B2(n15086), .A(n15085), .ZN(n15088) );
  INV_X1 U18393 ( .A(n15088), .ZN(n16249) );
  NAND2_X1 U18394 ( .A1(n15207), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15208) );
  NAND2_X1 U18395 ( .A1(n15208), .A2(n16244), .ZN(n15090) );
  NAND2_X1 U18396 ( .A1(n15090), .A2(n15089), .ZN(n16252) );
  OAI22_X1 U18397 ( .A1(n16239), .A2(n13174), .B1(n19886), .B2(n9722), .ZN(
        n15091) );
  AOI21_X1 U18398 ( .B1(n16227), .B2(n16108), .A(n15091), .ZN(n15093) );
  NAND2_X1 U18399 ( .A1(n16248), .A2(n19263), .ZN(n15092) );
  OAI211_X1 U18400 ( .C1(n16252), .C2(n16219), .A(n15093), .B(n15092), .ZN(
        n15094) );
  AOI21_X1 U18401 ( .B1(n16249), .B2(n19264), .A(n15094), .ZN(n15095) );
  INV_X1 U18402 ( .A(n15095), .ZN(P2_U2991) );
  OAI21_X1 U18403 ( .B1(n16239), .B2(n15097), .A(n15096), .ZN(n15098) );
  AOI21_X1 U18404 ( .B1(n16227), .B2(n15099), .A(n15098), .ZN(n15100) );
  OAI21_X1 U18405 ( .B1(n15101), .B2(n16214), .A(n15100), .ZN(n15102) );
  AOI21_X1 U18406 ( .B1(n15103), .B2(n19260), .A(n15102), .ZN(n15104) );
  OAI21_X1 U18407 ( .B1(n15105), .B2(n16220), .A(n15104), .ZN(P2_U2993) );
  NAND2_X1 U18408 ( .A1(n15107), .A2(n15106), .ZN(n15111) );
  NAND2_X1 U18409 ( .A1(n15109), .A2(n15108), .ZN(n15110) );
  XNOR2_X1 U18410 ( .A(n15111), .B(n15110), .ZN(n15240) );
  OAI21_X1 U18411 ( .B1(n15113), .B2(n15112), .A(n15229), .ZN(n15115) );
  AND2_X1 U18412 ( .A1(n15115), .A2(n15114), .ZN(n15238) );
  NOR2_X1 U18413 ( .A1(n9722), .A2(n15116), .ZN(n15231) );
  NOR2_X1 U18414 ( .A1(n15117), .A2(n19269), .ZN(n15118) );
  AOI211_X1 U18415 ( .C1(n19258), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15231), .B(n15118), .ZN(n15119) );
  OAI21_X1 U18416 ( .B1(n16214), .B2(n15235), .A(n15119), .ZN(n15120) );
  AOI21_X1 U18417 ( .B1(n15238), .B2(n19260), .A(n15120), .ZN(n15121) );
  OAI21_X1 U18418 ( .B1(n15240), .B2(n16220), .A(n15121), .ZN(P2_U2994) );
  XNOR2_X1 U18419 ( .A(n15123), .B(n15122), .ZN(n15257) );
  INV_X1 U18420 ( .A(n15241), .ZN(n18925) );
  NOR2_X1 U18421 ( .A1(n19877), .A2(n9722), .ZN(n15126) );
  AOI22_X1 U18422 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16227), .B2(n18920), .ZN(n15124) );
  INV_X1 U18423 ( .A(n15124), .ZN(n15125) );
  AOI211_X1 U18424 ( .C1(n19263), .C2(n18925), .A(n15126), .B(n15125), .ZN(
        n15130) );
  OR2_X2 U18425 ( .A1(n15330), .A2(n16259), .ZN(n15276) );
  NAND2_X1 U18426 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15242) );
  INV_X1 U18427 ( .A(n15127), .ZN(n15128) );
  OAI211_X1 U18428 ( .C1(n16142), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19260), .B(n15128), .ZN(n15129) );
  OAI211_X1 U18429 ( .C1(n15257), .C2(n16220), .A(n15130), .B(n15129), .ZN(
        P2_U2997) );
  XNOR2_X1 U18430 ( .A(n15132), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15133) );
  XNOR2_X1 U18431 ( .A(n15131), .B(n15133), .ZN(n16305) );
  INV_X1 U18432 ( .A(n16205), .ZN(n15138) );
  OAI21_X1 U18433 ( .B1(n15136), .B2(n15138), .A(n15135), .ZN(n15137) );
  OAI21_X1 U18434 ( .B1(n16206), .B2(n15138), .A(n15137), .ZN(n16302) );
  OAI22_X1 U18435 ( .A1(n16239), .A2(n15139), .B1(n19863), .B2(n9722), .ZN(
        n15140) );
  INV_X1 U18436 ( .A(n15140), .ZN(n15142) );
  NAND2_X1 U18437 ( .A1(n16227), .A2(n19025), .ZN(n15141) );
  OAI211_X1 U18438 ( .C1(n19029), .C2(n16214), .A(n15142), .B(n15141), .ZN(
        n15143) );
  AOI21_X1 U18439 ( .B1(n16302), .B2(n19264), .A(n15143), .ZN(n15144) );
  OAI21_X1 U18440 ( .B1(n16219), .B2(n16305), .A(n15144), .ZN(P2_U3007) );
  XNOR2_X1 U18441 ( .A(n15145), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15368) );
  XOR2_X1 U18442 ( .A(n15147), .B(n15146), .Z(n15366) );
  OAI22_X1 U18443 ( .A1(n19861), .A2(n9722), .B1(n19269), .B2(n19040), .ZN(
        n15151) );
  INV_X1 U18444 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15148) );
  OAI22_X1 U18445 ( .A1(n16214), .A2(n15149), .B1(n16239), .B2(n15148), .ZN(
        n15150) );
  AOI211_X1 U18446 ( .C1(n15366), .C2(n19264), .A(n15151), .B(n15150), .ZN(
        n15152) );
  OAI21_X1 U18447 ( .B1(n15368), .B2(n16219), .A(n15152), .ZN(P2_U3008) );
  NAND2_X1 U18448 ( .A1(n16281), .A2(n15153), .ZN(n15154) );
  OAI211_X1 U18449 ( .C1(n16058), .C2(n16283), .A(n15155), .B(n15154), .ZN(
        n15159) );
  NOR3_X1 U18450 ( .A1(n15157), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15156), .ZN(n15158) );
  NAND2_X1 U18451 ( .A1(n15161), .A2(n16274), .ZN(n15162) );
  OAI211_X1 U18452 ( .C1(n15164), .C2(n16315), .A(n15163), .B(n15162), .ZN(
        P2_U3017) );
  NAND3_X1 U18453 ( .A1(n15166), .A2(n16301), .A3(n15165), .ZN(n15176) );
  NOR2_X1 U18454 ( .A1(n15167), .A2(n15173), .ZN(n15172) );
  NAND2_X1 U18455 ( .A1(n16281), .A2(n15168), .ZN(n15169) );
  OAI211_X1 U18456 ( .C1(n16068), .C2(n16283), .A(n15170), .B(n15169), .ZN(
        n15171) );
  AOI211_X1 U18457 ( .C1(n15174), .C2(n15173), .A(n15172), .B(n15171), .ZN(
        n15175) );
  OAI211_X1 U18458 ( .C1(n15177), .C2(n16307), .A(n15176), .B(n15175), .ZN(
        P2_U3019) );
  XNOR2_X1 U18459 ( .A(n10038), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15178) );
  NAND2_X1 U18460 ( .A1(n15179), .A2(n15178), .ZN(n15183) );
  NOR2_X1 U18461 ( .A1(n16077), .A2(n16283), .ZN(n15180) );
  AOI211_X1 U18462 ( .C1(n16080), .C2(n16281), .A(n15181), .B(n15180), .ZN(
        n15182) );
  OAI211_X1 U18463 ( .C1(n15184), .C2(n10038), .A(n15183), .B(n15182), .ZN(
        n15185) );
  AOI21_X1 U18464 ( .B1(n15186), .B2(n16274), .A(n15185), .ZN(n15187) );
  OAI21_X1 U18465 ( .B1(n15188), .B2(n16315), .A(n15187), .ZN(P2_U3020) );
  INV_X1 U18466 ( .A(n16096), .ZN(n15195) );
  AOI221_X1 U18467 ( .B1(n15191), .B2(n15190), .C1(n15211), .C2(n15190), .A(
        n15189), .ZN(n15193) );
  NOR2_X1 U18468 ( .A1(n9722), .A2(n12555), .ZN(n15192) );
  AOI211_X1 U18469 ( .C1(n16281), .C2(n16095), .A(n15193), .B(n15192), .ZN(
        n15194) );
  OAI21_X1 U18470 ( .B1(n15195), .B2(n16283), .A(n15194), .ZN(n15196) );
  AOI21_X1 U18471 ( .B1(n15197), .B2(n16274), .A(n15196), .ZN(n15198) );
  OAI21_X1 U18472 ( .B1(n15199), .B2(n16315), .A(n15198), .ZN(P2_U3022) );
  NAND2_X1 U18473 ( .A1(n15201), .A2(n15200), .ZN(n15206) );
  NAND2_X1 U18474 ( .A1(n15204), .A2(n15203), .ZN(n15205) );
  INV_X1 U18475 ( .A(n15207), .ZN(n15210) );
  INV_X1 U18476 ( .A(n15208), .ZN(n15209) );
  AOI21_X1 U18477 ( .B1(n16242), .B2(n15210), .A(n15209), .ZN(n16136) );
  INV_X1 U18478 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15212) );
  OR2_X1 U18479 ( .A1(n15212), .A2(n15211), .ZN(n16241) );
  NOR2_X1 U18480 ( .A1(n15214), .A2(n15213), .ZN(n16245) );
  NAND2_X1 U18481 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n15077), .ZN(n15215) );
  OAI221_X1 U18482 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16241), 
        .C1(n16242), .C2(n16245), .A(n15215), .ZN(n15224) );
  INV_X1 U18483 ( .A(n15216), .ZN(n15218) );
  NAND2_X1 U18484 ( .A1(n15218), .A2(n15217), .ZN(n15220) );
  AND2_X1 U18485 ( .A1(n15220), .A2(n15219), .ZN(n16116) );
  INV_X1 U18486 ( .A(n16116), .ZN(n15221) );
  OAI22_X1 U18487 ( .A1(n15222), .A2(n16283), .B1(n16306), .B2(n15221), .ZN(
        n15223) );
  AOI211_X1 U18488 ( .C1(n16136), .C2(n16274), .A(n15224), .B(n15223), .ZN(
        n15225) );
  INV_X1 U18489 ( .A(n15226), .ZN(n15227) );
  AOI21_X1 U18490 ( .B1(n15228), .B2(n15227), .A(n15229), .ZN(n15237) );
  NAND3_X1 U18491 ( .A1(n16260), .A2(n15230), .A3(n15229), .ZN(n15234) );
  INV_X1 U18492 ( .A(n16125), .ZN(n15232) );
  AOI21_X1 U18493 ( .B1(n16281), .B2(n15232), .A(n15231), .ZN(n15233) );
  OAI211_X1 U18494 ( .C1(n15235), .C2(n16283), .A(n15234), .B(n15233), .ZN(
        n15236) );
  AOI211_X1 U18495 ( .C1(n15238), .C2(n16274), .A(n15237), .B(n15236), .ZN(
        n15239) );
  OAI21_X1 U18496 ( .B1(n15240), .B2(n16315), .A(n15239), .ZN(P2_U3026) );
  OAI22_X1 U18497 ( .A1(n16283), .A2(n15241), .B1(n19877), .B2(n9722), .ZN(
        n15244) );
  NOR2_X1 U18498 ( .A1(n15319), .A2(n16259), .ZN(n15288) );
  AOI21_X1 U18499 ( .B1(n16159), .B2(n16274), .A(n15288), .ZN(n15265) );
  NOR3_X1 U18500 ( .A1(n15265), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15242), .ZN(n15243) );
  AOI211_X1 U18501 ( .C1(n16281), .C2(n18926), .A(n15244), .B(n15243), .ZN(
        n15256) );
  AND2_X1 U18502 ( .A1(n16307), .A2(n15245), .ZN(n15246) );
  OR2_X1 U18503 ( .A1(n16142), .A2(n15246), .ZN(n15252) );
  AND2_X1 U18504 ( .A1(n15247), .A2(n16259), .ZN(n15248) );
  OR2_X1 U18505 ( .A1(n16255), .A2(n15248), .ZN(n15277) );
  NOR2_X1 U18506 ( .A1(n15249), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15250) );
  NOR2_X1 U18507 ( .A1(n15277), .A2(n15250), .ZN(n15251) );
  NAND2_X1 U18508 ( .A1(n15252), .A2(n15251), .ZN(n15268) );
  NOR2_X1 U18509 ( .A1(n15253), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15254) );
  OAI21_X1 U18510 ( .B1(n15268), .B2(n15254), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15255) );
  OAI211_X1 U18511 ( .C1(n15257), .C2(n16315), .A(n15256), .B(n15255), .ZN(
        P2_U3029) );
  OAI21_X1 U18512 ( .B1(n15260), .B2(n15259), .A(n15258), .ZN(n16144) );
  OAI21_X1 U18513 ( .B1(n15278), .B2(n15262), .A(n15261), .ZN(n15263) );
  INV_X1 U18514 ( .A(n15263), .ZN(n19109) );
  OAI22_X1 U18515 ( .A1(n16283), .A2(n18939), .B1(n15264), .B2(n9722), .ZN(
        n15267) );
  NOR3_X1 U18516 ( .A1(n15265), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15287), .ZN(n15266) );
  AOI211_X1 U18517 ( .C1(n16281), .C2(n19109), .A(n15267), .B(n15266), .ZN(
        n15270) );
  NAND2_X1 U18518 ( .A1(n15268), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15269) );
  OAI211_X1 U18519 ( .C1(n16144), .C2(n16315), .A(n15270), .B(n15269), .ZN(
        P2_U3030) );
  NAND2_X1 U18520 ( .A1(n15272), .A2(n15271), .ZN(n15275) );
  NAND2_X1 U18521 ( .A1(n15273), .A2(n16155), .ZN(n15274) );
  XOR2_X1 U18522 ( .A(n15275), .B(n15274), .Z(n16151) );
  XNOR2_X1 U18523 ( .A(n15276), .B(n15287), .ZN(n16150) );
  INV_X1 U18524 ( .A(n16150), .ZN(n15294) );
  NAND2_X1 U18525 ( .A1(n15277), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15292) );
  INV_X1 U18526 ( .A(n15278), .ZN(n15284) );
  INV_X1 U18527 ( .A(n15279), .ZN(n15282) );
  INV_X1 U18528 ( .A(n15280), .ZN(n15281) );
  NAND2_X1 U18529 ( .A1(n15282), .A2(n15281), .ZN(n15283) );
  NAND2_X1 U18530 ( .A1(n15284), .A2(n15283), .ZN(n19115) );
  INV_X1 U18531 ( .A(n19115), .ZN(n15286) );
  NOR2_X1 U18532 ( .A1(n18940), .A2(n9722), .ZN(n15285) );
  AOI21_X1 U18533 ( .B1(n16281), .B2(n15286), .A(n15285), .ZN(n15291) );
  NAND2_X1 U18534 ( .A1(n15288), .A2(n15287), .ZN(n15290) );
  NAND2_X1 U18535 ( .A1(n12589), .A2(n18952), .ZN(n15289) );
  NAND4_X1 U18536 ( .A1(n15292), .A2(n15291), .A3(n15290), .A4(n15289), .ZN(
        n15293) );
  AOI21_X1 U18537 ( .B1(n15294), .B2(n16274), .A(n15293), .ZN(n15295) );
  OAI21_X1 U18538 ( .B1(n16151), .B2(n16315), .A(n15295), .ZN(P2_U3031) );
  NAND2_X1 U18539 ( .A1(n15297), .A2(n15296), .ZN(n15298) );
  INV_X1 U18540 ( .A(n19119), .ZN(n15302) );
  NOR2_X1 U18541 ( .A1(n19871), .A2(n9722), .ZN(n15301) );
  AOI211_X1 U18542 ( .C1(n15320), .C2(n15299), .A(n16261), .B(n15319), .ZN(
        n15300) );
  AOI211_X1 U18543 ( .C1(n16281), .C2(n15302), .A(n15301), .B(n15300), .ZN(
        n15303) );
  OAI21_X1 U18544 ( .B1(n16283), .B2(n15304), .A(n15303), .ZN(n15306) );
  NOR2_X2 U18545 ( .A1(n15330), .A2(n15320), .ZN(n16173) );
  XNOR2_X1 U18546 ( .A(n16173), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16165) );
  NOR2_X1 U18547 ( .A1(n16165), .A2(n16307), .ZN(n15305) );
  AOI211_X1 U18548 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16255), .A(
        n15306), .B(n15305), .ZN(n15307) );
  OAI21_X1 U18549 ( .B1(n16315), .B2(n16164), .A(n15307), .ZN(P2_U3033) );
  OR2_X1 U18550 ( .A1(n15329), .A2(n15326), .ZN(n15309) );
  NAND2_X1 U18551 ( .A1(n15309), .A2(n15325), .ZN(n15313) );
  AND2_X1 U18552 ( .A1(n15311), .A2(n15310), .ZN(n15312) );
  XNOR2_X1 U18553 ( .A(n15313), .B(n15312), .ZN(n16171) );
  INV_X1 U18554 ( .A(n16171), .ZN(n15324) );
  AOI21_X1 U18555 ( .B1(n15315), .B2(n15334), .A(n15314), .ZN(n19120) );
  NAND2_X1 U18556 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n15077), .ZN(n15316) );
  OAI21_X1 U18557 ( .B1(n16283), .B2(n18977), .A(n15316), .ZN(n15317) );
  AOI21_X1 U18558 ( .B1(n16281), .B2(n19120), .A(n15317), .ZN(n15318) );
  OAI21_X1 U18559 ( .B1(n15319), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15318), .ZN(n15322) );
  AND2_X1 U18560 ( .A1(n15330), .A2(n15320), .ZN(n16172) );
  NOR3_X1 U18561 ( .A1(n16173), .A2(n16172), .A3(n16307), .ZN(n15321) );
  AOI211_X1 U18562 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16255), .A(
        n15322), .B(n15321), .ZN(n15323) );
  OAI21_X1 U18563 ( .B1(n16315), .B2(n15324), .A(n15323), .ZN(P2_U3034) );
  INV_X1 U18564 ( .A(n15325), .ZN(n15327) );
  NOR2_X1 U18565 ( .A1(n15327), .A2(n15326), .ZN(n15328) );
  XNOR2_X1 U18566 ( .A(n15329), .B(n15328), .ZN(n16180) );
  INV_X1 U18567 ( .A(n16192), .ZN(n15332) );
  INV_X1 U18568 ( .A(n15330), .ZN(n15331) );
  AOI21_X1 U18569 ( .B1(n15337), .B2(n15332), .A(n15331), .ZN(n16179) );
  OAI21_X1 U18570 ( .B1(n15335), .B2(n15333), .A(n15334), .ZN(n19122) );
  INV_X1 U18571 ( .A(n16269), .ZN(n15340) );
  NOR2_X1 U18572 ( .A1(n11291), .A2(n9722), .ZN(n15339) );
  NAND2_X1 U18573 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15351), .ZN(
        n16271) );
  AOI211_X1 U18574 ( .C1(n16270), .C2(n15337), .A(n15336), .B(n16271), .ZN(
        n15338) );
  AOI211_X1 U18575 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15340), .A(
        n15339), .B(n15338), .ZN(n15342) );
  NAND2_X1 U18576 ( .A1(n12589), .A2(n18986), .ZN(n15341) );
  OAI211_X1 U18577 ( .C1(n16306), .C2(n19122), .A(n15342), .B(n15341), .ZN(
        n15343) );
  AOI21_X1 U18578 ( .B1(n16179), .B2(n16274), .A(n15343), .ZN(n15344) );
  OAI21_X1 U18579 ( .B1(n16180), .B2(n16315), .A(n15344), .ZN(P2_U3035) );
  NOR2_X1 U18580 ( .A1(n15345), .A2(n10906), .ZN(n15347) );
  XOR2_X1 U18581 ( .A(n15347), .B(n15346), .Z(n16198) );
  OAI21_X1 U18582 ( .B1(n12591), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16190), .ZN(n16197) );
  NOR2_X1 U18583 ( .A1(n11264), .A2(n9722), .ZN(n15348) );
  AOI221_X1 U18584 ( .B1(n15351), .B2(n15350), .C1(n15349), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15348), .ZN(n15355) );
  OAI21_X1 U18585 ( .B1(n15352), .B2(n16279), .A(n16266), .ZN(n19126) );
  INV_X1 U18586 ( .A(n19126), .ZN(n15353) );
  AOI22_X1 U18587 ( .A1(n12589), .A2(n19009), .B1(n16281), .B2(n15353), .ZN(
        n15354) );
  OAI211_X1 U18588 ( .C1(n16197), .C2(n16307), .A(n15355), .B(n15354), .ZN(
        n15356) );
  INV_X1 U18589 ( .A(n15356), .ZN(n15357) );
  OAI21_X1 U18590 ( .B1(n16315), .B2(n16198), .A(n15357), .ZN(P2_U3037) );
  XNOR2_X1 U18591 ( .A(n15359), .B(n15358), .ZN(n19133) );
  NOR2_X1 U18592 ( .A1(n19861), .A2(n9722), .ZN(n15360) );
  AOI221_X1 U18593 ( .B1(n16299), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        n15362), .C2(n15361), .A(n15360), .ZN(n15364) );
  NAND2_X1 U18594 ( .A1(n12589), .A2(n19042), .ZN(n15363) );
  OAI211_X1 U18595 ( .C1(n16306), .C2(n19133), .A(n15364), .B(n15363), .ZN(
        n15365) );
  AOI21_X1 U18596 ( .B1(n15366), .B2(n16301), .A(n15365), .ZN(n15367) );
  OAI21_X1 U18597 ( .B1(n15368), .B2(n16307), .A(n15367), .ZN(P2_U3040) );
  MUX2_X1 U18598 ( .A(n11180), .B(n15370), .S(n15369), .Z(n15371) );
  AOI21_X1 U18599 ( .B1(n19094), .B2(n15386), .A(n15371), .ZN(n16325) );
  INV_X1 U18600 ( .A(n15372), .ZN(n15373) );
  OAI222_X1 U18601 ( .A1(n15390), .A2(n15375), .B1(n19916), .B2(n16325), .C1(
        n15374), .C2(n15373), .ZN(n15376) );
  MUX2_X1 U18602 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15376), .S(
        n15391), .Z(P2_U3601) );
  INV_X1 U18603 ( .A(n15377), .ZN(n15389) );
  OR2_X1 U18604 ( .A1(n15379), .A2(n15381), .ZN(n15383) );
  OAI21_X1 U18605 ( .B1(n10665), .B2(n15381), .A(n15380), .ZN(n15382) );
  OAI211_X1 U18606 ( .C1(n15378), .C2(n15384), .A(n15383), .B(n15382), .ZN(
        n15385) );
  AOI21_X1 U18607 ( .B1(n15387), .B2(n15386), .A(n15385), .ZN(n16317) );
  OAI222_X1 U18608 ( .A1(n19929), .A2(n15390), .B1(n15389), .B2(n15388), .C1(
        n19916), .C2(n16317), .ZN(n15392) );
  MUX2_X1 U18609 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15392), .S(
        n15391), .Z(P2_U3599) );
  INV_X1 U18610 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17038) );
  INV_X1 U18611 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17107) );
  NOR3_X1 U18612 ( .A1(n15394), .A2(n17321), .A3(n15393), .ZN(n15395) );
  AOI21_X1 U18613 ( .B1(n18635), .B2(n15396), .A(n15395), .ZN(n15692) );
  NAND2_X1 U18614 ( .A1(n18846), .A2(n16398), .ZN(n16381) );
  NAND4_X1 U18615 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .A3(P3_EBX_REG_0__SCAN_IN), .A4(P3_EBX_REG_1__SCAN_IN), .ZN(n17215) );
  NAND2_X1 U18616 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16980), .ZN(n16966) );
  NAND2_X1 U18617 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16971), .ZN(n15468) );
  NOR2_X1 U18618 ( .A1(n17321), .A2(n17227), .ZN(n17223) );
  NAND2_X1 U18619 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16955) );
  NOR2_X2 U18620 ( .A1(n18226), .A2(n17227), .ZN(n17228) );
  AOI22_X1 U18621 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15400) );
  AOI22_X1 U18622 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15399) );
  AOI22_X1 U18623 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15398) );
  AOI22_X1 U18624 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15397) );
  NAND4_X1 U18625 ( .A1(n15400), .A2(n15399), .A3(n15398), .A4(n15397), .ZN(
        n15406) );
  AOI22_X1 U18626 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15404) );
  AOI22_X1 U18627 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U18628 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15402) );
  AOI22_X1 U18629 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13276), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15401) );
  NAND4_X1 U18630 ( .A1(n15404), .A2(n15403), .A3(n15402), .A4(n15401), .ZN(
        n15405) );
  NOR2_X1 U18631 ( .A1(n15406), .A2(n15405), .ZN(n16962) );
  AOI22_X1 U18632 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U18633 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15409) );
  AOI22_X1 U18634 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15408) );
  AOI22_X1 U18635 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15407) );
  NAND4_X1 U18636 ( .A1(n15410), .A2(n15409), .A3(n15408), .A4(n15407), .ZN(
        n15416) );
  AOI22_X1 U18637 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15414) );
  AOI22_X1 U18638 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15413) );
  AOI22_X1 U18639 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15412) );
  AOI22_X1 U18640 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15411) );
  NAND4_X1 U18641 ( .A1(n15414), .A2(n15413), .A3(n15412), .A4(n15411), .ZN(
        n15415) );
  NOR2_X1 U18642 ( .A1(n15416), .A2(n15415), .ZN(n16972) );
  AOI22_X1 U18643 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15420) );
  AOI22_X1 U18644 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13276), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15419) );
  AOI22_X1 U18645 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U18646 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15417) );
  NAND4_X1 U18647 ( .A1(n15420), .A2(n15419), .A3(n15418), .A4(n15417), .ZN(
        n15426) );
  AOI22_X1 U18648 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15424) );
  AOI22_X1 U18649 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9728), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15423) );
  AOI22_X1 U18650 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U18651 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15421) );
  NAND4_X1 U18652 ( .A1(n15424), .A2(n15423), .A3(n15422), .A4(n15421), .ZN(
        n15425) );
  NOR2_X1 U18653 ( .A1(n15426), .A2(n15425), .ZN(n16983) );
  AOI22_X1 U18654 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17116), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15430) );
  AOI22_X1 U18655 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15429) );
  AOI22_X1 U18656 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15428) );
  AOI22_X1 U18657 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15427) );
  NAND4_X1 U18658 ( .A1(n15430), .A2(n15429), .A3(n15428), .A4(n15427), .ZN(
        n15436) );
  AOI22_X1 U18659 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15434) );
  AOI22_X1 U18660 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15433) );
  AOI22_X1 U18661 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15432) );
  AOI22_X1 U18662 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15431) );
  NAND4_X1 U18663 ( .A1(n15434), .A2(n15433), .A3(n15432), .A4(n15431), .ZN(
        n15435) );
  NOR2_X1 U18664 ( .A1(n15436), .A2(n15435), .ZN(n16982) );
  NOR2_X1 U18665 ( .A1(n16983), .A2(n16982), .ZN(n16978) );
  AOI22_X1 U18666 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17163), .ZN(n15447) );
  AOI22_X1 U18667 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15446) );
  AOI22_X1 U18668 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17183), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17173), .ZN(n15437) );
  OAI21_X1 U18669 ( .B1(n15438), .B2(n10125), .A(n15437), .ZN(n15444) );
  AOI22_X1 U18670 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17181), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17162), .ZN(n15442) );
  AOI22_X1 U18671 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17191), .ZN(n15441) );
  AOI22_X1 U18672 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9728), .ZN(n15440) );
  AOI22_X1 U18673 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17080), .ZN(n15439) );
  NAND4_X1 U18674 ( .A1(n15442), .A2(n15441), .A3(n15440), .A4(n15439), .ZN(
        n15443) );
  AOI211_X1 U18675 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n9725), .A(
        n15444), .B(n15443), .ZN(n15445) );
  NAND3_X1 U18676 ( .A1(n15447), .A2(n15446), .A3(n15445), .ZN(n16977) );
  NAND2_X1 U18677 ( .A1(n16978), .A2(n16977), .ZN(n16976) );
  NOR2_X1 U18678 ( .A1(n16972), .A2(n16976), .ZN(n16969) );
  AOI22_X1 U18679 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13276), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U18680 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15456) );
  AOI22_X1 U18681 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15448) );
  OAI21_X1 U18682 ( .B1(n15522), .B2(n17127), .A(n15448), .ZN(n15454) );
  AOI22_X1 U18683 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15452) );
  AOI22_X1 U18684 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U18685 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15450) );
  AOI22_X1 U18686 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15449) );
  NAND4_X1 U18687 ( .A1(n15452), .A2(n15451), .A3(n15450), .A4(n15449), .ZN(
        n15453) );
  AOI211_X1 U18688 ( .C1(n17184), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n15454), .B(n15453), .ZN(n15455) );
  NAND3_X1 U18689 ( .A1(n15457), .A2(n15456), .A3(n15455), .ZN(n16968) );
  NAND2_X1 U18690 ( .A1(n16969), .A2(n16968), .ZN(n16967) );
  NOR2_X1 U18691 ( .A1(n16962), .A2(n16967), .ZN(n16961) );
  AOI22_X1 U18692 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15461) );
  AOI22_X1 U18693 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9730), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15460) );
  AOI22_X1 U18694 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U18695 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15458) );
  NAND4_X1 U18696 ( .A1(n15461), .A2(n15460), .A3(n15459), .A4(n15458), .ZN(
        n15467) );
  AOI22_X1 U18697 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13276), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15465) );
  AOI22_X1 U18698 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15464) );
  AOI22_X1 U18699 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15463) );
  AOI22_X1 U18700 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15462) );
  NAND4_X1 U18701 ( .A1(n15465), .A2(n15464), .A3(n15463), .A4(n15462), .ZN(
        n15466) );
  NOR2_X1 U18702 ( .A1(n15467), .A2(n15466), .ZN(n16951) );
  XNOR2_X1 U18703 ( .A(n16961), .B(n16951), .ZN(n17249) );
  NAND3_X1 U18704 ( .A1(n18226), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17142), 
        .ZN(n17123) );
  NAND2_X1 U18705 ( .A1(n17225), .A2(n17095), .ZN(n15480) );
  AOI22_X1 U18706 ( .A1(n17085), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U18707 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U18708 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13276), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15469) );
  OAI21_X1 U18709 ( .B1(n15522), .B2(n17000), .A(n15469), .ZN(n15475) );
  AOI22_X1 U18710 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15473) );
  AOI22_X1 U18711 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U18712 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U18713 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15470) );
  NAND4_X1 U18714 ( .A1(n15473), .A2(n15472), .A3(n15471), .A4(n15470), .ZN(
        n15474) );
  AOI211_X1 U18715 ( .C1(n9730), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n15475), .B(n15474), .ZN(n15476) );
  NAND3_X1 U18716 ( .A1(n15478), .A2(n15477), .A3(n15476), .ZN(n17327) );
  NAND2_X1 U18717 ( .A1(n17228), .A2(n17327), .ZN(n15479) );
  OAI221_X1 U18718 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17123), .C1(n17107), 
        .C2(n15480), .A(n15479), .ZN(P3_U2690) );
  NAND2_X1 U18719 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18407) );
  AOI221_X1 U18720 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18407), .C1(n15482), 
        .C2(n18407), .A(n15481), .ZN(n18184) );
  NOR2_X1 U18721 ( .A1(n15483), .A2(n18672), .ZN(n15484) );
  OAI21_X1 U18722 ( .B1(n15484), .B2(n18543), .A(n18185), .ZN(n18182) );
  AOI22_X1 U18723 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18184), .B1(
        n18182), .B2(n18677), .ZN(P3_U2865) );
  INV_X1 U18724 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17983) );
  NOR2_X1 U18725 ( .A1(n15584), .A2(n17983), .ZN(n17982) );
  INV_X1 U18726 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17968) );
  INV_X1 U18727 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17624) );
  NOR2_X1 U18728 ( .A1(n17968), .A2(n17624), .ZN(n17952) );
  NAND3_X1 U18729 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17952), .ZN(n17595) );
  INV_X1 U18730 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17948) );
  NOR2_X1 U18731 ( .A1(n17595), .A2(n17948), .ZN(n15592) );
  NAND2_X1 U18732 ( .A1(n17982), .A2(n15592), .ZN(n17925) );
  NAND2_X1 U18733 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15486) );
  INV_X1 U18734 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18011) );
  INV_X1 U18735 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18074) );
  NOR2_X1 U18736 ( .A1(n18086), .A2(n18074), .ZN(n18068) );
  INV_X1 U18737 ( .A(n18068), .ZN(n18067) );
  INV_X1 U18738 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17739) );
  NOR2_X1 U18739 ( .A1(n18067), .A2(n17739), .ZN(n18055) );
  NAND3_X1 U18740 ( .A1(n18055), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18022) );
  INV_X1 U18741 ( .A(n18022), .ZN(n18021) );
  NAND2_X1 U18742 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18021), .ZN(
        n18009) );
  NOR2_X1 U18743 ( .A1(n18011), .A2(n18009), .ZN(n16453) );
  NAND3_X1 U18744 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18115) );
  NOR2_X1 U18745 ( .A1(n18150), .A2(n18115), .ZN(n18088) );
  INV_X1 U18746 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18092) );
  NAND2_X1 U18747 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18098) );
  NOR2_X1 U18748 ( .A1(n18092), .A2(n18098), .ZN(n18007) );
  AND2_X1 U18749 ( .A1(n18088), .A2(n18007), .ZN(n17997) );
  NAND2_X1 U18750 ( .A1(n16453), .A2(n17997), .ZN(n17932) );
  NOR3_X1 U18751 ( .A1(n17925), .A2(n15486), .A3(n17932), .ZN(n17897) );
  INV_X1 U18752 ( .A(n17925), .ZN(n17585) );
  NOR2_X1 U18753 ( .A1(n18115), .A2(n15485), .ZN(n18089) );
  AND2_X1 U18754 ( .A1(n18007), .A2(n18089), .ZN(n17998) );
  NAND2_X1 U18755 ( .A1(n16453), .A2(n17998), .ZN(n16454) );
  INV_X1 U18756 ( .A(n16454), .ZN(n17975) );
  NAND2_X1 U18757 ( .A1(n17585), .A2(n17975), .ZN(n17914) );
  NOR2_X1 U18758 ( .A1(n15486), .A2(n17914), .ZN(n17878) );
  AOI22_X1 U18759 ( .A1(n18664), .A2(n17897), .B1(n16452), .B2(n17878), .ZN(
        n17905) );
  NAND2_X1 U18760 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15593) );
  NOR2_X1 U18761 ( .A1(n17905), .A2(n15593), .ZN(n16435) );
  NAND2_X1 U18762 ( .A1(n18055), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18043) );
  AOI22_X1 U18763 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15496) );
  AOI22_X1 U18764 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15495) );
  AOI22_X1 U18765 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15487) );
  OAI21_X1 U18766 ( .B1(n9761), .B2(n17199), .A(n15487), .ZN(n15493) );
  AOI22_X1 U18767 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15491) );
  AOI22_X1 U18768 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15490) );
  AOI22_X1 U18769 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15508), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15489) );
  AOI22_X1 U18770 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15488) );
  NAND4_X1 U18771 ( .A1(n15491), .A2(n15490), .A3(n15489), .A4(n15488), .ZN(
        n15492) );
  AOI211_X1 U18772 ( .C1(n13289), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n15493), .B(n15492), .ZN(n15494) );
  AOI22_X1 U18773 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U18774 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15499) );
  AOI22_X1 U18775 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15508), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15498) );
  AOI22_X1 U18776 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15497) );
  NAND4_X1 U18777 ( .A1(n15500), .A2(n15499), .A3(n15498), .A4(n15497), .ZN(
        n15506) );
  AOI22_X1 U18778 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U18779 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15503) );
  AOI22_X1 U18780 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9725), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15502) );
  AOI22_X1 U18781 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15501) );
  NAND4_X1 U18782 ( .A1(n15504), .A2(n15503), .A3(n15502), .A4(n15501), .ZN(
        n15505) );
  NOR2_X1 U18783 ( .A1(n15507), .A2(n17364), .ZN(n15538) );
  AOI22_X1 U18784 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15520) );
  AOI22_X1 U18785 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15508), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15519) );
  AOI22_X1 U18786 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15509) );
  OAI21_X1 U18787 ( .B1(n15511), .B2(n15510), .A(n15509), .ZN(n15517) );
  AOI22_X1 U18788 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15515) );
  AOI22_X1 U18789 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15514) );
  AOI22_X1 U18790 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15513) );
  AOI22_X1 U18791 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15512) );
  NAND4_X1 U18792 ( .A1(n15515), .A2(n15514), .A3(n15513), .A4(n15512), .ZN(
        n15516) );
  AOI211_X1 U18793 ( .C1(n9725), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n15517), .B(n15516), .ZN(n15518) );
  NAND3_X1 U18794 ( .A1(n15520), .A2(n15519), .A3(n15518), .ZN(n15553) );
  NAND2_X1 U18795 ( .A1(n15538), .A2(n15553), .ZN(n15534) );
  NOR2_X1 U18796 ( .A1(n17356), .A2(n15534), .ZN(n15542) );
  AOI22_X1 U18797 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U18798 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15531) );
  AOI22_X1 U18799 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15521) );
  OAI21_X1 U18800 ( .B1(n15522), .B2(n17097), .A(n15521), .ZN(n15529) );
  AOI22_X1 U18801 ( .A1(n15508), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U18802 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15526) );
  AOI22_X1 U18803 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15525) );
  AOI22_X1 U18804 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15524) );
  NAND4_X1 U18805 ( .A1(n15527), .A2(n15526), .A3(n15525), .A4(n15524), .ZN(
        n15528) );
  AOI211_X1 U18806 ( .C1(n17175), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n15529), .B(n15528), .ZN(n15530) );
  NAND3_X1 U18807 ( .A1(n15532), .A2(n15531), .A3(n15530), .ZN(n15554) );
  NAND2_X1 U18808 ( .A1(n15542), .A2(n15554), .ZN(n15533) );
  NOR2_X1 U18809 ( .A1(n17349), .A2(n15533), .ZN(n15550) );
  XNOR2_X1 U18810 ( .A(n15533), .B(n16401), .ZN(n17798) );
  INV_X1 U18811 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18129) );
  XOR2_X1 U18812 ( .A(n15534), .B(n17356), .Z(n17821) );
  NAND2_X1 U18813 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15535), .ZN(
        n15537) );
  NAND2_X1 U18814 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15539), .ZN(
        n15540) );
  INV_X1 U18815 ( .A(n15553), .ZN(n17360) );
  XNOR2_X1 U18816 ( .A(n15538), .B(n17360), .ZN(n17836) );
  NAND2_X1 U18817 ( .A1(n17821), .A2(n17820), .ZN(n15541) );
  NOR2_X1 U18818 ( .A1(n17821), .A2(n17820), .ZN(n17819) );
  INV_X1 U18819 ( .A(n15554), .ZN(n17353) );
  XNOR2_X1 U18820 ( .A(n15542), .B(n17353), .ZN(n15544) );
  NAND2_X1 U18821 ( .A1(n15543), .A2(n15544), .ZN(n15545) );
  INV_X1 U18822 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18107) );
  NAND2_X1 U18823 ( .A1(n15550), .A2(n15546), .ZN(n15551) );
  INV_X1 U18824 ( .A(n15546), .ZN(n15549) );
  NAND2_X1 U18825 ( .A1(n17798), .A2(n17797), .ZN(n15548) );
  NAND2_X1 U18826 ( .A1(n15550), .A2(n15549), .ZN(n15547) );
  OAI211_X1 U18827 ( .C1(n15550), .C2(n15549), .A(n15548), .B(n15547), .ZN(
        n17779) );
  NAND2_X1 U18828 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17779), .ZN(
        n17778) );
  INV_X1 U18829 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17719) );
  INV_X1 U18830 ( .A(n15593), .ZN(n17879) );
  NAND3_X1 U18831 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n17879), .ZN(n15576) );
  NOR2_X1 U18832 ( .A1(n17925), .A2(n15576), .ZN(n15575) );
  INV_X1 U18833 ( .A(n15575), .ZN(n16455) );
  NAND2_X1 U18834 ( .A1(n15557), .A2(n15553), .ZN(n15556) );
  XNOR2_X1 U18835 ( .A(n17353), .B(n15555), .ZN(n15567) );
  XNOR2_X1 U18836 ( .A(n18122), .B(n15567), .ZN(n17806) );
  XOR2_X1 U18837 ( .A(n17356), .B(n15556), .Z(n15564) );
  XNOR2_X1 U18838 ( .A(n17360), .B(n15557), .ZN(n15558) );
  NAND2_X1 U18839 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15558), .ZN(
        n15563) );
  INV_X1 U18840 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18139) );
  XNOR2_X1 U18841 ( .A(n18139), .B(n15558), .ZN(n17831) );
  NAND2_X1 U18842 ( .A1(n15560), .A2(n15559), .ZN(n15562) );
  NAND2_X1 U18843 ( .A1(n15562), .A2(n15561), .ZN(n17830) );
  NAND2_X1 U18844 ( .A1(n17831), .A2(n17830), .ZN(n17829) );
  NAND2_X1 U18845 ( .A1(n15563), .A2(n17829), .ZN(n15565) );
  NAND2_X1 U18846 ( .A1(n15564), .A2(n15565), .ZN(n17815) );
  NAND2_X1 U18847 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17816), .ZN(
        n15566) );
  NAND2_X1 U18848 ( .A1(n17815), .A2(n15566), .ZN(n17805) );
  NAND2_X1 U18849 ( .A1(n17806), .A2(n17805), .ZN(n17804) );
  NAND2_X1 U18850 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15567), .ZN(
        n15568) );
  NAND2_X1 U18851 ( .A1(n17804), .A2(n15568), .ZN(n15570) );
  AOI21_X1 U18852 ( .B1(n17349), .B2(n16447), .A(n17786), .ZN(n15571) );
  XNOR2_X1 U18853 ( .A(n15570), .B(n15569), .ZN(n17792) );
  NAND2_X1 U18854 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17792), .ZN(
        n17791) );
  NAND2_X1 U18855 ( .A1(n15571), .A2(n15570), .ZN(n15572) );
  NAND2_X1 U18856 ( .A1(n17749), .A2(n16453), .ZN(n17939) );
  NOR2_X1 U18857 ( .A1(n16455), .A2(n17939), .ZN(n17880) );
  AOI22_X1 U18858 ( .A1(n18633), .A2(n17881), .B1(n17880), .B2(n18099), .ZN(
        n15573) );
  INV_X1 U18859 ( .A(n15573), .ZN(n15574) );
  INV_X1 U18860 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17529) );
  INV_X1 U18861 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17506) );
  NOR2_X1 U18862 ( .A1(n17529), .A2(n17506), .ZN(n16418) );
  OAI211_X1 U18863 ( .C1(n16435), .C2(n15574), .A(n18169), .B(n16418), .ZN(
        n15667) );
  INV_X1 U18864 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16430) );
  NAND2_X1 U18865 ( .A1(n18169), .A2(n18091), .ZN(n18134) );
  INV_X1 U18866 ( .A(n18134), .ZN(n18165) );
  NAND2_X1 U18867 ( .A1(n18668), .A2(n18144), .ZN(n18041) );
  INV_X1 U18868 ( .A(n18666), .ZN(n18651) );
  INV_X1 U18869 ( .A(n18145), .ZN(n17984) );
  INV_X1 U18870 ( .A(n17932), .ZN(n17976) );
  AOI21_X1 U18871 ( .B1(n15575), .B2(n17976), .A(n18144), .ZN(n17884) );
  AOI221_X1 U18872 ( .B1(n15576), .B2(n17984), .C1(n17914), .C2(n17984), .A(
        n17884), .ZN(n15577) );
  OAI211_X1 U18873 ( .C1(n18651), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15577), .B(n17974), .ZN(n15662) );
  AOI21_X1 U18874 ( .B1(n17529), .B2(n18041), .A(n15662), .ZN(n16450) );
  NAND2_X1 U18875 ( .A1(n16418), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15661) );
  INV_X1 U18876 ( .A(n15661), .ZN(n16436) );
  NAND2_X1 U18877 ( .A1(n17881), .A2(n16436), .ZN(n16417) );
  NAND2_X1 U18878 ( .A1(n16418), .A2(n17880), .ZN(n16443) );
  NOR2_X1 U18879 ( .A1(n16430), .A2(n16443), .ZN(n16419) );
  NOR3_X1 U18880 ( .A1(n16419), .A2(n16401), .A3(n18173), .ZN(n15578) );
  AOI211_X1 U18881 ( .C1(n18126), .C2(n16417), .A(n15578), .B(n18164), .ZN(
        n15670) );
  OAI21_X1 U18882 ( .B1(n16450), .B2(n18159), .A(n15670), .ZN(n15579) );
  AOI21_X1 U18883 ( .B1(n18165), .B2(n17506), .A(n15579), .ZN(n15600) );
  NAND3_X1 U18884 ( .A1(n16380), .A2(n18169), .A3(n16401), .ZN(n18080) );
  INV_X1 U18885 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17904) );
  NAND2_X1 U18886 ( .A1(n16453), .A2(n17784), .ZN(n15587) );
  INV_X1 U18887 ( .A(n15587), .ZN(n15585) );
  NOR2_X1 U18888 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17758) );
  NOR4_X1 U18889 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15581) );
  NAND4_X1 U18890 ( .A1(n17785), .A2(n17758), .A3(n15581), .A4(n18011), .ZN(
        n15582) );
  NAND2_X1 U18891 ( .A1(n17786), .A2(n15584), .ZN(n15583) );
  INV_X1 U18892 ( .A(n15586), .ZN(n17657) );
  NAND2_X1 U18893 ( .A1(n17657), .A2(n17983), .ZN(n17656) );
  NAND2_X1 U18894 ( .A1(n15588), .A2(n15587), .ZN(n17665) );
  INV_X1 U18895 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17917) );
  NOR2_X1 U18896 ( .A1(n17925), .A2(n17917), .ZN(n17912) );
  NOR2_X1 U18897 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17786), .ZN(
        n17648) );
  NAND2_X1 U18898 ( .A1(n17648), .A2(n17968), .ZN(n15589) );
  NOR2_X1 U18899 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15589), .ZN(
        n17611) );
  INV_X1 U18900 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17936) );
  NAND2_X1 U18901 ( .A1(n17611), .A2(n17936), .ZN(n17593) );
  NAND2_X1 U18902 ( .A1(n17982), .A2(n17665), .ZN(n17609) );
  NAND2_X1 U18903 ( .A1(n17622), .A2(n17609), .ZN(n17649) );
  NAND2_X1 U18904 ( .A1(n15592), .A2(n17649), .ZN(n17574) );
  OR2_X1 U18905 ( .A1(n17786), .A2(n17567), .ZN(n17545) );
  OAI221_X1 U18906 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17610), 
        .C1(n17904), .C2(n17546), .A(n17545), .ZN(n17534) );
  NOR2_X1 U18907 ( .A1(n17534), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17533) );
  NOR2_X1 U18908 ( .A1(n17546), .A2(n17610), .ZN(n15594) );
  NAND2_X1 U18909 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17786), .ZN(
        n16440) );
  NOR2_X2 U18910 ( .A1(n15596), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17520) );
  NAND2_X1 U18911 ( .A1(n17506), .A2(n17610), .ZN(n16441) );
  INV_X1 U18912 ( .A(n16441), .ZN(n15597) );
  OAI21_X1 U18913 ( .B1(n17521), .B2(n16440), .A(n15664), .ZN(n15598) );
  XNOR2_X1 U18914 ( .A(n15598), .B(n16430), .ZN(n16428) );
  AOI22_X1 U18915 ( .A1(n9724), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18096), 
        .B2(n16428), .ZN(n15599) );
  OAI221_X1 U18916 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15667), 
        .C1(n16430), .C2(n15600), .A(n15599), .ZN(P3_U2833) );
  AOI22_X1 U18917 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19081), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19058), .ZN(n15610) );
  INV_X1 U18918 ( .A(n15601), .ZN(n15602) );
  AOI22_X1 U18919 ( .A1(n15602), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n9707), .ZN(n15609) );
  AOI22_X1 U18920 ( .A1(n16137), .A2(n19093), .B1(n16116), .B2(n19019), .ZN(
        n15608) );
  AOI21_X1 U18921 ( .B1(n15605), .B2(n15604), .A(n15603), .ZN(n15606) );
  NAND2_X1 U18922 ( .A1(n19055), .A2(n15606), .ZN(n15607) );
  NAND4_X1 U18923 ( .A1(n15610), .A2(n15609), .A3(n15608), .A4(n15607), .ZN(
        P2_U2833) );
  INV_X1 U18924 ( .A(n15625), .ZN(n15623) );
  INV_X1 U18925 ( .A(n15621), .ZN(n15619) );
  AOI211_X1 U18926 ( .C1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n15612), .A(
        n20628), .B(n15611), .ZN(n15617) );
  INV_X1 U18927 ( .A(n15617), .ZN(n15615) );
  OAI211_X1 U18928 ( .C1(n15615), .C2(n20587), .A(n15614), .B(n15613), .ZN(
        n15616) );
  OAI21_X1 U18929 ( .B1(n15617), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15616), .ZN(n15618) );
  AOI21_X1 U18930 ( .B1(n15619), .B2(n12247), .A(n15618), .ZN(n15620) );
  AOI21_X1 U18931 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15621), .A(
        n15620), .ZN(n15622) );
  OAI21_X1 U18932 ( .B1(n15623), .B2(n20549), .A(n15622), .ZN(n15624) );
  OAI21_X1 U18933 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15625), .A(
        n15624), .ZN(n15637) );
  NAND2_X1 U18934 ( .A1(n19998), .A2(n13394), .ZN(n15632) );
  OAI21_X1 U18935 ( .B1(n15628), .B2(n15627), .A(n15626), .ZN(n15631) );
  INV_X1 U18936 ( .A(n15629), .ZN(n15630) );
  AOI211_X1 U18937 ( .C1(n15633), .C2(n15632), .A(n15631), .B(n15630), .ZN(
        n15635) );
  NAND2_X1 U18938 ( .A1(n15635), .A2(n15634), .ZN(n15636) );
  AOI21_X1 U18939 ( .B1(n15637), .B2(n20188), .A(n15636), .ZN(n15654) );
  INV_X1 U18940 ( .A(n15654), .ZN(n15645) );
  NAND4_X1 U18941 ( .A1(n15639), .A2(n12214), .A3(n15638), .A4(n20633), .ZN(
        n15643) );
  OAI21_X1 U18942 ( .B1(n20864), .B2(n15641), .A(n15640), .ZN(n15642) );
  OAI21_X1 U18943 ( .B1(n15644), .B2(n15643), .A(n15642), .ZN(n16018) );
  AOI221_X1 U18944 ( .B1(n20761), .B2(n20760), .C1(n15645), .C2(n20760), .A(
        n16018), .ZN(n16020) );
  NOR2_X1 U18945 ( .A1(n15646), .A2(n16015), .ZN(n15647) );
  NOR2_X1 U18946 ( .A1(n16020), .A2(n15647), .ZN(n15652) );
  INV_X1 U18947 ( .A(n16015), .ZN(n15648) );
  AOI211_X1 U18948 ( .C1(n15671), .C2(n20764), .A(n15649), .B(n15648), .ZN(
        n15650) );
  NAND2_X1 U18949 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15650), .ZN(n15651) );
  OAI22_X1 U18950 ( .A1(n15652), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n16020), 
        .B2(n15651), .ZN(n15653) );
  OAI21_X1 U18951 ( .B1(n15654), .B2(n19992), .A(n15653), .ZN(P1_U3161) );
  AOI22_X1 U18952 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15861), .B1(
        n16000), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15660) );
  INV_X1 U18953 ( .A(n15655), .ZN(n15658) );
  INV_X1 U18954 ( .A(n15656), .ZN(n15657) );
  AOI22_X1 U18955 ( .A1(n15658), .A2(n20182), .B1(n15999), .B2(n15657), .ZN(
        n15659) );
  OAI211_X1 U18956 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15862), .A(
        n15660), .B(n15659), .ZN(P1_U3010) );
  OAI211_X1 U18957 ( .C1(n15662), .C2(n15661), .A(n18091), .B(n18169), .ZN(
        n16432) );
  NOR2_X1 U18958 ( .A1(n17521), .A2(n16440), .ZN(n15663) );
  NAND2_X1 U18959 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15663), .ZN(
        n16384) );
  INV_X1 U18960 ( .A(n16384), .ZN(n15665) );
  NOR2_X1 U18961 ( .A1(n15665), .A2(n16382), .ZN(n15666) );
  XNOR2_X1 U18962 ( .A(n15666), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16411) );
  NOR2_X1 U18963 ( .A1(n18162), .A2(n18794), .ZN(n16409) );
  NOR3_X1 U18964 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16430), .A3(
        n15667), .ZN(n15668) );
  AOI211_X1 U18965 ( .C1(n18096), .C2(n16411), .A(n16409), .B(n15668), .ZN(
        n15669) );
  OAI221_X1 U18966 ( .B1(n16413), .B2(n15670), .C1(n16413), .C2(n16432), .A(
        n15669), .ZN(P3_U2832) );
  NAND2_X1 U18967 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15671), .ZN(n20771) );
  INV_X1 U18968 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20781) );
  NAND3_X1 U18969 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .A3(n20781), .ZN(
        n15673) );
  INV_X1 U18970 ( .A(HOLD), .ZN(n20773) );
  OAI211_X1 U18971 ( .C1(n20781), .C2(n20773), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15672) );
  NAND4_X1 U18972 ( .A1(n15674), .A2(n20771), .A3(n15673), .A4(n15672), .ZN(
        P1_U3195) );
  INV_X1 U18973 ( .A(n20144), .ZN(n20135) );
  INV_X1 U18974 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16541) );
  NOR2_X1 U18975 ( .A1(n20135), .A2(n16541), .ZN(P1_U2905) );
  INV_X1 U18976 ( .A(n15675), .ZN(n15676) );
  NAND3_X1 U18977 ( .A1(n14744), .A2(n15676), .A3(n15874), .ZN(n15677) );
  NAND2_X1 U18978 ( .A1(n15678), .A2(n15677), .ZN(n15680) );
  XNOR2_X1 U18979 ( .A(n15680), .B(n15679), .ZN(n15776) );
  INV_X1 U18980 ( .A(n15681), .ZN(n15684) );
  AOI22_X1 U18981 ( .A1(n15874), .A2(n15928), .B1(n15682), .B2(n20175), .ZN(
        n15683) );
  OAI211_X1 U18982 ( .C1(n15966), .C2(n15684), .A(n15946), .B(n15683), .ZN(
        n15873) );
  INV_X1 U18983 ( .A(n15873), .ZN(n15686) );
  INV_X1 U18984 ( .A(n15878), .ZN(n15931) );
  NOR2_X1 U18985 ( .A1(n20172), .A2(n15931), .ZN(n15915) );
  AOI22_X1 U18986 ( .A1(n20175), .A2(n15917), .B1(n15685), .B2(n15915), .ZN(
        n15930) );
  AOI221_X1 U18987 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15686), 
        .C1(n15930), .C2(n15686), .A(n15679), .ZN(n15687) );
  NOR2_X1 U18988 ( .A1(n20177), .A2(n20817), .ZN(n15774) );
  AOI211_X1 U18989 ( .C1(n15776), .C2(n20182), .A(n15687), .B(n15774), .ZN(
        n15689) );
  NAND3_X1 U18990 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15875), .A3(
        n15679), .ZN(n15688) );
  OAI211_X1 U18991 ( .C1(n15721), .C2(n20179), .A(n15689), .B(n15688), .ZN(
        P1_U3011) );
  NOR3_X1 U18992 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15690) );
  NOR3_X1 U18993 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19969), .A3(n19822), 
        .ZN(n16365) );
  NOR4_X1 U18994 ( .A1(n15690), .A2(n19975), .A3(n15691), .A4(n16365), .ZN(
        P2_U3178) );
  AOI221_X1 U18995 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15691), .C1(n19956), .C2(
        n15691), .A(n19768), .ZN(n19951) );
  INV_X1 U18996 ( .A(n19951), .ZN(n19948) );
  NOR2_X1 U18997 ( .A1(n16336), .A2(n19948), .ZN(P2_U3047) );
  OR3_X1 U18998 ( .A1(n15692), .A2(n17387), .A3(n16398), .ZN(n15693) );
  AOI21_X2 U18999 ( .B1(n15694), .B2(n15693), .A(n18697), .ZN(n17231) );
  NAND2_X1 U19000 ( .A1(n18226), .A2(n17231), .ZN(n17379) );
  INV_X1 U19001 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17452) );
  NAND2_X1 U19002 ( .A1(n18667), .A2(n17231), .ZN(n17372) );
  AOI22_X1 U19003 ( .A1(n17378), .A2(BUF2_REG_0__SCAN_IN), .B1(n17377), .B2(
        n17862), .ZN(n15695) );
  OAI221_X1 U19004 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17379), .C1(n17452), 
        .C2(n17231), .A(n15695), .ZN(P3_U2735) );
  INV_X1 U19005 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15703) );
  NAND2_X1 U19006 ( .A1(n15696), .A2(n20824), .ZN(n15697) );
  OAI22_X1 U19007 ( .A1(n15707), .A2(n20824), .B1(n15698), .B2(n15697), .ZN(
        n15699) );
  AOI21_X1 U19008 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n20093), .A(n15699), .ZN(
        n15702) );
  OAI22_X1 U19009 ( .A1(n15853), .A2(n20081), .B1(n15766), .B2(n20088), .ZN(
        n15700) );
  AOI21_X1 U19010 ( .B1(n15763), .B2(n20051), .A(n15700), .ZN(n15701) );
  OAI211_X1 U19011 ( .C1(n15703), .C2(n20064), .A(n15702), .B(n15701), .ZN(
        P1_U2816) );
  AOI22_X1 U19012 ( .A1(n15704), .A2(n20102), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n20093), .ZN(n15712) );
  NOR3_X1 U19013 ( .A1(n20091), .A2(n20814), .A3(n15705), .ZN(n15720) );
  AND2_X1 U19014 ( .A1(n15706), .A2(n15720), .ZN(n15717) );
  AOI21_X1 U19015 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15717), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15708) );
  OAI22_X1 U19016 ( .A1(n15709), .A2(n20029), .B1(n15708), .B2(n15707), .ZN(
        n15710) );
  AOI21_X1 U19017 ( .B1(n20099), .B2(n15856), .A(n15710), .ZN(n15711) );
  OAI211_X1 U19018 ( .C1(n15713), .C2(n20064), .A(n15712), .B(n15711), .ZN(
        P1_U2817) );
  AOI22_X1 U19019 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20092), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(n20093), .ZN(n15719) );
  INV_X1 U19020 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20821) );
  OAI21_X1 U19021 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n20091), .A(n15722), 
        .ZN(n15716) );
  OAI22_X1 U19022 ( .A1(n15714), .A2(n20029), .B1(n20081), .B2(n15868), .ZN(
        n15715) );
  AOI221_X1 U19023 ( .B1(n15717), .B2(n20821), .C1(n15716), .C2(
        P1_REIP_REG_22__SCAN_IN), .A(n15715), .ZN(n15718) );
  OAI211_X1 U19024 ( .C1(n15773), .C2(n20088), .A(n15719), .B(n15718), .ZN(
        P1_U2818) );
  AOI22_X1 U19025 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20092), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(n20093), .ZN(n15726) );
  NOR2_X1 U19026 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15720), .ZN(n15723) );
  OAI22_X1 U19027 ( .A1(n15723), .A2(n15722), .B1(n15721), .B2(n20081), .ZN(
        n15724) );
  AOI21_X1 U19028 ( .B1(n15775), .B2(n20051), .A(n15724), .ZN(n15725) );
  OAI211_X1 U19029 ( .C1(n15779), .C2(n20088), .A(n15726), .B(n15725), .ZN(
        P1_U2820) );
  NAND2_X1 U19030 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n20092), .ZN(
        n15727) );
  OAI211_X1 U19031 ( .C1(n20024), .C2(n15728), .A(n20177), .B(n15727), .ZN(
        n15729) );
  AOI211_X1 U19032 ( .C1(n20102), .C2(n15731), .A(n15730), .B(n15729), .ZN(
        n15735) );
  AOI22_X1 U19033 ( .A1(n15733), .A2(n20051), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n15732), .ZN(n15734) );
  OAI211_X1 U19034 ( .C1(n20081), .C2(n15882), .A(n15735), .B(n15734), .ZN(
        P1_U2822) );
  NAND2_X1 U19035 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15738) );
  AOI21_X1 U19036 ( .B1(n15738), .B2(n15737), .A(n15736), .ZN(n15747) );
  AOI22_X1 U19037 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n20093), .B1(n20099), 
        .B2(n15933), .ZN(n15739) );
  OAI211_X1 U19038 ( .C1(n20064), .C2(n15740), .A(n15739), .B(n20177), .ZN(
        n15744) );
  OAI22_X1 U19039 ( .A1(n15742), .A2(n20029), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n15741), .ZN(n15743) );
  AOI211_X1 U19040 ( .C1(n15745), .C2(n20102), .A(n15744), .B(n15743), .ZN(
        n15746) );
  OAI21_X1 U19041 ( .B1(n15747), .B2(n20804), .A(n15746), .ZN(P1_U2827) );
  NAND2_X1 U19042 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15756), .ZN(n15748) );
  AOI21_X1 U19043 ( .B1(n20802), .B2(n15748), .A(n15747), .ZN(n15751) );
  AOI22_X1 U19044 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20092), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(n20093), .ZN(n15749) );
  OAI211_X1 U19045 ( .C1(n15956), .C2(n20081), .A(n15749), .B(n20177), .ZN(
        n15750) );
  AOI211_X1 U19046 ( .C1(n20102), .C2(n15808), .A(n15751), .B(n15750), .ZN(
        n15752) );
  OAI21_X1 U19047 ( .B1(n20029), .B2(n15812), .A(n15752), .ZN(P1_U2828) );
  OAI21_X1 U19048 ( .B1(n20064), .B2(n11936), .A(n20177), .ZN(n15755) );
  INV_X1 U19049 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15753) );
  OAI22_X1 U19050 ( .A1(n15819), .A2(n20088), .B1(n15753), .B2(n20024), .ZN(
        n15754) );
  AOI211_X1 U19051 ( .C1(n20099), .C2(n15958), .A(n15755), .B(n15754), .ZN(
        n15758) );
  AOI22_X1 U19052 ( .A1(n15816), .A2(n20051), .B1(n15756), .B2(n20800), .ZN(
        n15757) );
  OAI211_X1 U19053 ( .C1(n15759), .C2(n20800), .A(n15758), .B(n15757), .ZN(
        P1_U2829) );
  AOI22_X1 U19054 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n15765) );
  AOI22_X1 U19055 ( .A1(n15849), .A2(n20167), .B1(n15799), .B2(n15763), .ZN(
        n15764) );
  OAI211_X1 U19056 ( .C1(n20157), .C2(n15766), .A(n15765), .B(n15764), .ZN(
        P1_U2975) );
  AOI22_X1 U19057 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15772) );
  NAND2_X1 U19058 ( .A1(n15767), .A2(n15768), .ZN(n15769) );
  XOR2_X1 U19059 ( .A(n12357), .B(n15769), .Z(n15865) );
  AOI22_X1 U19060 ( .A1(n15865), .A2(n20167), .B1(n15799), .B2(n15770), .ZN(
        n15771) );
  OAI211_X1 U19061 ( .C1(n20157), .C2(n15773), .A(n15772), .B(n15771), .ZN(
        P1_U2977) );
  AOI21_X1 U19062 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20165), .A(
        n15774), .ZN(n15778) );
  AOI22_X1 U19063 ( .A1(n15776), .A2(n20167), .B1(n15799), .B2(n15775), .ZN(
        n15777) );
  OAI211_X1 U19064 ( .C1(n20157), .C2(n15779), .A(n15778), .B(n15777), .ZN(
        P1_U2979) );
  AOI22_X1 U19065 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15788) );
  INV_X1 U19066 ( .A(n15780), .ZN(n15782) );
  AOI21_X1 U19067 ( .B1(n15783), .B2(n15782), .A(n15781), .ZN(n15785) );
  XNOR2_X1 U19068 ( .A(n15785), .B(n15784), .ZN(n15904) );
  AOI22_X1 U19069 ( .A1(n15786), .A2(n15799), .B1(n20167), .B2(n15904), .ZN(
        n15787) );
  OAI211_X1 U19070 ( .C1(n20157), .C2(n15789), .A(n15788), .B(n15787), .ZN(
        P1_U2983) );
  MUX2_X1 U19071 ( .A(n12689), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .S(
        n9712), .Z(n15797) );
  AOI21_X1 U19072 ( .B1(n14183), .B2(n15792), .A(n15791), .ZN(n15795) );
  INV_X1 U19073 ( .A(n15793), .ZN(n15794) );
  NOR2_X1 U19074 ( .A1(n15795), .A2(n15794), .ZN(n15796) );
  XOR2_X1 U19075 ( .A(n15797), .B(n15796), .Z(n15922) );
  AOI22_X1 U19076 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15802) );
  AOI22_X1 U19077 ( .A1(n15800), .A2(n15799), .B1(n15809), .B2(n15798), .ZN(
        n15801) );
  OAI211_X1 U19078 ( .C1(n15922), .C2(n20158), .A(n15802), .B(n15801), .ZN(
        P1_U2985) );
  AOI22_X1 U19079 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15811) );
  AND2_X1 U19080 ( .A1(n15804), .A2(n15803), .ZN(n15806) );
  OAI21_X1 U19081 ( .B1(n15807), .B2(n15806), .A(n15805), .ZN(n15953) );
  AOI22_X1 U19082 ( .A1(n20167), .A2(n15953), .B1(n15809), .B2(n15808), .ZN(
        n15810) );
  OAI211_X1 U19083 ( .C1(n20191), .C2(n15812), .A(n15811), .B(n15810), .ZN(
        P1_U2987) );
  AOI22_X1 U19084 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15818) );
  NOR3_X1 U19085 ( .A1(n14183), .A2(n9757), .A3(n15976), .ZN(n15814) );
  NOR2_X1 U19086 ( .A1(n15814), .A2(n15813), .ZN(n15815) );
  XNOR2_X1 U19087 ( .A(n15815), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15960) );
  AOI22_X1 U19088 ( .A1(n20167), .A2(n15960), .B1(n15799), .B2(n15816), .ZN(
        n15817) );
  OAI211_X1 U19089 ( .C1(n20157), .C2(n15819), .A(n15818), .B(n15817), .ZN(
        P1_U2988) );
  AOI22_X1 U19090 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15825) );
  XNOR2_X1 U19091 ( .A(n15821), .B(n15997), .ZN(n15822) );
  XNOR2_X1 U19092 ( .A(n15823), .B(n15822), .ZN(n15993) );
  AOI22_X1 U19093 ( .A1(n15993), .A2(n20167), .B1(n15799), .B2(n20044), .ZN(
        n15824) );
  OAI211_X1 U19094 ( .C1(n20157), .C2(n20047), .A(n15825), .B(n15824), .ZN(
        P1_U2992) );
  AOI22_X1 U19095 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16000), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15832) );
  NAND2_X1 U19096 ( .A1(n15829), .A2(n15828), .ZN(n15830) );
  XNOR2_X1 U19097 ( .A(n15827), .B(n15830), .ZN(n16002) );
  AOI22_X1 U19098 ( .A1(n16002), .A2(n20167), .B1(n15799), .B2(n20052), .ZN(
        n15831) );
  OAI211_X1 U19099 ( .C1(n20157), .C2(n20058), .A(n15832), .B(n15831), .ZN(
        P1_U2993) );
  INV_X1 U19100 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20065) );
  OAI222_X1 U19101 ( .A1(n20157), .A2(n20074), .B1(n15833), .B2(n20158), .C1(
        n20191), .C2(n20068), .ZN(n15834) );
  INV_X1 U19102 ( .A(n15834), .ZN(n15836) );
  OAI211_X1 U19103 ( .C1(n20065), .C2(n15837), .A(n15836), .B(n15835), .ZN(
        P1_U2994) );
  INV_X1 U19104 ( .A(n15838), .ZN(n15839) );
  AOI22_X1 U19105 ( .A1(n15840), .A2(n20182), .B1(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15839), .ZN(n15845) );
  NAND2_X1 U19106 ( .A1(n16000), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15844) );
  NAND2_X1 U19107 ( .A1(n15999), .A2(n15841), .ZN(n15842) );
  NAND4_X1 U19108 ( .A1(n15845), .A2(n15844), .A3(n15843), .A4(n15842), .ZN(
        P1_U3006) );
  INV_X1 U19109 ( .A(n15846), .ZN(n15847) );
  NOR3_X1 U19110 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14726), .A3(
        n15847), .ZN(n15848) );
  NOR2_X1 U19111 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15863), .ZN(
        n15854) );
  OAI221_X1 U19112 ( .B1(n15851), .B2(n15850), .C1(n15851), .C2(n15854), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15852) );
  INV_X1 U19113 ( .A(n15862), .ZN(n15855) );
  AOI22_X1 U19114 ( .A1(n16000), .A2(P1_REIP_REG_23__SCAN_IN), .B1(n15855), 
        .B2(n15854), .ZN(n15859) );
  AOI22_X1 U19115 ( .A1(n15857), .A2(n20182), .B1(n15999), .B2(n15856), .ZN(
        n15858) );
  OAI211_X1 U19116 ( .C1(n15860), .C2(n14726), .A(n15859), .B(n15858), .ZN(
        P1_U3008) );
  AOI22_X1 U19117 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15861), .B1(
        n16000), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15867) );
  AOI21_X1 U19118 ( .B1(n12701), .B2(n12357), .A(n15862), .ZN(n15864) );
  AOI22_X1 U19119 ( .A1(n15865), .A2(n20182), .B1(n15864), .B2(n15863), .ZN(
        n15866) );
  OAI211_X1 U19120 ( .C1(n20179), .C2(n15868), .A(n15867), .B(n15866), .ZN(
        P1_U3009) );
  INV_X1 U19121 ( .A(n15869), .ZN(n15871) );
  AOI22_X1 U19122 ( .A1(n15871), .A2(n20182), .B1(n15999), .B2(n15870), .ZN(
        n15877) );
  NOR2_X1 U19123 ( .A1(n20177), .A2(n20814), .ZN(n15872) );
  AOI221_X1 U19124 ( .B1(n15875), .B2(n15874), .C1(n15873), .C2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15872), .ZN(n15876) );
  NAND2_X1 U19125 ( .A1(n15877), .A2(n15876), .ZN(P1_U3012) );
  NOR2_X1 U19126 ( .A1(n15937), .A2(n12689), .ZN(n15880) );
  NAND2_X1 U19127 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15878), .ZN(
        n15920) );
  INV_X1 U19128 ( .A(n15946), .ZN(n15967) );
  AOI221_X1 U19129 ( .B1(n12689), .B2(n15943), .C1(n15920), .C2(n15943), .A(
        n15967), .ZN(n15879) );
  OAI221_X1 U19130 ( .B1(n15916), .B2(n15880), .C1(n15916), .C2(n15917), .A(
        n15879), .ZN(n15908) );
  AOI21_X1 U19131 ( .B1(n15985), .B2(n15881), .A(n15908), .ZN(n15897) );
  NOR2_X1 U19132 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15881), .ZN(
        n15885) );
  INV_X1 U19133 ( .A(n15939), .ZN(n15957) );
  NAND3_X1 U19134 ( .A1(n15917), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15957), .ZN(n15927) );
  NOR2_X1 U19135 ( .A1(n12689), .A2(n15927), .ZN(n15899) );
  OAI22_X1 U19136 ( .A1(n15883), .A2(n15988), .B1(n20179), .B2(n15882), .ZN(
        n15884) );
  AOI21_X1 U19137 ( .B1(n15885), .B2(n15899), .A(n15884), .ZN(n15887) );
  NAND2_X1 U19138 ( .A1(n16000), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15886) );
  OAI211_X1 U19139 ( .C1(n15897), .C2(n15888), .A(n15887), .B(n15886), .ZN(
        P1_U3013) );
  NOR2_X1 U19140 ( .A1(n15898), .A2(n15889), .ZN(n15890) );
  AOI21_X1 U19141 ( .B1(n15890), .B2(n15899), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15896) );
  INV_X1 U19142 ( .A(n15891), .ZN(n15893) );
  AOI22_X1 U19143 ( .A1(n15893), .A2(n20182), .B1(n15999), .B2(n15892), .ZN(
        n15895) );
  NAND2_X1 U19144 ( .A1(n16000), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15894) );
  OAI211_X1 U19145 ( .C1(n15897), .C2(n15896), .A(n15895), .B(n15894), .ZN(
        P1_U3014) );
  INV_X1 U19146 ( .A(n15899), .ZN(n15913) );
  NOR2_X1 U19147 ( .A1(n15898), .A2(n15913), .ZN(n15902) );
  AOI21_X1 U19148 ( .B1(n15899), .B2(n15898), .A(n15908), .ZN(n15900) );
  INV_X1 U19149 ( .A(n15900), .ZN(n15901) );
  MUX2_X1 U19150 ( .A(n15902), .B(n15901), .S(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(n15903) );
  AOI21_X1 U19151 ( .B1(n15904), .B2(n20182), .A(n15903), .ZN(n15906) );
  NAND2_X1 U19152 ( .A1(n16000), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15905) );
  OAI211_X1 U19153 ( .C1(n20179), .C2(n15907), .A(n15906), .B(n15905), .ZN(
        P1_U3015) );
  AOI22_X1 U19154 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15908), .B1(
        n16000), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15912) );
  AOI22_X1 U19155 ( .A1(n15910), .A2(n20182), .B1(n15999), .B2(n15909), .ZN(
        n15911) );
  OAI211_X1 U19156 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15913), .A(
        n15912), .B(n15911), .ZN(P1_U3016) );
  OAI22_X1 U19157 ( .A1(n15917), .A2(n15916), .B1(n15915), .B2(n15914), .ZN(
        n15918) );
  AOI211_X1 U19158 ( .C1(n15928), .C2(n15920), .A(n15919), .B(n15918), .ZN(
        n15938) );
  OAI21_X1 U19159 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15930), .A(
        n15938), .ZN(n15925) );
  NOR2_X1 U19160 ( .A1(n20177), .A2(n20805), .ZN(n15924) );
  OAI22_X1 U19161 ( .A1(n15922), .A2(n15988), .B1(n20179), .B2(n15921), .ZN(
        n15923) );
  AOI211_X1 U19162 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15925), .A(
        n15924), .B(n15923), .ZN(n15926) );
  OAI21_X1 U19163 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15927), .A(
        n15926), .ZN(P1_U3017) );
  INV_X1 U19164 ( .A(n15928), .ZN(n15929) );
  AOI221_X1 U19165 ( .B1(n15931), .B2(n15930), .C1(n15929), .C2(n15930), .A(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15932) );
  AOI21_X1 U19166 ( .B1(n16000), .B2(P1_REIP_REG_13__SCAN_IN), .A(n15932), 
        .ZN(n15936) );
  AOI22_X1 U19167 ( .A1(n15934), .A2(n20182), .B1(n15999), .B2(n15933), .ZN(
        n15935) );
  OAI211_X1 U19168 ( .C1(n15938), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        P1_U3018) );
  NOR2_X1 U19169 ( .A1(n15939), .A2(n15944), .ZN(n15951) );
  NAND2_X1 U19170 ( .A1(n15941), .A2(n15940), .ZN(n15963) );
  INV_X1 U19171 ( .A(n15963), .ZN(n15947) );
  AOI22_X1 U19172 ( .A1(n20175), .A2(n15944), .B1(n15943), .B2(n15942), .ZN(
        n15945) );
  NAND2_X1 U19173 ( .A1(n15946), .A2(n15945), .ZN(n15959) );
  AOI21_X1 U19174 ( .B1(n15948), .B2(n15947), .A(n15959), .ZN(n15949) );
  INV_X1 U19175 ( .A(n15949), .ZN(n15950) );
  MUX2_X1 U19176 ( .A(n15951), .B(n15950), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n15952) );
  AOI21_X1 U19177 ( .B1(n15953), .B2(n20182), .A(n15952), .ZN(n15955) );
  NAND2_X1 U19178 ( .A1(n16000), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15954) );
  OAI211_X1 U19179 ( .C1(n20179), .C2(n15956), .A(n15955), .B(n15954), .ZN(
        P1_U3019) );
  NAND2_X1 U19180 ( .A1(n15965), .A2(n15957), .ZN(n16005) );
  AOI22_X1 U19181 ( .A1(n16000), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n15999), 
        .B2(n15958), .ZN(n15962) );
  AOI22_X1 U19182 ( .A1(n15960), .A2(n20182), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15959), .ZN(n15961) );
  OAI211_X1 U19183 ( .C1(n16005), .C2(n15963), .A(n15962), .B(n15961), .ZN(
        P1_U3020) );
  AOI21_X1 U19184 ( .B1(n15966), .B2(n15965), .A(n15964), .ZN(n15969) );
  AOI221_X1 U19185 ( .B1(n15969), .B2(n15985), .C1(n15968), .C2(n15985), .A(
        n15967), .ZN(n15984) );
  NOR2_X1 U19186 ( .A1(n15986), .A2(n16005), .ZN(n15994) );
  NAND3_X1 U19187 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n15994), .ZN(n15978) );
  AOI221_X1 U19188 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n15976), .C2(n15983), .A(
        n15978), .ZN(n15970) );
  AOI21_X1 U19189 ( .B1(n16000), .B2(P1_REIP_REG_10__SCAN_IN), .A(n15970), 
        .ZN(n15971) );
  OAI21_X1 U19190 ( .B1(n20179), .B2(n15972), .A(n15971), .ZN(n15973) );
  AOI21_X1 U19191 ( .B1(n15974), .B2(n20182), .A(n15973), .ZN(n15975) );
  OAI21_X1 U19192 ( .B1(n15984), .B2(n15976), .A(n15975), .ZN(P1_U3021) );
  INV_X1 U19193 ( .A(n15977), .ZN(n20014) );
  NOR2_X1 U19194 ( .A1(n20177), .A2(n20796), .ZN(n15981) );
  OAI22_X1 U19195 ( .A1(n15979), .A2(n15988), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15978), .ZN(n15980) );
  AOI211_X1 U19196 ( .C1(n15999), .C2(n20014), .A(n15981), .B(n15980), .ZN(
        n15982) );
  OAI21_X1 U19197 ( .B1(n15984), .B2(n15983), .A(n15982), .ZN(P1_U3022) );
  AOI21_X1 U19198 ( .B1(n15986), .B2(n15985), .A(n16001), .ZN(n15998) );
  INV_X1 U19199 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20793) );
  OAI222_X1 U19200 ( .A1(n20036), .A2(n20179), .B1(n20177), .B2(n20793), .C1(
        n15988), .C2(n15987), .ZN(n15989) );
  INV_X1 U19201 ( .A(n15989), .ZN(n15991) );
  OAI221_X1 U19202 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15992), .C2(n15997), .A(
        n15994), .ZN(n15990) );
  OAI211_X1 U19203 ( .C1(n15998), .C2(n15992), .A(n15991), .B(n15990), .ZN(
        P1_U3023) );
  AOI22_X1 U19204 ( .A1(n16000), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n15999), 
        .B2(n20038), .ZN(n15996) );
  AOI22_X1 U19205 ( .A1(n15994), .A2(n15997), .B1(n20182), .B2(n15993), .ZN(
        n15995) );
  OAI211_X1 U19206 ( .C1(n15998), .C2(n15997), .A(n15996), .B(n15995), .ZN(
        P1_U3024) );
  AOI22_X1 U19207 ( .A1(n16000), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n15999), 
        .B2(n20049), .ZN(n16004) );
  AOI22_X1 U19208 ( .A1(n16002), .A2(n20182), .B1(n16001), .B2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16003) );
  OAI211_X1 U19209 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16005), .A(
        n16004), .B(n16003), .ZN(P1_U3025) );
  INV_X1 U19210 ( .A(n16006), .ZN(n16009) );
  NAND3_X1 U19211 ( .A1(n16009), .A2(n16008), .A3(n16007), .ZN(n16010) );
  OAI21_X1 U19212 ( .B1(n16011), .B2(n13674), .A(n16010), .ZN(P1_U3468) );
  NAND4_X1 U19213 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20764), .A4(n20864), .ZN(n16012) );
  NAND2_X1 U19214 ( .A1(n16013), .A2(n16012), .ZN(n20762) );
  INV_X1 U19215 ( .A(n20867), .ZN(n16016) );
  OAI21_X1 U19216 ( .B1(n16020), .B2(n20761), .A(n20760), .ZN(n16014) );
  OAI211_X1 U19217 ( .C1(n16016), .C2(n20864), .A(n16015), .B(n16014), .ZN(
        n16017) );
  AOI221_X1 U19218 ( .B1(n16019), .B2(n16018), .C1(n20762), .C2(n16018), .A(
        n16017), .ZN(P1_U3162) );
  NOR2_X1 U19219 ( .A1(n16020), .A2(n20761), .ZN(n16022) );
  OAI22_X1 U19220 ( .A1(n20593), .A2(n16022), .B1(n16021), .B2(n20761), .ZN(
        P1_U3466) );
  OR3_X1 U19221 ( .A1(n16023), .A2(P2_EBX_REG_30__SCAN_IN), .A3(n19063), .ZN(
        n16025) );
  NAND2_X1 U19222 ( .A1(n19081), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n16024) );
  OAI211_X1 U19223 ( .C1(n16026), .C2(n14876), .A(n16025), .B(n16024), .ZN(
        n16027) );
  AOI21_X1 U19224 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n9707), .A(
        n16027), .ZN(n16032) );
  INV_X1 U19225 ( .A(n16028), .ZN(n16034) );
  NOR2_X1 U19226 ( .A1(n19069), .A2(n16029), .ZN(n16053) );
  OAI211_X1 U19227 ( .C1(n16033), .C2(n19075), .A(n16032), .B(n16031), .ZN(
        P2_U2824) );
  AOI21_X1 U19228 ( .B1(n16035), .B2(n16034), .A(n19825), .ZN(n16045) );
  NAND2_X1 U19229 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n9707), .ZN(
        n16038) );
  AOI22_X1 U19230 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n19081), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n19058), .ZN(n16037) );
  OAI211_X1 U19231 ( .C1(n16039), .C2(n19063), .A(n16038), .B(n16037), .ZN(
        n16040) );
  AOI21_X1 U19232 ( .B1(n16041), .B2(n19019), .A(n16040), .ZN(n16042) );
  INV_X1 U19233 ( .A(n16042), .ZN(n16043) );
  AOI21_X1 U19234 ( .B1(n16045), .B2(n16044), .A(n16043), .ZN(n16046) );
  OAI21_X1 U19235 ( .B1(n16047), .B2(n19075), .A(n16046), .ZN(P2_U2825) );
  AOI22_X1 U19236 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19081), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19058), .ZN(n16050) );
  AOI22_X1 U19237 ( .A1(n16048), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n9707), .ZN(n16049) );
  OAI211_X1 U19238 ( .C1(n16051), .C2(n19083), .A(n16050), .B(n16049), .ZN(
        n16056) );
  AOI211_X1 U19239 ( .C1(n16054), .C2(n16053), .A(n16052), .B(n19825), .ZN(
        n16055) );
  NOR2_X1 U19240 ( .A1(n16056), .A2(n16055), .ZN(n16057) );
  OAI21_X1 U19241 ( .B1(n16058), .B2(n19075), .A(n16057), .ZN(P2_U2826) );
  AOI22_X1 U19242 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n19081), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n19058), .ZN(n16061) );
  AOI22_X1 U19243 ( .A1(n16059), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n9707), .ZN(n16060) );
  OAI211_X1 U19244 ( .C1(n16062), .C2(n19083), .A(n16061), .B(n16060), .ZN(
        n16066) );
  AOI211_X1 U19245 ( .C1(n16064), .C2(n16063), .A(n9852), .B(n19825), .ZN(
        n16065) );
  NOR2_X1 U19246 ( .A1(n16066), .A2(n16065), .ZN(n16067) );
  OAI21_X1 U19247 ( .B1(n16068), .B2(n19075), .A(n16067), .ZN(P2_U2828) );
  AOI211_X1 U19248 ( .C1(n16071), .C2(n16070), .A(n16069), .B(n19825), .ZN(
        n16079) );
  AOI22_X1 U19249 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19081), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19058), .ZN(n16076) );
  INV_X1 U19250 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16072) );
  OAI22_X1 U19251 ( .A1(n16073), .A2(n19063), .B1(n16072), .B2(n19079), .ZN(
        n16074) );
  INV_X1 U19252 ( .A(n16074), .ZN(n16075) );
  OAI211_X1 U19253 ( .C1(n16077), .C2(n19075), .A(n16076), .B(n16075), .ZN(
        n16078) );
  AOI211_X1 U19254 ( .C1(n19019), .C2(n16080), .A(n16079), .B(n16078), .ZN(
        n16081) );
  INV_X1 U19255 ( .A(n16081), .ZN(P2_U2829) );
  AOI211_X1 U19256 ( .C1(n16084), .C2(n16082), .A(n16083), .B(n19825), .ZN(
        n16092) );
  AOI22_X1 U19257 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19081), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19058), .ZN(n16089) );
  OAI22_X1 U19258 ( .A1(n16086), .A2(n19063), .B1(n16085), .B2(n19079), .ZN(
        n16087) );
  INV_X1 U19259 ( .A(n16087), .ZN(n16088) );
  OAI211_X1 U19260 ( .C1(n16090), .C2(n19083), .A(n16089), .B(n16088), .ZN(
        n16091) );
  AOI211_X1 U19261 ( .C1(n19093), .C2(n16093), .A(n16092), .B(n16091), .ZN(
        n16094) );
  INV_X1 U19262 ( .A(n16094), .ZN(P2_U2830) );
  AOI22_X1 U19263 ( .A1(n16096), .A2(n19093), .B1(n16095), .B2(n19019), .ZN(
        n16105) );
  AOI211_X1 U19264 ( .C1(n16099), .C2(n16098), .A(n16097), .B(n19825), .ZN(
        n16103) );
  AOI22_X1 U19265 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n9707), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n19058), .ZN(n16100) );
  OAI21_X1 U19266 ( .B1(n16101), .B2(n19063), .A(n16100), .ZN(n16102) );
  AOI211_X1 U19267 ( .C1(n19081), .C2(P2_REIP_REG_24__SCAN_IN), .A(n16103), 
        .B(n16102), .ZN(n16104) );
  NAND2_X1 U19268 ( .A1(n16105), .A2(n16104), .ZN(P2_U2831) );
  AOI211_X1 U19269 ( .C1(n16108), .C2(n16107), .A(n16106), .B(n19825), .ZN(
        n16113) );
  AOI22_X1 U19270 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19081), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n19058), .ZN(n16111) );
  AOI22_X1 U19271 ( .A1(n16109), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n9707), .ZN(n16110) );
  OAI211_X1 U19272 ( .C1(n16243), .C2(n19083), .A(n16111), .B(n16110), .ZN(
        n16112) );
  AOI211_X1 U19273 ( .C1(n19093), .C2(n16248), .A(n16113), .B(n16112), .ZN(
        n16114) );
  INV_X1 U19274 ( .A(n16114), .ZN(P2_U2832) );
  OAI22_X1 U19275 ( .A1(n16122), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16121), .ZN(n19306) );
  INV_X1 U19276 ( .A(n19306), .ZN(n16115) );
  AOI22_X1 U19277 ( .A1(n19105), .A2(n16115), .B1(n19157), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16120) );
  AOI22_X1 U19278 ( .A1(n19107), .A2(BUF2_REG_22__SCAN_IN), .B1(n19106), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16119) );
  AOI22_X1 U19279 ( .A1(n16117), .A2(n19146), .B1(n19158), .B2(n16116), .ZN(
        n16118) );
  NAND3_X1 U19280 ( .A1(n16120), .A2(n16119), .A3(n16118), .ZN(P2_U2897) );
  OAI22_X1 U19281 ( .A1(n16122), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16121), .ZN(n19296) );
  INV_X1 U19282 ( .A(n19296), .ZN(n16123) );
  AOI22_X1 U19283 ( .A1(n19105), .A2(n16123), .B1(n19157), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16130) );
  AOI22_X1 U19284 ( .A1(n19107), .A2(BUF2_REG_20__SCAN_IN), .B1(n19106), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16129) );
  NOR2_X1 U19285 ( .A1(n16125), .A2(n16124), .ZN(n16126) );
  AOI21_X1 U19286 ( .B1(n16127), .B2(n19146), .A(n16126), .ZN(n16128) );
  NAND3_X1 U19287 ( .A1(n16130), .A2(n16129), .A3(n16128), .ZN(P2_U2899) );
  AOI22_X1 U19288 ( .A1(n19105), .A2(n16131), .B1(n19157), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16135) );
  AOI22_X1 U19289 ( .A1(n19107), .A2(BUF2_REG_18__SCAN_IN), .B1(n19106), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16134) );
  AOI22_X1 U19290 ( .A1(n16132), .A2(n19146), .B1(n19158), .B2(n18913), .ZN(
        n16133) );
  NAND3_X1 U19291 ( .A1(n16135), .A2(n16134), .A3(n16133), .ZN(P2_U2901) );
  AOI22_X1 U19292 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n15077), .ZN(n16140) );
  AOI222_X1 U19293 ( .A1(n16138), .A2(n19264), .B1(n19263), .B2(n16137), .C1(
        n19260), .C2(n16136), .ZN(n16139) );
  OAI211_X1 U19294 ( .C1(n19269), .C2(n16141), .A(n16140), .B(n16139), .ZN(
        P2_U2992) );
  AOI22_X1 U19295 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n15077), .ZN(n16149) );
  INV_X1 U19296 ( .A(n18939), .ZN(n16147) );
  AOI21_X1 U19297 ( .B1(n16159), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16143) );
  NOR3_X1 U19298 ( .A1(n16143), .A2(n16142), .A3(n16219), .ZN(n16146) );
  NOR2_X1 U19299 ( .A1(n16144), .A2(n16220), .ZN(n16145) );
  AOI211_X1 U19300 ( .C1(n19263), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        n16148) );
  OAI211_X1 U19301 ( .C1(n19269), .C2(n18935), .A(n16149), .B(n16148), .ZN(
        P2_U2998) );
  AOI22_X1 U19302 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n12404), .B1(n16227), 
        .B2(n18949), .ZN(n16154) );
  OAI22_X1 U19303 ( .A1(n16151), .A2(n16220), .B1(n16219), .B2(n16150), .ZN(
        n16152) );
  AOI21_X1 U19304 ( .B1(n19263), .B2(n18952), .A(n16152), .ZN(n16153) );
  OAI211_X1 U19305 ( .C1(n16239), .C2(n18941), .A(n16154), .B(n16153), .ZN(
        P2_U2999) );
  AOI22_X1 U19306 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n12404), .ZN(n16162) );
  NAND2_X1 U19307 ( .A1(n16156), .A2(n16155), .ZN(n16157) );
  XNOR2_X1 U19308 ( .A(n16158), .B(n16157), .ZN(n16258) );
  INV_X1 U19309 ( .A(n18966), .ZN(n16257) );
  AOI21_X1 U19310 ( .B1(n16173), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16160) );
  NOR2_X1 U19311 ( .A1(n16160), .A2(n16159), .ZN(n16256) );
  AOI222_X1 U19312 ( .A1(n16258), .A2(n19264), .B1(n19263), .B2(n16257), .C1(
        n19260), .C2(n16256), .ZN(n16161) );
  AOI22_X1 U19313 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n12404), .B1(n16227), 
        .B2(n16163), .ZN(n16169) );
  OAI22_X1 U19314 ( .A1(n16165), .A2(n16219), .B1(n16164), .B2(n16220), .ZN(
        n16166) );
  AOI21_X1 U19315 ( .B1(n19263), .B2(n16167), .A(n16166), .ZN(n16168) );
  OAI211_X1 U19316 ( .C1(n16239), .C2(n16170), .A(n16169), .B(n16168), .ZN(
        P2_U3001) );
  AOI22_X1 U19317 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n15077), .ZN(n16178) );
  NAND2_X1 U19318 ( .A1(n16171), .A2(n19264), .ZN(n16175) );
  OR3_X1 U19319 ( .A1(n16173), .A2(n16172), .A3(n16219), .ZN(n16174) );
  OAI211_X1 U19320 ( .C1(n16214), .C2(n18977), .A(n16175), .B(n16174), .ZN(
        n16176) );
  INV_X1 U19321 ( .A(n16176), .ZN(n16177) );
  OAI211_X1 U19322 ( .C1(n19269), .C2(n18972), .A(n16178), .B(n16177), .ZN(
        P2_U3002) );
  AOI22_X1 U19323 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n12404), .B1(n16227), 
        .B2(n18984), .ZN(n16184) );
  INV_X1 U19324 ( .A(n16179), .ZN(n16181) );
  OAI22_X1 U19325 ( .A1(n16181), .A2(n16219), .B1(n16180), .B2(n16220), .ZN(
        n16182) );
  AOI21_X1 U19326 ( .B1(n19263), .B2(n18986), .A(n16182), .ZN(n16183) );
  OAI211_X1 U19327 ( .C1(n16239), .C2(n18978), .A(n16184), .B(n16183), .ZN(
        P2_U3003) );
  AOI22_X1 U19328 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n12404), .ZN(n16196) );
  NAND2_X1 U19329 ( .A1(n16186), .A2(n16185), .ZN(n16189) );
  NOR2_X1 U19330 ( .A1(n16187), .A2(n10084), .ZN(n16188) );
  XNOR2_X1 U19331 ( .A(n16189), .B(n16188), .ZN(n16278) );
  INV_X1 U19332 ( .A(n16278), .ZN(n16194) );
  AND2_X1 U19333 ( .A1(n16190), .A2(n16270), .ZN(n16191) );
  NOR2_X1 U19334 ( .A1(n16192), .A2(n16191), .ZN(n16275) );
  AOI222_X1 U19335 ( .A1(n16194), .A2(n19264), .B1(n19263), .B2(n16193), .C1(
        n19260), .C2(n16275), .ZN(n16195) );
  OAI211_X1 U19336 ( .C1(n19269), .C2(n18994), .A(n16196), .B(n16195), .ZN(
        P2_U3004) );
  AOI22_X1 U19337 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n12404), .B1(n16227), 
        .B2(n19007), .ZN(n16201) );
  OAI22_X1 U19338 ( .A1(n16198), .A2(n16220), .B1(n16219), .B2(n16197), .ZN(
        n16199) );
  AOI21_X1 U19339 ( .B1(n19263), .B2(n19009), .A(n16199), .ZN(n16200) );
  OAI211_X1 U19340 ( .C1(n16239), .C2(n19001), .A(n16201), .B(n16200), .ZN(
        P2_U3005) );
  AOI22_X1 U19341 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n15077), .ZN(n16217) );
  INV_X1 U19342 ( .A(n16202), .ZN(n16203) );
  XNOR2_X1 U19343 ( .A(n16204), .B(n16203), .ZN(n16282) );
  NAND2_X1 U19344 ( .A1(n16282), .A2(n19260), .ZN(n16213) );
  NAND2_X1 U19345 ( .A1(n16206), .A2(n16205), .ZN(n16211) );
  INV_X1 U19346 ( .A(n16207), .ZN(n16208) );
  NOR2_X1 U19347 ( .A1(n16209), .A2(n16208), .ZN(n16210) );
  XNOR2_X1 U19348 ( .A(n16211), .B(n16210), .ZN(n16286) );
  NAND2_X1 U19349 ( .A1(n16286), .A2(n19264), .ZN(n16212) );
  OAI211_X1 U19350 ( .C1(n16214), .C2(n19023), .A(n16213), .B(n16212), .ZN(
        n16215) );
  INV_X1 U19351 ( .A(n16215), .ZN(n16216) );
  OAI211_X1 U19352 ( .C1(n19269), .C2(n19017), .A(n16217), .B(n16216), .ZN(
        P2_U3006) );
  AOI22_X1 U19353 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n12404), .B1(n16227), 
        .B2(n19052), .ZN(n16224) );
  OAI22_X1 U19354 ( .A1(n16221), .A2(n16220), .B1(n16219), .B2(n16218), .ZN(
        n16222) );
  AOI21_X1 U19355 ( .B1(n19263), .B2(n19053), .A(n16222), .ZN(n16223) );
  OAI211_X1 U19356 ( .C1(n16239), .C2(n16225), .A(n16224), .B(n16223), .ZN(
        P2_U3009) );
  AOI22_X1 U19357 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n12404), .B1(n16227), 
        .B2(n16226), .ZN(n16238) );
  OAI21_X1 U19358 ( .B1(n16230), .B2(n16229), .A(n16228), .ZN(n16308) );
  INV_X1 U19359 ( .A(n16308), .ZN(n16236) );
  XNOR2_X1 U19360 ( .A(n16232), .B(n16231), .ZN(n16233) );
  XNOR2_X1 U19361 ( .A(n9718), .B(n16233), .ZN(n16316) );
  INV_X1 U19362 ( .A(n16316), .ZN(n16235) );
  AOI222_X1 U19363 ( .A1(n10640), .A2(n19263), .B1(n19260), .B2(n16236), .C1(
        n16235), .C2(n19264), .ZN(n16237) );
  OAI211_X1 U19364 ( .C1(n16240), .C2(n16239), .A(n16238), .B(n16237), .ZN(
        P2_U3011) );
  AOI221_X1 U19365 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C1(n16244), .C2(n16242), .A(
        n16241), .ZN(n16247) );
  OAI22_X1 U19366 ( .A1(n16245), .A2(n16244), .B1(n16306), .B2(n16243), .ZN(
        n16246) );
  AOI211_X1 U19367 ( .C1(n15077), .C2(P2_REIP_REG_23__SCAN_IN), .A(n16247), 
        .B(n16246), .ZN(n16251) );
  AOI22_X1 U19368 ( .A1(n16249), .A2(n16301), .B1(n12589), .B2(n16248), .ZN(
        n16250) );
  OAI211_X1 U19369 ( .C1(n16307), .C2(n16252), .A(n16251), .B(n16250), .ZN(
        P2_U3023) );
  AOI21_X1 U19370 ( .B1(n16254), .B2(n16253), .A(n15280), .ZN(n19116) );
  AOI22_X1 U19371 ( .A1(n16255), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16281), .B2(n19116), .ZN(n16265) );
  AOI222_X1 U19372 ( .A1(n16258), .A2(n16301), .B1(n12589), .B2(n16257), .C1(
        n16274), .C2(n16256), .ZN(n16264) );
  NAND2_X1 U19373 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n12404), .ZN(n16263) );
  OAI211_X1 U19374 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16261), .A(
        n16260), .B(n16259), .ZN(n16262) );
  NAND4_X1 U19375 ( .A1(n16265), .A2(n16264), .A3(n16263), .A4(n16262), .ZN(
        P2_U3032) );
  AOI21_X1 U19376 ( .B1(n16267), .B2(n16266), .A(n15333), .ZN(n19123) );
  NAND2_X1 U19377 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n15077), .ZN(n16268) );
  OAI221_X1 U19378 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16271), 
        .C1(n16270), .C2(n16269), .A(n16268), .ZN(n16272) );
  AOI21_X1 U19379 ( .B1(n16281), .B2(n19123), .A(n16272), .ZN(n16277) );
  NOR2_X1 U19380 ( .A1(n16283), .A2(n18999), .ZN(n16273) );
  AOI21_X1 U19381 ( .B1(n16275), .B2(n16274), .A(n16273), .ZN(n16276) );
  OAI211_X1 U19382 ( .C1(n16278), .C2(n16315), .A(n16277), .B(n16276), .ZN(
        P2_U3036) );
  AOI21_X1 U19383 ( .B1(n16280), .B2(n16293), .A(n16279), .ZN(n19127) );
  AOI22_X1 U19384 ( .A1(n16299), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16281), .B2(n19127), .ZN(n16292) );
  INV_X1 U19385 ( .A(n16282), .ZN(n16284) );
  OAI22_X1 U19386 ( .A1(n16284), .A2(n16307), .B1(n16283), .B2(n19023), .ZN(
        n16285) );
  AOI21_X1 U19387 ( .B1(n16301), .B2(n16286), .A(n16285), .ZN(n16291) );
  NAND2_X1 U19388 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n15077), .ZN(n16290) );
  INV_X1 U19389 ( .A(n16287), .ZN(n16298) );
  OAI211_X1 U19390 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16298), .B(n16288), .ZN(n16289) );
  NAND4_X1 U19391 ( .A1(n16292), .A2(n16291), .A3(n16290), .A4(n16289), .ZN(
        P2_U3038) );
  OAI21_X1 U19392 ( .B1(n16295), .B2(n16294), .A(n16293), .ZN(n19131) );
  OAI22_X1 U19393 ( .A1(n19131), .A2(n16306), .B1(n19863), .B2(n9722), .ZN(
        n16296) );
  AOI221_X1 U19394 ( .B1(n16299), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n16298), .C2(n16297), .A(n16296), .ZN(n16304) );
  INV_X1 U19395 ( .A(n19029), .ZN(n16300) );
  AOI22_X1 U19396 ( .A1(n16302), .A2(n16301), .B1(n12589), .B2(n16300), .ZN(
        n16303) );
  OAI211_X1 U19397 ( .C1(n16307), .C2(n16305), .A(n16304), .B(n16303), .ZN(
        P2_U3039) );
  OAI22_X1 U19398 ( .A1(n19923), .A2(n16306), .B1(n11214), .B2(n9722), .ZN(
        n16310) );
  NOR2_X1 U19399 ( .A1(n16308), .A2(n16307), .ZN(n16309) );
  AOI211_X1 U19400 ( .C1(n12589), .C2(n10640), .A(n16310), .B(n16309), .ZN(
        n16314) );
  OAI21_X1 U19401 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16312), .A(
        n16311), .ZN(n16313) );
  OAI211_X1 U19402 ( .C1(n16316), .C2(n16315), .A(n16314), .B(n16313), .ZN(
        P2_U3043) );
  NAND2_X1 U19403 ( .A1(n16317), .A2(n16359), .ZN(n16320) );
  INV_X1 U19404 ( .A(n16359), .ZN(n16322) );
  NAND2_X1 U19405 ( .A1(n16322), .A2(n16318), .ZN(n16319) );
  NAND2_X1 U19406 ( .A1(n16320), .A2(n16319), .ZN(n16338) );
  NOR2_X1 U19407 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19382) );
  INV_X1 U19408 ( .A(n19382), .ZN(n19349) );
  OR2_X1 U19409 ( .A1(n16321), .A2(n16322), .ZN(n16324) );
  NAND2_X1 U19410 ( .A1(n16322), .A2(n10470), .ZN(n16323) );
  NAND2_X1 U19411 ( .A1(n16324), .A2(n16323), .ZN(n16333) );
  NAND2_X1 U19412 ( .A1(n16333), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16332) );
  NAND2_X1 U19413 ( .A1(n16325), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16329) );
  NAND2_X1 U19414 ( .A1(n16329), .A2(n19943), .ZN(n16327) );
  NAND2_X1 U19415 ( .A1(n16327), .A2(n16326), .ZN(n16328) );
  OAI211_X1 U19416 ( .C1(n19943), .C2(n16329), .A(n16328), .B(n16359), .ZN(
        n16330) );
  AOI21_X1 U19417 ( .B1(n16338), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16330), .ZN(n16331) );
  NAND2_X1 U19418 ( .A1(n16332), .A2(n16331), .ZN(n16335) );
  INV_X1 U19419 ( .A(n16333), .ZN(n16362) );
  NAND2_X1 U19420 ( .A1(n16362), .A2(n19926), .ZN(n16334) );
  OAI211_X1 U19421 ( .C1(n16338), .C2(n19349), .A(n16335), .B(n16334), .ZN(
        n16337) );
  NAND2_X1 U19422 ( .A1(n16337), .A2(n16336), .ZN(n16364) );
  INV_X1 U19423 ( .A(n16338), .ZN(n16361) );
  INV_X1 U19424 ( .A(n16339), .ZN(n16340) );
  AOI22_X1 U19425 ( .A1(n16344), .A2(n16341), .B1(n11186), .B2(n16340), .ZN(
        n16342) );
  OAI21_X1 U19426 ( .B1(n16344), .B2(n16343), .A(n16342), .ZN(n19959) );
  INV_X1 U19427 ( .A(n19959), .ZN(n16357) );
  NOR2_X1 U19428 ( .A1(n16346), .A2(n16345), .ZN(n16347) );
  AND2_X1 U19429 ( .A1(n16348), .A2(n16347), .ZN(n18874) );
  INV_X1 U19430 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n16349) );
  NAND2_X1 U19431 ( .A1(n18876), .A2(n16349), .ZN(n16355) );
  NAND2_X1 U19432 ( .A1(n19283), .A2(n16350), .ZN(n16352) );
  OAI22_X1 U19433 ( .A1(n9710), .A2(n16352), .B1(n10982), .B2(n16351), .ZN(
        n16354) );
  AOI21_X1 U19434 ( .B1(n18874), .B2(n16355), .A(n16354), .ZN(n16356) );
  OAI211_X1 U19435 ( .C1(n16359), .C2(n16358), .A(n16357), .B(n16356), .ZN(
        n16360) );
  AOI21_X1 U19436 ( .B1(n16362), .B2(n16361), .A(n16360), .ZN(n16363) );
  NAND2_X1 U19437 ( .A1(n16364), .A2(n16363), .ZN(n16371) );
  AOI211_X1 U19438 ( .C1(n16367), .C2(n16371), .A(n16366), .B(n16365), .ZN(
        n16376) );
  OR2_X1 U19439 ( .A1(n19963), .A2(n19973), .ZN(n16368) );
  AOI21_X1 U19440 ( .B1(n10553), .B2(n16369), .A(n16368), .ZN(n16372) );
  INV_X1 U19441 ( .A(n19822), .ZN(n19974) );
  AOI22_X1 U19442 ( .A1(n16370), .A2(n19975), .B1(n16372), .B2(n19974), .ZN(
        n16374) );
  OAI21_X1 U19443 ( .B1(n16371), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16373) );
  AND2_X1 U19444 ( .A1(n16373), .A2(n16372), .ZN(n19824) );
  INV_X1 U19445 ( .A(n19824), .ZN(n19821) );
  NAND2_X1 U19446 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19821), .ZN(n16377) );
  OAI21_X1 U19447 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16374), .A(n16377), 
        .ZN(n16375) );
  OAI211_X1 U19448 ( .C1(n19956), .C2(n16378), .A(n16376), .B(n16375), .ZN(
        P2_U3176) );
  INV_X1 U19449 ( .A(n16377), .ZN(n16379) );
  OAI21_X1 U19450 ( .B1(n16379), .B2(n19533), .A(n16378), .ZN(P2_U3593) );
  NOR2_X1 U19451 ( .A1(n16391), .A2(n16381), .ZN(n16400) );
  NAND2_X1 U19452 ( .A1(n16400), .A2(n16401), .ZN(n17756) );
  NOR2_X1 U19453 ( .A1(n17786), .A2(n16382), .ZN(n16390) );
  OAI21_X1 U19454 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17786), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16383) );
  OAI221_X1 U19455 ( .B1(n16413), .B2(n16384), .C1(n17786), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16383), .ZN(n16389) );
  OAI21_X1 U19456 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16413), .A(
        n16384), .ZN(n16387) );
  NAND2_X1 U19457 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17786), .ZN(
        n16385) );
  OAI22_X1 U19458 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17786), .B1(
        n16385), .B2(n16413), .ZN(n16386) );
  OAI21_X1 U19459 ( .B1(n16390), .B2(n16387), .A(n16386), .ZN(n16388) );
  OAI21_X1 U19460 ( .B1(n16390), .B2(n16389), .A(n16388), .ZN(n16439) );
  INV_X1 U19461 ( .A(n16791), .ZN(n16869) );
  NOR2_X1 U19462 ( .A1(n18162), .A2(n18792), .ZN(n16437) );
  NAND2_X1 U19463 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17639) );
  NAND2_X1 U19464 ( .A1(n17655), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17638) );
  NOR2_X1 U19465 ( .A1(n17639), .A2(n17638), .ZN(n17617) );
  NAND2_X1 U19466 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17617), .ZN(
        n17590) );
  NOR3_X1 U19467 ( .A1(n17600), .A2(n9872), .A3(n17590), .ZN(n17548) );
  NAND3_X1 U19468 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(n17548), .ZN(n17536) );
  NOR2_X1 U19469 ( .A1(n17537), .A2(n17536), .ZN(n17514) );
  NAND3_X1 U19470 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(n17514), .ZN(n16424) );
  NOR2_X1 U19471 ( .A1(n16392), .A2(n16424), .ZN(n16393) );
  NOR2_X1 U19472 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18862), .ZN(n17712) );
  INV_X1 U19473 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17867) );
  OAI21_X1 U19474 ( .B1(n17618), .B2(n17867), .A(n18221), .ZN(n17707) );
  NAND2_X1 U19475 ( .A1(n16393), .A2(n17707), .ZN(n16406) );
  INV_X1 U19476 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16395) );
  XOR2_X1 U19477 ( .A(n16395), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16396) );
  NOR2_X1 U19478 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17618), .ZN(
        n16421) );
  INV_X1 U19479 ( .A(n17712), .ZN(n17668) );
  OR2_X1 U19480 ( .A1(n18221), .A2(n16393), .ZN(n16425) );
  OAI211_X1 U19481 ( .C1(n16394), .C2(n17668), .A(n16425), .B(n17872), .ZN(
        n16420) );
  NOR2_X1 U19482 ( .A1(n16421), .A2(n16420), .ZN(n16407) );
  OAI22_X1 U19483 ( .A1(n16406), .A2(n16396), .B1(n16407), .B2(n16395), .ZN(
        n16397) );
  AOI211_X1 U19484 ( .C1(n16869), .C2(n17729), .A(n16437), .B(n16397), .ZN(
        n16404) );
  NOR2_X2 U19485 ( .A1(n16398), .A2(n16555), .ZN(n17824) );
  INV_X1 U19486 ( .A(n16417), .ZN(n16410) );
  NAND2_X1 U19487 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16410), .ZN(
        n16399) );
  XNOR2_X1 U19488 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16399), .ZN(
        n16434) );
  NAND2_X1 U19489 ( .A1(n16419), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16402) );
  XNOR2_X1 U19490 ( .A(n16402), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16433) );
  AOI22_X1 U19491 ( .A1(n17824), .A2(n16434), .B1(n17788), .B2(n16433), .ZN(
        n16403) );
  OAI211_X1 U19492 ( .C1(n17756), .C2(n16439), .A(n16404), .B(n16403), .ZN(
        P3_U2799) );
  INV_X1 U19493 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16405) );
  AOI22_X1 U19494 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16407), .B1(
        n16406), .B2(n16405), .ZN(n16408) );
  AOI211_X1 U19495 ( .C1(n17729), .C2(n16573), .A(n16409), .B(n16408), .ZN(
        n16416) );
  OAI22_X1 U19496 ( .A1(n16410), .A2(n17877), .B1(n16419), .B2(n17748), .ZN(
        n16412) );
  AOI22_X1 U19497 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16412), .B1(
        n17787), .B2(n16411), .ZN(n16415) );
  INV_X1 U19498 ( .A(n17749), .ZN(n18062) );
  OAI22_X1 U19499 ( .A1(n18063), .A2(n17877), .B1(n17748), .B2(n18062), .ZN(
        n17722) );
  NAND2_X1 U19500 ( .A1(n16453), .A2(n17722), .ZN(n17613) );
  NOR2_X1 U19501 ( .A1(n16455), .A2(n17613), .ZN(n17530) );
  NAND3_X1 U19502 ( .A1(n16436), .A2(n17530), .A3(n16413), .ZN(n16414) );
  NAND3_X1 U19503 ( .A1(n16416), .A2(n16415), .A3(n16414), .ZN(P3_U2800) );
  NAND2_X1 U19504 ( .A1(n17824), .A2(n16417), .ZN(n16431) );
  NAND2_X1 U19505 ( .A1(n17881), .A2(n16418), .ZN(n16444) );
  AOI211_X1 U19506 ( .C1(n16430), .C2(n16443), .A(n16419), .B(n17748), .ZN(
        n16427) );
  AOI22_X1 U19507 ( .A1(n9724), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16420), .ZN(n16423) );
  OAI21_X1 U19508 ( .B1(n17729), .B2(n16421), .A(n16582), .ZN(n16422) );
  OAI211_X1 U19509 ( .C1(n16425), .C2(n16424), .A(n16423), .B(n16422), .ZN(
        n16426) );
  AOI211_X1 U19510 ( .C1(n17787), .C2(n16428), .A(n16427), .B(n16426), .ZN(
        n16429) );
  OAI221_X1 U19511 ( .B1(n16431), .B2(n16430), .C1(n16431), .C2(n16444), .A(
        n16429), .ZN(P3_U2801) );
  OAI211_X1 U19512 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18134), .A(
        n16432), .B(n18133), .ZN(n16438) );
  INV_X1 U19513 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18808) );
  AOI21_X1 U19514 ( .B1(n17786), .B2(n17521), .A(n17520), .ZN(n17510) );
  NAND2_X1 U19515 ( .A1(n16441), .A2(n16440), .ZN(n17509) );
  NOR2_X1 U19516 ( .A1(n17510), .A2(n17509), .ZN(n17508) );
  NOR3_X1 U19517 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17508), .A3(
        n16447), .ZN(n16442) );
  OAI221_X1 U19518 ( .B1(n16442), .B2(n17520), .C1(n16442), .C2(n17509), .A(
        n18096), .ZN(n16458) );
  AOI22_X1 U19519 ( .A1(n18633), .A2(n16444), .B1(n18099), .B2(n16443), .ZN(
        n16449) );
  NOR2_X1 U19520 ( .A1(n17349), .A2(n18639), .ZN(n16446) );
  INV_X1 U19521 ( .A(n17508), .ZN(n16445) );
  OAI211_X1 U19522 ( .C1(n17521), .C2(n16447), .A(n16446), .B(n16445), .ZN(
        n16448) );
  NAND4_X1 U19523 ( .A1(n18169), .A2(n16450), .A3(n16449), .A4(n16448), .ZN(
        n16451) );
  NAND3_X1 U19524 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n13328), .A3(
        n16451), .ZN(n16457) );
  NAND2_X1 U19525 ( .A1(n9724), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17517) );
  INV_X1 U19526 ( .A(n16452), .ZN(n18146) );
  INV_X1 U19527 ( .A(n16453), .ZN(n17938) );
  AOI22_X1 U19528 ( .A1(n18633), .A2(n17747), .B1(n17749), .B2(n18099), .ZN(
        n18035) );
  OAI222_X1 U19529 ( .A1(n18146), .A2(n16454), .B1(n17938), .B2(n18035), .C1(
        n18144), .C2(n17932), .ZN(n17924) );
  NAND2_X1 U19530 ( .A1(n18169), .A2(n17924), .ZN(n17985) );
  NOR2_X1 U19531 ( .A1(n16455), .A2(n17985), .ZN(n17886) );
  NAND3_X1 U19532 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17886), .A3(
        n17506), .ZN(n16456) );
  NAND4_X1 U19533 ( .A1(n16458), .A2(n16457), .A3(n17517), .A4(n16456), .ZN(
        P3_U2834) );
  NOR3_X1 U19534 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16460) );
  NOR4_X1 U19535 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16459) );
  NAND4_X1 U19536 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16460), .A3(n16459), .A4(
        U215), .ZN(U213) );
  INV_X1 U19537 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19167) );
  INV_X2 U19538 ( .A(U214), .ZN(n16509) );
  NOR2_X2 U19539 ( .A1(n16509), .A2(n16461), .ZN(n16502) );
  OAI222_X1 U19540 ( .A1(U212), .A2(n19167), .B1(n16511), .B2(n16462), .C1(
        U214), .C2(n16541), .ZN(U216) );
  AOI222_X1 U19541 ( .A1(n16508), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16502), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16509), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n16463) );
  INV_X1 U19542 ( .A(n16463), .ZN(U217) );
  INV_X1 U19543 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16465) );
  AOI22_X1 U19544 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16508), .ZN(n16464) );
  OAI21_X1 U19545 ( .B1(n16465), .B2(n16511), .A(n16464), .ZN(U218) );
  INV_X1 U19546 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n16467) );
  OAI222_X1 U19547 ( .A1(U214), .A2(n16467), .B1(n16511), .B2(n16466), .C1(
        U212), .C2(n16537), .ZN(U219) );
  AOI22_X1 U19548 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16508), .ZN(n16468) );
  OAI21_X1 U19549 ( .B1(n16469), .B2(n16511), .A(n16468), .ZN(U220) );
  INV_X1 U19550 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n16471) );
  OAI222_X1 U19551 ( .A1(U214), .A2(n16471), .B1(n16511), .B2(n16470), .C1(
        U212), .C2(n19172), .ZN(U221) );
  INV_X1 U19552 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16473) );
  AOI22_X1 U19553 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16508), .ZN(n16472) );
  OAI21_X1 U19554 ( .B1(n16473), .B2(n16511), .A(n16472), .ZN(U222) );
  AOI22_X1 U19555 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16508), .ZN(n16474) );
  OAI21_X1 U19556 ( .B1(n16475), .B2(n16511), .A(n16474), .ZN(U223) );
  AOI222_X1 U19557 ( .A1(n16509), .A2(P1_DATAO_REG_23__SCAN_IN), .B1(n16502), 
        .B2(BUF1_REG_23__SCAN_IN), .C1(n16508), .C2(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n16476) );
  INV_X1 U19558 ( .A(n16476), .ZN(U224) );
  AOI22_X1 U19559 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16508), .ZN(n16477) );
  OAI21_X1 U19560 ( .B1(n14643), .B2(n16511), .A(n16477), .ZN(U225) );
  AOI222_X1 U19561 ( .A1(n16509), .A2(P1_DATAO_REG_21__SCAN_IN), .B1(n16502), 
        .B2(BUF1_REG_21__SCAN_IN), .C1(n16508), .C2(P2_DATAO_REG_21__SCAN_IN), 
        .ZN(n16478) );
  INV_X1 U19562 ( .A(n16478), .ZN(U226) );
  AOI22_X1 U19563 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16508), .ZN(n16479) );
  OAI21_X1 U19564 ( .B1(n16480), .B2(n16511), .A(n16479), .ZN(U227) );
  INV_X1 U19565 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U19566 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16508), .ZN(n16481) );
  OAI21_X1 U19567 ( .B1(n16482), .B2(n16511), .A(n16481), .ZN(U228) );
  AOI222_X1 U19568 ( .A1(n16509), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n16502), 
        .B2(BUF1_REG_18__SCAN_IN), .C1(n16508), .C2(P2_DATAO_REG_18__SCAN_IN), 
        .ZN(n16483) );
  INV_X1 U19569 ( .A(n16483), .ZN(U229) );
  INV_X1 U19570 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16485) );
  AOI22_X1 U19571 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16508), .ZN(n16484) );
  OAI21_X1 U19572 ( .B1(n16485), .B2(n16511), .A(n16484), .ZN(U230) );
  AOI22_X1 U19573 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16508), .ZN(n16486) );
  OAI21_X1 U19574 ( .B1(n14672), .B2(n16511), .A(n16486), .ZN(U231) );
  AOI22_X1 U19575 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16502), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16509), .ZN(n16487) );
  OAI21_X1 U19576 ( .B1(n19178), .B2(U212), .A(n16487), .ZN(U232) );
  INV_X1 U19577 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16524) );
  AOI22_X1 U19578 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16502), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16509), .ZN(n16488) );
  OAI21_X1 U19579 ( .B1(n16524), .B2(U212), .A(n16488), .ZN(U233) );
  AOI22_X1 U19580 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16508), .ZN(n16489) );
  OAI21_X1 U19581 ( .B1(n16490), .B2(n16511), .A(n16489), .ZN(U234) );
  INV_X1 U19582 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16522) );
  AOI22_X1 U19583 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16502), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16509), .ZN(n16491) );
  OAI21_X1 U19584 ( .B1(n16522), .B2(U212), .A(n16491), .ZN(U235) );
  OAI222_X1 U19585 ( .A1(U212), .A2(n19187), .B1(n16511), .B2(n14969), .C1(
        U214), .C2(n20122), .ZN(U236) );
  AOI222_X1 U19586 ( .A1(n16509), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n16502), 
        .B2(BUF1_REG_10__SCAN_IN), .C1(n16508), .C2(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n16492) );
  INV_X1 U19587 ( .A(n16492), .ZN(U237) );
  INV_X1 U19588 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16521) );
  AOI22_X1 U19589 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16502), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16509), .ZN(n16493) );
  OAI21_X1 U19590 ( .B1(n16521), .B2(U212), .A(n16493), .ZN(U238) );
  INV_X1 U19591 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16495) );
  AOI22_X1 U19592 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16508), .ZN(n16494) );
  OAI21_X1 U19593 ( .B1(n16495), .B2(n16511), .A(n16494), .ZN(U239) );
  INV_X1 U19594 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16519) );
  AOI22_X1 U19595 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16502), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16509), .ZN(n16496) );
  OAI21_X1 U19596 ( .B1(n16519), .B2(U212), .A(n16496), .ZN(U240) );
  INV_X1 U19597 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16498) );
  AOI22_X1 U19598 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16508), .ZN(n16497) );
  OAI21_X1 U19599 ( .B1(n16498), .B2(n16511), .A(n16497), .ZN(U241) );
  AOI22_X1 U19600 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16502), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16508), .ZN(n16499) );
  OAI21_X1 U19601 ( .B1(n20134), .B2(U214), .A(n16499), .ZN(U242) );
  INV_X1 U19602 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16501) );
  AOI22_X1 U19603 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16508), .ZN(n16500) );
  OAI21_X1 U19604 ( .B1(n16501), .B2(n16511), .A(n16500), .ZN(U243) );
  AOI22_X1 U19605 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16502), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16509), .ZN(n16503) );
  OAI21_X1 U19606 ( .B1(n19206), .B2(U212), .A(n16503), .ZN(U244) );
  AOI22_X1 U19607 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16508), .ZN(n16504) );
  OAI21_X1 U19608 ( .B1(n16505), .B2(n16511), .A(n16504), .ZN(U245) );
  AOI22_X1 U19609 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16508), .ZN(n16506) );
  OAI21_X1 U19610 ( .B1(n16507), .B2(n16511), .A(n16506), .ZN(U246) );
  AOI22_X1 U19611 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16509), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16508), .ZN(n16510) );
  OAI21_X1 U19612 ( .B1(n16512), .B2(n16511), .A(n16510), .ZN(U247) );
  INV_X1 U19613 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16513) );
  AOI22_X1 U19614 ( .A1(n16540), .A2(n16513), .B1(n18186), .B2(U215), .ZN(U251) );
  OAI22_X1 U19615 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16540), .ZN(n16514) );
  INV_X1 U19616 ( .A(n16514), .ZN(U252) );
  INV_X1 U19617 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16515) );
  AOI22_X1 U19618 ( .A1(n16540), .A2(n16515), .B1(n18198), .B2(U215), .ZN(U253) );
  INV_X1 U19619 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18203) );
  AOI22_X1 U19620 ( .A1(n16540), .A2(n19206), .B1(n18203), .B2(U215), .ZN(U254) );
  INV_X1 U19621 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16516) );
  INV_X1 U19622 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18207) );
  AOI22_X1 U19623 ( .A1(n16540), .A2(n16516), .B1(n18207), .B2(U215), .ZN(U255) );
  INV_X1 U19624 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16517) );
  INV_X1 U19625 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18212) );
  AOI22_X1 U19626 ( .A1(n16540), .A2(n16517), .B1(n18212), .B2(U215), .ZN(U256) );
  INV_X1 U19627 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16518) );
  INV_X1 U19628 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U19629 ( .A1(n16540), .A2(n16518), .B1(n18216), .B2(U215), .ZN(U257) );
  AOI22_X1 U19630 ( .A1(n16540), .A2(n16519), .B1(n18223), .B2(U215), .ZN(U258) );
  INV_X1 U19631 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16520) );
  INV_X1 U19632 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U19633 ( .A1(n16534), .A2(n16520), .B1(n17484), .B2(U215), .ZN(U259) );
  AOI22_X1 U19634 ( .A1(n16540), .A2(n16521), .B1(n17486), .B2(U215), .ZN(U260) );
  AOI22_X1 U19635 ( .A1(n16534), .A2(n19190), .B1(n17488), .B2(U215), .ZN(U261) );
  AOI22_X1 U19636 ( .A1(n16534), .A2(n19187), .B1(n17490), .B2(U215), .ZN(U262) );
  INV_X1 U19637 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U19638 ( .A1(n16540), .A2(n16522), .B1(n17492), .B2(U215), .ZN(U263) );
  OAI22_X1 U19639 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16534), .ZN(n16523) );
  INV_X1 U19640 ( .A(n16523), .ZN(U264) );
  INV_X1 U19641 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U19642 ( .A1(n16534), .A2(n16524), .B1(n17498), .B2(U215), .ZN(U265) );
  INV_X1 U19643 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n16525) );
  AOI22_X1 U19644 ( .A1(n16540), .A2(n19178), .B1(n16525), .B2(U215), .ZN(U266) );
  OAI22_X1 U19645 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16540), .ZN(n16526) );
  INV_X1 U19646 ( .A(n16526), .ZN(U267) );
  OAI22_X1 U19647 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16540), .ZN(n16527) );
  INV_X1 U19648 ( .A(n16527), .ZN(U268) );
  INV_X1 U19649 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18197) );
  AOI22_X1 U19650 ( .A1(n16534), .A2(n19175), .B1(n18197), .B2(U215), .ZN(U269) );
  INV_X1 U19651 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16528) );
  AOI22_X1 U19652 ( .A1(n16540), .A2(n16528), .B1(n18202), .B2(U215), .ZN(U270) );
  OAI22_X1 U19653 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16540), .ZN(n16529) );
  INV_X1 U19654 ( .A(n16529), .ZN(U271) );
  INV_X1 U19655 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18211) );
  AOI22_X1 U19656 ( .A1(n16534), .A2(n16530), .B1(n18211), .B2(U215), .ZN(U272) );
  INV_X1 U19657 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16531) );
  INV_X1 U19658 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n17279) );
  AOI22_X1 U19659 ( .A1(n16534), .A2(n16531), .B1(n17279), .B2(U215), .ZN(U273) );
  AOI22_X1 U19660 ( .A1(n16540), .A2(n16532), .B1(n18222), .B2(U215), .ZN(U274) );
  OAI22_X1 U19661 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16534), .ZN(n16533) );
  INV_X1 U19662 ( .A(n16533), .ZN(U275) );
  OAI22_X1 U19663 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16534), .ZN(n16535) );
  INV_X1 U19664 ( .A(n16535), .ZN(U276) );
  INV_X1 U19665 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18196) );
  AOI22_X1 U19666 ( .A1(n16540), .A2(n19172), .B1(n18196), .B2(U215), .ZN(U277) );
  OAI22_X1 U19667 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16540), .ZN(n16536) );
  INV_X1 U19668 ( .A(n16536), .ZN(U278) );
  INV_X1 U19669 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17253) );
  AOI22_X1 U19670 ( .A1(n16540), .A2(n16537), .B1(n17253), .B2(U215), .ZN(U279) );
  OAI22_X1 U19671 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16540), .ZN(n16538) );
  INV_X1 U19672 ( .A(n16538), .ZN(U280) );
  OAI22_X1 U19673 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16540), .ZN(n16539) );
  INV_X1 U19674 ( .A(n16539), .ZN(U281) );
  INV_X1 U19675 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18220) );
  AOI22_X1 U19676 ( .A1(n16540), .A2(n19167), .B1(n18220), .B2(U215), .ZN(U282) );
  INV_X1 U19677 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17386) );
  AOI222_X1 U19678 ( .A1(n16541), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19167), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17386), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16542) );
  INV_X2 U19679 ( .A(n16544), .ZN(n16543) );
  INV_X1 U19680 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18748) );
  INV_X1 U19681 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U19682 ( .A1(n16543), .A2(n18748), .B1(n19868), .B2(n16544), .ZN(
        U347) );
  INV_X1 U19683 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18746) );
  INV_X1 U19684 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19867) );
  AOI22_X1 U19685 ( .A1(n16543), .A2(n18746), .B1(n19867), .B2(n16544), .ZN(
        U348) );
  INV_X1 U19686 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18744) );
  AOI22_X1 U19687 ( .A1(n16543), .A2(n18744), .B1(n19866), .B2(n16544), .ZN(
        U349) );
  INV_X1 U19688 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18742) );
  INV_X1 U19689 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U19690 ( .A1(n16543), .A2(n18742), .B1(n19864), .B2(n16544), .ZN(
        U350) );
  INV_X1 U19691 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18740) );
  INV_X1 U19692 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19862) );
  AOI22_X1 U19693 ( .A1(n16543), .A2(n18740), .B1(n19862), .B2(n16544), .ZN(
        U351) );
  INV_X1 U19694 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18738) );
  INV_X1 U19695 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19860) );
  AOI22_X1 U19696 ( .A1(n16543), .A2(n18738), .B1(n19860), .B2(n16544), .ZN(
        U352) );
  INV_X1 U19697 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18736) );
  INV_X1 U19698 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19858) );
  AOI22_X1 U19699 ( .A1(n16543), .A2(n18736), .B1(n19858), .B2(n16544), .ZN(
        U353) );
  INV_X1 U19700 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18734) );
  AOI22_X1 U19701 ( .A1(n16543), .A2(n18734), .B1(n19857), .B2(n16544), .ZN(
        U354) );
  INV_X1 U19702 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18793) );
  INV_X1 U19703 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19899) );
  AOI22_X1 U19704 ( .A1(n16543), .A2(n18793), .B1(n19899), .B2(n16544), .ZN(
        U355) );
  INV_X1 U19705 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18789) );
  INV_X1 U19706 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U19707 ( .A1(n16543), .A2(n18789), .B1(n19897), .B2(n16544), .ZN(
        U356) );
  INV_X1 U19708 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18784) );
  INV_X1 U19709 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19895) );
  AOI22_X1 U19710 ( .A1(n16543), .A2(n18784), .B1(n19895), .B2(n16544), .ZN(
        U357) );
  INV_X1 U19711 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18783) );
  INV_X1 U19712 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19892) );
  AOI22_X1 U19713 ( .A1(n16543), .A2(n18783), .B1(n19892), .B2(n16544), .ZN(
        U358) );
  INV_X1 U19714 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18781) );
  INV_X1 U19715 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U19716 ( .A1(n16543), .A2(n18781), .B1(n19891), .B2(n16544), .ZN(
        U359) );
  INV_X1 U19717 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U19718 ( .A1(n16543), .A2(n18779), .B1(n19890), .B2(n16544), .ZN(
        U360) );
  INV_X1 U19719 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18777) );
  INV_X1 U19720 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19888) );
  AOI22_X1 U19721 ( .A1(n16543), .A2(n18777), .B1(n19888), .B2(n16544), .ZN(
        U361) );
  INV_X1 U19722 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18775) );
  INV_X1 U19723 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U19724 ( .A1(n16543), .A2(n18775), .B1(n19887), .B2(n16544), .ZN(
        U362) );
  INV_X1 U19725 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18773) );
  INV_X1 U19726 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U19727 ( .A1(n16543), .A2(n18773), .B1(n19885), .B2(n16544), .ZN(
        U363) );
  INV_X1 U19728 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18770) );
  INV_X1 U19729 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U19730 ( .A1(n16543), .A2(n18770), .B1(n19884), .B2(n16544), .ZN(
        U364) );
  INV_X1 U19731 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19856) );
  AOI22_X1 U19732 ( .A1(n16543), .A2(n18732), .B1(n19856), .B2(n16544), .ZN(
        U365) );
  INV_X1 U19733 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19882) );
  AOI22_X1 U19734 ( .A1(n16543), .A2(n18768), .B1(n19882), .B2(n16544), .ZN(
        U366) );
  INV_X1 U19735 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18767) );
  INV_X1 U19736 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U19737 ( .A1(n16543), .A2(n18767), .B1(n19881), .B2(n16544), .ZN(
        U367) );
  INV_X1 U19738 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18765) );
  INV_X1 U19739 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U19740 ( .A1(n16543), .A2(n18765), .B1(n19879), .B2(n16544), .ZN(
        U368) );
  INV_X1 U19741 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18762) );
  INV_X1 U19742 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19878) );
  AOI22_X1 U19743 ( .A1(n16543), .A2(n18762), .B1(n19878), .B2(n16544), .ZN(
        U369) );
  INV_X1 U19744 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18760) );
  INV_X1 U19745 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19876) );
  AOI22_X1 U19746 ( .A1(n16543), .A2(n18760), .B1(n19876), .B2(n16544), .ZN(
        U370) );
  INV_X1 U19747 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18759) );
  INV_X1 U19748 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19875) );
  AOI22_X1 U19749 ( .A1(n16543), .A2(n18759), .B1(n19875), .B2(n16544), .ZN(
        U371) );
  INV_X1 U19750 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18756) );
  INV_X1 U19751 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U19752 ( .A1(n16543), .A2(n18756), .B1(n19874), .B2(n16544), .ZN(
        U372) );
  INV_X1 U19753 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18754) );
  AOI22_X1 U19754 ( .A1(n16543), .A2(n18754), .B1(n19872), .B2(n16544), .ZN(
        U373) );
  INV_X1 U19755 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18752) );
  INV_X1 U19756 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19870) );
  AOI22_X1 U19757 ( .A1(n16543), .A2(n18752), .B1(n19870), .B2(n16544), .ZN(
        U374) );
  INV_X1 U19758 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18750) );
  INV_X1 U19759 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19869) );
  AOI22_X1 U19760 ( .A1(n16543), .A2(n18750), .B1(n19869), .B2(n16544), .ZN(
        U375) );
  INV_X1 U19761 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18731) );
  INV_X1 U19762 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19854) );
  AOI22_X1 U19763 ( .A1(n16543), .A2(n18731), .B1(n19854), .B2(n16544), .ZN(
        U376) );
  INV_X1 U19764 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16545) );
  NOR2_X1 U19765 ( .A1(n18716), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18719) );
  OAI22_X1 U19766 ( .A1(n18728), .A2(n18719), .B1(n18716), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18711) );
  INV_X1 U19767 ( .A(n18711), .ZN(n18800) );
  OAI21_X1 U19768 ( .B1(n18728), .B2(n16545), .A(n18713), .ZN(P3_U2633) );
  NOR2_X1 U19769 ( .A1(n17454), .A2(n16546), .ZN(n16552) );
  INV_X1 U19770 ( .A(n17453), .ZN(n16547) );
  OAI21_X1 U19771 ( .B1(n16552), .B2(n16547), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16548) );
  OAI21_X1 U19772 ( .B1(n16549), .B2(n18700), .A(n16548), .ZN(P3_U2634) );
  AOI21_X1 U19773 ( .B1(n18728), .B2(n18730), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16550) );
  AOI22_X1 U19774 ( .A1(n18788), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16550), 
        .B2(n18841), .ZN(P3_U2635) );
  INV_X1 U19775 ( .A(n16551), .ZN(n18714) );
  OAI21_X1 U19776 ( .B1(n18714), .B2(BS16), .A(n18800), .ZN(n18798) );
  OAI21_X1 U19777 ( .B1(n18800), .B2(n18849), .A(n18798), .ZN(P3_U2636) );
  NOR3_X1 U19778 ( .A1(n16554), .A2(n16553), .A3(n16552), .ZN(n18640) );
  NOR2_X1 U19779 ( .A1(n18640), .A2(n18697), .ZN(n18843) );
  OAI21_X1 U19780 ( .B1(n18843), .B2(n18180), .A(n16555), .ZN(P3_U2637) );
  INV_X1 U19781 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18839) );
  NOR4_X1 U19782 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n16559) );
  NOR4_X1 U19783 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n16558) );
  NOR4_X1 U19784 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16557) );
  NOR4_X1 U19785 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_23__SCAN_IN), .A3(P3_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16556) );
  NAND4_X1 U19786 ( .A1(n16559), .A2(n16558), .A3(n16557), .A4(n16556), .ZN(
        n16565) );
  NOR4_X1 U19787 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16563) );
  AOI211_X1 U19788 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_25__SCAN_IN), .B(
        P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(n16562) );
  NOR4_X1 U19789 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n16561) );
  NOR4_X1 U19790 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16560) );
  NAND4_X1 U19791 ( .A1(n16563), .A2(n16562), .A3(n16561), .A4(n16560), .ZN(
        n16564) );
  NOR2_X1 U19792 ( .A1(n16565), .A2(n16564), .ZN(n18834) );
  INV_X1 U19793 ( .A(n18834), .ZN(n18838) );
  INV_X1 U19794 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18799) );
  NOR2_X1 U19795 ( .A1(n18838), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18840) );
  AND3_X1 U19796 ( .A1(n16566), .A2(n18799), .A3(n18840), .ZN(n16568) );
  AOI21_X1 U19797 ( .B1(P3_BYTEENABLE_REG_1__SCAN_IN), .B2(n18838), .A(n16568), 
        .ZN(n16567) );
  OAI21_X1 U19798 ( .B1(n18839), .B2(n18838), .A(n16567), .ZN(P3_U2638) );
  NAND2_X1 U19799 ( .A1(n18834), .A2(n18839), .ZN(n18836) );
  AOI21_X1 U19800 ( .B1(P3_BYTEENABLE_REG_3__SCAN_IN), .B2(n18838), .A(n16568), 
        .ZN(n16569) );
  OAI21_X1 U19801 ( .B1(P3_DATAWIDTH_REG_1__SCAN_IN), .B2(n18836), .A(n16569), 
        .ZN(P3_U2639) );
  OAI21_X1 U19802 ( .B1(n16579), .B2(n16925), .A(n16570), .ZN(n16578) );
  AOI211_X1 U19803 ( .C1(n16573), .C2(n16572), .A(n16571), .B(n16808), .ZN(
        n16575) );
  OAI22_X1 U19804 ( .A1(n18794), .A2(n16584), .B1(n16925), .B2(n16910), .ZN(
        n16574) );
  AOI211_X1 U19805 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16575), .B(n16574), .ZN(n16577) );
  OAI211_X1 U19806 ( .C1(n16911), .C2(n16578), .A(n16577), .B(n16576), .ZN(
        P3_U2641) );
  AOI211_X1 U19807 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16589), .A(n16579), .B(
        n16911), .ZN(n16588) );
  AOI211_X1 U19808 ( .C1(n16582), .C2(n16581), .A(n16580), .B(n16808), .ZN(
        n16587) );
  AOI22_X1 U19809 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16898), .B1(
        P3_EBX_REG_29__SCAN_IN), .B2(n16871), .ZN(n16583) );
  OAI221_X1 U19810 ( .B1(P3_REIP_REG_29__SCAN_IN), .B2(n16585), .C1(n18787), 
        .C2(n16584), .A(n16583), .ZN(n16586) );
  OR3_X1 U19811 ( .A1(n16588), .A2(n16587), .A3(n16586), .ZN(P3_U2642) );
  OAI21_X1 U19812 ( .B1(n16602), .B2(n16593), .A(n16589), .ZN(n16598) );
  AOI211_X1 U19813 ( .C1(n17505), .C2(n16591), .A(n16590), .B(n16808), .ZN(
        n16595) );
  NAND2_X1 U19814 ( .A1(n16912), .A2(n16592), .ZN(n16610) );
  OAI22_X1 U19815 ( .A1(n18785), .A2(n16610), .B1(n16593), .B2(n16910), .ZN(
        n16594) );
  AOI211_X1 U19816 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16595), .B(n16594), .ZN(n16597) );
  INV_X1 U19817 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18782) );
  OAI221_X1 U19818 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(P3_REIP_REG_27__SCAN_IN), .C1(n18785), .C2(n18782), .A(n16605), .ZN(n16596) );
  OAI211_X1 U19819 ( .C1(n16598), .C2(n16911), .A(n16597), .B(n16596), .ZN(
        P3_U2643) );
  AOI22_X1 U19820 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16898), .B1(
        P3_EBX_REG_27__SCAN_IN), .B2(n16871), .ZN(n16607) );
  AOI211_X1 U19821 ( .C1(n16601), .C2(n16600), .A(n16599), .B(n16808), .ZN(
        n16604) );
  AOI211_X1 U19822 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16613), .A(n16602), .B(
        n16911), .ZN(n16603) );
  AOI211_X1 U19823 ( .C1(n16605), .C2(n18782), .A(n16604), .B(n16603), .ZN(
        n16606) );
  OAI211_X1 U19824 ( .C1(n18782), .C2(n16610), .A(n16607), .B(n16606), .ZN(
        P3_U2644) );
  AOI211_X1 U19825 ( .C1(n17540), .C2(n16609), .A(n16608), .B(n16808), .ZN(
        n16612) );
  OAI22_X1 U19826 ( .A1(n18780), .A2(n16610), .B1(n16956), .B2(n16910), .ZN(
        n16611) );
  AOI211_X1 U19827 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16612), .B(n16611), .ZN(n16615) );
  OAI211_X1 U19828 ( .C1(n16618), .C2(n16956), .A(n16906), .B(n16613), .ZN(
        n16614) );
  OAI211_X1 U19829 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16616), .A(n16615), 
        .B(n16614), .ZN(P3_U2645) );
  INV_X1 U19830 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16628) );
  INV_X1 U19831 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18778) );
  AOI22_X1 U19832 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16898), .B1(
        n16617), .B2(n18778), .ZN(n16627) );
  OAI21_X1 U19833 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16902), .A(n16638), 
        .ZN(n16625) );
  AOI211_X1 U19834 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16619), .A(n16618), .B(
        n16911), .ZN(n16624) );
  AOI211_X1 U19835 ( .C1(n16622), .C2(n16621), .A(n16620), .B(n18704), .ZN(
        n16623) );
  AOI211_X1 U19836 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16625), .A(n16624), 
        .B(n16623), .ZN(n16626) );
  OAI211_X1 U19837 ( .C1(n16628), .C2(n16910), .A(n16627), .B(n16626), .ZN(
        P3_U2646) );
  AOI211_X1 U19838 ( .C1(n17559), .C2(n16630), .A(n16629), .B(n16808), .ZN(
        n16633) );
  NOR3_X1 U19839 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16631), .A3(n16902), 
        .ZN(n16632) );
  AOI211_X1 U19840 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16633), .B(n16632), .ZN(n16637) );
  XNOR2_X1 U19841 ( .A(P3_EBX_REG_24__SCAN_IN), .B(n16634), .ZN(n16635) );
  AOI22_X1 U19842 ( .A1(n16906), .A2(n16635), .B1(P3_EBX_REG_24__SCAN_IN), 
        .B2(n16871), .ZN(n16636) );
  OAI211_X1 U19843 ( .C1(n16638), .C2(n18776), .A(n16637), .B(n16636), .ZN(
        P3_U2647) );
  AOI22_X1 U19844 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16898), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n16871), .ZN(n16649) );
  AOI21_X1 U19845 ( .B1(n16639), .B2(n16888), .A(n16894), .ZN(n16670) );
  INV_X1 U19846 ( .A(n16670), .ZN(n16657) );
  NOR3_X1 U19847 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16639), .A3(n16902), 
        .ZN(n16650) );
  AOI211_X1 U19848 ( .C1(n17591), .C2(n16641), .A(n16640), .B(n18704), .ZN(
        n16642) );
  AOI221_X1 U19849 ( .B1(n16657), .B2(P3_REIP_REG_22__SCAN_IN), .C1(n16650), 
        .C2(P3_REIP_REG_22__SCAN_IN), .A(n16642), .ZN(n16648) );
  OAI211_X1 U19850 ( .C1(n16651), .C2(n16644), .A(n16906), .B(n16643), .ZN(
        n16647) );
  INV_X1 U19851 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18772) );
  NAND3_X1 U19852 ( .A1(n16645), .A2(n16888), .A3(n18772), .ZN(n16646) );
  NAND4_X1 U19853 ( .A1(n16649), .A2(n16648), .A3(n16647), .A4(n16646), .ZN(
        P3_U2649) );
  AOI21_X1 U19854 ( .B1(n16871), .B2(P3_EBX_REG_21__SCAN_IN), .A(n16650), .ZN(
        n16659) );
  AOI211_X1 U19855 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16666), .A(n16651), .B(
        n16911), .ZN(n16656) );
  AOI211_X1 U19856 ( .C1(n16654), .C2(n16653), .A(n16652), .B(n18704), .ZN(
        n16655) );
  AOI211_X1 U19857 ( .C1(n16657), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16656), 
        .B(n16655), .ZN(n16658) );
  OAI211_X1 U19858 ( .C1(n17607), .C2(n16891), .A(n16659), .B(n16658), .ZN(
        P3_U2650) );
  AOI21_X1 U19859 ( .B1(n16660), .B2(n16888), .A(P3_REIP_REG_20__SCAN_IN), 
        .ZN(n16671) );
  AOI211_X1 U19860 ( .C1(n17620), .C2(n16662), .A(n16661), .B(n18704), .ZN(
        n16665) );
  INV_X1 U19861 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16663) );
  OAI22_X1 U19862 ( .A1(n16663), .A2(n16891), .B1(n16667), .B2(n16910), .ZN(
        n16664) );
  NOR2_X1 U19863 ( .A1(n16665), .A2(n16664), .ZN(n16669) );
  OAI211_X1 U19864 ( .C1(n16682), .C2(n16667), .A(n16906), .B(n16666), .ZN(
        n16668) );
  OAI211_X1 U19865 ( .C1(n16671), .C2(n16670), .A(n16669), .B(n16668), .ZN(
        P3_U2651) );
  INV_X1 U19866 ( .A(n16672), .ZN(n16675) );
  INV_X1 U19867 ( .A(n16673), .ZN(n16674) );
  NAND2_X1 U19868 ( .A1(n16914), .A2(n16674), .ZN(n16735) );
  OAI21_X1 U19869 ( .B1(n16675), .B2(n16735), .A(n16912), .ZN(n16701) );
  INV_X1 U19870 ( .A(n16701), .ZN(n16696) );
  NAND2_X1 U19871 ( .A1(n16674), .A2(n16888), .ZN(n16716) );
  NOR3_X1 U19872 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16675), .A3(n16716), 
        .ZN(n16695) );
  NOR2_X1 U19873 ( .A1(n16696), .A2(n16695), .ZN(n16687) );
  NOR3_X1 U19874 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16676), .A3(n16716), 
        .ZN(n16677) );
  AOI211_X1 U19875 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16871), .A(n9724), .B(
        n16677), .ZN(n16686) );
  NOR2_X1 U19876 ( .A1(n16698), .A2(n17646), .ZN(n16679) );
  INV_X1 U19877 ( .A(n16679), .ZN(n16688) );
  AOI21_X1 U19878 ( .B1(n16678), .B2(n16688), .A(n9740), .ZN(n17631) );
  AOI21_X1 U19879 ( .B1(n16679), .B2(n16883), .A(n16843), .ZN(n16681) );
  NOR2_X1 U19880 ( .A1(n17631), .A2(n16681), .ZN(n16680) );
  AOI211_X1 U19881 ( .C1(n17631), .C2(n16681), .A(n18704), .B(n16680), .ZN(
        n16684) );
  AOI211_X1 U19882 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16691), .A(n16682), .B(
        n16911), .ZN(n16683) );
  AOI211_X1 U19883 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16684), .B(n16683), .ZN(n16685) );
  OAI211_X1 U19884 ( .C1(n16687), .C2(n18766), .A(n16686), .B(n16685), .ZN(
        P3_U2652) );
  INV_X1 U19885 ( .A(n16698), .ZN(n17630) );
  OAI21_X1 U19886 ( .B1(n17630), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16688), .ZN(n17643) );
  OAI21_X1 U19887 ( .B1(n17638), .B2(n16757), .A(n16869), .ZN(n16690) );
  AOI21_X1 U19888 ( .B1(n17643), .B2(n16690), .A(n16808), .ZN(n16689) );
  OAI21_X1 U19889 ( .B1(n17643), .B2(n16690), .A(n16689), .ZN(n16693) );
  OAI211_X1 U19890 ( .C1(n16703), .C2(n17053), .A(n16906), .B(n16691), .ZN(
        n16692) );
  OAI211_X1 U19891 ( .C1(n16891), .C2(n17646), .A(n16693), .B(n16692), .ZN(
        n16694) );
  AOI211_X1 U19892 ( .C1(n16696), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16695), 
        .B(n16694), .ZN(n16697) );
  OAI211_X1 U19893 ( .C1(n17053), .C2(n16910), .A(n16697), .B(n13328), .ZN(
        P3_U2653) );
  OAI21_X1 U19894 ( .B1(n16699), .B2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16698), .ZN(n17660) );
  OAI21_X1 U19895 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16710), .A(
        n16869), .ZN(n16700) );
  XNOR2_X1 U19896 ( .A(n17660), .B(n16700), .ZN(n16708) );
  AOI21_X1 U19897 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16871), .A(n9724), .ZN(
        n16707) );
  AOI221_X1 U19898 ( .B1(n16702), .B2(n18763), .C1(n16716), .C2(n18763), .A(
        n16701), .ZN(n16705) );
  AOI211_X1 U19899 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16713), .A(n16703), .B(
        n16911), .ZN(n16704) );
  AOI211_X1 U19900 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16705), .B(n16704), .ZN(n16706) );
  OAI211_X1 U19901 ( .C1(n16808), .C2(n16708), .A(n16707), .B(n16706), .ZN(
        P3_U2654) );
  NOR2_X1 U19902 ( .A1(n16709), .A2(n16843), .ZN(n16712) );
  NOR2_X1 U19903 ( .A1(n17679), .A2(n17867), .ZN(n17669) );
  INV_X1 U19904 ( .A(n17669), .ZN(n16731) );
  NOR2_X1 U19905 ( .A1(n17685), .A2(n16731), .ZN(n16711) );
  OAI21_X1 U19906 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16711), .A(
        n16710), .ZN(n17674) );
  XOR2_X1 U19907 ( .A(n16712), .B(n17674), .Z(n16720) );
  AOI22_X1 U19908 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16898), .B1(
        P3_EBX_REG_16__SCAN_IN), .B2(n16871), .ZN(n16719) );
  NAND2_X1 U19909 ( .A1(n16912), .A2(n16735), .ZN(n16729) );
  INV_X1 U19910 ( .A(n16729), .ZN(n16740) );
  NOR2_X1 U19911 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16716), .ZN(n16721) );
  INV_X1 U19912 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18761) );
  NAND2_X1 U19913 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n18761), .ZN(n16715) );
  OAI211_X1 U19914 ( .C1(n16724), .C2(n17039), .A(n16906), .B(n16713), .ZN(
        n16714) );
  OAI211_X1 U19915 ( .C1(n16716), .C2(n16715), .A(n18162), .B(n16714), .ZN(
        n16717) );
  AOI221_X1 U19916 ( .B1(n16740), .B2(P3_REIP_REG_16__SCAN_IN), .C1(n16721), 
        .C2(P3_REIP_REG_16__SCAN_IN), .A(n16717), .ZN(n16718) );
  OAI211_X1 U19917 ( .C1(n16808), .C2(n16720), .A(n16719), .B(n16718), .ZN(
        P3_U2655) );
  INV_X1 U19918 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18758) );
  AOI211_X1 U19919 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16871), .A(n9724), .B(
        n16721), .ZN(n16728) );
  AOI22_X1 U19920 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16731), .B1(
        n17669), .B2(n17685), .ZN(n17681) );
  OAI21_X1 U19921 ( .B1(n17679), .B2(n16757), .A(n16869), .ZN(n16723) );
  NOR2_X1 U19922 ( .A1(n17681), .A2(n16723), .ZN(n16722) );
  AOI211_X1 U19923 ( .C1(n17681), .C2(n16723), .A(n18704), .B(n16722), .ZN(
        n16726) );
  AOI211_X1 U19924 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16741), .A(n16724), .B(
        n16911), .ZN(n16725) );
  AOI211_X1 U19925 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16726), .B(n16725), .ZN(n16727) );
  OAI211_X1 U19926 ( .C1(n18758), .C2(n16729), .A(n16728), .B(n16727), .ZN(
        P3_U2656) );
  INV_X1 U19927 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16744) );
  INV_X1 U19928 ( .A(n17708), .ZN(n16730) );
  NAND2_X1 U19929 ( .A1(n17709), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17711) );
  NOR2_X1 U19930 ( .A1(n16730), .A2(n17711), .ZN(n16732) );
  INV_X1 U19931 ( .A(n16732), .ZN(n16745) );
  OAI21_X1 U19932 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16745), .A(
        n16869), .ZN(n16734) );
  OAI21_X1 U19933 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16732), .A(
        n16731), .ZN(n17698) );
  NOR2_X1 U19934 ( .A1(n16734), .A2(n17698), .ZN(n16733) );
  AOI211_X1 U19935 ( .C1(n16734), .C2(n17698), .A(n18704), .B(n16733), .ZN(
        n16739) );
  NAND3_X1 U19936 ( .A1(n16888), .A2(n16736), .A3(n16735), .ZN(n16737) );
  OAI211_X1 U19937 ( .C1(n17111), .C2(n16910), .A(n18162), .B(n16737), .ZN(
        n16738) );
  AOI211_X1 U19938 ( .C1(n16740), .C2(P3_REIP_REG_14__SCAN_IN), .A(n16739), 
        .B(n16738), .ZN(n16743) );
  OAI211_X1 U19939 ( .C1(n16749), .C2(n17111), .A(n16906), .B(n16741), .ZN(
        n16742) );
  OAI211_X1 U19940 ( .C1(n16891), .C2(n16744), .A(n16743), .B(n16742), .ZN(
        P3_U2657) );
  NOR2_X1 U19941 ( .A1(n17724), .A2(n17711), .ZN(n16756) );
  OAI21_X1 U19942 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16756), .A(
        n16745), .ZN(n16746) );
  INV_X1 U19943 ( .A(n16746), .ZN(n17716) );
  AOI21_X1 U19944 ( .B1(n16756), .B2(n16883), .A(n16843), .ZN(n16747) );
  XNOR2_X1 U19945 ( .A(n17716), .B(n16747), .ZN(n16755) );
  NOR3_X1 U19946 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16748), .A3(n16902), 
        .ZN(n16752) );
  AOI211_X1 U19947 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16764), .A(n16749), .B(
        n16911), .ZN(n16751) );
  OAI22_X1 U19948 ( .A1(n17713), .A2(n16891), .B1(n17107), .B2(n16910), .ZN(
        n16750) );
  NOR4_X1 U19949 ( .A1(n9724), .A2(n16752), .A3(n16751), .A4(n16750), .ZN(
        n16754) );
  NOR2_X1 U19950 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16902), .ZN(n16759) );
  OAI21_X1 U19951 ( .B1(n16760), .B2(n16902), .A(n16914), .ZN(n16769) );
  OAI21_X1 U19952 ( .B1(n16759), .B2(n16769), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16753) );
  OAI211_X1 U19953 ( .C1(n16755), .C2(n16808), .A(n16754), .B(n16753), .ZN(
        P3_U2658) );
  AOI21_X1 U19954 ( .B1(n17724), .B2(n17711), .A(n16756), .ZN(n17728) );
  INV_X1 U19955 ( .A(n16757), .ZN(n16886) );
  AOI21_X1 U19956 ( .B1(n17709), .B2(n16886), .A(n16843), .ZN(n16758) );
  XNOR2_X1 U19957 ( .A(n17728), .B(n16758), .ZN(n16762) );
  AOI22_X1 U19958 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16871), .B1(n16760), 
        .B2(n16759), .ZN(n16761) );
  OAI211_X1 U19959 ( .C1(n18704), .C2(n16762), .A(n16761), .B(n18162), .ZN(
        n16763) );
  AOI21_X1 U19960 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16769), .A(n16763), 
        .ZN(n16767) );
  OAI211_X1 U19961 ( .C1(n16768), .C2(n16765), .A(n16906), .B(n16764), .ZN(
        n16766) );
  OAI211_X1 U19962 ( .C1(n16891), .C2(n17724), .A(n16767), .B(n16766), .ZN(
        P3_U2659) );
  AOI211_X1 U19963 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n16787), .A(n16768), .B(
        n16911), .ZN(n16776) );
  INV_X1 U19964 ( .A(n16769), .ZN(n16774) );
  INV_X1 U19965 ( .A(n16786), .ZN(n16770) );
  NOR2_X1 U19966 ( .A1(n16778), .A2(n16902), .ZN(n16795) );
  AOI21_X1 U19967 ( .B1(n16770), .B2(n16795), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16773) );
  NAND2_X1 U19968 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17741) );
  NAND2_X1 U19969 ( .A1(n9814), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16829) );
  NOR2_X1 U19970 ( .A1(n17794), .A2(n16829), .ZN(n16817) );
  NAND2_X1 U19971 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16817), .ZN(
        n16805) );
  NOR2_X1 U19972 ( .A1(n17741), .A2(n16805), .ZN(n16779) );
  AOI21_X1 U19973 ( .B1(n16779), .B2(n16883), .A(n16843), .ZN(n16771) );
  OAI21_X1 U19974 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16779), .A(
        n17711), .ZN(n17742) );
  XOR2_X1 U19975 ( .A(n16771), .B(n17742), .Z(n16772) );
  OAI22_X1 U19976 ( .A1(n16774), .A2(n16773), .B1(n16808), .B2(n16772), .ZN(
        n16775) );
  AOI211_X1 U19977 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16776), .B(n16775), .ZN(n16777) );
  OAI211_X1 U19978 ( .C1(n17138), .C2(n16910), .A(n16777), .B(n13328), .ZN(
        P3_U2660) );
  AOI21_X1 U19979 ( .B1(n16778), .B2(n16888), .A(n16894), .ZN(n16809) );
  INV_X1 U19980 ( .A(n16809), .ZN(n16785) );
  INV_X1 U19981 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16782) );
  INV_X1 U19982 ( .A(n16805), .ZN(n16793) );
  NAND2_X1 U19983 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16793), .ZN(
        n16792) );
  AOI21_X1 U19984 ( .B1(n16782), .B2(n16792), .A(n16779), .ZN(n17761) );
  INV_X1 U19985 ( .A(n16792), .ZN(n16780) );
  AOI21_X1 U19986 ( .B1(n16780), .B2(n16883), .A(n16843), .ZN(n16799) );
  NOR2_X1 U19987 ( .A1(n17761), .A2(n16799), .ZN(n16781) );
  AOI211_X1 U19988 ( .C1(n17761), .C2(n16799), .A(n18704), .B(n16781), .ZN(
        n16784) );
  OAI22_X1 U19989 ( .A1(n16782), .A2(n16891), .B1(n17155), .B2(n16910), .ZN(
        n16783) );
  AOI211_X1 U19990 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n16785), .A(n16784), 
        .B(n16783), .ZN(n16790) );
  OAI211_X1 U19991 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(P3_REIP_REG_10__SCAN_IN), 
        .A(n16795), .B(n16786), .ZN(n16789) );
  OAI211_X1 U19992 ( .C1(n16794), .C2(n17155), .A(n16906), .B(n16787), .ZN(
        n16788) );
  NAND4_X1 U19993 ( .A1(n16790), .A2(n13328), .A3(n16789), .A4(n16788), .ZN(
        P3_U2661) );
  NAND2_X1 U19994 ( .A1(n16830), .A2(n16791), .ZN(n16882) );
  OAI21_X1 U19995 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16793), .A(
        n16792), .ZN(n17770) );
  AOI211_X1 U19996 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16812), .A(n16794), .B(
        n16911), .ZN(n16798) );
  INV_X1 U19997 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18747) );
  AOI22_X1 U19998 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16898), .B1(
        n16795), .B2(n18747), .ZN(n16796) );
  OAI211_X1 U19999 ( .C1(n18747), .C2(n16809), .A(n16796), .B(n18162), .ZN(
        n16797) );
  AOI211_X1 U20000 ( .C1(n16871), .C2(P3_EBX_REG_9__SCAN_IN), .A(n16798), .B(
        n16797), .ZN(n16802) );
  NOR2_X1 U20001 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16805), .ZN(
        n16800) );
  OAI211_X1 U20002 ( .C1(n16800), .C2(n17770), .A(n16830), .B(n16799), .ZN(
        n16801) );
  OAI211_X1 U20003 ( .C1(n16882), .C2(n17770), .A(n16802), .B(n16801), .ZN(
        P3_U2662) );
  AOI21_X1 U20004 ( .B1(n16803), .B2(n16888), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n16810) );
  NOR2_X1 U20005 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16829), .ZN(
        n16804) );
  AOI21_X1 U20006 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16804), .A(
        n16843), .ZN(n16806) );
  OAI21_X1 U20007 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16817), .A(
        n16805), .ZN(n17782) );
  XOR2_X1 U20008 ( .A(n16806), .B(n17782), .Z(n16807) );
  OAI22_X1 U20009 ( .A1(n16810), .A2(n16809), .B1(n16808), .B2(n16807), .ZN(
        n16811) );
  AOI211_X1 U20010 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16871), .A(n9724), .B(
        n16811), .ZN(n16815) );
  OAI211_X1 U20011 ( .C1(n16818), .C2(n16813), .A(n16906), .B(n16812), .ZN(
        n16814) );
  OAI211_X1 U20012 ( .C1(n16891), .C2(n16816), .A(n16815), .B(n16814), .ZN(
        P3_U2663) );
  AOI21_X1 U20013 ( .B1(n17794), .B2(n16829), .A(n16817), .ZN(n17800) );
  OAI21_X1 U20014 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16829), .A(
        n16869), .ZN(n16832) );
  XOR2_X1 U20015 ( .A(n17800), .B(n16832), .Z(n16827) );
  AOI211_X1 U20016 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16833), .A(n16818), .B(
        n16911), .ZN(n16819) );
  AOI211_X1 U20017 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16871), .A(n9724), .B(
        n16819), .ZN(n16826) );
  INV_X1 U20018 ( .A(n16821), .ZN(n16820) );
  AOI21_X1 U20019 ( .B1(n16888), .B2(n16820), .A(n16894), .ZN(n16845) );
  INV_X1 U20020 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18741) );
  NAND3_X1 U20021 ( .A1(n16821), .A2(n16888), .A3(n18741), .ZN(n16835) );
  AOI21_X1 U20022 ( .B1(n16845), .B2(n16835), .A(n18743), .ZN(n16824) );
  NOR3_X1 U20023 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16822), .A3(n16902), .ZN(
        n16823) );
  AOI211_X1 U20024 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16824), .B(n16823), .ZN(n16825) );
  OAI211_X1 U20025 ( .C1(n18704), .C2(n16827), .A(n16826), .B(n16825), .ZN(
        P3_U2664) );
  NOR2_X1 U20026 ( .A1(n16828), .A2(n17867), .ZN(n16841) );
  OAI21_X1 U20027 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16841), .A(
        n16829), .ZN(n17810) );
  OAI21_X1 U20028 ( .B1(n16843), .B2(n16883), .A(n16830), .ZN(n16909) );
  AOI211_X1 U20029 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16869), .A(
        n17810), .B(n16909), .ZN(n16839) );
  NAND2_X1 U20030 ( .A1(n16830), .A2(n17810), .ZN(n16831) );
  OAI22_X1 U20031 ( .A1(n9874), .A2(n16891), .B1(n16832), .B2(n16831), .ZN(
        n16838) );
  OAI211_X1 U20032 ( .C1(n16847), .C2(n16836), .A(n16906), .B(n16833), .ZN(
        n16834) );
  OAI211_X1 U20033 ( .C1(n16910), .C2(n16836), .A(n16835), .B(n16834), .ZN(
        n16837) );
  NOR4_X1 U20034 ( .A1(n9724), .A2(n16839), .A3(n16838), .A4(n16837), .ZN(
        n16840) );
  OAI21_X1 U20035 ( .B1(n18741), .B2(n16845), .A(n16840), .ZN(P3_U2665) );
  INV_X1 U20036 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16842) );
  NAND2_X1 U20037 ( .A1(n17814), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16853) );
  AOI21_X1 U20038 ( .B1(n16842), .B2(n16853), .A(n16841), .ZN(n17823) );
  INV_X1 U20039 ( .A(n16853), .ZN(n16844) );
  AOI21_X1 U20040 ( .B1(n16844), .B2(n16883), .A(n16843), .ZN(n16859) );
  XNOR2_X1 U20041 ( .A(n17823), .B(n16859), .ZN(n16852) );
  AOI21_X1 U20042 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n16871), .A(n9724), .ZN(
        n16851) );
  AOI221_X1 U20043 ( .B1(n16846), .B2(n18739), .C1(n16902), .C2(n18739), .A(
        n16845), .ZN(n16849) );
  AOI211_X1 U20044 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n16854), .A(n16847), .B(
        n16911), .ZN(n16848) );
  AOI211_X1 U20045 ( .C1(n16898), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16849), .B(n16848), .ZN(n16850) );
  OAI211_X1 U20046 ( .C1(n18704), .C2(n16852), .A(n16851), .B(n16850), .ZN(
        P3_U2666) );
  NOR2_X1 U20047 ( .A1(n16858), .A2(n17867), .ZN(n16867) );
  OAI21_X1 U20048 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16867), .A(
        n16853), .ZN(n17837) );
  NOR2_X1 U20049 ( .A1(n17387), .A2(n18859), .ZN(n16880) );
  AOI221_X1 U20050 ( .B1(n17163), .B2(n16880), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n16880), .A(n9724), .ZN(
        n16866) );
  OAI211_X1 U20051 ( .C1(n16873), .C2(n16857), .A(n16906), .B(n16854), .ZN(
        n16856) );
  INV_X1 U20052 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18737) );
  NAND3_X1 U20053 ( .A1(n16860), .A2(n16888), .A3(n18737), .ZN(n16855) );
  OAI211_X1 U20054 ( .C1(n16910), .C2(n16857), .A(n16856), .B(n16855), .ZN(
        n16864) );
  NOR2_X1 U20055 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16858), .ZN(
        n17832) );
  AOI22_X1 U20056 ( .A1(n16886), .A2(n17832), .B1(n16859), .B2(n17837), .ZN(
        n16862) );
  INV_X1 U20057 ( .A(n16860), .ZN(n16861) );
  AOI21_X1 U20058 ( .B1(n16888), .B2(n16861), .A(n16894), .ZN(n16874) );
  OAI22_X1 U20059 ( .A1(n16862), .A2(n18704), .B1(n18737), .B2(n16874), .ZN(
        n16863) );
  AOI211_X1 U20060 ( .C1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n16898), .A(
        n16864), .B(n16863), .ZN(n16865) );
  OAI211_X1 U20061 ( .C1(n17837), .C2(n16882), .A(n16866), .B(n16865), .ZN(
        P3_U2667) );
  INV_X1 U20062 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17859) );
  NOR2_X1 U20063 ( .A1(n17859), .A2(n17867), .ZN(n16884) );
  INV_X1 U20064 ( .A(n16867), .ZN(n16868) );
  OAI21_X1 U20065 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16884), .A(
        n16868), .ZN(n17849) );
  INV_X1 U20066 ( .A(n16884), .ZN(n16881) );
  OAI21_X1 U20067 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16881), .A(
        n16869), .ZN(n16870) );
  XNOR2_X1 U20068 ( .A(n17849), .B(n16870), .ZN(n16879) );
  AOI22_X1 U20069 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16898), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(n16871), .ZN(n16878) );
  NOR2_X1 U20070 ( .A1(n18817), .A2(n18825), .ZN(n18652) );
  NAND2_X1 U20071 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18652), .ZN(
        n18650) );
  AOI21_X1 U20072 ( .B1(n18650), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n17191), .ZN(n16872) );
  INV_X1 U20073 ( .A(n16872), .ZN(n18804) );
  AOI211_X1 U20074 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16895), .A(n16873), .B(
        n16911), .ZN(n16876) );
  AOI221_X1 U20075 ( .B1(n16887), .B2(n18735), .C1(n16902), .C2(n18735), .A(
        n16874), .ZN(n16875) );
  AOI211_X1 U20076 ( .C1(n16880), .C2(n18804), .A(n16876), .B(n16875), .ZN(
        n16877) );
  OAI211_X1 U20077 ( .C1(n18704), .C2(n16879), .A(n16878), .B(n16877), .ZN(
        P3_U2668) );
  NAND2_X1 U20078 ( .A1(n18817), .A2(n18657), .ZN(n18654) );
  NAND2_X1 U20079 ( .A1(n18654), .A2(n18650), .ZN(n18811) );
  INV_X1 U20080 ( .A(n16880), .ZN(n16917) );
  OAI21_X1 U20081 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16881), .ZN(n17856) );
  OAI22_X1 U20082 ( .A1(n18811), .A2(n16917), .B1(n17856), .B2(n16882), .ZN(
        n16893) );
  NAND2_X1 U20083 ( .A1(n16884), .A2(n16883), .ZN(n16885) );
  OAI211_X1 U20084 ( .C1(n16886), .C2(n17856), .A(n16899), .B(n16885), .ZN(
        n16890) );
  OAI211_X1 U20085 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16888), .B(n16887), .ZN(n16889) );
  OAI211_X1 U20086 ( .C1(n16891), .C2(n17859), .A(n16890), .B(n16889), .ZN(
        n16892) );
  AOI211_X1 U20087 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n16894), .A(n16893), .B(
        n16892), .ZN(n16897) );
  OAI211_X1 U20088 ( .C1(n16900), .C2(n17213), .A(n16906), .B(n16895), .ZN(
        n16896) );
  OAI211_X1 U20089 ( .C1(n16910), .C2(n17213), .A(n16897), .B(n16896), .ZN(
        P3_U2669) );
  AOI21_X1 U20090 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16899), .A(
        n16898), .ZN(n16908) );
  AOI21_X1 U20091 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n16900), .ZN(n17222) );
  INV_X1 U20092 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n16901) );
  OAI22_X1 U20093 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16902), .B1(n16901), 
        .B2(n16910), .ZN(n16905) );
  NAND2_X1 U20094 ( .A1(n16903), .A2(n18657), .ZN(n18818) );
  OAI22_X1 U20095 ( .A1(n18839), .A2(n16914), .B1(n18818), .B2(n16917), .ZN(
        n16904) );
  AOI211_X1 U20096 ( .C1(n16906), .C2(n17222), .A(n16905), .B(n16904), .ZN(
        n16907) );
  OAI221_X1 U20097 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16909), .C1(
        n17867), .C2(n16908), .A(n16907), .ZN(P3_U2670) );
  NAND2_X1 U20098 ( .A1(n16911), .A2(n16910), .ZN(n16913) );
  AOI22_X1 U20099 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16913), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16912), .ZN(n16916) );
  NAND3_X1 U20100 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18813), .A3(
        n16914), .ZN(n16915) );
  OAI211_X1 U20101 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n16917), .A(
        n16916), .B(n16915), .ZN(P3_U2671) );
  NOR2_X1 U20102 ( .A1(n16956), .A2(n16955), .ZN(n16921) );
  NAND2_X1 U20103 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .ZN(n16918) );
  NOR4_X1 U20104 ( .A1(n16919), .A2(n16975), .A3(n16998), .A4(n16918), .ZN(
        n16920) );
  NAND4_X1 U20105 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16921), .A4(n16920), .ZN(n16924) );
  NAND2_X1 U20106 ( .A1(n17225), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16923) );
  NAND2_X1 U20107 ( .A1(n16950), .A2(n18226), .ZN(n16922) );
  OAI22_X1 U20108 ( .A1(n16950), .A2(n16923), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16922), .ZN(P3_U2672) );
  NAND2_X1 U20109 ( .A1(n16925), .A2(n16924), .ZN(n16926) );
  NAND2_X1 U20110 ( .A1(n16926), .A2(n17225), .ZN(n16949) );
  AOI22_X1 U20111 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16930) );
  AOI22_X1 U20112 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U20113 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16928) );
  AOI22_X1 U20114 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16927) );
  NAND4_X1 U20115 ( .A1(n16930), .A2(n16929), .A3(n16928), .A4(n16927), .ZN(
        n16936) );
  AOI22_X1 U20116 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U20117 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U20118 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20119 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13290), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16931) );
  NAND4_X1 U20120 ( .A1(n16934), .A2(n16933), .A3(n16932), .A4(n16931), .ZN(
        n16935) );
  NOR2_X1 U20121 ( .A1(n16936), .A2(n16935), .ZN(n16948) );
  AOI22_X1 U20122 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20123 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20124 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16938) );
  AOI22_X1 U20125 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16937) );
  NAND4_X1 U20126 ( .A1(n16940), .A2(n16939), .A3(n16938), .A4(n16937), .ZN(
        n16946) );
  AOI22_X1 U20127 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16944) );
  AOI22_X1 U20128 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13290), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20129 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20130 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16941) );
  NAND4_X1 U20131 ( .A1(n16944), .A2(n16943), .A3(n16942), .A4(n16941), .ZN(
        n16945) );
  NOR2_X1 U20132 ( .A1(n16946), .A2(n16945), .ZN(n16953) );
  INV_X1 U20133 ( .A(n16961), .ZN(n16952) );
  NOR3_X1 U20134 ( .A1(n16953), .A2(n16952), .A3(n16951), .ZN(n16947) );
  XOR2_X1 U20135 ( .A(n16948), .B(n16947), .Z(n17242) );
  OAI22_X1 U20136 ( .A1(n16950), .A2(n16949), .B1(n17242), .B2(n17225), .ZN(
        P3_U2673) );
  INV_X1 U20137 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16959) );
  NOR2_X1 U20138 ( .A1(n16952), .A2(n16951), .ZN(n16954) );
  XNOR2_X1 U20139 ( .A(n16954), .B(n16953), .ZN(n17246) );
  NOR4_X1 U20140 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16956), .A3(n16966), .A4(
        n16955), .ZN(n16957) );
  AOI21_X1 U20141 ( .B1(n17228), .B2(n17246), .A(n16957), .ZN(n16958) );
  OAI21_X1 U20142 ( .B1(n16960), .B2(n16959), .A(n16958), .ZN(P3_U2674) );
  INV_X1 U20143 ( .A(n16971), .ZN(n16965) );
  AOI21_X1 U20144 ( .B1(n16962), .B2(n16967), .A(n16961), .ZN(n17254) );
  AOI22_X1 U20145 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16963), .B1(n17228), 
        .B2(n17254), .ZN(n16964) );
  OAI21_X1 U20146 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16965), .A(n16964), .ZN(
        P3_U2676) );
  INV_X1 U20147 ( .A(n16966), .ZN(n16974) );
  AOI21_X1 U20148 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17225), .A(n16974), .ZN(
        n16970) );
  OAI21_X1 U20149 ( .B1(n16969), .B2(n16968), .A(n16967), .ZN(n17262) );
  OAI22_X1 U20150 ( .A1(n16971), .A2(n16970), .B1(n17225), .B2(n17262), .ZN(
        P3_U2677) );
  AOI21_X1 U20151 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17225), .A(n16980), .ZN(
        n16973) );
  XNOR2_X1 U20152 ( .A(n16972), .B(n16976), .ZN(n17267) );
  OAI22_X1 U20153 ( .A1(n16974), .A2(n16973), .B1(n17225), .B2(n17267), .ZN(
        P3_U2678) );
  NOR2_X1 U20154 ( .A1(n16975), .A2(n16981), .ZN(n16985) );
  AOI21_X1 U20155 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17225), .A(n16985), .ZN(
        n16979) );
  OAI21_X1 U20156 ( .B1(n16978), .B2(n16977), .A(n16976), .ZN(n17272) );
  OAI22_X1 U20157 ( .A1(n16980), .A2(n16979), .B1(n17225), .B2(n17272), .ZN(
        P3_U2679) );
  INV_X1 U20158 ( .A(n16981), .ZN(n16997) );
  AOI21_X1 U20159 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17225), .A(n16997), .ZN(
        n16984) );
  XNOR2_X1 U20160 ( .A(n16983), .B(n16982), .ZN(n17277) );
  OAI22_X1 U20161 ( .A1(n16985), .A2(n16984), .B1(n17225), .B2(n17277), .ZN(
        P3_U2680) );
  AOI22_X1 U20162 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17225), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n9780), .ZN(n16996) );
  AOI22_X1 U20163 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20164 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20165 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20166 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16986) );
  NAND4_X1 U20167 ( .A1(n16989), .A2(n16988), .A3(n16987), .A4(n16986), .ZN(
        n16995) );
  AOI22_X1 U20168 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20169 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16992) );
  AOI22_X1 U20170 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13290), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16991) );
  AOI22_X1 U20171 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16990) );
  NAND4_X1 U20172 ( .A1(n16993), .A2(n16992), .A3(n16991), .A4(n16990), .ZN(
        n16994) );
  NOR2_X1 U20173 ( .A1(n16995), .A2(n16994), .ZN(n17280) );
  OAI22_X1 U20174 ( .A1(n16997), .A2(n16996), .B1(n17280), .B2(n17225), .ZN(
        P3_U2681) );
  NAND2_X1 U20175 ( .A1(n17225), .A2(n16998), .ZN(n17023) );
  AOI22_X1 U20176 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20177 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20178 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16999) );
  OAI21_X1 U20179 ( .B1(n13277), .B2(n17000), .A(n16999), .ZN(n17006) );
  AOI22_X1 U20180 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20181 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20182 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20183 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13290), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17001) );
  NAND4_X1 U20184 ( .A1(n17004), .A2(n17003), .A3(n17002), .A4(n17001), .ZN(
        n17005) );
  AOI211_X1 U20185 ( .C1(n9729), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n17006), .B(n17005), .ZN(n17008) );
  NAND3_X1 U20186 ( .A1(n17010), .A2(n17009), .A3(n17008), .ZN(n17284) );
  AOI22_X1 U20187 ( .A1(n17228), .A2(n17284), .B1(n9780), .B2(n9925), .ZN(
        n17011) );
  OAI21_X1 U20188 ( .B1(n9925), .B2(n17023), .A(n17011), .ZN(P3_U2682) );
  AOI22_X1 U20189 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20190 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20191 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20192 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17012) );
  NAND4_X1 U20193 ( .A1(n17015), .A2(n17014), .A3(n17013), .A4(n17012), .ZN(
        n17021) );
  AOI22_X1 U20194 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9730), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20195 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20196 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U20197 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13290), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17016) );
  NAND4_X1 U20198 ( .A1(n17019), .A2(n17018), .A3(n17017), .A4(n17016), .ZN(
        n17020) );
  NOR2_X1 U20199 ( .A1(n17021), .A2(n17020), .ZN(n17292) );
  NOR2_X1 U20200 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17022), .ZN(n17024) );
  OAI22_X1 U20201 ( .A1(n17292), .A2(n17225), .B1(n17024), .B2(n17023), .ZN(
        P3_U2683) );
  NAND2_X1 U20202 ( .A1(n17225), .A2(n17035), .ZN(n17052) );
  AOI22_X1 U20203 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20204 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20205 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17025) );
  OAI21_X1 U20206 ( .B1(n9756), .B2(n17127), .A(n17025), .ZN(n17031) );
  AOI22_X1 U20207 ( .A1(n15523), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20208 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20209 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20210 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17026) );
  NAND4_X1 U20211 ( .A1(n17029), .A2(n17028), .A3(n17027), .A4(n17026), .ZN(
        n17030) );
  AOI211_X1 U20212 ( .C1(n17175), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17031), .B(n17030), .ZN(n17032) );
  NAND3_X1 U20213 ( .A1(n17034), .A2(n17033), .A3(n17032), .ZN(n17293) );
  NOR3_X1 U20214 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17321), .A3(n17035), .ZN(
        n17036) );
  AOI21_X1 U20215 ( .B1(n17228), .B2(n17293), .A(n17036), .ZN(n17037) );
  OAI21_X1 U20216 ( .B1(n17038), .B2(n17052), .A(n17037), .ZN(P3_U2684) );
  NOR3_X1 U20217 ( .A1(n17321), .A2(n17039), .A3(n17092), .ZN(n17065) );
  NAND2_X1 U20218 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17065), .ZN(n17064) );
  AOI22_X1 U20219 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13290), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17050) );
  AOI22_X1 U20220 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20221 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17040) );
  OAI21_X1 U20222 ( .B1(n17180), .B2(n17220), .A(n17040), .ZN(n17047) );
  AOI22_X1 U20223 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20224 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20225 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20226 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17042) );
  NAND4_X1 U20227 ( .A1(n17045), .A2(n17044), .A3(n17043), .A4(n17042), .ZN(
        n17046) );
  AOI211_X1 U20228 ( .C1(n17173), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n17047), .B(n17046), .ZN(n17048) );
  NAND3_X1 U20229 ( .A1(n17050), .A2(n17049), .A3(n17048), .ZN(n17298) );
  NAND2_X1 U20230 ( .A1(n17228), .A2(n17298), .ZN(n17051) );
  OAI221_X1 U20231 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17064), .C1(n17053), 
        .C2(n17052), .A(n17051), .ZN(P3_U2685) );
  AOI22_X1 U20232 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20233 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17163), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20234 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9730), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20235 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17080), .ZN(n17054) );
  NAND4_X1 U20236 ( .A1(n17057), .A2(n17056), .A3(n17055), .A4(n17054), .ZN(
        n17063) );
  AOI22_X1 U20237 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17177), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20238 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17182), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U20239 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17191), .ZN(n17059) );
  AOI22_X1 U20240 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17162), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17058) );
  NAND4_X1 U20241 ( .A1(n17061), .A2(n17060), .A3(n17059), .A4(n17058), .ZN(
        n17062) );
  NOR2_X1 U20242 ( .A1(n17063), .A2(n17062), .ZN(n17309) );
  OAI211_X1 U20243 ( .C1(n17065), .C2(P3_EBX_REG_17__SCAN_IN), .A(n17225), .B(
        n17064), .ZN(n17066) );
  OAI21_X1 U20244 ( .B1(n17309), .B2(n17225), .A(n17066), .ZN(P3_U2686) );
  INV_X1 U20245 ( .A(n17092), .ZN(n17067) );
  OAI21_X1 U20246 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17067), .A(n17225), .ZN(
        n17078) );
  AOI22_X1 U20247 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20248 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20249 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20250 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17068) );
  NAND4_X1 U20251 ( .A1(n17071), .A2(n17070), .A3(n17069), .A4(n17068), .ZN(
        n17077) );
  AOI22_X1 U20252 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U20253 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13290), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20254 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9730), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20255 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17072) );
  NAND4_X1 U20256 ( .A1(n17075), .A2(n17074), .A3(n17073), .A4(n17072), .ZN(
        n17076) );
  NOR2_X1 U20257 ( .A1(n17077), .A2(n17076), .ZN(n17315) );
  OAI22_X1 U20258 ( .A1(n17079), .A2(n17078), .B1(n17315), .B2(n17225), .ZN(
        P3_U2687) );
  AOI22_X1 U20259 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20260 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20261 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13290), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20262 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17081) );
  NAND4_X1 U20263 ( .A1(n17084), .A2(n17083), .A3(n17082), .A4(n17081), .ZN(
        n17091) );
  AOI22_X1 U20264 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17089) );
  AOI22_X1 U20265 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20266 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U20267 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17085), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17086) );
  NAND4_X1 U20268 ( .A1(n17089), .A2(n17088), .A3(n17087), .A4(n17086), .ZN(
        n17090) );
  NOR2_X1 U20269 ( .A1(n17091), .A2(n17090), .ZN(n17320) );
  OAI21_X1 U20270 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17093), .A(n17092), .ZN(
        n17094) );
  AOI22_X1 U20271 ( .A1(n17228), .A2(n17320), .B1(n17094), .B2(n17225), .ZN(
        P3_U2688) );
  AOI22_X1 U20272 ( .A1(n17223), .A2(n17107), .B1(n17225), .B2(n17095), .ZN(
        n17110) );
  AOI22_X1 U20273 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20274 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U20275 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17096) );
  OAI21_X1 U20276 ( .B1(n13277), .B2(n17097), .A(n17096), .ZN(n17103) );
  AOI22_X1 U20277 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20278 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20279 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20280 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17098) );
  NAND4_X1 U20281 ( .A1(n17101), .A2(n17100), .A3(n17099), .A4(n17098), .ZN(
        n17102) );
  AOI211_X1 U20282 ( .C1(n17184), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17103), .B(n17102), .ZN(n17104) );
  NAND3_X1 U20283 ( .A1(n17106), .A2(n17105), .A3(n17104), .ZN(n17323) );
  NOR3_X1 U20284 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17107), .A3(n17123), .ZN(
        n17108) );
  AOI21_X1 U20285 ( .B1(n17228), .B2(n17323), .A(n17108), .ZN(n17109) );
  OAI21_X1 U20286 ( .B1(n17111), .B2(n17110), .A(n17109), .ZN(P3_U2689) );
  AOI22_X1 U20287 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20288 ( .A1(n10107), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20289 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20290 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9725), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17112) );
  NAND4_X1 U20291 ( .A1(n17115), .A2(n17114), .A3(n17113), .A4(n17112), .ZN(
        n17122) );
  AOI22_X1 U20292 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U20293 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20294 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20295 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13290), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17117) );
  NAND4_X1 U20296 ( .A1(n17120), .A2(n17119), .A3(n17118), .A4(n17117), .ZN(
        n17121) );
  NOR2_X1 U20297 ( .A1(n17122), .A2(n17121), .ZN(n17332) );
  OAI21_X1 U20298 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17142), .A(n17123), .ZN(
        n17124) );
  AOI22_X1 U20299 ( .A1(n17228), .A2(n17332), .B1(n17124), .B2(n17225), .ZN(
        P3_U2691) );
  AOI22_X1 U20300 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20301 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17116), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20302 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17126) );
  OAI21_X1 U20303 ( .B1(n17128), .B2(n17127), .A(n17126), .ZN(n17134) );
  AOI22_X1 U20304 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20305 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20306 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20307 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17129) );
  NAND4_X1 U20308 ( .A1(n17132), .A2(n17131), .A3(n17130), .A4(n17129), .ZN(
        n17133) );
  AOI211_X1 U20309 ( .C1(n9725), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n17134), .B(n17133), .ZN(n17135) );
  NAND3_X1 U20310 ( .A1(n17137), .A2(n17136), .A3(n17135), .ZN(n17335) );
  NAND3_X1 U20311 ( .A1(n17225), .A2(n17139), .A3(n17138), .ZN(n17140) );
  OAI21_X1 U20312 ( .B1(n17225), .B2(n17335), .A(n17140), .ZN(n17141) );
  AOI21_X1 U20313 ( .B1(n18226), .B2(n17142), .A(n17141), .ZN(P3_U2692) );
  AOI22_X1 U20314 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17153) );
  AOI22_X1 U20315 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20316 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17143) );
  OAI21_X1 U20317 ( .B1(n17144), .B2(n17220), .A(n17143), .ZN(n17150) );
  AOI22_X1 U20318 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20319 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20320 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U20321 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17145) );
  NAND4_X1 U20322 ( .A1(n17148), .A2(n17147), .A3(n17146), .A4(n17145), .ZN(
        n17149) );
  AOI211_X1 U20323 ( .C1(n17174), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17150), .B(n17149), .ZN(n17151) );
  NAND3_X1 U20324 ( .A1(n17153), .A2(n17152), .A3(n17151), .ZN(n17338) );
  OAI33_X1 U20325 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17170), .A3(n17321), 
        .B1(n17155), .B2(n17228), .B3(n17154), .ZN(n17156) );
  AOI21_X1 U20326 ( .B1(n17228), .B2(n17338), .A(n17156), .ZN(n17157) );
  INV_X1 U20327 ( .A(n17157), .ZN(P3_U2693) );
  AOI22_X1 U20328 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20329 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17181), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17125), .ZN(n17160) );
  AOI22_X1 U20330 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17177), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20331 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17158) );
  NAND4_X1 U20332 ( .A1(n17161), .A2(n17160), .A3(n17159), .A4(n17158), .ZN(
        n17169) );
  AOI22_X1 U20333 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17183), .ZN(n17167) );
  AOI22_X1 U20334 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17173), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20335 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17174), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17162), .ZN(n17165) );
  AOI22_X1 U20336 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17175), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17163), .ZN(n17164) );
  NAND4_X1 U20337 ( .A1(n17167), .A2(n17166), .A3(n17165), .A4(n17164), .ZN(
        n17168) );
  NOR2_X1 U20338 ( .A1(n17169), .A2(n17168), .ZN(n17342) );
  OAI211_X1 U20339 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n17171), .A(n17170), .B(
        n17225), .ZN(n17172) );
  OAI21_X1 U20340 ( .B1(n17342), .B2(n17225), .A(n17172), .ZN(P3_U2694) );
  AOI22_X1 U20341 ( .A1(n9730), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20342 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20343 ( .A1(n17177), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17178) );
  OAI21_X1 U20344 ( .B1(n17180), .B2(n17179), .A(n17178), .ZN(n17190) );
  AOI22_X1 U20345 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20346 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20347 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9725), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17186) );
  AOI22_X1 U20348 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17080), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17185) );
  NAND4_X1 U20349 ( .A1(n17188), .A2(n17187), .A3(n17186), .A4(n17185), .ZN(
        n17189) );
  AOI211_X1 U20350 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n17190), .B(n17189), .ZN(n17192) );
  NAND3_X1 U20351 ( .A1(n17194), .A2(n17193), .A3(n17192), .ZN(n17345) );
  INV_X1 U20352 ( .A(n17345), .ZN(n17197) );
  OAI21_X1 U20353 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17201), .A(n17195), .ZN(
        n17196) );
  AOI22_X1 U20354 ( .A1(n17228), .A2(n17197), .B1(n17196), .B2(n17225), .ZN(
        P3_U2695) );
  OAI21_X1 U20355 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17198), .A(n17225), .ZN(
        n17200) );
  OAI22_X1 U20356 ( .A1(n17201), .A2(n17200), .B1(n17199), .B2(n17225), .ZN(
        P3_U2696) );
  NAND2_X1 U20357 ( .A1(n18226), .A2(n17202), .ZN(n17204) );
  NOR2_X1 U20358 ( .A1(n17228), .A2(n17202), .ZN(n17205) );
  AOI22_X1 U20359 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17228), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17205), .ZN(n17203) );
  OAI21_X1 U20360 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17204), .A(n17203), .ZN(
        P3_U2697) );
  INV_X1 U20361 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17208) );
  OAI21_X1 U20362 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17206), .A(n17205), .ZN(
        n17207) );
  OAI21_X1 U20363 ( .B1(n17225), .B2(n17208), .A(n17207), .ZN(P3_U2698) );
  INV_X1 U20364 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17212) );
  OAI21_X1 U20365 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17210), .A(n17209), .ZN(
        n17211) );
  AOI22_X1 U20366 ( .A1(n17228), .A2(n17212), .B1(n17211), .B2(n17225), .ZN(
        P3_U2699) );
  NAND3_X1 U20367 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(n17223), .ZN(n17221) );
  NOR2_X1 U20368 ( .A1(n17213), .A2(n17221), .ZN(n17214) );
  AOI21_X1 U20369 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17225), .A(n17214), .ZN(
        n17218) );
  INV_X1 U20370 ( .A(n17223), .ZN(n17230) );
  NOR2_X1 U20371 ( .A1(n17215), .A2(n17230), .ZN(n17217) );
  INV_X1 U20372 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17216) );
  OAI22_X1 U20373 ( .A1(n17218), .A2(n17217), .B1(n17216), .B2(n17225), .ZN(
        P3_U2700) );
  NAND3_X1 U20374 ( .A1(n17221), .A2(P3_EBX_REG_2__SCAN_IN), .A3(n17225), .ZN(
        n17219) );
  OAI221_X1 U20375 ( .B1(n17221), .B2(P3_EBX_REG_2__SCAN_IN), .C1(n17225), 
        .C2(n17220), .A(n17219), .ZN(P3_U2701) );
  INV_X1 U20376 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20377 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n17227), .B1(n17223), .B2(
        n17222), .ZN(n17224) );
  OAI21_X1 U20378 ( .B1(n17226), .B2(n17225), .A(n17224), .ZN(P3_U2702) );
  AOI22_X1 U20379 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17228), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17227), .ZN(n17229) );
  OAI21_X1 U20380 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17230), .A(n17229), .ZN(
        P3_U2703) );
  INV_X1 U20381 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17472) );
  INV_X1 U20382 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17394) );
  INV_X1 U20383 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17398) );
  INV_X1 U20384 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17503) );
  NAND2_X1 U20385 ( .A1(n17231), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n17380) );
  NAND4_X1 U20386 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17232) );
  NOR2_X1 U20387 ( .A1(n17380), .A2(n17232), .ZN(n17233) );
  NAND4_X1 U20388 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .A4(n17233), .ZN(n17346) );
  NAND4_X1 U20389 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n17322)
         );
  NOR2_X1 U20390 ( .A1(n17346), .A2(n17322), .ZN(n17234) );
  NAND4_X1 U20391 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(n17234), .ZN(n17324) );
  NAND2_X1 U20392 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n17278) );
  NAND4_X1 U20393 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n17235)
         );
  NOR3_X2 U20394 ( .A1(n17312), .A2(n17278), .A3(n17235), .ZN(n17274) );
  NAND2_X1 U20395 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17274), .ZN(n17273) );
  NOR2_X2 U20396 ( .A1(n17321), .A2(n17273), .ZN(n17269) );
  NOR2_X2 U20397 ( .A1(n17398), .A2(n17268), .ZN(n17263) );
  NAND2_X1 U20398 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17255), .ZN(n17250) );
  NAND2_X1 U20399 ( .A1(n17243), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17239) );
  NOR2_X2 U20400 ( .A1(n18217), .A2(n17363), .ZN(n17310) );
  OAI22_X1 U20401 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17379), .B1(n17317), 
        .B2(n17243), .ZN(n17236) );
  AOI22_X1 U20402 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17310), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17236), .ZN(n17237) );
  OAI21_X1 U20403 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17239), .A(n17237), .ZN(
        P3_U2704) );
  NOR2_X2 U20404 ( .A1(n17238), .A2(n17363), .ZN(n17311) );
  AOI22_X1 U20405 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17311), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17310), .ZN(n17241) );
  OAI211_X1 U20406 ( .C1(n17243), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17363), .B(
        n17239), .ZN(n17240) );
  OAI211_X1 U20407 ( .C1(n17242), .C2(n17372), .A(n17241), .B(n17240), .ZN(
        P3_U2705) );
  INV_X1 U20408 ( .A(n17243), .ZN(n17245) );
  OAI21_X1 U20409 ( .B1(n17317), .B2(n17472), .A(n17250), .ZN(n17244) );
  AOI22_X1 U20410 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n17310), .B1(n17245), .B2(
        n17244), .ZN(n17248) );
  AOI22_X1 U20411 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17311), .B1(n17246), .B2(
        n17377), .ZN(n17247) );
  NAND2_X1 U20412 ( .A1(n17248), .A2(n17247), .ZN(P3_U2706) );
  INV_X1 U20413 ( .A(n17310), .ZN(n17297) );
  AOI22_X1 U20414 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17311), .B1(n17249), .B2(
        n17377), .ZN(n17252) );
  OAI211_X1 U20415 ( .C1(n17255), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17363), .B(
        n17250), .ZN(n17251) );
  OAI211_X1 U20416 ( .C1(n17297), .C2(n17253), .A(n17252), .B(n17251), .ZN(
        P3_U2707) );
  INV_X1 U20417 ( .A(n17311), .ZN(n17303) );
  AOI22_X1 U20418 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n17310), .B1(n17254), .B2(
        n17377), .ZN(n17258) );
  AOI211_X1 U20419 ( .C1(n17394), .C2(n17259), .A(n17255), .B(n17317), .ZN(
        n17256) );
  INV_X1 U20420 ( .A(n17256), .ZN(n17257) );
  OAI211_X1 U20421 ( .C1(n17303), .C2(n17490), .A(n17258), .B(n17257), .ZN(
        P3_U2708) );
  AOI22_X1 U20422 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17311), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17310), .ZN(n17261) );
  OAI211_X1 U20423 ( .C1(n17263), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17363), .B(
        n17259), .ZN(n17260) );
  OAI211_X1 U20424 ( .C1(n17372), .C2(n17262), .A(n17261), .B(n17260), .ZN(
        P3_U2709) );
  AOI22_X1 U20425 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17311), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17310), .ZN(n17266) );
  AOI211_X1 U20426 ( .C1(n17398), .C2(n17268), .A(n17263), .B(n17317), .ZN(
        n17264) );
  INV_X1 U20427 ( .A(n17264), .ZN(n17265) );
  OAI211_X1 U20428 ( .C1(n17372), .C2(n17267), .A(n17266), .B(n17265), .ZN(
        P3_U2710) );
  AOI22_X1 U20429 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17311), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17310), .ZN(n17271) );
  OAI211_X1 U20430 ( .C1(n17269), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17363), .B(
        n17268), .ZN(n17270) );
  OAI211_X1 U20431 ( .C1(n17372), .C2(n17272), .A(n17271), .B(n17270), .ZN(
        P3_U2711) );
  AOI22_X1 U20432 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17311), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17310), .ZN(n17276) );
  OAI211_X1 U20433 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17274), .A(n17273), .B(
        n17363), .ZN(n17275) );
  OAI211_X1 U20434 ( .C1(n17372), .C2(n17277), .A(n17276), .B(n17275), .ZN(
        P3_U2712) );
  INV_X1 U20435 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17408) );
  NOR3_X1 U20436 ( .A1(n17321), .A2(n17312), .A3(n17278), .ZN(n17299) );
  NAND2_X1 U20437 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17299), .ZN(n17294) );
  NAND2_X1 U20438 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17288), .ZN(n17285) );
  NAND2_X1 U20439 ( .A1(n17285), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17283) );
  OAI22_X1 U20440 ( .A1(n17280), .A2(n17372), .B1(n17279), .B2(n17297), .ZN(
        n17281) );
  AOI21_X1 U20441 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17311), .A(n17281), .ZN(
        n17282) );
  OAI221_X1 U20442 ( .B1(n17285), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17283), 
        .C2(n17317), .A(n17282), .ZN(P3_U2713) );
  AOI22_X1 U20443 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17311), .B1(n17377), .B2(
        n17284), .ZN(n17287) );
  OAI211_X1 U20444 ( .C1(n17288), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17363), .B(
        n17285), .ZN(n17286) );
  OAI211_X1 U20445 ( .C1(n17297), .C2(n18211), .A(n17287), .B(n17286), .ZN(
        P3_U2714) );
  AOI22_X1 U20446 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17311), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17310), .ZN(n17291) );
  AOI211_X1 U20447 ( .C1(n17408), .C2(n17294), .A(n17288), .B(n17317), .ZN(
        n17289) );
  INV_X1 U20448 ( .A(n17289), .ZN(n17290) );
  OAI211_X1 U20449 ( .C1(n17292), .C2(n17372), .A(n17291), .B(n17290), .ZN(
        P3_U2715) );
  AOI22_X1 U20450 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17311), .B1(n17377), .B2(
        n17293), .ZN(n17296) );
  OAI211_X1 U20451 ( .C1(n17299), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17363), .B(
        n17294), .ZN(n17295) );
  OAI211_X1 U20452 ( .C1(n17297), .C2(n18202), .A(n17296), .B(n17295), .ZN(
        P3_U2716) );
  AOI22_X1 U20453 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17310), .B1(n17377), .B2(
        n17298), .ZN(n17302) );
  INV_X1 U20454 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17458) );
  NOR2_X1 U20455 ( .A1(n17312), .A2(n17458), .ZN(n17304) );
  INV_X1 U20456 ( .A(n17299), .ZN(n17300) );
  OAI211_X1 U20457 ( .C1(n17304), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17363), .B(
        n17300), .ZN(n17301) );
  OAI211_X1 U20458 ( .C1(n17303), .C2(n18198), .A(n17302), .B(n17301), .ZN(
        P3_U2717) );
  AOI22_X1 U20459 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17311), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17310), .ZN(n17308) );
  INV_X1 U20460 ( .A(n17312), .ZN(n17306) );
  INV_X1 U20461 ( .A(n17304), .ZN(n17305) );
  OAI211_X1 U20462 ( .C1(n17306), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17363), .B(
        n17305), .ZN(n17307) );
  OAI211_X1 U20463 ( .C1(n17309), .C2(n17372), .A(n17308), .B(n17307), .ZN(
        P3_U2718) );
  AOI22_X1 U20464 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17311), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17310), .ZN(n17314) );
  OAI211_X1 U20465 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17316), .A(n17369), .B(
        n17312), .ZN(n17313) );
  OAI211_X1 U20466 ( .C1(n17315), .C2(n17372), .A(n17314), .B(n17313), .ZN(
        P3_U2719) );
  AOI211_X1 U20467 ( .C1(n17503), .C2(n17324), .A(n17317), .B(n17316), .ZN(
        n17318) );
  AOI21_X1 U20468 ( .B1(n17378), .B2(BUF2_REG_15__SCAN_IN), .A(n17318), .ZN(
        n17319) );
  OAI21_X1 U20469 ( .B1(n17320), .B2(n17372), .A(n17319), .ZN(P3_U2720) );
  NOR2_X1 U20470 ( .A1(n17321), .A2(n17346), .ZN(n17351) );
  NAND3_X1 U20471 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n17351), .ZN(n17340) );
  NOR2_X1 U20472 ( .A1(n17322), .A2(n17340), .ZN(n17330) );
  INV_X1 U20473 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17419) );
  AOI22_X1 U20474 ( .A1(n17377), .A2(n17323), .B1(n17330), .B2(n17419), .ZN(
        n17326) );
  NAND3_X1 U20475 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17369), .A3(n17324), 
        .ZN(n17325) );
  OAI211_X1 U20476 ( .C1(n17375), .C2(n17498), .A(n17326), .B(n17325), .ZN(
        P3_U2721) );
  INV_X1 U20477 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17426) );
  NOR3_X1 U20478 ( .A1(n17424), .A2(n17426), .A3(n17340), .ZN(n17331) );
  AND2_X1 U20479 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17331), .ZN(n17334) );
  AOI21_X1 U20480 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17369), .A(n17334), .ZN(
        n17329) );
  AOI22_X1 U20481 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17378), .B1(n17377), .B2(
        n17327), .ZN(n17328) );
  OAI21_X1 U20482 ( .B1(n17330), .B2(n17329), .A(n17328), .ZN(P3_U2722) );
  AOI21_X1 U20483 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17369), .A(n17331), .ZN(
        n17333) );
  OAI222_X1 U20484 ( .A1(n17375), .A2(n17492), .B1(n17334), .B2(n17333), .C1(
        n17372), .C2(n17332), .ZN(P3_U2723) );
  INV_X1 U20485 ( .A(n17340), .ZN(n17344) );
  NAND2_X1 U20486 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17344), .ZN(n17337) );
  OAI21_X1 U20487 ( .B1(n17426), .B2(n17340), .A(n17363), .ZN(n17341) );
  AOI22_X1 U20488 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17378), .B1(n17377), .B2(
        n17335), .ZN(n17336) );
  OAI221_X1 U20489 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17337), .C1(n17424), 
        .C2(n17341), .A(n17336), .ZN(P3_U2724) );
  AOI22_X1 U20490 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17378), .B1(n17377), .B2(
        n17338), .ZN(n17339) );
  OAI221_X1 U20491 ( .B1(n17341), .B2(n17426), .C1(n17341), .C2(n17340), .A(
        n17339), .ZN(P3_U2725) );
  AOI22_X1 U20492 ( .A1(n17351), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17363), .ZN(n17343) );
  OAI222_X1 U20493 ( .A1(n17375), .A2(n17486), .B1(n17344), .B2(n17343), .C1(
        n17372), .C2(n17342), .ZN(P3_U2726) );
  INV_X1 U20494 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20495 ( .A1(n17377), .A2(n17345), .B1(n17351), .B2(n17430), .ZN(
        n17348) );
  NAND3_X1 U20496 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17369), .A3(n17346), .ZN(
        n17347) );
  OAI211_X1 U20497 ( .C1(n17375), .C2(n17484), .A(n17348), .B(n17347), .ZN(
        P3_U2727) );
  INV_X1 U20498 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17434) );
  INV_X1 U20499 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17439) );
  INV_X1 U20500 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17445) );
  NOR2_X1 U20501 ( .A1(n17452), .A2(n17379), .ZN(n17382) );
  NAND2_X1 U20502 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17382), .ZN(n17367) );
  NOR2_X1 U20503 ( .A1(n17445), .A2(n17367), .ZN(n17374) );
  NAND2_X1 U20504 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17374), .ZN(n17359) );
  NOR2_X1 U20505 ( .A1(n17439), .A2(n17359), .ZN(n17362) );
  NAND2_X1 U20506 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17362), .ZN(n17352) );
  NOR2_X1 U20507 ( .A1(n17434), .A2(n17352), .ZN(n17355) );
  AOI21_X1 U20508 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17369), .A(n17355), .ZN(
        n17350) );
  OAI222_X1 U20509 ( .A1(n17375), .A2(n18223), .B1(n17351), .B2(n17350), .C1(
        n17372), .C2(n17349), .ZN(P3_U2728) );
  INV_X1 U20510 ( .A(n17352), .ZN(n17358) );
  AOI21_X1 U20511 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17369), .A(n17358), .ZN(
        n17354) );
  OAI222_X1 U20512 ( .A1(n17375), .A2(n18216), .B1(n17355), .B2(n17354), .C1(
        n17372), .C2(n17353), .ZN(P3_U2729) );
  AOI21_X1 U20513 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17369), .A(n17362), .ZN(
        n17357) );
  OAI222_X1 U20514 ( .A1(n17375), .A2(n18212), .B1(n17358), .B2(n17357), .C1(
        n17372), .C2(n17356), .ZN(P3_U2730) );
  INV_X1 U20515 ( .A(n17359), .ZN(n17366) );
  AOI21_X1 U20516 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17363), .A(n17366), .ZN(
        n17361) );
  OAI222_X1 U20517 ( .A1(n17375), .A2(n18207), .B1(n17362), .B2(n17361), .C1(
        n17372), .C2(n17360), .ZN(P3_U2731) );
  AOI21_X1 U20518 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17363), .A(n17374), .ZN(
        n17365) );
  OAI222_X1 U20519 ( .A1(n17375), .A2(n18203), .B1(n17366), .B2(n17365), .C1(
        n17372), .C2(n17364), .ZN(P3_U2732) );
  INV_X1 U20520 ( .A(n17367), .ZN(n17368) );
  AOI21_X1 U20521 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17369), .A(n17368), .ZN(
        n17373) );
  INV_X1 U20522 ( .A(n17370), .ZN(n17371) );
  OAI222_X1 U20523 ( .A1(n18198), .A2(n17375), .B1(n17374), .B2(n17373), .C1(
        n17372), .C2(n17371), .ZN(P3_U2733) );
  AOI22_X1 U20524 ( .A1(n17378), .A2(BUF2_REG_1__SCAN_IN), .B1(n17377), .B2(
        n17376), .ZN(n17384) );
  NOR2_X1 U20525 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17379), .ZN(n17381) );
  OAI22_X1 U20526 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17382), .B1(n17381), .B2(
        n17380), .ZN(n17383) );
  NAND2_X1 U20527 ( .A1(n17384), .A2(n17383), .ZN(P3_U2734) );
  OR2_X1 U20528 ( .A1(n18810), .A2(n17668), .ZN(n17436) );
  NOR2_X1 U20529 ( .A1(n17442), .A2(n17386), .ZN(P3_U2736) );
  INV_X1 U20530 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17389) );
  NAND2_X1 U20531 ( .A1(n17440), .A2(n17387), .ZN(n17416) );
  INV_X2 U20532 ( .A(n17436), .ZN(n17449) );
  AOI22_X1 U20533 ( .A1(n17449), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17388) );
  OAI21_X1 U20534 ( .B1(n17389), .B2(n17416), .A(n17388), .ZN(P3_U2737) );
  AOI22_X1 U20535 ( .A1(n17449), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20536 ( .B1(n17472), .B2(n17416), .A(n17390), .ZN(P3_U2738) );
  INV_X1 U20537 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20538 ( .A1(n17449), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U20539 ( .B1(n17392), .B2(n17416), .A(n17391), .ZN(P3_U2739) );
  AOI22_X1 U20540 ( .A1(n17449), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17393) );
  OAI21_X1 U20541 ( .B1(n17394), .B2(n17416), .A(n17393), .ZN(P3_U2740) );
  INV_X1 U20542 ( .A(n17416), .ZN(n17411) );
  AOI22_X1 U20543 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17411), .B1(n17449), 
        .B2(P3_UWORD_REG_10__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20544 ( .B1(n17396), .B2(n17442), .A(n17395), .ZN(P3_U2741) );
  AOI22_X1 U20545 ( .A1(n17449), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17397) );
  OAI21_X1 U20546 ( .B1(n17398), .B2(n17416), .A(n17397), .ZN(P3_U2742) );
  AOI22_X1 U20547 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17411), .B1(n17449), 
        .B2(P3_UWORD_REG_8__SCAN_IN), .ZN(n17399) );
  OAI21_X1 U20548 ( .B1(n17400), .B2(n17442), .A(n17399), .ZN(P3_U2743) );
  AOI22_X1 U20549 ( .A1(P3_DATAO_REG_23__SCAN_IN), .A2(n17448), .B1(n17449), 
        .B2(P3_UWORD_REG_7__SCAN_IN), .ZN(n17401) );
  OAI21_X1 U20550 ( .B1(n17402), .B2(n17416), .A(n17401), .ZN(P3_U2744) );
  INV_X1 U20551 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17404) );
  AOI22_X1 U20552 ( .A1(n17449), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20553 ( .B1(n17404), .B2(n17416), .A(n17403), .ZN(P3_U2745) );
  INV_X1 U20554 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U20555 ( .A1(n17449), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20556 ( .B1(n17406), .B2(n17416), .A(n17405), .ZN(P3_U2746) );
  AOI22_X1 U20557 ( .A1(n17449), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17407) );
  OAI21_X1 U20558 ( .B1(n17408), .B2(n17416), .A(n17407), .ZN(P3_U2747) );
  INV_X1 U20559 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U20560 ( .A1(n17449), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20561 ( .B1(n17410), .B2(n17416), .A(n17409), .ZN(P3_U2748) );
  AOI22_X1 U20562 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17411), .B1(n17449), 
        .B2(P3_UWORD_REG_2__SCAN_IN), .ZN(n17412) );
  OAI21_X1 U20563 ( .B1(n17413), .B2(n17442), .A(n17412), .ZN(P3_U2749) );
  AOI22_X1 U20564 ( .A1(n17449), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17414) );
  OAI21_X1 U20565 ( .B1(n17458), .B2(n17416), .A(n17414), .ZN(P3_U2750) );
  INV_X1 U20566 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U20567 ( .A1(n17449), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17415) );
  OAI21_X1 U20568 ( .B1(n17456), .B2(n17416), .A(n17415), .ZN(P3_U2751) );
  AOI22_X1 U20569 ( .A1(n17449), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17417) );
  OAI21_X1 U20570 ( .B1(n17503), .B2(n17451), .A(n17417), .ZN(P3_U2752) );
  AOI22_X1 U20571 ( .A1(n17449), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U20572 ( .B1(n17419), .B2(n17451), .A(n17418), .ZN(P3_U2753) );
  INV_X1 U20573 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U20574 ( .A1(n17449), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17420) );
  OAI21_X1 U20575 ( .B1(n17494), .B2(n17451), .A(n17420), .ZN(P3_U2754) );
  INV_X1 U20576 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20577 ( .A1(n17449), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17446), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17421) );
  OAI21_X1 U20578 ( .B1(n17422), .B2(n17451), .A(n17421), .ZN(P3_U2755) );
  AOI22_X1 U20579 ( .A1(n17449), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17446), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17423) );
  OAI21_X1 U20580 ( .B1(n17424), .B2(n17451), .A(n17423), .ZN(P3_U2756) );
  AOI22_X1 U20581 ( .A1(n17449), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17446), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17425) );
  OAI21_X1 U20582 ( .B1(n17426), .B2(n17451), .A(n17425), .ZN(P3_U2757) );
  INV_X1 U20583 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20584 ( .A1(n17449), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17446), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17427) );
  OAI21_X1 U20585 ( .B1(n17428), .B2(n17451), .A(n17427), .ZN(P3_U2758) );
  AOI22_X1 U20586 ( .A1(n17449), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17446), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17429) );
  OAI21_X1 U20587 ( .B1(n17430), .B2(n17451), .A(n17429), .ZN(P3_U2759) );
  AOI22_X1 U20588 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17440), .B1(n17449), .B2(
        P3_LWORD_REG_7__SCAN_IN), .ZN(n17431) );
  OAI21_X1 U20589 ( .B1(n17432), .B2(n17442), .A(n17431), .ZN(P3_U2760) );
  AOI22_X1 U20590 ( .A1(P3_LWORD_REG_6__SCAN_IN), .A2(n17449), .B1(n17448), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17433) );
  OAI21_X1 U20591 ( .B1(n17434), .B2(n17451), .A(n17433), .ZN(P3_U2761) );
  AOI22_X1 U20592 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17440), .B1(n17448), .B2(
        P3_DATAO_REG_5__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20593 ( .B1(n17437), .B2(n17436), .A(n17435), .ZN(P3_U2762) );
  AOI22_X1 U20594 ( .A1(n17449), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17446), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17438) );
  OAI21_X1 U20595 ( .B1(n17439), .B2(n17451), .A(n17438), .ZN(P3_U2763) );
  AOI22_X1 U20596 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17440), .B1(n17449), .B2(
        P3_LWORD_REG_3__SCAN_IN), .ZN(n17441) );
  OAI21_X1 U20597 ( .B1(n17443), .B2(n17442), .A(n17441), .ZN(P3_U2764) );
  AOI22_X1 U20598 ( .A1(n17449), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17446), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17444) );
  OAI21_X1 U20599 ( .B1(n17445), .B2(n17451), .A(n17444), .ZN(P3_U2765) );
  INV_X1 U20600 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20601 ( .A1(n17449), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17446), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20602 ( .B1(n17476), .B2(n17451), .A(n17447), .ZN(P3_U2766) );
  AOI22_X1 U20603 ( .A1(n17449), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17448), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17450) );
  OAI21_X1 U20604 ( .B1(n17452), .B2(n17451), .A(n17450), .ZN(P3_U2767) );
  NAND3_X1 U20605 ( .A1(n18850), .A2(n17454), .A3(n17453), .ZN(n17502) );
  AOI22_X1 U20606 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17500), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17499), .ZN(n17455) );
  OAI21_X1 U20607 ( .B1(n17456), .B2(n17502), .A(n17455), .ZN(P3_U2768) );
  AOI22_X1 U20608 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17500), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17499), .ZN(n17457) );
  OAI21_X1 U20609 ( .B1(n17458), .B2(n17502), .A(n17457), .ZN(P3_U2769) );
  AOI22_X1 U20610 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17499), .ZN(n17459) );
  OAI21_X1 U20611 ( .B1(n18198), .B2(n17497), .A(n17459), .ZN(P3_U2770) );
  AOI22_X1 U20612 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17469), .ZN(n17460) );
  OAI21_X1 U20613 ( .B1(n18203), .B2(n17497), .A(n17460), .ZN(P3_U2771) );
  AOI22_X1 U20614 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17469), .ZN(n17461) );
  OAI21_X1 U20615 ( .B1(n18207), .B2(n17497), .A(n17461), .ZN(P3_U2772) );
  AOI22_X1 U20616 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17469), .ZN(n17462) );
  OAI21_X1 U20617 ( .B1(n18212), .B2(n17497), .A(n17462), .ZN(P3_U2773) );
  AOI22_X1 U20618 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17469), .ZN(n17463) );
  OAI21_X1 U20619 ( .B1(n18216), .B2(n17497), .A(n17463), .ZN(P3_U2774) );
  AOI22_X1 U20620 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17469), .ZN(n17464) );
  OAI21_X1 U20621 ( .B1(n18223), .B2(n17497), .A(n17464), .ZN(P3_U2775) );
  AOI22_X1 U20622 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17469), .ZN(n17465) );
  OAI21_X1 U20623 ( .B1(n17484), .B2(n17497), .A(n17465), .ZN(P3_U2776) );
  AOI22_X1 U20624 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17469), .ZN(n17466) );
  OAI21_X1 U20625 ( .B1(n17486), .B2(n17497), .A(n17466), .ZN(P3_U2777) );
  AOI22_X1 U20626 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17469), .ZN(n17467) );
  OAI21_X1 U20627 ( .B1(n17488), .B2(n17497), .A(n17467), .ZN(P3_U2778) );
  AOI22_X1 U20628 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17469), .ZN(n17468) );
  OAI21_X1 U20629 ( .B1(n17490), .B2(n17497), .A(n17468), .ZN(P3_U2779) );
  AOI22_X1 U20630 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17469), .ZN(n17470) );
  OAI21_X1 U20631 ( .B1(n17492), .B2(n17497), .A(n17470), .ZN(P3_U2780) );
  AOI22_X1 U20632 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17500), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17499), .ZN(n17471) );
  OAI21_X1 U20633 ( .B1(n17472), .B2(n17502), .A(n17471), .ZN(P3_U2781) );
  AOI22_X1 U20634 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17495), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17499), .ZN(n17473) );
  OAI21_X1 U20635 ( .B1(n17498), .B2(n17497), .A(n17473), .ZN(P3_U2782) );
  AOI22_X1 U20636 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17499), .ZN(n17474) );
  OAI21_X1 U20637 ( .B1(n18186), .B2(n17497), .A(n17474), .ZN(P3_U2783) );
  AOI22_X1 U20638 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17500), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17499), .ZN(n17475) );
  OAI21_X1 U20639 ( .B1(n17476), .B2(n17502), .A(n17475), .ZN(P3_U2784) );
  AOI22_X1 U20640 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17499), .ZN(n17477) );
  OAI21_X1 U20641 ( .B1(n18198), .B2(n17497), .A(n17477), .ZN(P3_U2785) );
  AOI22_X1 U20642 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17499), .ZN(n17478) );
  OAI21_X1 U20643 ( .B1(n18203), .B2(n17497), .A(n17478), .ZN(P3_U2786) );
  AOI22_X1 U20644 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17499), .ZN(n17479) );
  OAI21_X1 U20645 ( .B1(n18207), .B2(n17497), .A(n17479), .ZN(P3_U2787) );
  AOI22_X1 U20646 ( .A1(P3_LWORD_REG_5__SCAN_IN), .A2(n17499), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n17495), .ZN(n17480) );
  OAI21_X1 U20647 ( .B1(n18212), .B2(n17497), .A(n17480), .ZN(P3_U2788) );
  AOI22_X1 U20648 ( .A1(P3_LWORD_REG_6__SCAN_IN), .A2(n17499), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17495), .ZN(n17481) );
  OAI21_X1 U20649 ( .B1(n18216), .B2(n17497), .A(n17481), .ZN(P3_U2789) );
  AOI22_X1 U20650 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17499), .ZN(n17482) );
  OAI21_X1 U20651 ( .B1(n18223), .B2(n17497), .A(n17482), .ZN(P3_U2790) );
  AOI22_X1 U20652 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17499), .ZN(n17483) );
  OAI21_X1 U20653 ( .B1(n17484), .B2(n17497), .A(n17483), .ZN(P3_U2791) );
  AOI22_X1 U20654 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17499), .ZN(n17485) );
  OAI21_X1 U20655 ( .B1(n17486), .B2(n17497), .A(n17485), .ZN(P3_U2792) );
  AOI22_X1 U20656 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17499), .ZN(n17487) );
  OAI21_X1 U20657 ( .B1(n17488), .B2(n17497), .A(n17487), .ZN(P3_U2793) );
  AOI22_X1 U20658 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17499), .ZN(n17489) );
  OAI21_X1 U20659 ( .B1(n17490), .B2(n17497), .A(n17489), .ZN(P3_U2794) );
  AOI22_X1 U20660 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17499), .ZN(n17491) );
  OAI21_X1 U20661 ( .B1(n17492), .B2(n17497), .A(n17491), .ZN(P3_U2795) );
  AOI22_X1 U20662 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17500), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17499), .ZN(n17493) );
  OAI21_X1 U20663 ( .B1(n17494), .B2(n17502), .A(n17493), .ZN(P3_U2796) );
  AOI22_X1 U20664 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17495), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17499), .ZN(n17496) );
  OAI21_X1 U20665 ( .B1(n17498), .B2(n17497), .A(n17496), .ZN(P3_U2797) );
  AOI22_X1 U20666 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17500), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17499), .ZN(n17501) );
  OAI21_X1 U20667 ( .B1(n17503), .B2(n17502), .A(n17501), .ZN(P3_U2798) );
  OAI21_X1 U20668 ( .B1(n17514), .B2(n17846), .A(n17872), .ZN(n17504) );
  AOI21_X1 U20669 ( .B1(n17712), .B2(n9805), .A(n17504), .ZN(n17535) );
  OAI21_X1 U20670 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17618), .A(
        n17535), .ZN(n17526) );
  AOI22_X1 U20671 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17526), .B1(
        n17729), .B2(n17505), .ZN(n17519) );
  NOR2_X1 U20672 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17529), .ZN(
        n17513) );
  NOR2_X1 U20673 ( .A1(n17824), .A2(n17788), .ZN(n17596) );
  OAI22_X1 U20674 ( .A1(n17881), .A2(n17877), .B1(n17880), .B2(n17748), .ZN(
        n17543) );
  NOR2_X1 U20675 ( .A1(n17529), .A2(n17543), .ZN(n17507) );
  NOR3_X1 U20676 ( .A1(n17596), .A2(n17507), .A3(n17506), .ZN(n17512) );
  AOI211_X1 U20677 ( .C1(n17510), .C2(n17509), .A(n17508), .B(n17756), .ZN(
        n17511) );
  AOI211_X1 U20678 ( .C1(n17530), .C2(n17513), .A(n17512), .B(n17511), .ZN(
        n17518) );
  AND2_X1 U20679 ( .A1(n17707), .A2(n17514), .ZN(n17528) );
  NAND2_X1 U20680 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17515) );
  OAI211_X1 U20681 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17528), .B(n17515), .ZN(n17516) );
  NAND4_X1 U20682 ( .A1(n17519), .A2(n17518), .A3(n17517), .A4(n17516), .ZN(
        P3_U2802) );
  INV_X1 U20683 ( .A(n17520), .ZN(n17522) );
  NAND2_X1 U20684 ( .A1(n17522), .A2(n17521), .ZN(n17523) );
  XNOR2_X1 U20685 ( .A(n17786), .B(n17523), .ZN(n17889) );
  INV_X1 U20686 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17527) );
  OAI22_X1 U20687 ( .A1(n18162), .A2(n18782), .B1(n17682), .B2(n17524), .ZN(
        n17525) );
  AOI221_X1 U20688 ( .B1(n17528), .B2(n17527), .C1(n17526), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17525), .ZN(n17532) );
  AOI22_X1 U20689 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17543), .B1(
        n17530), .B2(n17529), .ZN(n17531) );
  OAI211_X1 U20690 ( .C1(n17889), .C2(n17756), .A(n17532), .B(n17531), .ZN(
        P3_U2803) );
  INV_X1 U20691 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17891) );
  NAND3_X1 U20692 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n17891), .ZN(n17890) );
  INV_X2 U20693 ( .A(n17613), .ZN(n17677) );
  NAND2_X1 U20694 ( .A1(n17912), .A2(n17677), .ZN(n17569) );
  AOI21_X1 U20695 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17534), .A(
        n17533), .ZN(n17896) );
  INV_X1 U20696 ( .A(n17618), .ZN(n17539) );
  AOI221_X1 U20697 ( .B1(n18221), .B2(n17537), .C1(n17536), .C2(n17537), .A(
        n17535), .ZN(n17538) );
  AOI221_X1 U20698 ( .B1(n17729), .B2(n17540), .C1(n17539), .C2(n17540), .A(
        n17538), .ZN(n17541) );
  NAND2_X1 U20699 ( .A1(n9724), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17894) );
  OAI211_X1 U20700 ( .C1(n17896), .C2(n17756), .A(n17541), .B(n17894), .ZN(
        n17542) );
  AOI21_X1 U20701 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17543), .A(
        n17542), .ZN(n17544) );
  OAI21_X1 U20702 ( .B1(n17890), .B2(n17569), .A(n17544), .ZN(P3_U2804) );
  OAI21_X1 U20703 ( .B1(n17610), .B2(n17546), .A(n17545), .ZN(n17547) );
  XNOR2_X1 U20704 ( .A(n17547), .B(n17904), .ZN(n17909) );
  INV_X1 U20705 ( .A(n17548), .ZN(n17550) );
  INV_X1 U20706 ( .A(n17872), .ZN(n17860) );
  AOI21_X1 U20707 ( .B1(n18577), .B2(n17550), .A(n17860), .ZN(n17577) );
  OAI21_X1 U20708 ( .B1(n17549), .B2(n17668), .A(n17577), .ZN(n17561) );
  INV_X1 U20709 ( .A(n17707), .ZN(n17680) );
  NOR2_X1 U20710 ( .A1(n17680), .A2(n17550), .ZN(n17563) );
  OAI211_X1 U20711 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17563), .B(n17551), .ZN(n17552) );
  NAND2_X1 U20712 ( .A1(n9724), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17907) );
  OAI211_X1 U20713 ( .C1(n17682), .C2(n17553), .A(n17552), .B(n17907), .ZN(
        n17554) );
  AOI21_X1 U20714 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17561), .A(
        n17554), .ZN(n17558) );
  NAND3_X1 U20715 ( .A1(n18010), .A2(n17912), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17555) );
  XNOR2_X1 U20716 ( .A(n17555), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17901) );
  INV_X1 U20717 ( .A(n17912), .ZN(n17564) );
  NOR2_X1 U20718 ( .A1(n17939), .A2(n17564), .ZN(n17916) );
  NAND2_X1 U20719 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17916), .ZN(
        n17556) );
  XNOR2_X1 U20720 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17556), .ZN(
        n17900) );
  AOI22_X1 U20721 ( .A1(n17824), .A2(n17901), .B1(n17788), .B2(n17900), .ZN(
        n17557) );
  OAI211_X1 U20722 ( .C1(n17756), .C2(n17909), .A(n17558), .B(n17557), .ZN(
        P3_U2805) );
  INV_X1 U20723 ( .A(n17559), .ZN(n17573) );
  NOR2_X1 U20724 ( .A1(n18162), .A2(n18776), .ZN(n17560) );
  AOI221_X1 U20725 ( .B1(n17563), .B2(n17562), .C1(n17561), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17560), .ZN(n17572) );
  NOR2_X1 U20726 ( .A1(n17565), .A2(n17564), .ZN(n17566) );
  OAI22_X1 U20727 ( .A1(n17566), .A2(n17877), .B1(n17916), .B2(n17748), .ZN(
        n17584) );
  AOI21_X1 U20728 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17568), .A(
        n17567), .ZN(n17923) );
  OAI22_X1 U20729 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17569), .B1(
        n17923), .B2(n17756), .ZN(n17570) );
  AOI21_X1 U20730 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17584), .A(
        n17570), .ZN(n17571) );
  OAI211_X1 U20731 ( .C1(n17682), .C2(n17573), .A(n17572), .B(n17571), .ZN(
        P3_U2806) );
  AOI22_X1 U20732 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17610), .B1(
        n17574), .B2(n17593), .ZN(n17575) );
  NAND2_X1 U20733 ( .A1(n17622), .A2(n17575), .ZN(n17576) );
  XNOR2_X1 U20734 ( .A(n17576), .B(n17917), .ZN(n17930) );
  AOI221_X1 U20735 ( .B1(n17578), .B2(n17577), .C1(n17668), .C2(n17577), .A(
        n9872), .ZN(n17583) );
  NAND2_X1 U20736 ( .A1(n9724), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17928) );
  NOR2_X1 U20737 ( .A1(n17680), .A2(n17590), .ZN(n17608) );
  NAND3_X1 U20738 ( .A1(n17579), .A2(n17608), .A3(n9872), .ZN(n17580) );
  OAI211_X1 U20739 ( .C1(n17682), .C2(n17581), .A(n17928), .B(n17580), .ZN(
        n17582) );
  AOI211_X1 U20740 ( .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17584), .A(
        n17583), .B(n17582), .ZN(n17587) );
  NAND3_X1 U20741 ( .A1(n17585), .A2(n17677), .A3(n17917), .ZN(n17586) );
  OAI211_X1 U20742 ( .C1(n17930), .C2(n17756), .A(n17587), .B(n17586), .ZN(
        P3_U2807) );
  OAI21_X1 U20743 ( .B1(n9740), .B2(n17668), .A(n17872), .ZN(n17589) );
  AOI21_X1 U20744 ( .B1(n17667), .B2(n17590), .A(n17589), .ZN(n17629) );
  OAI21_X1 U20745 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17618), .A(
        n17629), .ZN(n17606) );
  AOI22_X1 U20746 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17606), .B1(
        n17729), .B2(n17591), .ZN(n17603) );
  INV_X1 U20747 ( .A(n17622), .ZN(n17592) );
  AOI221_X1 U20748 ( .B1(n17595), .B2(n17593), .C1(n17609), .C2(n17593), .A(
        n17592), .ZN(n17594) );
  XNOR2_X1 U20749 ( .A(n17594), .B(n17948), .ZN(n17945) );
  INV_X1 U20750 ( .A(n17982), .ZN(n17651) );
  OR2_X1 U20751 ( .A1(n17651), .A2(n17595), .ZN(n17940) );
  NOR2_X1 U20752 ( .A1(n17613), .A2(n17940), .ZN(n17598) );
  INV_X1 U20753 ( .A(n17596), .ZN(n17621) );
  NAND2_X1 U20754 ( .A1(n17788), .A2(n17939), .ZN(n17694) );
  OAI21_X1 U20755 ( .B1(n18010), .B2(n17877), .A(n17694), .ZN(n17676) );
  AOI21_X1 U20756 ( .B1(n17621), .B2(n17940), .A(n17676), .ZN(n17616) );
  INV_X1 U20757 ( .A(n17616), .ZN(n17597) );
  MUX2_X1 U20758 ( .A(n17598), .B(n17597), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17599) );
  AOI21_X1 U20759 ( .B1(n17787), .B2(n17945), .A(n17599), .ZN(n17602) );
  NAND2_X1 U20760 ( .A1(n9724), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17946) );
  OAI211_X1 U20761 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17608), .B(n17600), .ZN(n17601) );
  NAND4_X1 U20762 ( .A1(n17603), .A2(n17602), .A3(n17946), .A4(n17601), .ZN(
        P3_U2808) );
  OAI22_X1 U20763 ( .A1(n18162), .A2(n18771), .B1(n17682), .B2(n17604), .ZN(
        n17605) );
  AOI221_X1 U20764 ( .B1(n17608), .B2(n17607), .C1(n17606), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17605), .ZN(n17615) );
  NOR3_X1 U20765 ( .A1(n17654), .A2(n17610), .A3(n17609), .ZN(n17632) );
  INV_X1 U20766 ( .A(n17649), .ZN(n17633) );
  AOI22_X1 U20767 ( .A1(n17952), .A2(n17632), .B1(n17633), .B2(n17611), .ZN(
        n17612) );
  XNOR2_X1 U20768 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17612), .ZN(
        n17956) );
  INV_X1 U20769 ( .A(n17952), .ZN(n17937) );
  NOR2_X1 U20770 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17937), .ZN(
        n17955) );
  NAND2_X1 U20771 ( .A1(n17982), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17954) );
  NOR2_X1 U20772 ( .A1(n17613), .A2(n17954), .ZN(n17637) );
  AOI22_X1 U20773 ( .A1(n17787), .A2(n17956), .B1(n17955), .B2(n17637), .ZN(
        n17614) );
  OAI211_X1 U20774 ( .C1(n17616), .C2(n17936), .A(n17615), .B(n17614), .ZN(
        P3_U2809) );
  AOI21_X1 U20775 ( .B1(n18577), .B2(n17617), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17628) );
  INV_X1 U20776 ( .A(n17857), .ZN(n17619) );
  AOI22_X1 U20777 ( .A1(n9724), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17620), 
        .B2(n17619), .ZN(n17627) );
  NOR2_X1 U20778 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17968), .ZN(
        n17959) );
  NOR2_X1 U20779 ( .A1(n17968), .A2(n17954), .ZN(n17934) );
  INV_X1 U20780 ( .A(n17934), .ZN(n17962) );
  AOI21_X1 U20781 ( .B1(n17621), .B2(n17962), .A(n17676), .ZN(n17635) );
  OAI221_X1 U20782 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17648), 
        .C1(n17968), .C2(n17632), .A(n17622), .ZN(n17623) );
  XNOR2_X1 U20783 ( .A(n17624), .B(n17623), .ZN(n17967) );
  OAI22_X1 U20784 ( .A1(n17635), .A2(n17624), .B1(n17756), .B2(n17967), .ZN(
        n17625) );
  AOI21_X1 U20785 ( .B1(n17959), .B2(n17637), .A(n17625), .ZN(n17626) );
  OAI211_X1 U20786 ( .C1(n17629), .C2(n17628), .A(n17627), .B(n17626), .ZN(
        P3_U2810) );
  AOI21_X1 U20787 ( .B1(n17667), .B2(n17638), .A(n17860), .ZN(n17663) );
  OAI21_X1 U20788 ( .B1(n17630), .B2(n17668), .A(n17663), .ZN(n17645) );
  AOI22_X1 U20789 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17645), .B1(
        n17729), .B2(n17631), .ZN(n17642) );
  AOI21_X1 U20790 ( .B1(n17633), .B2(n17648), .A(n17632), .ZN(n17634) );
  XNOR2_X1 U20791 ( .A(n17634), .B(n17968), .ZN(n17973) );
  OAI22_X1 U20792 ( .A1(n17973), .A2(n17756), .B1(n17635), .B2(n17968), .ZN(
        n17636) );
  AOI21_X1 U20793 ( .B1(n17637), .B2(n17968), .A(n17636), .ZN(n17641) );
  NAND2_X1 U20794 ( .A1(n9724), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17971) );
  NOR2_X1 U20795 ( .A1(n17680), .A2(n17638), .ZN(n17647) );
  OAI211_X1 U20796 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17647), .B(n17639), .ZN(n17640) );
  NAND4_X1 U20797 ( .A1(n17642), .A2(n17641), .A3(n17971), .A4(n17640), .ZN(
        P3_U2811) );
  AOI21_X1 U20798 ( .B1(n17677), .B2(n17651), .A(n17676), .ZN(n17659) );
  INV_X1 U20799 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18764) );
  OAI22_X1 U20800 ( .A1(n18162), .A2(n18764), .B1(n17682), .B2(n17643), .ZN(
        n17644) );
  AOI221_X1 U20801 ( .B1(n17647), .B2(n17646), .C1(n17645), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17644), .ZN(n17653) );
  AOI21_X1 U20802 ( .B1(n17786), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17648), .ZN(n17650) );
  XNOR2_X1 U20803 ( .A(n17650), .B(n17649), .ZN(n17987) );
  NOR2_X1 U20804 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17651), .ZN(
        n17986) );
  AOI22_X1 U20805 ( .A1(n17787), .A2(n17987), .B1(n17677), .B2(n17986), .ZN(
        n17652) );
  OAI211_X1 U20806 ( .C1(n17659), .C2(n17654), .A(n17653), .B(n17652), .ZN(
        P3_U2812) );
  AOI21_X1 U20807 ( .B1(n17655), .B2(n18577), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17664) );
  OAI21_X1 U20808 ( .B1(n17657), .B2(n17983), .A(n17656), .ZN(n17991) );
  AOI21_X1 U20809 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17677), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17658) );
  OAI22_X1 U20810 ( .A1(n17857), .A2(n17660), .B1(n17659), .B2(n17658), .ZN(
        n17661) );
  AOI21_X1 U20811 ( .B1(n17787), .B2(n17991), .A(n17661), .ZN(n17662) );
  NAND2_X1 U20812 ( .A1(n9724), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17994) );
  OAI211_X1 U20813 ( .C1(n17664), .C2(n17663), .A(n17662), .B(n17994), .ZN(
        P3_U2813) );
  NAND2_X1 U20814 ( .A1(n17786), .A2(n17784), .ZN(n17766) );
  OAI22_X1 U20815 ( .A1(n17786), .A2(n17665), .B1(n17766), .B2(n17938), .ZN(
        n17666) );
  XNOR2_X1 U20816 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17666), .ZN(
        n18005) );
  AOI21_X1 U20817 ( .B1(n17667), .B2(n17679), .A(n17860), .ZN(n17700) );
  OAI21_X1 U20818 ( .B1(n17669), .B2(n17668), .A(n17700), .ZN(n17684) );
  INV_X1 U20819 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17670) );
  AOI211_X1 U20820 ( .C1(n17670), .C2(n17685), .A(n17680), .B(n17679), .ZN(
        n17672) );
  AOI22_X1 U20821 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17684), .B1(
        n17672), .B2(n17671), .ZN(n17673) );
  NAND2_X1 U20822 ( .A1(n9724), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18003) );
  OAI211_X1 U20823 ( .C1(n17682), .C2(n17674), .A(n17673), .B(n18003), .ZN(
        n17675) );
  AOI221_X1 U20824 ( .B1(n17677), .B2(n15584), .C1(n17676), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17675), .ZN(n17678) );
  OAI21_X1 U20825 ( .B1(n18005), .B2(n17756), .A(n17678), .ZN(P3_U2814) );
  NAND3_X1 U20826 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17749), .A3(
        n18021), .ZN(n17701) );
  NAND2_X1 U20827 ( .A1(n18011), .A2(n17701), .ZN(n18015) );
  INV_X1 U20828 ( .A(n18015), .ZN(n17695) );
  NOR2_X1 U20829 ( .A1(n17680), .A2(n17679), .ZN(n17686) );
  NAND2_X1 U20830 ( .A1(n9724), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18018) );
  OAI21_X1 U20831 ( .B1(n17682), .B2(n17681), .A(n18018), .ZN(n17683) );
  AOI221_X1 U20832 ( .B1(n17686), .B2(n17685), .C1(n17684), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17683), .ZN(n17693) );
  INV_X1 U20833 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18033) );
  INV_X1 U20834 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17731) );
  NAND3_X1 U20835 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18055), .A3(
        n17784), .ZN(n17687) );
  NAND4_X1 U20836 ( .A1(n17754), .A2(n17758), .A3(n18092), .A4(n17739), .ZN(
        n17730) );
  AOI22_X1 U20837 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17687), .B1(
        n17730), .B2(n17719), .ZN(n17688) );
  OAI221_X1 U20838 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18033), 
        .C1(n17731), .C2(n17786), .A(n17688), .ZN(n17689) );
  XNOR2_X1 U20839 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17689), .ZN(
        n18017) );
  NOR2_X1 U20840 ( .A1(n18010), .A2(n17877), .ZN(n17691) );
  NAND2_X1 U20841 ( .A1(n18012), .A2(n18011), .ZN(n17690) );
  AOI22_X1 U20842 ( .A1(n17787), .A2(n18017), .B1(n17691), .B2(n17690), .ZN(
        n17692) );
  OAI211_X1 U20843 ( .C1(n17695), .C2(n17694), .A(n17693), .B(n17692), .ZN(
        P3_U2815) );
  OAI21_X1 U20844 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17696), .A(
        n18012), .ZN(n18027) );
  NAND3_X1 U20845 ( .A1(n17803), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18577), .ZN(n17740) );
  NOR2_X1 U20846 ( .A1(n17697), .A2(n17740), .ZN(n17744) );
  AOI21_X1 U20847 ( .B1(n17708), .B2(n17744), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17699) );
  OAI22_X1 U20848 ( .A1(n17700), .A2(n17699), .B1(n17857), .B2(n17698), .ZN(
        n17705) );
  NOR2_X1 U20849 ( .A1(n18062), .A2(n18022), .ZN(n17702) );
  OAI21_X1 U20850 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17702), .A(
        n17701), .ZN(n18026) );
  OAI22_X1 U20851 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17730), .B1(
        n17766), .B2(n18043), .ZN(n17718) );
  OAI221_X1 U20852 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17731), 
        .C1(n17719), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17718), .ZN(
        n17703) );
  XNOR2_X1 U20853 ( .A(n18033), .B(n17703), .ZN(n18028) );
  OAI22_X1 U20854 ( .A1(n17748), .A2(n18026), .B1(n17756), .B2(n18028), .ZN(
        n17704) );
  AOI211_X1 U20855 ( .C1(n9724), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17705), .B(
        n17704), .ZN(n17706) );
  OAI21_X1 U20856 ( .B1(n17877), .B2(n18027), .A(n17706), .ZN(P3_U2816) );
  INV_X1 U20857 ( .A(n17722), .ZN(n17777) );
  OR2_X1 U20858 ( .A1(n18043), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18049) );
  NAND2_X1 U20859 ( .A1(n17709), .A2(n17707), .ZN(n17725) );
  AOI211_X1 U20860 ( .C1(n17713), .C2(n17724), .A(n17708), .B(n17725), .ZN(
        n17715) );
  OAI21_X1 U20861 ( .B1(n17709), .B2(n17846), .A(n17872), .ZN(n17710) );
  AOI21_X1 U20862 ( .B1(n17712), .B2(n17711), .A(n17710), .ZN(n17723) );
  NAND2_X1 U20863 ( .A1(n9724), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18047) );
  OAI21_X1 U20864 ( .B1(n17723), .B2(n17713), .A(n18047), .ZN(n17714) );
  AOI211_X1 U20865 ( .C1(n17729), .C2(n17716), .A(n17715), .B(n17714), .ZN(
        n17721) );
  NOR2_X1 U20866 ( .A1(n18043), .A2(n18062), .ZN(n18040) );
  OAI22_X1 U20867 ( .A1(n17717), .A2(n17877), .B1(n18040), .B2(n17748), .ZN(
        n17733) );
  XNOR2_X1 U20868 ( .A(n17719), .B(n17718), .ZN(n18045) );
  AOI22_X1 U20869 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17733), .B1(
        n17787), .B2(n18045), .ZN(n17720) );
  OAI211_X1 U20870 ( .C1(n17777), .C2(n18049), .A(n17721), .B(n17720), .ZN(
        P3_U2817) );
  AND3_X1 U20871 ( .A1(n17731), .A2(n17722), .A3(n18055), .ZN(n17727) );
  NAND2_X1 U20872 ( .A1(n9724), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18057) );
  OAI221_X1 U20873 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17725), .C1(
        n17724), .C2(n17723), .A(n18057), .ZN(n17726) );
  AOI211_X1 U20874 ( .C1(n17729), .C2(n17728), .A(n17727), .B(n17726), .ZN(
        n17735) );
  OR2_X1 U20875 ( .A1(n18067), .A2(n17766), .ZN(n17736) );
  OAI21_X1 U20876 ( .B1(n17739), .B2(n17736), .A(n17730), .ZN(n17732) );
  XNOR2_X1 U20877 ( .A(n17732), .B(n17731), .ZN(n18056) );
  AOI22_X1 U20878 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17733), .B1(
        n17787), .B2(n18056), .ZN(n17734) );
  NAND2_X1 U20879 ( .A1(n17735), .A2(n17734), .ZN(P3_U2818) );
  NAND2_X1 U20880 ( .A1(n18068), .A2(n17739), .ZN(n18073) );
  NAND3_X1 U20881 ( .A1(n17754), .A2(n17758), .A3(n18092), .ZN(n17737) );
  NAND2_X1 U20882 ( .A1(n17737), .A2(n17736), .ZN(n17738) );
  XNOR2_X1 U20883 ( .A(n17739), .B(n17738), .ZN(n18061) );
  NOR2_X1 U20884 ( .A1(n18162), .A2(n18751), .ZN(n17746) );
  INV_X1 U20885 ( .A(n17740), .ZN(n17795) );
  NAND2_X1 U20886 ( .A1(n17781), .A2(n17795), .ZN(n17752) );
  NOR2_X1 U20887 ( .A1(n17741), .A2(n17752), .ZN(n17764) );
  AOI21_X1 U20888 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17868), .A(
        n17764), .ZN(n17743) );
  OAI22_X1 U20889 ( .A1(n17744), .A2(n17743), .B1(n17857), .B2(n17742), .ZN(
        n17745) );
  AOI211_X1 U20890 ( .C1(n17787), .C2(n18061), .A(n17746), .B(n17745), .ZN(
        n17751) );
  NOR2_X1 U20891 ( .A1(n18068), .A2(n17777), .ZN(n17753) );
  OAI22_X1 U20892 ( .A1(n17749), .A2(n17748), .B1(n17877), .B2(n17747), .ZN(
        n17765) );
  OAI21_X1 U20893 ( .B1(n17753), .B2(n17765), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17750) );
  OAI211_X1 U20894 ( .C1(n17777), .C2(n18073), .A(n17751), .B(n17750), .ZN(
        P3_U2819) );
  INV_X1 U20895 ( .A(n17752), .ZN(n17769) );
  AND2_X1 U20896 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17769), .ZN(
        n17772) );
  AOI21_X1 U20897 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17868), .A(
        n17772), .ZN(n17763) );
  INV_X1 U20898 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18749) );
  NOR2_X1 U20899 ( .A1(n18162), .A2(n18749), .ZN(n17760) );
  AOI21_X1 U20900 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17765), .A(
        n17753), .ZN(n17757) );
  NAND2_X1 U20901 ( .A1(n17754), .A2(n18092), .ZN(n17767) );
  AOI22_X1 U20902 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17766), .B1(
        n17767), .B2(n18086), .ZN(n17755) );
  XNOR2_X1 U20903 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17755), .ZN(
        n18081) );
  OAI22_X1 U20904 ( .A1(n17758), .A2(n17757), .B1(n18081), .B2(n17756), .ZN(
        n17759) );
  AOI211_X1 U20905 ( .C1(n17761), .C2(n17619), .A(n17760), .B(n17759), .ZN(
        n17762) );
  OAI21_X1 U20906 ( .B1(n17764), .B2(n17763), .A(n17762), .ZN(P3_U2820) );
  INV_X1 U20907 ( .A(n17765), .ZN(n17776) );
  NAND2_X1 U20908 ( .A1(n17767), .A2(n17766), .ZN(n17768) );
  XNOR2_X1 U20909 ( .A(n17768), .B(n18086), .ZN(n18083) );
  NOR2_X1 U20910 ( .A1(n18162), .A2(n18747), .ZN(n17774) );
  AOI21_X1 U20911 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17868), .A(
        n17769), .ZN(n17771) );
  OAI22_X1 U20912 ( .A1(n17772), .A2(n17771), .B1(n17857), .B2(n17770), .ZN(
        n17773) );
  AOI211_X1 U20913 ( .C1(n17787), .C2(n18083), .A(n17774), .B(n17773), .ZN(
        n17775) );
  OAI221_X1 U20914 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17777), .C1(
        n18086), .C2(n17776), .A(n17775), .ZN(P3_U2821) );
  OAI21_X1 U20915 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17779), .A(
        n17778), .ZN(n18104) );
  OAI21_X1 U20916 ( .B1(n9814), .B2(n17846), .A(n17872), .ZN(n17793) );
  INV_X1 U20917 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18745) );
  NOR2_X1 U20918 ( .A1(n18162), .A2(n18745), .ZN(n18094) );
  OAI211_X1 U20919 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n9814), .B(n18577), .ZN(n17780)
         );
  OAI22_X1 U20920 ( .A1(n17857), .A2(n17782), .B1(n17781), .B2(n17780), .ZN(
        n17783) );
  AOI211_X1 U20921 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17793), .A(
        n18094), .B(n17783), .ZN(n17790) );
  NOR2_X1 U20922 ( .A1(n17785), .A2(n17784), .ZN(n18100) );
  XNOR2_X1 U20923 ( .A(n17786), .B(n18100), .ZN(n18095) );
  AOI22_X1 U20924 ( .A1(n17788), .A2(n18100), .B1(n17787), .B2(n18095), .ZN(
        n17789) );
  OAI211_X1 U20925 ( .C1(n17877), .C2(n18104), .A(n17790), .B(n17789), .ZN(
        P3_U2822) );
  OAI21_X1 U20926 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17792), .A(
        n17791), .ZN(n18113) );
  NOR2_X1 U20927 ( .A1(n18162), .A2(n18743), .ZN(n18105) );
  AOI221_X1 U20928 ( .B1(n17795), .B2(n17794), .C1(n17793), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18105), .ZN(n17802) );
  AOI21_X1 U20929 ( .B1(n17798), .B2(n17797), .A(n17796), .ZN(n17799) );
  XNOR2_X1 U20930 ( .A(n17799), .B(n18107), .ZN(n18106) );
  AOI22_X1 U20931 ( .A1(n17824), .A2(n18106), .B1(n17800), .B2(n17619), .ZN(
        n17801) );
  OAI211_X1 U20932 ( .C1(n17876), .C2(n18113), .A(n17802), .B(n17801), .ZN(
        P3_U2823) );
  NAND2_X1 U20933 ( .A1(n17803), .A2(n18577), .ZN(n17807) );
  NAND2_X1 U20934 ( .A1(n17868), .A2(n17807), .ZN(n17827) );
  OAI21_X1 U20935 ( .B1(n17806), .B2(n17805), .A(n17804), .ZN(n18116) );
  OAI22_X1 U20936 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17807), .B1(
        n17876), .B2(n18116), .ZN(n17812) );
  OAI21_X1 U20937 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17809), .A(
        n17808), .ZN(n18117) );
  OAI22_X1 U20938 ( .A1(n17857), .A2(n17810), .B1(n17877), .B2(n18117), .ZN(
        n17811) );
  AOI211_X1 U20939 ( .C1(n9724), .C2(P3_REIP_REG_6__SCAN_IN), .A(n17812), .B(
        n17811), .ZN(n17813) );
  OAI21_X1 U20940 ( .B1(n9874), .B2(n17827), .A(n17813), .ZN(P3_U2824) );
  AOI21_X1 U20941 ( .B1(n17814), .B2(n17872), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17828) );
  NAND2_X1 U20942 ( .A1(n17816), .A2(n17815), .ZN(n17817) );
  XOR2_X1 U20943 ( .A(n17817), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18132) );
  OAI22_X1 U20944 ( .A1(n17876), .A2(n18132), .B1(n13328), .B2(n18739), .ZN(
        n17818) );
  INV_X1 U20945 ( .A(n17818), .ZN(n17826) );
  AOI21_X1 U20946 ( .B1(n17821), .B2(n17820), .A(n17819), .ZN(n17822) );
  XNOR2_X1 U20947 ( .A(n17822), .B(n18129), .ZN(n18125) );
  AOI22_X1 U20948 ( .A1(n17824), .A2(n18125), .B1(n17823), .B2(n17619), .ZN(
        n17825) );
  OAI211_X1 U20949 ( .C1(n17828), .C2(n17827), .A(n17826), .B(n17825), .ZN(
        P3_U2825) );
  OAI21_X1 U20950 ( .B1(n17831), .B2(n17830), .A(n17829), .ZN(n18136) );
  AOI22_X1 U20951 ( .A1(n9724), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18577), .B2(
        n17832), .ZN(n17840) );
  OAI21_X1 U20952 ( .B1(n17833), .B2(n17846), .A(n17872), .ZN(n17845) );
  OAI21_X1 U20953 ( .B1(n17836), .B2(n17835), .A(n17834), .ZN(n18142) );
  OAI22_X1 U20954 ( .A1(n17857), .A2(n17837), .B1(n17877), .B2(n18142), .ZN(
        n17838) );
  AOI21_X1 U20955 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17845), .A(
        n17838), .ZN(n17839) );
  OAI211_X1 U20956 ( .C1(n17876), .C2(n18136), .A(n17840), .B(n17839), .ZN(
        P3_U2826) );
  OAI22_X1 U20957 ( .A1(n17877), .A2(n17842), .B1(n17876), .B2(n17841), .ZN(
        n17843) );
  AOI211_X1 U20958 ( .C1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n17845), .A(
        n17844), .B(n17843), .ZN(n17848) );
  OR4_X1 U20959 ( .A1(n17859), .A2(n17846), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(n17860), .ZN(n17847) );
  OAI211_X1 U20960 ( .C1(n17857), .C2(n17849), .A(n17848), .B(n17847), .ZN(
        P3_U2827) );
  OAI21_X1 U20961 ( .B1(n17852), .B2(n17851), .A(n17850), .ZN(n18158) );
  OAI21_X1 U20962 ( .B1(n17855), .B2(n17854), .A(n17853), .ZN(n18154) );
  OAI22_X1 U20963 ( .A1(n17857), .A2(n17856), .B1(n17877), .B2(n18154), .ZN(
        n17858) );
  AOI221_X1 U20964 ( .B1(n17860), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18577), .C2(n17859), .A(n17858), .ZN(n17861) );
  NAND2_X1 U20965 ( .A1(n9724), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18156) );
  OAI211_X1 U20966 ( .C1(n17876), .C2(n18158), .A(n17861), .B(n18156), .ZN(
        P3_U2828) );
  NOR2_X1 U20967 ( .A1(n17862), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17863) );
  XNOR2_X1 U20968 ( .A(n17863), .B(n17865), .ZN(n18168) );
  OAI21_X1 U20969 ( .B1(n17865), .B2(n17870), .A(n17864), .ZN(n18161) );
  OAI22_X1 U20970 ( .A1(n17876), .A2(n18161), .B1(n13328), .B2(n18839), .ZN(
        n17866) );
  AOI221_X1 U20971 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17868), .C1(
        n17867), .C2(n17619), .A(n17866), .ZN(n17869) );
  OAI21_X1 U20972 ( .B1(n18168), .B2(n17877), .A(n17869), .ZN(P3_U2829) );
  AOI21_X1 U20973 ( .B1(n17871), .B2(n18828), .A(n17870), .ZN(n18176) );
  INV_X1 U20974 ( .A(n18176), .ZN(n18174) );
  OAI21_X1 U20975 ( .B1(n17873), .B2(n18853), .A(n17872), .ZN(n17874) );
  AOI22_X1 U20976 ( .A1(n9724), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17874), .ZN(n17875) );
  OAI221_X1 U20977 ( .B1(n18176), .B2(n17877), .C1(n18174), .C2(n17876), .A(
        n17875), .ZN(P3_U2830) );
  AOI22_X1 U20978 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18164), .B1(
        n9724), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n17888) );
  AOI21_X1 U20979 ( .B1(n17878), .B2(n17974), .A(n18145), .ZN(n17898) );
  OAI22_X1 U20980 ( .A1(n18668), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18651), .B2(n17879), .ZN(n17883) );
  OAI22_X1 U20981 ( .A1(n17881), .A2(n18153), .B1(n17880), .B2(n18039), .ZN(
        n17882) );
  NOR4_X1 U20982 ( .A1(n17884), .A2(n17898), .A3(n17883), .A4(n17882), .ZN(
        n17892) );
  OAI211_X1 U20983 ( .C1(n18668), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17892), .ZN(n17885) );
  OAI211_X1 U20984 ( .C1(n17886), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18169), .B(n17885), .ZN(n17887) );
  OAI211_X1 U20985 ( .C1(n17889), .C2(n18080), .A(n17888), .B(n17887), .ZN(
        P3_U2835) );
  NAND2_X1 U20986 ( .A1(n17912), .A2(n17924), .ZN(n17910) );
  OAI22_X1 U20987 ( .A1(n17892), .A2(n17891), .B1(n17910), .B2(n17890), .ZN(
        n17893) );
  AOI22_X1 U20988 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18164), .B1(
        n18169), .B2(n17893), .ZN(n17895) );
  OAI211_X1 U20989 ( .C1(n17896), .C2(n18080), .A(n17895), .B(n17894), .ZN(
        P3_U2836) );
  INV_X1 U20990 ( .A(n17897), .ZN(n17899) );
  AOI21_X1 U20991 ( .B1(n18664), .B2(n17899), .A(n17898), .ZN(n17903) );
  AOI22_X1 U20992 ( .A1(n18633), .A2(n17901), .B1(n18099), .B2(n17900), .ZN(
        n17902) );
  OAI221_X1 U20993 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17905), 
        .C1(n17904), .C2(n17903), .A(n17902), .ZN(n17906) );
  AOI22_X1 U20994 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18164), .B1(
        n18169), .B2(n17906), .ZN(n17908) );
  OAI211_X1 U20995 ( .C1(n17909), .C2(n18080), .A(n17908), .B(n17907), .ZN(
        P3_U2837) );
  NOR3_X1 U20996 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18159), .A3(
        n17910), .ZN(n17911) );
  AOI21_X1 U20997 ( .B1(n9724), .B2(P3_REIP_REG_24__SCAN_IN), .A(n17911), .ZN(
        n17922) );
  AOI21_X1 U20998 ( .B1(n18010), .B2(n17912), .A(n18153), .ZN(n17913) );
  AOI211_X1 U20999 ( .C1(n17984), .C2(n17914), .A(n17913), .B(n18149), .ZN(
        n17915) );
  OAI211_X1 U21000 ( .C1(n17916), .C2(n18039), .A(n17915), .B(n18133), .ZN(
        n17920) );
  INV_X1 U21001 ( .A(n17920), .ZN(n17919) );
  AOI221_X1 U21002 ( .B1(n17925), .B2(n18664), .C1(n17932), .C2(n18664), .A(
        n17917), .ZN(n17918) );
  AOI21_X1 U21003 ( .B1(n17919), .B2(n17918), .A(n9724), .ZN(n17926) );
  OAI211_X1 U21004 ( .C1(n18091), .C2(n17920), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17926), .ZN(n17921) );
  OAI211_X1 U21005 ( .C1(n17923), .C2(n18080), .A(n17922), .B(n17921), .ZN(
        P3_U2838) );
  INV_X1 U21006 ( .A(n17924), .ZN(n17931) );
  NOR3_X1 U21007 ( .A1(n18164), .A2(n17931), .A3(n17925), .ZN(n17927) );
  OAI21_X1 U21008 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17927), .A(
        n17926), .ZN(n17929) );
  OAI211_X1 U21009 ( .C1(n18080), .C2(n17930), .A(n17929), .B(n17928), .ZN(
        P3_U2839) );
  AOI221_X1 U21010 ( .B1(n17931), .B2(n17948), .C1(n17940), .C2(n17948), .A(
        n18159), .ZN(n17944) );
  NAND2_X1 U21011 ( .A1(n18153), .A2(n18039), .ZN(n18066) );
  NOR2_X1 U21012 ( .A1(n18668), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17935) );
  OAI21_X1 U21013 ( .B1(n17932), .B2(n17954), .A(n18664), .ZN(n17933) );
  OAI221_X1 U21014 ( .B1(n18668), .B2(n17975), .C1(n18668), .C2(n17934), .A(
        n17933), .ZN(n17961) );
  AOI211_X1 U21015 ( .C1(n18066), .C2(n17940), .A(n17935), .B(n17961), .ZN(
        n17951) );
  AOI22_X1 U21016 ( .A1(n18664), .A2(n17937), .B1(n17936), .B2(n18041), .ZN(
        n17942) );
  NAND2_X1 U21017 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17998), .ZN(
        n18042) );
  NOR2_X1 U21018 ( .A1(n17938), .A2(n18042), .ZN(n17996) );
  INV_X1 U21019 ( .A(n17996), .ZN(n17949) );
  NAND2_X1 U21020 ( .A1(n18099), .A2(n17939), .ZN(n18006) );
  OAI21_X1 U21021 ( .B1(n18010), .B2(n18153), .A(n18006), .ZN(n17977) );
  AOI221_X1 U21022 ( .B1(n17949), .B2(n18666), .C1(n17940), .C2(n18666), .A(
        n17977), .ZN(n17941) );
  NAND4_X1 U21023 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17951), .A3(
        n17942), .A4(n17941), .ZN(n17943) );
  AOI22_X1 U21024 ( .A1(n18096), .A2(n17945), .B1(n17944), .B2(n17943), .ZN(
        n17947) );
  OAI211_X1 U21025 ( .C1(n18133), .C2(n17948), .A(n17947), .B(n17946), .ZN(
        P3_U2840) );
  NOR2_X1 U21026 ( .A1(n18159), .A2(n17977), .ZN(n18000) );
  OAI21_X1 U21027 ( .B1(n17954), .B2(n17949), .A(n18666), .ZN(n17950) );
  NAND2_X1 U21028 ( .A1(n18000), .A2(n17950), .ZN(n17960) );
  NOR2_X1 U21029 ( .A1(n18664), .A2(n18666), .ZN(n18160) );
  OAI21_X1 U21030 ( .B1(n17952), .B2(n18160), .A(n17951), .ZN(n17953) );
  OAI21_X1 U21031 ( .B1(n17960), .B2(n17953), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17958) );
  NOR2_X1 U21032 ( .A1(n17985), .A2(n17954), .ZN(n17969) );
  AOI22_X1 U21033 ( .A1(n18096), .A2(n17956), .B1(n17969), .B2(n17955), .ZN(
        n17957) );
  OAI221_X1 U21034 ( .B1(n9724), .B2(n17958), .C1(n13328), .C2(n18771), .A(
        n17957), .ZN(P3_U2841) );
  AOI22_X1 U21035 ( .A1(n9724), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17969), 
        .B2(n17959), .ZN(n17966) );
  AOI211_X1 U21036 ( .C1(n17962), .C2(n18066), .A(n17961), .B(n17960), .ZN(
        n17963) );
  NOR2_X1 U21037 ( .A1(n9724), .A2(n17963), .ZN(n17970) );
  NOR3_X1 U21038 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18160), .A3(
        n18862), .ZN(n17964) );
  OAI21_X1 U21039 ( .B1(n17970), .B2(n17964), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17965) );
  OAI211_X1 U21040 ( .C1(n17967), .C2(n18080), .A(n17966), .B(n17965), .ZN(
        P3_U2842) );
  AOI22_X1 U21041 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17970), .B1(
        n17969), .B2(n17968), .ZN(n17972) );
  OAI211_X1 U21042 ( .C1(n17973), .C2(n18080), .A(n17972), .B(n17971), .ZN(
        P3_U2843) );
  INV_X1 U21043 ( .A(n18066), .ZN(n17981) );
  NAND3_X1 U21044 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17975), .A3(
        n17974), .ZN(n17979) );
  AOI21_X1 U21045 ( .B1(n17982), .B2(n17976), .A(n18144), .ZN(n17978) );
  AOI211_X1 U21046 ( .C1(n17984), .C2(n17979), .A(n17978), .B(n17977), .ZN(
        n17980) );
  OAI211_X1 U21047 ( .C1(n17982), .C2(n17981), .A(n17980), .B(n18133), .ZN(
        n17992) );
  OAI221_X1 U21048 ( .B1(n17992), .B2(n17984), .C1(n17992), .C2(n17983), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17989) );
  INV_X1 U21049 ( .A(n17985), .ZN(n18001) );
  AOI22_X1 U21050 ( .A1(n18096), .A2(n17987), .B1(n18001), .B2(n17986), .ZN(
        n17988) );
  OAI221_X1 U21051 ( .B1(n9724), .B2(n17989), .C1(n13328), .C2(n18764), .A(
        n17988), .ZN(P3_U2844) );
  NOR2_X1 U21052 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n15584), .ZN(
        n17990) );
  AOI22_X1 U21053 ( .A1(n18096), .A2(n17991), .B1(n18001), .B2(n17990), .ZN(
        n17995) );
  NAND3_X1 U21054 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18162), .A3(
        n17992), .ZN(n17993) );
  NAND3_X1 U21055 ( .A1(n17995), .A2(n17994), .A3(n17993), .ZN(P3_U2845) );
  AOI21_X1 U21056 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18651), .A(
        n17996), .ZN(n17999) );
  OAI22_X1 U21057 ( .A1(n18668), .A2(n17998), .B1(n17997), .B2(n18144), .ZN(
        n18036) );
  AOI211_X1 U21058 ( .C1(n18009), .C2(n18041), .A(n17999), .B(n18036), .ZN(
        n18008) );
  AOI221_X1 U21059 ( .B1(n18076), .B2(n18000), .C1(n18008), .C2(n18000), .A(
        n9724), .ZN(n18002) );
  AOI22_X1 U21060 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18002), .B1(
        n18001), .B2(n15584), .ZN(n18004) );
  OAI211_X1 U21061 ( .C1(n18005), .C2(n18080), .A(n18004), .B(n18003), .ZN(
        P3_U2846) );
  INV_X1 U21062 ( .A(n18006), .ZN(n18016) );
  NOR2_X1 U21063 ( .A1(n18128), .A2(n18115), .ZN(n18110) );
  NAND2_X1 U21064 ( .A1(n18007), .A2(n18110), .ZN(n18034) );
  AOI221_X1 U21065 ( .B1(n18009), .B2(n18011), .C1(n18034), .C2(n18011), .A(
        n18008), .ZN(n18014) );
  AOI211_X1 U21066 ( .C1(n18012), .C2(n18011), .A(n18010), .B(n18153), .ZN(
        n18013) );
  AOI211_X1 U21067 ( .C1(n18016), .C2(n18015), .A(n18014), .B(n18013), .ZN(
        n18020) );
  AOI22_X1 U21068 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18164), .B1(
        n18096), .B2(n18017), .ZN(n18019) );
  OAI211_X1 U21069 ( .C1(n18020), .C2(n18159), .A(n18019), .B(n18018), .ZN(
        P3_U2847) );
  AOI21_X1 U21070 ( .B1(n18666), .B2(n18042), .A(n18036), .ZN(n18065) );
  OAI21_X1 U21071 ( .B1(n18076), .B2(n18021), .A(n18065), .ZN(n18024) );
  OAI21_X1 U21072 ( .B1(n18022), .B2(n18034), .A(n18033), .ZN(n18023) );
  OAI21_X1 U21073 ( .B1(n18033), .B2(n18024), .A(n18023), .ZN(n18025) );
  OAI21_X1 U21074 ( .B1(n18039), .B2(n18026), .A(n18025), .ZN(n18030) );
  OAI22_X1 U21075 ( .A1(n18080), .A2(n18028), .B1(n18175), .B2(n18027), .ZN(
        n18029) );
  AOI21_X1 U21076 ( .B1(n18169), .B2(n18030), .A(n18029), .ZN(n18032) );
  NAND2_X1 U21077 ( .A1(n9724), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n18031) );
  OAI211_X1 U21078 ( .C1(n18133), .C2(n18033), .A(n18032), .B(n18031), .ZN(
        P3_U2848) );
  NAND2_X1 U21079 ( .A1(n18035), .A2(n18034), .ZN(n18054) );
  NAND2_X1 U21080 ( .A1(n18169), .A2(n18054), .ZN(n18087) );
  OAI21_X1 U21081 ( .B1(n18668), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18051) );
  OAI22_X1 U21082 ( .A1(n18668), .A2(n18068), .B1(n18055), .B2(n18144), .ZN(
        n18070) );
  AOI211_X1 U21083 ( .C1(n18633), .C2(n18037), .A(n18036), .B(n18070), .ZN(
        n18038) );
  OAI21_X1 U21084 ( .B1(n18040), .B2(n18039), .A(n18038), .ZN(n18052) );
  AOI211_X1 U21085 ( .C1(n18041), .C2(n18051), .A(n18159), .B(n18052), .ZN(
        n18044) );
  NOR2_X1 U21086 ( .A1(n18043), .A2(n18042), .ZN(n18050) );
  AOI221_X1 U21087 ( .B1(n18651), .B2(n18044), .C1(n18050), .C2(n18044), .A(
        n9724), .ZN(n18046) );
  AOI22_X1 U21088 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18046), .B1(
        n18096), .B2(n18045), .ZN(n18048) );
  OAI211_X1 U21089 ( .C1(n18087), .C2(n18049), .A(n18048), .B(n18047), .ZN(
        P3_U2849) );
  INV_X1 U21090 ( .A(n18050), .ZN(n18053) );
  AOI211_X1 U21091 ( .C1(n18053), .C2(n18666), .A(n18052), .B(n18051), .ZN(
        n18060) );
  OAI221_X1 U21092 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18055), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18054), .A(n18169), .ZN(
        n18059) );
  AOI22_X1 U21093 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18164), .B1(
        n18096), .B2(n18056), .ZN(n18058) );
  OAI211_X1 U21094 ( .C1(n18060), .C2(n18059), .A(n18058), .B(n18057), .ZN(
        P3_U2850) );
  AOI22_X1 U21095 ( .A1(n9724), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18096), 
        .B2(n18061), .ZN(n18072) );
  AOI22_X1 U21096 ( .A1(n18633), .A2(n18063), .B1(n18099), .B2(n18062), .ZN(
        n18064) );
  NAND3_X1 U21097 ( .A1(n18169), .A2(n18065), .A3(n18064), .ZN(n18082) );
  AOI21_X1 U21098 ( .B1(n18067), .B2(n18066), .A(n18082), .ZN(n18075) );
  OAI21_X1 U21099 ( .B1(n18651), .B2(n18068), .A(n18075), .ZN(n18069) );
  OAI211_X1 U21100 ( .C1(n18070), .C2(n18069), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n13328), .ZN(n18071) );
  OAI211_X1 U21101 ( .C1(n18073), .C2(n18087), .A(n18072), .B(n18071), .ZN(
        P3_U2851) );
  AOI221_X1 U21102 ( .B1(n18076), .B2(n18075), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18075), .A(n18074), .ZN(
        n18078) );
  NOR3_X1 U21103 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18086), .A3(
        n18087), .ZN(n18077) );
  AOI221_X1 U21104 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n9724), .C1(n18078), 
        .C2(n18162), .A(n18077), .ZN(n18079) );
  OAI21_X1 U21105 ( .B1(n18081), .B2(n18080), .A(n18079), .ZN(P3_U2852) );
  NAND2_X1 U21106 ( .A1(n13328), .A2(n18082), .ZN(n18085) );
  AOI22_X1 U21107 ( .A1(n9724), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18096), .B2(
        n18083), .ZN(n18084) );
  OAI221_X1 U21108 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18087), .C1(
        n18086), .C2(n18085), .A(n18084), .ZN(P3_U2853) );
  OAI22_X1 U21109 ( .A1(n18145), .A2(n18089), .B1(n18088), .B2(n18144), .ZN(
        n18090) );
  OR2_X1 U21110 ( .A1(n18149), .A2(n18090), .ZN(n18114) );
  AOI21_X1 U21111 ( .B1(n18091), .B2(n18098), .A(n18114), .ZN(n18108) );
  AOI221_X1 U21112 ( .B1(n18108), .B2(n18133), .C1(n18134), .C2(n18133), .A(
        n18092), .ZN(n18093) );
  AOI211_X1 U21113 ( .C1(n18096), .C2(n18095), .A(n18094), .B(n18093), .ZN(
        n18103) );
  INV_X1 U21114 ( .A(n18110), .ZN(n18097) );
  NOR3_X1 U21115 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18098), .A3(
        n18097), .ZN(n18101) );
  OAI221_X1 U21116 ( .B1(n18101), .B2(n18100), .C1(n18101), .C2(n18099), .A(
        n18169), .ZN(n18102) );
  OAI211_X1 U21117 ( .C1(n18104), .C2(n18175), .A(n18103), .B(n18102), .ZN(
        P3_U2854) );
  AOI21_X1 U21118 ( .B1(n18106), .B2(n18126), .A(n18105), .ZN(n18112) );
  OAI22_X1 U21119 ( .A1(n18108), .A2(n18159), .B1(n18107), .B2(n18133), .ZN(
        n18109) );
  OAI221_X1 U21120 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18110), .A(n18109), .ZN(
        n18111) );
  OAI211_X1 U21121 ( .C1(n18113), .C2(n18173), .A(n18112), .B(n18111), .ZN(
        P3_U2855) );
  AOI21_X1 U21122 ( .B1(n18169), .B2(n18114), .A(n18164), .ZN(n18123) );
  NOR4_X1 U21123 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18128), .A3(
        n18159), .A4(n18115), .ZN(n18119) );
  OAI22_X1 U21124 ( .A1(n18175), .A2(n18117), .B1(n18173), .B2(n18116), .ZN(
        n18118) );
  NOR2_X1 U21125 ( .A1(n18119), .A2(n18118), .ZN(n18121) );
  NAND2_X1 U21126 ( .A1(n9724), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18120) );
  OAI211_X1 U21127 ( .C1(n18123), .C2(n18122), .A(n18121), .B(n18120), .ZN(
        P3_U2856) );
  OAI22_X1 U21128 ( .A1(n18123), .A2(n18129), .B1(n13328), .B2(n18739), .ZN(
        n18124) );
  AOI21_X1 U21129 ( .B1(n18126), .B2(n18125), .A(n18124), .ZN(n18131) );
  NOR3_X1 U21130 ( .A1(n18128), .A2(n18159), .A3(n18127), .ZN(n18140) );
  NAND3_X1 U21131 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18140), .A3(
        n18129), .ZN(n18130) );
  OAI211_X1 U21132 ( .C1(n18132), .C2(n18173), .A(n18131), .B(n18130), .ZN(
        P3_U2857) );
  OAI21_X1 U21133 ( .B1(n18135), .B2(n18134), .A(n18133), .ZN(n18138) );
  OAI22_X1 U21134 ( .A1(n18162), .A2(n18737), .B1(n18173), .B2(n18136), .ZN(
        n18137) );
  AOI221_X1 U21135 ( .B1(n18140), .B2(n18139), .C1(n18138), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18137), .ZN(n18141) );
  OAI21_X1 U21136 ( .B1(n18175), .B2(n18142), .A(n18141), .ZN(P3_U2858) );
  NAND2_X1 U21137 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18143) );
  OAI22_X1 U21138 ( .A1(n18145), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n18144), .B2(n18143), .ZN(n18148) );
  INV_X1 U21139 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18809) );
  NOR3_X1 U21140 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18809), .A3(
        n18146), .ZN(n18147) );
  AOI221_X1 U21141 ( .B1(n18149), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18148), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n18147), .ZN(
        n18152) );
  NAND2_X1 U21142 ( .A1(n18664), .A2(n18150), .ZN(n18151) );
  OAI211_X1 U21143 ( .C1(n18154), .C2(n18153), .A(n18152), .B(n18151), .ZN(
        n18155) );
  AOI22_X1 U21144 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18164), .B1(
        n18169), .B2(n18155), .ZN(n18157) );
  OAI211_X1 U21145 ( .C1(n18173), .C2(n18158), .A(n18157), .B(n18156), .ZN(
        P3_U2860) );
  NOR3_X1 U21146 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18160), .A3(
        n18159), .ZN(n18170) );
  OAI22_X1 U21147 ( .A1(n18162), .A2(n18839), .B1(n18173), .B2(n18161), .ZN(
        n18163) );
  AOI221_X1 U21148 ( .B1(n18164), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18170), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n18163), .ZN(
        n18167) );
  OAI211_X1 U21149 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18658), .A(
        n18165), .B(n18809), .ZN(n18166) );
  OAI211_X1 U21150 ( .C1(n18168), .C2(n18175), .A(n18167), .B(n18166), .ZN(
        P3_U2861) );
  AOI21_X1 U21151 ( .B1(n18668), .B2(n18169), .A(n18828), .ZN(n18171) );
  AOI221_X1 U21152 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n9724), .C1(n18171), 
        .C2(n13328), .A(n18170), .ZN(n18172) );
  OAI221_X1 U21153 ( .B1(n18176), .B2(n18175), .C1(n18174), .C2(n18173), .A(
        n18172), .ZN(P3_U2862) );
  INV_X1 U21154 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18483) );
  INV_X1 U21155 ( .A(n18177), .ZN(n18178) );
  AOI21_X1 U21156 ( .B1(n18180), .B2(n18179), .A(n18178), .ZN(n18692) );
  OAI21_X1 U21157 ( .B1(n18692), .B2(n18230), .A(n18185), .ZN(n18181) );
  OAI221_X1 U21158 ( .B1(n18483), .B2(n18845), .C1(n18483), .C2(n18185), .A(
        n18181), .ZN(P3_U2863) );
  NOR2_X1 U21159 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18677), .ZN(
        n18361) );
  INV_X1 U21160 ( .A(n18361), .ZN(n18363) );
  NAND2_X1 U21161 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18677), .ZN(
        n18457) );
  INV_X1 U21162 ( .A(n18457), .ZN(n18459) );
  NAND2_X1 U21163 ( .A1(n18543), .A2(n18459), .ZN(n18484) );
  AND2_X1 U21164 ( .A1(n18363), .A2(n18484), .ZN(n18183) );
  OAI22_X1 U21165 ( .A1(n18184), .A2(n18680), .B1(n18183), .B2(n18182), .ZN(
        P3_U2866) );
  NOR2_X1 U21166 ( .A1(n18681), .A2(n18185), .ZN(P3_U2867) );
  NAND2_X1 U21167 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18187) );
  NOR2_X1 U21168 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18187), .ZN(
        n18576) );
  NAND2_X1 U21169 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18576), .ZN(
        n18526) );
  NAND2_X1 U21170 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18577), .ZN(n18581) );
  AND2_X1 U21171 ( .A1(n18577), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18573) );
  NAND2_X1 U21172 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18483), .ZN(
        n18250) );
  NOR2_X2 U21173 ( .A1(n18187), .A2(n18250), .ZN(n18566) );
  NOR2_X2 U21174 ( .A1(n18231), .A2(n18186), .ZN(n18572) );
  NAND2_X1 U21175 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18671) );
  NOR2_X2 U21176 ( .A1(n18671), .A2(n18187), .ZN(n18625) );
  NAND2_X1 U21177 ( .A1(n18672), .A2(n18483), .ZN(n18673) );
  NAND2_X1 U21178 ( .A1(n18677), .A2(n18680), .ZN(n18316) );
  NOR2_X2 U21179 ( .A1(n18673), .A2(n18316), .ZN(n18279) );
  NOR2_X1 U21180 ( .A1(n18625), .A2(n18279), .ZN(n18188) );
  NOR2_X1 U21181 ( .A1(n9706), .A2(n18188), .ZN(n18224) );
  AOI22_X1 U21182 ( .A1(n18573), .A2(n18566), .B1(n18572), .B2(n18224), .ZN(
        n18193) );
  INV_X1 U21183 ( .A(n18250), .ZN(n18430) );
  NOR2_X1 U21184 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18483), .ZN(
        n18406) );
  NOR2_X1 U21185 ( .A1(n18430), .A2(n18406), .ZN(n18485) );
  NOR2_X1 U21186 ( .A1(n18485), .A2(n18187), .ZN(n18544) );
  AOI21_X1 U21187 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18231), .ZN(n18541) );
  INV_X1 U21188 ( .A(n18188), .ZN(n18251) );
  AOI22_X1 U21189 ( .A1(n18577), .A2(n18544), .B1(n18541), .B2(n18251), .ZN(
        n18227) );
  NAND2_X1 U21190 ( .A1(n18190), .A2(n18189), .ZN(n18225) );
  NOR2_X1 U21191 ( .A1(n18191), .A2(n18225), .ZN(n18578) );
  AOI22_X1 U21192 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18227), .B1(
        n18279), .B2(n18578), .ZN(n18192) );
  OAI211_X1 U21193 ( .C1(n18526), .C2(n18581), .A(n18193), .B(n18192), .ZN(
        P3_U2868) );
  NAND2_X1 U21194 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18577), .ZN(n18495) );
  AND2_X1 U21195 ( .A1(n18577), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18584) );
  AND2_X1 U21196 ( .A1(n18487), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18582) );
  AOI22_X1 U21197 ( .A1(n18566), .A2(n18584), .B1(n18224), .B2(n18582), .ZN(
        n18195) );
  NOR2_X1 U21198 ( .A1(n18850), .A2(n18225), .ZN(n18492) );
  AOI22_X1 U21199 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18227), .B1(
        n18279), .B2(n18492), .ZN(n18194) );
  OAI211_X1 U21200 ( .C1(n18526), .C2(n18495), .A(n18195), .B(n18194), .ZN(
        P3_U2869) );
  NOR2_X1 U21201 ( .A1(n18196), .A2(n18221), .ZN(n18465) );
  INV_X1 U21202 ( .A(n18465), .ZN(n18593) );
  NOR2_X2 U21203 ( .A1(n18221), .A2(n18197), .ZN(n18589) );
  NOR2_X2 U21204 ( .A1(n18231), .A2(n18198), .ZN(n18588) );
  AOI22_X1 U21205 ( .A1(n18566), .A2(n18589), .B1(n18224), .B2(n18588), .ZN(
        n18201) );
  NOR2_X1 U21206 ( .A1(n18199), .A2(n18225), .ZN(n18590) );
  AOI22_X1 U21207 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18227), .B1(
        n18279), .B2(n18590), .ZN(n18200) );
  OAI211_X1 U21208 ( .C1(n18526), .C2(n18593), .A(n18201), .B(n18200), .ZN(
        P3_U2870) );
  NAND2_X1 U21209 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18577), .ZN(n18554) );
  NOR2_X2 U21210 ( .A1(n18202), .A2(n18221), .ZN(n18596) );
  NOR2_X2 U21211 ( .A1(n18203), .A2(n18231), .ZN(n18594) );
  AOI22_X1 U21212 ( .A1(n18566), .A2(n18596), .B1(n18224), .B2(n18594), .ZN(
        n18206) );
  NOR2_X1 U21213 ( .A1(n18204), .A2(n18225), .ZN(n18551) );
  AOI22_X1 U21214 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18227), .B1(
        n18279), .B2(n18551), .ZN(n18205) );
  OAI211_X1 U21215 ( .C1(n18526), .C2(n18554), .A(n18206), .B(n18205), .ZN(
        P3_U2871) );
  NAND2_X1 U21216 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18577), .ZN(n18445) );
  AND2_X1 U21217 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18577), .ZN(n18602) );
  NOR2_X2 U21218 ( .A1(n18207), .A2(n18231), .ZN(n18600) );
  AOI22_X1 U21219 ( .A1(n18566), .A2(n18602), .B1(n18224), .B2(n18600), .ZN(
        n18210) );
  NOR2_X1 U21220 ( .A1(n18208), .A2(n18225), .ZN(n18442) );
  AOI22_X1 U21221 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18227), .B1(
        n18279), .B2(n18442), .ZN(n18209) );
  OAI211_X1 U21222 ( .C1(n18526), .C2(n18445), .A(n18210), .B(n18209), .ZN(
        P3_U2872) );
  NAND2_X1 U21223 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18577), .ZN(n18562) );
  NOR2_X2 U21224 ( .A1(n18211), .A2(n18221), .ZN(n18609) );
  NOR2_X2 U21225 ( .A1(n18212), .A2(n18231), .ZN(n18606) );
  AOI22_X1 U21226 ( .A1(n18566), .A2(n18609), .B1(n18224), .B2(n18606), .ZN(
        n18215) );
  NOR2_X1 U21227 ( .A1(n18213), .A2(n18225), .ZN(n18559) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18227), .B1(
        n18279), .B2(n18559), .ZN(n18214) );
  OAI211_X1 U21229 ( .C1(n18526), .C2(n18562), .A(n18215), .B(n18214), .ZN(
        P3_U2873) );
  INV_X1 U21230 ( .A(n18566), .ZN(n18558) );
  NAND2_X1 U21231 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18577), .ZN(n18533) );
  INV_X1 U21232 ( .A(n18526), .ZN(n18623) );
  NAND2_X1 U21233 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18577), .ZN(n18619) );
  INV_X1 U21234 ( .A(n18619), .ZN(n18530) );
  NOR2_X2 U21235 ( .A1(n18216), .A2(n18231), .ZN(n18614) );
  AOI22_X1 U21236 ( .A1(n18623), .A2(n18530), .B1(n18224), .B2(n18614), .ZN(
        n18219) );
  NOR2_X2 U21237 ( .A1(n18217), .A2(n18225), .ZN(n18616) );
  AOI22_X1 U21238 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18227), .B1(
        n18279), .B2(n18616), .ZN(n18218) );
  OAI211_X1 U21239 ( .C1(n18558), .C2(n18533), .A(n18219), .B(n18218), .ZN(
        P3_U2874) );
  NOR2_X1 U21240 ( .A1(n18220), .A2(n18221), .ZN(n18509) );
  INV_X1 U21241 ( .A(n18509), .ZN(n18630) );
  NOR2_X2 U21242 ( .A1(n18223), .A2(n18231), .ZN(n18621) );
  AOI22_X1 U21243 ( .A1(n18566), .A2(n18622), .B1(n18224), .B2(n18621), .ZN(
        n18229) );
  NOR2_X2 U21244 ( .A1(n18226), .A2(n18225), .ZN(n18624) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18227), .B1(
        n18279), .B2(n18624), .ZN(n18228) );
  OAI211_X1 U21246 ( .C1(n18526), .C2(n18630), .A(n18229), .B(n18228), .ZN(
        P3_U2875) );
  INV_X1 U21247 ( .A(n18578), .ZN(n18491) );
  INV_X1 U21248 ( .A(n18316), .ZN(n18272) );
  NAND2_X1 U21249 ( .A1(n18272), .A2(n18406), .ZN(n18310) );
  INV_X1 U21250 ( .A(n18581), .ZN(n18488) );
  AOI22_X1 U21251 ( .A1(n18488), .A2(n18566), .B1(n18572), .B2(n18246), .ZN(
        n18233) );
  NOR2_X1 U21252 ( .A1(n18680), .A2(n18407), .ZN(n18574) );
  NOR2_X1 U21253 ( .A1(n18231), .A2(n18230), .ZN(n18575) );
  INV_X1 U21254 ( .A(n18575), .ZN(n18271) );
  NOR2_X1 U21255 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18271), .ZN(
        n18317) );
  AOI22_X1 U21256 ( .A1(n18577), .A2(n18574), .B1(n18272), .B2(n18317), .ZN(
        n18247) );
  AOI22_X1 U21257 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18247), .B1(
        n18625), .B2(n18573), .ZN(n18232) );
  OAI211_X1 U21258 ( .C1(n18491), .C2(n18310), .A(n18233), .B(n18232), .ZN(
        P3_U2876) );
  INV_X1 U21259 ( .A(n18492), .ZN(n18587) );
  INV_X1 U21260 ( .A(n18495), .ZN(n18583) );
  AOI22_X1 U21261 ( .A1(n18566), .A2(n18583), .B1(n18582), .B2(n18246), .ZN(
        n18235) );
  AOI22_X1 U21262 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18247), .B1(
        n18625), .B2(n18584), .ZN(n18234) );
  OAI211_X1 U21263 ( .C1(n18587), .C2(n18310), .A(n18235), .B(n18234), .ZN(
        P3_U2877) );
  INV_X1 U21264 ( .A(n18590), .ZN(n18468) );
  AOI22_X1 U21265 ( .A1(n18566), .A2(n18465), .B1(n18588), .B2(n18246), .ZN(
        n18237) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18247), .B1(
        n18625), .B2(n18589), .ZN(n18236) );
  OAI211_X1 U21267 ( .C1(n18468), .C2(n18310), .A(n18237), .B(n18236), .ZN(
        P3_U2878) );
  AOI22_X1 U21268 ( .A1(n18625), .A2(n18596), .B1(n18594), .B2(n18246), .ZN(
        n18239) );
  INV_X1 U21269 ( .A(n18310), .ZN(n18312) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18247), .B1(
        n18551), .B2(n18312), .ZN(n18238) );
  OAI211_X1 U21271 ( .C1(n18558), .C2(n18554), .A(n18239), .B(n18238), .ZN(
        P3_U2879) );
  AOI22_X1 U21272 ( .A1(n18625), .A2(n18602), .B1(n18600), .B2(n18246), .ZN(
        n18241) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18247), .B1(
        n18442), .B2(n18312), .ZN(n18240) );
  OAI211_X1 U21274 ( .C1(n18558), .C2(n18445), .A(n18241), .B(n18240), .ZN(
        P3_U2880) );
  AOI22_X1 U21275 ( .A1(n18625), .A2(n18609), .B1(n18606), .B2(n18246), .ZN(
        n18243) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18247), .B1(
        n18559), .B2(n18312), .ZN(n18242) );
  OAI211_X1 U21277 ( .C1(n18558), .C2(n18562), .A(n18243), .B(n18242), .ZN(
        P3_U2881) );
  INV_X1 U21278 ( .A(n18625), .ZN(n18613) );
  AOI22_X1 U21279 ( .A1(n18566), .A2(n18530), .B1(n18614), .B2(n18246), .ZN(
        n18245) );
  AOI22_X1 U21280 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18247), .B1(
        n18616), .B2(n18312), .ZN(n18244) );
  OAI211_X1 U21281 ( .C1(n18613), .C2(n18533), .A(n18245), .B(n18244), .ZN(
        P3_U2882) );
  INV_X1 U21282 ( .A(n18622), .ZN(n18513) );
  AOI22_X1 U21283 ( .A1(n18566), .A2(n18509), .B1(n18621), .B2(n18246), .ZN(
        n18249) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18247), .B1(
        n18624), .B2(n18312), .ZN(n18248) );
  OAI211_X1 U21285 ( .C1(n18613), .C2(n18513), .A(n18249), .B(n18248), .ZN(
        P3_U2883) );
  NOR2_X2 U21286 ( .A1(n18316), .A2(n18250), .ZN(n18331) );
  NOR2_X1 U21287 ( .A1(n18312), .A2(n18331), .ZN(n18294) );
  NOR2_X1 U21288 ( .A1(n9706), .A2(n18294), .ZN(n18267) );
  AOI22_X1 U21289 ( .A1(n18279), .A2(n18573), .B1(n18572), .B2(n18267), .ZN(
        n18254) );
  INV_X1 U21290 ( .A(n18294), .ZN(n18252) );
  OAI221_X1 U21291 ( .B1(n18252), .B2(n18543), .C1(n18252), .C2(n18251), .A(
        n18541), .ZN(n18268) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18268), .B1(
        n18578), .B2(n18331), .ZN(n18253) );
  OAI211_X1 U21293 ( .C1(n18613), .C2(n18581), .A(n18254), .B(n18253), .ZN(
        P3_U2884) );
  INV_X1 U21294 ( .A(n18331), .ZN(n18338) );
  AOI22_X1 U21295 ( .A1(n18625), .A2(n18583), .B1(n18582), .B2(n18267), .ZN(
        n18256) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18268), .B1(
        n18279), .B2(n18584), .ZN(n18255) );
  OAI211_X1 U21297 ( .C1(n18587), .C2(n18338), .A(n18256), .B(n18255), .ZN(
        P3_U2885) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18268), .B1(
        n18588), .B2(n18267), .ZN(n18258) );
  AOI22_X1 U21299 ( .A1(n18279), .A2(n18589), .B1(n18590), .B2(n18331), .ZN(
        n18257) );
  OAI211_X1 U21300 ( .C1(n18613), .C2(n18593), .A(n18258), .B(n18257), .ZN(
        P3_U2886) );
  INV_X1 U21301 ( .A(n18551), .ZN(n18599) );
  INV_X1 U21302 ( .A(n18554), .ZN(n18595) );
  AOI22_X1 U21303 ( .A1(n18625), .A2(n18595), .B1(n18594), .B2(n18267), .ZN(
        n18260) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18268), .B1(
        n18279), .B2(n18596), .ZN(n18259) );
  OAI211_X1 U21305 ( .C1(n18599), .C2(n18338), .A(n18260), .B(n18259), .ZN(
        P3_U2887) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18268), .B1(
        n18600), .B2(n18267), .ZN(n18262) );
  AOI22_X1 U21307 ( .A1(n18279), .A2(n18602), .B1(n18442), .B2(n18331), .ZN(
        n18261) );
  OAI211_X1 U21308 ( .C1(n18613), .C2(n18445), .A(n18262), .B(n18261), .ZN(
        P3_U2888) );
  INV_X1 U21309 ( .A(n18559), .ZN(n18612) );
  INV_X1 U21310 ( .A(n18562), .ZN(n18608) );
  AOI22_X1 U21311 ( .A1(n18625), .A2(n18608), .B1(n18606), .B2(n18267), .ZN(
        n18264) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18268), .B1(
        n18279), .B2(n18609), .ZN(n18263) );
  OAI211_X1 U21313 ( .C1(n18612), .C2(n18338), .A(n18264), .B(n18263), .ZN(
        P3_U2889) );
  INV_X1 U21314 ( .A(n18279), .ZN(n18292) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18268), .B1(
        n18614), .B2(n18267), .ZN(n18266) );
  AOI22_X1 U21316 ( .A1(n18625), .A2(n18530), .B1(n18616), .B2(n18331), .ZN(
        n18265) );
  OAI211_X1 U21317 ( .C1(n18292), .C2(n18533), .A(n18266), .B(n18265), .ZN(
        P3_U2890) );
  AOI22_X1 U21318 ( .A1(n18279), .A2(n18622), .B1(n18621), .B2(n18267), .ZN(
        n18270) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18268), .B1(
        n18624), .B2(n18331), .ZN(n18269) );
  OAI211_X1 U21320 ( .C1(n18613), .C2(n18630), .A(n18270), .B(n18269), .ZN(
        P3_U2891) );
  INV_X1 U21321 ( .A(n18671), .ZN(n18456) );
  NAND2_X1 U21322 ( .A1(n18456), .A2(n18272), .ZN(n18360) );
  AOI22_X1 U21323 ( .A1(n18279), .A2(n18488), .B1(n18572), .B2(n18288), .ZN(
        n18274) );
  INV_X1 U21324 ( .A(n18543), .ZN(n18431) );
  AOI21_X1 U21325 ( .B1(n18672), .B2(n18431), .A(n18271), .ZN(n18362) );
  NAND2_X1 U21326 ( .A1(n18272), .A2(n18362), .ZN(n18289) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18289), .B1(
        n18573), .B2(n18312), .ZN(n18273) );
  OAI211_X1 U21328 ( .C1(n18491), .C2(n18360), .A(n18274), .B(n18273), .ZN(
        P3_U2892) );
  AOI22_X1 U21329 ( .A1(n18279), .A2(n18583), .B1(n18582), .B2(n18288), .ZN(
        n18276) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18289), .B1(
        n18584), .B2(n18312), .ZN(n18275) );
  OAI211_X1 U21331 ( .C1(n18587), .C2(n18360), .A(n18276), .B(n18275), .ZN(
        P3_U2893) );
  AOI22_X1 U21332 ( .A1(n18588), .A2(n18288), .B1(n18589), .B2(n18312), .ZN(
        n18278) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18289), .B1(
        n18279), .B2(n18465), .ZN(n18277) );
  OAI211_X1 U21334 ( .C1(n18468), .C2(n18360), .A(n18278), .B(n18277), .ZN(
        P3_U2894) );
  AOI22_X1 U21335 ( .A1(n18596), .A2(n18312), .B1(n18594), .B2(n18288), .ZN(
        n18281) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18289), .B1(
        n18279), .B2(n18595), .ZN(n18280) );
  OAI211_X1 U21337 ( .C1(n18599), .C2(n18360), .A(n18281), .B(n18280), .ZN(
        P3_U2895) );
  AOI22_X1 U21338 ( .A1(n18602), .A2(n18312), .B1(n18600), .B2(n18288), .ZN(
        n18283) );
  INV_X1 U21339 ( .A(n18360), .ZN(n18353) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18289), .B1(
        n18442), .B2(n18353), .ZN(n18282) );
  OAI211_X1 U21341 ( .C1(n18292), .C2(n18445), .A(n18283), .B(n18282), .ZN(
        P3_U2896) );
  AOI22_X1 U21342 ( .A1(n18609), .A2(n18312), .B1(n18606), .B2(n18288), .ZN(
        n18285) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18289), .B1(
        n18559), .B2(n18353), .ZN(n18284) );
  OAI211_X1 U21344 ( .C1(n18292), .C2(n18562), .A(n18285), .B(n18284), .ZN(
        P3_U2897) );
  INV_X1 U21345 ( .A(n18533), .ZN(n18615) );
  AOI22_X1 U21346 ( .A1(n18615), .A2(n18312), .B1(n18614), .B2(n18288), .ZN(
        n18287) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18289), .B1(
        n18616), .B2(n18353), .ZN(n18286) );
  OAI211_X1 U21348 ( .C1(n18292), .C2(n18619), .A(n18287), .B(n18286), .ZN(
        P3_U2898) );
  AOI22_X1 U21349 ( .A1(n18622), .A2(n18312), .B1(n18621), .B2(n18288), .ZN(
        n18291) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18289), .B1(
        n18624), .B2(n18353), .ZN(n18290) );
  OAI211_X1 U21351 ( .C1(n18292), .C2(n18630), .A(n18291), .B(n18290), .ZN(
        P3_U2899) );
  INV_X1 U21352 ( .A(n18673), .ZN(n18293) );
  NAND2_X1 U21353 ( .A1(n18293), .A2(n18361), .ZN(n18383) );
  AOI21_X1 U21354 ( .B1(n18360), .B2(n18383), .A(n9706), .ZN(n18311) );
  AOI22_X1 U21355 ( .A1(n18573), .A2(n18331), .B1(n18572), .B2(n18311), .ZN(
        n18297) );
  INV_X1 U21356 ( .A(n18383), .ZN(n18372) );
  AOI221_X1 U21357 ( .B1(n18294), .B2(n18360), .C1(n18431), .C2(n18360), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18295) );
  OAI21_X1 U21358 ( .B1(n18372), .B2(n18295), .A(n18487), .ZN(n18313) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18313), .B1(
        n18578), .B2(n18372), .ZN(n18296) );
  OAI211_X1 U21360 ( .C1(n18581), .C2(n18310), .A(n18297), .B(n18296), .ZN(
        P3_U2900) );
  AOI22_X1 U21361 ( .A1(n18583), .A2(n18312), .B1(n18582), .B2(n18311), .ZN(
        n18299) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18313), .B1(
        n18584), .B2(n18331), .ZN(n18298) );
  OAI211_X1 U21363 ( .C1(n18587), .C2(n18383), .A(n18299), .B(n18298), .ZN(
        P3_U2901) );
  AOI22_X1 U21364 ( .A1(n18588), .A2(n18311), .B1(n18589), .B2(n18331), .ZN(
        n18301) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18313), .B1(
        n18590), .B2(n18372), .ZN(n18300) );
  OAI211_X1 U21366 ( .C1(n18593), .C2(n18310), .A(n18301), .B(n18300), .ZN(
        P3_U2902) );
  AOI22_X1 U21367 ( .A1(n18596), .A2(n18331), .B1(n18594), .B2(n18311), .ZN(
        n18303) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18313), .B1(
        n18551), .B2(n18372), .ZN(n18302) );
  OAI211_X1 U21369 ( .C1(n18554), .C2(n18310), .A(n18303), .B(n18302), .ZN(
        P3_U2903) );
  AOI22_X1 U21370 ( .A1(n18602), .A2(n18331), .B1(n18600), .B2(n18311), .ZN(
        n18305) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18313), .B1(
        n18442), .B2(n18372), .ZN(n18304) );
  OAI211_X1 U21372 ( .C1(n18445), .C2(n18310), .A(n18305), .B(n18304), .ZN(
        P3_U2904) );
  AOI22_X1 U21373 ( .A1(n18609), .A2(n18331), .B1(n18606), .B2(n18311), .ZN(
        n18307) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18313), .B1(
        n18559), .B2(n18372), .ZN(n18306) );
  OAI211_X1 U21375 ( .C1(n18562), .C2(n18310), .A(n18307), .B(n18306), .ZN(
        P3_U2905) );
  AOI22_X1 U21376 ( .A1(n18615), .A2(n18331), .B1(n18614), .B2(n18311), .ZN(
        n18309) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18313), .B1(
        n18616), .B2(n18372), .ZN(n18308) );
  OAI211_X1 U21378 ( .C1(n18619), .C2(n18310), .A(n18309), .B(n18308), .ZN(
        P3_U2906) );
  AOI22_X1 U21379 ( .A1(n18509), .A2(n18312), .B1(n18621), .B2(n18311), .ZN(
        n18315) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18313), .B1(
        n18624), .B2(n18372), .ZN(n18314) );
  OAI211_X1 U21381 ( .C1(n18513), .C2(n18338), .A(n18315), .B(n18314), .ZN(
        P3_U2907) );
  NAND2_X1 U21382 ( .A1(n18406), .A2(n18361), .ZN(n18405) );
  AOI22_X1 U21383 ( .A1(n18573), .A2(n18353), .B1(n18572), .B2(n18334), .ZN(
        n18320) );
  NOR2_X1 U21384 ( .A1(n18672), .A2(n18316), .ZN(n18318) );
  AOI22_X1 U21385 ( .A1(n18577), .A2(n18318), .B1(n18317), .B2(n18361), .ZN(
        n18335) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18335), .B1(
        n18488), .B2(n18331), .ZN(n18319) );
  OAI211_X1 U21387 ( .C1(n18491), .C2(n18405), .A(n18320), .B(n18319), .ZN(
        P3_U2908) );
  AOI22_X1 U21388 ( .A1(n18582), .A2(n18334), .B1(n18584), .B2(n18353), .ZN(
        n18322) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18335), .B1(
        n18583), .B2(n18331), .ZN(n18321) );
  OAI211_X1 U21390 ( .C1(n18587), .C2(n18405), .A(n18322), .B(n18321), .ZN(
        P3_U2909) );
  AOI22_X1 U21391 ( .A1(n18588), .A2(n18334), .B1(n18589), .B2(n18353), .ZN(
        n18324) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18335), .B1(
        n18465), .B2(n18331), .ZN(n18323) );
  OAI211_X1 U21393 ( .C1(n18468), .C2(n18405), .A(n18324), .B(n18323), .ZN(
        P3_U2910) );
  AOI22_X1 U21394 ( .A1(n18595), .A2(n18331), .B1(n18594), .B2(n18334), .ZN(
        n18326) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18335), .B1(
        n18596), .B2(n18353), .ZN(n18325) );
  OAI211_X1 U21396 ( .C1(n18599), .C2(n18405), .A(n18326), .B(n18325), .ZN(
        P3_U2911) );
  INV_X1 U21397 ( .A(n18442), .ZN(n18605) );
  INV_X1 U21398 ( .A(n18445), .ZN(n18601) );
  AOI22_X1 U21399 ( .A1(n18601), .A2(n18331), .B1(n18600), .B2(n18334), .ZN(
        n18328) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18335), .B1(
        n18602), .B2(n18353), .ZN(n18327) );
  OAI211_X1 U21401 ( .C1(n18605), .C2(n18405), .A(n18328), .B(n18327), .ZN(
        P3_U2912) );
  AOI22_X1 U21402 ( .A1(n18609), .A2(n18353), .B1(n18606), .B2(n18334), .ZN(
        n18330) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18335), .B1(
        n18608), .B2(n18331), .ZN(n18329) );
  OAI211_X1 U21404 ( .C1(n18612), .C2(n18405), .A(n18330), .B(n18329), .ZN(
        P3_U2913) );
  AOI22_X1 U21405 ( .A1(n18530), .A2(n18331), .B1(n18614), .B2(n18334), .ZN(
        n18333) );
  INV_X1 U21406 ( .A(n18405), .ZN(n18390) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18335), .B1(
        n18616), .B2(n18390), .ZN(n18332) );
  OAI211_X1 U21408 ( .C1(n18533), .C2(n18360), .A(n18333), .B(n18332), .ZN(
        P3_U2914) );
  AOI22_X1 U21409 ( .A1(n18622), .A2(n18353), .B1(n18621), .B2(n18334), .ZN(
        n18337) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18335), .B1(
        n18624), .B2(n18390), .ZN(n18336) );
  OAI211_X1 U21411 ( .C1(n18630), .C2(n18338), .A(n18337), .B(n18336), .ZN(
        P3_U2915) );
  NAND2_X1 U21412 ( .A1(n18430), .A2(n18361), .ZN(n18424) );
  INV_X1 U21413 ( .A(n18424), .ZN(n18426) );
  NOR2_X1 U21414 ( .A1(n18390), .A2(n18426), .ZN(n18384) );
  NOR2_X1 U21415 ( .A1(n9706), .A2(n18384), .ZN(n18356) );
  AOI22_X1 U21416 ( .A1(n18488), .A2(n18353), .B1(n18572), .B2(n18356), .ZN(
        n18342) );
  NOR2_X1 U21417 ( .A1(n18353), .A2(n18372), .ZN(n18339) );
  OAI21_X1 U21418 ( .B1(n18339), .B2(n18431), .A(n18384), .ZN(n18340) );
  OAI211_X1 U21419 ( .C1(n18426), .C2(n18803), .A(n18487), .B(n18340), .ZN(
        n18357) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18357), .B1(
        n18573), .B2(n18372), .ZN(n18341) );
  OAI211_X1 U21421 ( .C1(n18491), .C2(n18424), .A(n18342), .B(n18341), .ZN(
        P3_U2916) );
  AOI22_X1 U21422 ( .A1(n18582), .A2(n18356), .B1(n18584), .B2(n18372), .ZN(
        n18344) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18357), .B1(
        n18492), .B2(n18426), .ZN(n18343) );
  OAI211_X1 U21424 ( .C1(n18495), .C2(n18360), .A(n18344), .B(n18343), .ZN(
        P3_U2917) );
  AOI22_X1 U21425 ( .A1(n18465), .A2(n18353), .B1(n18588), .B2(n18356), .ZN(
        n18346) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18357), .B1(
        n18589), .B2(n18372), .ZN(n18345) );
  OAI211_X1 U21427 ( .C1(n18468), .C2(n18424), .A(n18346), .B(n18345), .ZN(
        P3_U2918) );
  AOI22_X1 U21428 ( .A1(n18595), .A2(n18353), .B1(n18594), .B2(n18356), .ZN(
        n18348) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18357), .B1(
        n18596), .B2(n18372), .ZN(n18347) );
  OAI211_X1 U21430 ( .C1(n18599), .C2(n18424), .A(n18348), .B(n18347), .ZN(
        P3_U2919) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18357), .B1(
        n18600), .B2(n18356), .ZN(n18350) );
  AOI22_X1 U21432 ( .A1(n18442), .A2(n18426), .B1(n18602), .B2(n18372), .ZN(
        n18349) );
  OAI211_X1 U21433 ( .C1(n18445), .C2(n18360), .A(n18350), .B(n18349), .ZN(
        P3_U2920) );
  AOI22_X1 U21434 ( .A1(n18608), .A2(n18353), .B1(n18606), .B2(n18356), .ZN(
        n18352) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18357), .B1(
        n18609), .B2(n18372), .ZN(n18351) );
  OAI211_X1 U21436 ( .C1(n18612), .C2(n18424), .A(n18352), .B(n18351), .ZN(
        P3_U2921) );
  AOI22_X1 U21437 ( .A1(n18530), .A2(n18353), .B1(n18614), .B2(n18356), .ZN(
        n18355) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18357), .B1(
        n18616), .B2(n18426), .ZN(n18354) );
  OAI211_X1 U21439 ( .C1(n18533), .C2(n18383), .A(n18355), .B(n18354), .ZN(
        P3_U2922) );
  AOI22_X1 U21440 ( .A1(n18622), .A2(n18372), .B1(n18621), .B2(n18356), .ZN(
        n18359) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18357), .B1(
        n18624), .B2(n18426), .ZN(n18358) );
  OAI211_X1 U21442 ( .C1(n18630), .C2(n18360), .A(n18359), .B(n18358), .ZN(
        P3_U2923) );
  AOI22_X1 U21443 ( .A1(n18573), .A2(n18390), .B1(n18572), .B2(n18379), .ZN(
        n18365) );
  NAND2_X1 U21444 ( .A1(n18362), .A2(n18361), .ZN(n18380) );
  NOR2_X2 U21445 ( .A1(n18671), .A2(n18363), .ZN(n18448) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18380), .B1(
        n18578), .B2(n18448), .ZN(n18364) );
  OAI211_X1 U21447 ( .C1(n18581), .C2(n18383), .A(n18365), .B(n18364), .ZN(
        P3_U2924) );
  INV_X1 U21448 ( .A(n18448), .ZN(n18455) );
  AOI22_X1 U21449 ( .A1(n18583), .A2(n18372), .B1(n18582), .B2(n18379), .ZN(
        n18367) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18380), .B1(
        n18584), .B2(n18390), .ZN(n18366) );
  OAI211_X1 U21451 ( .C1(n18587), .C2(n18455), .A(n18367), .B(n18366), .ZN(
        P3_U2925) );
  AOI22_X1 U21452 ( .A1(n18465), .A2(n18372), .B1(n18588), .B2(n18379), .ZN(
        n18369) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18380), .B1(
        n18589), .B2(n18390), .ZN(n18368) );
  OAI211_X1 U21454 ( .C1(n18468), .C2(n18455), .A(n18369), .B(n18368), .ZN(
        P3_U2926) );
  AOI22_X1 U21455 ( .A1(n18596), .A2(n18390), .B1(n18594), .B2(n18379), .ZN(
        n18371) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18380), .B1(
        n18551), .B2(n18448), .ZN(n18370) );
  OAI211_X1 U21457 ( .C1(n18554), .C2(n18383), .A(n18371), .B(n18370), .ZN(
        P3_U2927) );
  AOI22_X1 U21458 ( .A1(n18601), .A2(n18372), .B1(n18600), .B2(n18379), .ZN(
        n18374) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18380), .B1(
        n18602), .B2(n18390), .ZN(n18373) );
  OAI211_X1 U21460 ( .C1(n18605), .C2(n18455), .A(n18374), .B(n18373), .ZN(
        P3_U2928) );
  AOI22_X1 U21461 ( .A1(n18609), .A2(n18390), .B1(n18606), .B2(n18379), .ZN(
        n18376) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18380), .B1(
        n18559), .B2(n18448), .ZN(n18375) );
  OAI211_X1 U21463 ( .C1(n18562), .C2(n18383), .A(n18376), .B(n18375), .ZN(
        P3_U2929) );
  AOI22_X1 U21464 ( .A1(n18615), .A2(n18390), .B1(n18614), .B2(n18379), .ZN(
        n18378) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18380), .B1(
        n18616), .B2(n18448), .ZN(n18377) );
  OAI211_X1 U21466 ( .C1(n18619), .C2(n18383), .A(n18378), .B(n18377), .ZN(
        P3_U2930) );
  AOI22_X1 U21467 ( .A1(n18622), .A2(n18390), .B1(n18621), .B2(n18379), .ZN(
        n18382) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18380), .B1(
        n18624), .B2(n18448), .ZN(n18381) );
  OAI211_X1 U21469 ( .C1(n18630), .C2(n18383), .A(n18382), .B(n18381), .ZN(
        P3_U2931) );
  NOR2_X1 U21470 ( .A1(n18673), .A2(n18457), .ZN(n18464) );
  CLKBUF_X1 U21471 ( .A(n18464), .Z(n18473) );
  NOR2_X1 U21472 ( .A1(n18448), .A2(n18473), .ZN(n18432) );
  NOR2_X1 U21473 ( .A1(n9706), .A2(n18432), .ZN(n18401) );
  AOI22_X1 U21474 ( .A1(n18573), .A2(n18426), .B1(n18572), .B2(n18401), .ZN(
        n18387) );
  OAI21_X1 U21475 ( .B1(n18384), .B2(n18431), .A(n18432), .ZN(n18385) );
  OAI211_X1 U21476 ( .C1(n18473), .C2(n18803), .A(n18487), .B(n18385), .ZN(
        n18402) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18402), .B1(
        n18578), .B2(n18464), .ZN(n18386) );
  OAI211_X1 U21478 ( .C1(n18581), .C2(n18405), .A(n18387), .B(n18386), .ZN(
        P3_U2932) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18402), .B1(
        n18582), .B2(n18401), .ZN(n18389) );
  AOI22_X1 U21480 ( .A1(n18492), .A2(n18473), .B1(n18584), .B2(n18426), .ZN(
        n18388) );
  OAI211_X1 U21481 ( .C1(n18495), .C2(n18405), .A(n18389), .B(n18388), .ZN(
        P3_U2933) );
  INV_X1 U21482 ( .A(n18464), .ZN(n18482) );
  AOI22_X1 U21483 ( .A1(n18465), .A2(n18390), .B1(n18588), .B2(n18401), .ZN(
        n18392) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18402), .B1(
        n18589), .B2(n18426), .ZN(n18391) );
  OAI211_X1 U21485 ( .C1(n18468), .C2(n18482), .A(n18392), .B(n18391), .ZN(
        P3_U2934) );
  AOI22_X1 U21486 ( .A1(n18596), .A2(n18426), .B1(n18594), .B2(n18401), .ZN(
        n18394) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18402), .B1(
        n18551), .B2(n18464), .ZN(n18393) );
  OAI211_X1 U21488 ( .C1(n18554), .C2(n18405), .A(n18394), .B(n18393), .ZN(
        P3_U2935) );
  AOI22_X1 U21489 ( .A1(n18602), .A2(n18426), .B1(n18600), .B2(n18401), .ZN(
        n18396) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18402), .B1(
        n18442), .B2(n18473), .ZN(n18395) );
  OAI211_X1 U21491 ( .C1(n18445), .C2(n18405), .A(n18396), .B(n18395), .ZN(
        P3_U2936) );
  AOI22_X1 U21492 ( .A1(n18609), .A2(n18426), .B1(n18606), .B2(n18401), .ZN(
        n18398) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18402), .B1(
        n18559), .B2(n18464), .ZN(n18397) );
  OAI211_X1 U21494 ( .C1(n18562), .C2(n18405), .A(n18398), .B(n18397), .ZN(
        P3_U2937) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18402), .B1(
        n18614), .B2(n18401), .ZN(n18400) );
  AOI22_X1 U21496 ( .A1(n18615), .A2(n18426), .B1(n18616), .B2(n18473), .ZN(
        n18399) );
  OAI211_X1 U21497 ( .C1(n18619), .C2(n18405), .A(n18400), .B(n18399), .ZN(
        P3_U2938) );
  AOI22_X1 U21498 ( .A1(n18622), .A2(n18426), .B1(n18621), .B2(n18401), .ZN(
        n18404) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18402), .B1(
        n18624), .B2(n18464), .ZN(n18403) );
  OAI211_X1 U21500 ( .C1(n18630), .C2(n18405), .A(n18404), .B(n18403), .ZN(
        P3_U2939) );
  NAND2_X1 U21501 ( .A1(n18406), .A2(n18459), .ZN(n18506) );
  AOI22_X1 U21502 ( .A1(n18573), .A2(n18448), .B1(n18572), .B2(n18425), .ZN(
        n18411) );
  NOR2_X1 U21503 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18407), .ZN(
        n18409) );
  NOR2_X1 U21504 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18457), .ZN(
        n18408) );
  AOI22_X1 U21505 ( .A1(n18577), .A2(n18409), .B1(n18575), .B2(n18408), .ZN(
        n18427) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18427), .B1(
        n18488), .B2(n18426), .ZN(n18410) );
  OAI211_X1 U21507 ( .C1(n18491), .C2(n18506), .A(n18411), .B(n18410), .ZN(
        P3_U2940) );
  AOI22_X1 U21508 ( .A1(n18582), .A2(n18425), .B1(n18584), .B2(n18448), .ZN(
        n18413) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18427), .B1(
        n18583), .B2(n18426), .ZN(n18412) );
  OAI211_X1 U21510 ( .C1(n18587), .C2(n18506), .A(n18413), .B(n18412), .ZN(
        P3_U2941) );
  AOI22_X1 U21511 ( .A1(n18465), .A2(n18426), .B1(n18588), .B2(n18425), .ZN(
        n18415) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18427), .B1(
        n18589), .B2(n18448), .ZN(n18414) );
  OAI211_X1 U21513 ( .C1(n18468), .C2(n18506), .A(n18415), .B(n18414), .ZN(
        P3_U2942) );
  AOI22_X1 U21514 ( .A1(n18595), .A2(n18426), .B1(n18594), .B2(n18425), .ZN(
        n18417) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18427), .B1(
        n18596), .B2(n18448), .ZN(n18416) );
  OAI211_X1 U21516 ( .C1(n18599), .C2(n18506), .A(n18417), .B(n18416), .ZN(
        P3_U2943) );
  AOI22_X1 U21517 ( .A1(n18602), .A2(n18448), .B1(n18600), .B2(n18425), .ZN(
        n18419) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18427), .B1(
        n18601), .B2(n18426), .ZN(n18418) );
  OAI211_X1 U21519 ( .C1(n18605), .C2(n18506), .A(n18419), .B(n18418), .ZN(
        P3_U2944) );
  AOI22_X1 U21520 ( .A1(n18609), .A2(n18448), .B1(n18606), .B2(n18425), .ZN(
        n18421) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18427), .B1(
        n18608), .B2(n18426), .ZN(n18420) );
  OAI211_X1 U21522 ( .C1(n18612), .C2(n18506), .A(n18421), .B(n18420), .ZN(
        P3_U2945) );
  AOI22_X1 U21523 ( .A1(n18615), .A2(n18448), .B1(n18614), .B2(n18425), .ZN(
        n18423) );
  INV_X1 U21524 ( .A(n18506), .ZN(n18508) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18427), .B1(
        n18616), .B2(n18508), .ZN(n18422) );
  OAI211_X1 U21526 ( .C1(n18619), .C2(n18424), .A(n18423), .B(n18422), .ZN(
        P3_U2946) );
  AOI22_X1 U21527 ( .A1(n18509), .A2(n18426), .B1(n18621), .B2(n18425), .ZN(
        n18429) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18427), .B1(
        n18624), .B2(n18508), .ZN(n18428) );
  OAI211_X1 U21529 ( .C1(n18513), .C2(n18455), .A(n18429), .B(n18428), .ZN(
        P3_U2947) );
  NAND2_X1 U21530 ( .A1(n18430), .A2(n18459), .ZN(n18538) );
  AOI21_X1 U21531 ( .B1(n18506), .B2(n18538), .A(n9706), .ZN(n18451) );
  AOI22_X1 U21532 ( .A1(n18573), .A2(n18473), .B1(n18572), .B2(n18451), .ZN(
        n18435) );
  OAI211_X1 U21533 ( .C1(n18432), .C2(n18431), .A(n18506), .B(n18538), .ZN(
        n18433) );
  NAND2_X1 U21534 ( .A1(n18541), .A2(n18433), .ZN(n18452) );
  INV_X1 U21535 ( .A(n18538), .ZN(n18529) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18452), .B1(
        n18578), .B2(n18529), .ZN(n18434) );
  OAI211_X1 U21537 ( .C1(n18581), .C2(n18455), .A(n18435), .B(n18434), .ZN(
        P3_U2948) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18452), .B1(
        n18582), .B2(n18451), .ZN(n18437) );
  AOI22_X1 U21539 ( .A1(n18492), .A2(n18529), .B1(n18584), .B2(n18473), .ZN(
        n18436) );
  OAI211_X1 U21540 ( .C1(n18495), .C2(n18455), .A(n18437), .B(n18436), .ZN(
        P3_U2949) );
  AOI22_X1 U21541 ( .A1(n18465), .A2(n18448), .B1(n18588), .B2(n18451), .ZN(
        n18439) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18452), .B1(
        n18589), .B2(n18464), .ZN(n18438) );
  OAI211_X1 U21543 ( .C1(n18468), .C2(n18538), .A(n18439), .B(n18438), .ZN(
        P3_U2950) );
  AOI22_X1 U21544 ( .A1(n18596), .A2(n18464), .B1(n18594), .B2(n18451), .ZN(
        n18441) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18452), .B1(
        n18551), .B2(n18529), .ZN(n18440) );
  OAI211_X1 U21546 ( .C1(n18554), .C2(n18455), .A(n18441), .B(n18440), .ZN(
        P3_U2951) );
  AOI22_X1 U21547 ( .A1(n18602), .A2(n18473), .B1(n18600), .B2(n18451), .ZN(
        n18444) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18452), .B1(
        n18442), .B2(n18529), .ZN(n18443) );
  OAI211_X1 U21549 ( .C1(n18445), .C2(n18455), .A(n18444), .B(n18443), .ZN(
        P3_U2952) );
  AOI22_X1 U21550 ( .A1(n18608), .A2(n18448), .B1(n18606), .B2(n18451), .ZN(
        n18447) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18452), .B1(
        n18609), .B2(n18464), .ZN(n18446) );
  OAI211_X1 U21552 ( .C1(n18612), .C2(n18538), .A(n18447), .B(n18446), .ZN(
        P3_U2953) );
  AOI22_X1 U21553 ( .A1(n18530), .A2(n18448), .B1(n18614), .B2(n18451), .ZN(
        n18450) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18452), .B1(
        n18616), .B2(n18529), .ZN(n18449) );
  OAI211_X1 U21555 ( .C1(n18533), .C2(n18482), .A(n18450), .B(n18449), .ZN(
        P3_U2954) );
  AOI22_X1 U21556 ( .A1(n18622), .A2(n18464), .B1(n18621), .B2(n18451), .ZN(
        n18454) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18452), .B1(
        n18624), .B2(n18529), .ZN(n18453) );
  OAI211_X1 U21558 ( .C1(n18630), .C2(n18455), .A(n18454), .B(n18453), .ZN(
        P3_U2955) );
  NAND2_X1 U21559 ( .A1(n18456), .A2(n18459), .ZN(n18570) );
  NOR2_X1 U21560 ( .A1(n18672), .A2(n18457), .ZN(n18515) );
  INV_X1 U21561 ( .A(n18515), .ZN(n18458) );
  NOR2_X1 U21562 ( .A1(n9706), .A2(n18458), .ZN(n18478) );
  AOI22_X1 U21563 ( .A1(n18488), .A2(n18473), .B1(n18572), .B2(n18478), .ZN(
        n18461) );
  OAI211_X1 U21564 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18577), .A(
        n18575), .B(n18459), .ZN(n18479) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18479), .B1(
        n18573), .B2(n18508), .ZN(n18460) );
  OAI211_X1 U21566 ( .C1(n18491), .C2(n18570), .A(n18461), .B(n18460), .ZN(
        P3_U2956) );
  AOI22_X1 U21567 ( .A1(n18582), .A2(n18478), .B1(n18584), .B2(n18508), .ZN(
        n18463) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18479), .B1(
        n18583), .B2(n18464), .ZN(n18462) );
  OAI211_X1 U21569 ( .C1(n18587), .C2(n18570), .A(n18463), .B(n18462), .ZN(
        P3_U2957) );
  AOI22_X1 U21570 ( .A1(n18588), .A2(n18478), .B1(n18589), .B2(n18508), .ZN(
        n18467) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18479), .B1(
        n18465), .B2(n18464), .ZN(n18466) );
  OAI211_X1 U21572 ( .C1(n18468), .C2(n18570), .A(n18467), .B(n18466), .ZN(
        P3_U2958) );
  AOI22_X1 U21573 ( .A1(n18595), .A2(n18473), .B1(n18594), .B2(n18478), .ZN(
        n18470) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18479), .B1(
        n18596), .B2(n18508), .ZN(n18469) );
  OAI211_X1 U21575 ( .C1(n18599), .C2(n18570), .A(n18470), .B(n18469), .ZN(
        P3_U2959) );
  AOI22_X1 U21576 ( .A1(n18602), .A2(n18508), .B1(n18600), .B2(n18478), .ZN(
        n18472) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18479), .B1(
        n18601), .B2(n18473), .ZN(n18471) );
  OAI211_X1 U21578 ( .C1(n18605), .C2(n18570), .A(n18472), .B(n18471), .ZN(
        P3_U2960) );
  AOI22_X1 U21579 ( .A1(n18609), .A2(n18508), .B1(n18606), .B2(n18478), .ZN(
        n18475) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18479), .B1(
        n18608), .B2(n18473), .ZN(n18474) );
  OAI211_X1 U21581 ( .C1(n18612), .C2(n18570), .A(n18475), .B(n18474), .ZN(
        P3_U2961) );
  AOI22_X1 U21582 ( .A1(n18615), .A2(n18508), .B1(n18614), .B2(n18478), .ZN(
        n18477) );
  INV_X1 U21583 ( .A(n18570), .ZN(n18555) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18479), .B1(
        n18616), .B2(n18555), .ZN(n18476) );
  OAI211_X1 U21585 ( .C1(n18619), .C2(n18482), .A(n18477), .B(n18476), .ZN(
        P3_U2962) );
  AOI22_X1 U21586 ( .A1(n18622), .A2(n18508), .B1(n18621), .B2(n18478), .ZN(
        n18481) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18479), .B1(
        n18624), .B2(n18555), .ZN(n18480) );
  OAI211_X1 U21588 ( .C1(n18630), .C2(n18482), .A(n18481), .B(n18480), .ZN(
        P3_U2963) );
  NAND2_X1 U21589 ( .A1(n18576), .A2(n18483), .ZN(n18629) );
  INV_X1 U21590 ( .A(n18629), .ZN(n18607) );
  NOR2_X1 U21591 ( .A1(n18555), .A2(n18607), .ZN(n18540) );
  NOR2_X1 U21592 ( .A1(n9706), .A2(n18540), .ZN(n18507) );
  AOI22_X1 U21593 ( .A1(n18573), .A2(n18529), .B1(n18572), .B2(n18507), .ZN(
        n18490) );
  OAI21_X1 U21594 ( .B1(n18485), .B2(n18484), .A(n18540), .ZN(n18486) );
  OAI211_X1 U21595 ( .C1(n18607), .C2(n18803), .A(n18487), .B(n18486), .ZN(
        n18510) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18510), .B1(
        n18488), .B2(n18508), .ZN(n18489) );
  OAI211_X1 U21597 ( .C1(n18491), .C2(n18629), .A(n18490), .B(n18489), .ZN(
        P3_U2964) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18510), .B1(
        n18582), .B2(n18507), .ZN(n18494) );
  AOI22_X1 U21599 ( .A1(n18492), .A2(n18607), .B1(n18584), .B2(n18529), .ZN(
        n18493) );
  OAI211_X1 U21600 ( .C1(n18495), .C2(n18506), .A(n18494), .B(n18493), .ZN(
        P3_U2965) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18510), .B1(
        n18588), .B2(n18507), .ZN(n18497) );
  AOI22_X1 U21602 ( .A1(n18590), .A2(n18607), .B1(n18589), .B2(n18529), .ZN(
        n18496) );
  OAI211_X1 U21603 ( .C1(n18593), .C2(n18506), .A(n18497), .B(n18496), .ZN(
        P3_U2966) );
  AOI22_X1 U21604 ( .A1(n18595), .A2(n18508), .B1(n18594), .B2(n18507), .ZN(
        n18499) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18510), .B1(
        n18596), .B2(n18529), .ZN(n18498) );
  OAI211_X1 U21606 ( .C1(n18599), .C2(n18629), .A(n18499), .B(n18498), .ZN(
        P3_U2967) );
  AOI22_X1 U21607 ( .A1(n18601), .A2(n18508), .B1(n18600), .B2(n18507), .ZN(
        n18501) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18510), .B1(
        n18602), .B2(n18529), .ZN(n18500) );
  OAI211_X1 U21609 ( .C1(n18605), .C2(n18629), .A(n18501), .B(n18500), .ZN(
        P3_U2968) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18510), .B1(
        n18606), .B2(n18507), .ZN(n18503) );
  AOI22_X1 U21611 ( .A1(n18559), .A2(n18607), .B1(n18609), .B2(n18529), .ZN(
        n18502) );
  OAI211_X1 U21612 ( .C1(n18562), .C2(n18506), .A(n18503), .B(n18502), .ZN(
        P3_U2969) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18510), .B1(
        n18614), .B2(n18507), .ZN(n18505) );
  AOI22_X1 U21614 ( .A1(n18615), .A2(n18529), .B1(n18616), .B2(n18607), .ZN(
        n18504) );
  OAI211_X1 U21615 ( .C1(n18619), .C2(n18506), .A(n18505), .B(n18504), .ZN(
        P3_U2970) );
  AOI22_X1 U21616 ( .A1(n18509), .A2(n18508), .B1(n18621), .B2(n18507), .ZN(
        n18512) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18510), .B1(
        n18624), .B2(n18607), .ZN(n18511) );
  OAI211_X1 U21618 ( .C1(n18513), .C2(n18538), .A(n18512), .B(n18511), .ZN(
        P3_U2971) );
  INV_X1 U21619 ( .A(n18576), .ZN(n18514) );
  NOR2_X1 U21620 ( .A1(n9706), .A2(n18514), .ZN(n18534) );
  AOI22_X1 U21621 ( .A1(n18573), .A2(n18555), .B1(n18572), .B2(n18534), .ZN(
        n18517) );
  AOI22_X1 U21622 ( .A1(n18577), .A2(n18515), .B1(n18576), .B2(n18575), .ZN(
        n18535) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18535), .B1(
        n18623), .B2(n18578), .ZN(n18516) );
  OAI211_X1 U21624 ( .C1(n18581), .C2(n18538), .A(n18517), .B(n18516), .ZN(
        P3_U2972) );
  AOI22_X1 U21625 ( .A1(n18583), .A2(n18529), .B1(n18582), .B2(n18534), .ZN(
        n18519) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18535), .B1(
        n18584), .B2(n18555), .ZN(n18518) );
  OAI211_X1 U21627 ( .C1(n18526), .C2(n18587), .A(n18519), .B(n18518), .ZN(
        P3_U2973) );
  AOI22_X1 U21628 ( .A1(n18588), .A2(n18534), .B1(n18589), .B2(n18555), .ZN(
        n18521) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18535), .B1(
        n18623), .B2(n18590), .ZN(n18520) );
  OAI211_X1 U21630 ( .C1(n18593), .C2(n18538), .A(n18521), .B(n18520), .ZN(
        P3_U2974) );
  AOI22_X1 U21631 ( .A1(n18596), .A2(n18555), .B1(n18594), .B2(n18534), .ZN(
        n18523) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18535), .B1(
        n18623), .B2(n18551), .ZN(n18522) );
  OAI211_X1 U21633 ( .C1(n18554), .C2(n18538), .A(n18523), .B(n18522), .ZN(
        P3_U2975) );
  AOI22_X1 U21634 ( .A1(n18601), .A2(n18529), .B1(n18600), .B2(n18534), .ZN(
        n18525) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18535), .B1(
        n18602), .B2(n18555), .ZN(n18524) );
  OAI211_X1 U21636 ( .C1(n18526), .C2(n18605), .A(n18525), .B(n18524), .ZN(
        P3_U2976) );
  AOI22_X1 U21637 ( .A1(n18609), .A2(n18555), .B1(n18606), .B2(n18534), .ZN(
        n18528) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18535), .B1(
        n18623), .B2(n18559), .ZN(n18527) );
  OAI211_X1 U21639 ( .C1(n18562), .C2(n18538), .A(n18528), .B(n18527), .ZN(
        P3_U2977) );
  AOI22_X1 U21640 ( .A1(n18530), .A2(n18529), .B1(n18614), .B2(n18534), .ZN(
        n18532) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18535), .B1(
        n18623), .B2(n18616), .ZN(n18531) );
  OAI211_X1 U21642 ( .C1(n18533), .C2(n18570), .A(n18532), .B(n18531), .ZN(
        P3_U2978) );
  AOI22_X1 U21643 ( .A1(n18622), .A2(n18555), .B1(n18621), .B2(n18534), .ZN(
        n18537) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18535), .B1(
        n18623), .B2(n18624), .ZN(n18536) );
  OAI211_X1 U21645 ( .C1(n18630), .C2(n18538), .A(n18537), .B(n18536), .ZN(
        P3_U2979) );
  INV_X1 U21646 ( .A(n18544), .ZN(n18539) );
  NOR2_X1 U21647 ( .A1(n9706), .A2(n18539), .ZN(n18565) );
  AOI22_X1 U21648 ( .A1(n18573), .A2(n18607), .B1(n18572), .B2(n18565), .ZN(
        n18546) );
  INV_X1 U21649 ( .A(n18540), .ZN(n18542) );
  OAI221_X1 U21650 ( .B1(n18544), .B2(n18543), .C1(n18544), .C2(n18542), .A(
        n18541), .ZN(n18567) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18567), .B1(
        n18578), .B2(n18566), .ZN(n18545) );
  OAI211_X1 U21652 ( .C1(n18581), .C2(n18570), .A(n18546), .B(n18545), .ZN(
        P3_U2980) );
  AOI22_X1 U21653 ( .A1(n18583), .A2(n18555), .B1(n18582), .B2(n18565), .ZN(
        n18548) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18567), .B1(
        n18584), .B2(n18607), .ZN(n18547) );
  OAI211_X1 U21655 ( .C1(n18558), .C2(n18587), .A(n18548), .B(n18547), .ZN(
        P3_U2981) );
  AOI22_X1 U21656 ( .A1(n18588), .A2(n18565), .B1(n18589), .B2(n18607), .ZN(
        n18550) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18567), .B1(
        n18566), .B2(n18590), .ZN(n18549) );
  OAI211_X1 U21658 ( .C1(n18593), .C2(n18570), .A(n18550), .B(n18549), .ZN(
        P3_U2982) );
  AOI22_X1 U21659 ( .A1(n18596), .A2(n18607), .B1(n18594), .B2(n18565), .ZN(
        n18553) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18567), .B1(
        n18566), .B2(n18551), .ZN(n18552) );
  OAI211_X1 U21661 ( .C1(n18554), .C2(n18570), .A(n18553), .B(n18552), .ZN(
        P3_U2983) );
  AOI22_X1 U21662 ( .A1(n18601), .A2(n18555), .B1(n18600), .B2(n18565), .ZN(
        n18557) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18567), .B1(
        n18602), .B2(n18607), .ZN(n18556) );
  OAI211_X1 U21664 ( .C1(n18558), .C2(n18605), .A(n18557), .B(n18556), .ZN(
        P3_U2984) );
  AOI22_X1 U21665 ( .A1(n18609), .A2(n18607), .B1(n18606), .B2(n18565), .ZN(
        n18561) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18567), .B1(
        n18566), .B2(n18559), .ZN(n18560) );
  OAI211_X1 U21667 ( .C1(n18562), .C2(n18570), .A(n18561), .B(n18560), .ZN(
        P3_U2985) );
  AOI22_X1 U21668 ( .A1(n18615), .A2(n18607), .B1(n18614), .B2(n18565), .ZN(
        n18564) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18567), .B1(
        n18566), .B2(n18616), .ZN(n18563) );
  OAI211_X1 U21670 ( .C1(n18619), .C2(n18570), .A(n18564), .B(n18563), .ZN(
        P3_U2986) );
  AOI22_X1 U21671 ( .A1(n18622), .A2(n18607), .B1(n18621), .B2(n18565), .ZN(
        n18569) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18567), .B1(
        n18566), .B2(n18624), .ZN(n18568) );
  OAI211_X1 U21673 ( .C1(n18630), .C2(n18570), .A(n18569), .B(n18568), .ZN(
        P3_U2987) );
  INV_X1 U21674 ( .A(n18574), .ZN(n18571) );
  NOR2_X1 U21675 ( .A1(n9706), .A2(n18571), .ZN(n18620) );
  AOI22_X1 U21676 ( .A1(n18623), .A2(n18573), .B1(n18572), .B2(n18620), .ZN(
        n18580) );
  AOI22_X1 U21677 ( .A1(n18577), .A2(n18576), .B1(n18575), .B2(n18574), .ZN(
        n18626) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n18578), .ZN(n18579) );
  OAI211_X1 U21679 ( .C1(n18581), .C2(n18629), .A(n18580), .B(n18579), .ZN(
        P3_U2988) );
  AOI22_X1 U21680 ( .A1(n18583), .A2(n18607), .B1(n18582), .B2(n18620), .ZN(
        n18586) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18626), .B1(
        n18623), .B2(n18584), .ZN(n18585) );
  OAI211_X1 U21682 ( .C1(n18613), .C2(n18587), .A(n18586), .B(n18585), .ZN(
        P3_U2989) );
  AOI22_X1 U21683 ( .A1(n18623), .A2(n18589), .B1(n18588), .B2(n18620), .ZN(
        n18592) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n18590), .ZN(n18591) );
  OAI211_X1 U21685 ( .C1(n18593), .C2(n18629), .A(n18592), .B(n18591), .ZN(
        P3_U2990) );
  AOI22_X1 U21686 ( .A1(n18595), .A2(n18607), .B1(n18594), .B2(n18620), .ZN(
        n18598) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18626), .B1(
        n18623), .B2(n18596), .ZN(n18597) );
  OAI211_X1 U21688 ( .C1(n18613), .C2(n18599), .A(n18598), .B(n18597), .ZN(
        P3_U2991) );
  AOI22_X1 U21689 ( .A1(n18601), .A2(n18607), .B1(n18600), .B2(n18620), .ZN(
        n18604) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18626), .B1(
        n18623), .B2(n18602), .ZN(n18603) );
  OAI211_X1 U21691 ( .C1(n18613), .C2(n18605), .A(n18604), .B(n18603), .ZN(
        P3_U2992) );
  AOI22_X1 U21692 ( .A1(n18608), .A2(n18607), .B1(n18606), .B2(n18620), .ZN(
        n18611) );
  AOI22_X1 U21693 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18626), .B1(
        n18623), .B2(n18609), .ZN(n18610) );
  OAI211_X1 U21694 ( .C1(n18613), .C2(n18612), .A(n18611), .B(n18610), .ZN(
        P3_U2993) );
  AOI22_X1 U21695 ( .A1(n18623), .A2(n18615), .B1(n18614), .B2(n18620), .ZN(
        n18618) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n18616), .ZN(n18617) );
  OAI211_X1 U21697 ( .C1(n18619), .C2(n18629), .A(n18618), .B(n18617), .ZN(
        P3_U2994) );
  AOI22_X1 U21698 ( .A1(n18623), .A2(n18622), .B1(n18621), .B2(n18620), .ZN(
        n18628) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n18624), .ZN(n18627) );
  OAI211_X1 U21700 ( .C1(n18630), .C2(n18629), .A(n18628), .B(n18627), .ZN(
        P3_U2995) );
  NOR2_X1 U21701 ( .A1(n18632), .A2(n18631), .ZN(n18636) );
  NOR2_X1 U21702 ( .A1(n18664), .A2(n18633), .ZN(n18634) );
  OAI222_X1 U21703 ( .A1(n18639), .A2(n18638), .B1(n18637), .B2(n18636), .C1(
        n18635), .C2(n18634), .ZN(n18844) );
  OAI21_X1 U21704 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n18640), .ZN(n18642) );
  OAI211_X1 U21705 ( .C1(n18665), .C2(n18643), .A(n18642), .B(n18641), .ZN(
        n18686) );
  INV_X1 U21706 ( .A(n18665), .ZN(n18675) );
  OAI21_X1 U21707 ( .B1(n18646), .B2(n18645), .A(n18644), .ZN(n18659) );
  AOI21_X1 U21708 ( .B1(n18648), .B2(n18647), .A(n18652), .ZN(n18649) );
  AOI211_X1 U21709 ( .C1(n18659), .C2(n18650), .A(n18649), .B(n18807), .ZN(
        n18655) );
  OAI21_X1 U21710 ( .B1(n18651), .B2(n18831), .A(n18668), .ZN(n18656) );
  AOI22_X1 U21711 ( .A1(n18664), .A2(n18654), .B1(n18652), .B2(n18656), .ZN(
        n18653) );
  AOI22_X1 U21712 ( .A1(n18655), .A2(n18654), .B1(n18653), .B2(n18807), .ZN(
        n18805) );
  AOI22_X1 U21713 ( .A1(n18675), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18805), .B2(n18665), .ZN(n18684) );
  INV_X1 U21714 ( .A(n18656), .ZN(n18669) );
  NOR2_X1 U21715 ( .A1(n18825), .A2(n18669), .ZN(n18662) );
  OAI221_X1 U21716 ( .B1(n18659), .B2(n18825), .C1(n18659), .C2(n18658), .A(
        n18657), .ZN(n18660) );
  INV_X1 U21717 ( .A(n18660), .ZN(n18661) );
  MUX2_X1 U21718 ( .A(n18662), .B(n18661), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n18663) );
  AOI21_X1 U21719 ( .B1(n18664), .B2(n18811), .A(n18663), .ZN(n18814) );
  AOI22_X1 U21720 ( .A1(n18675), .A2(n18817), .B1(n18814), .B2(n18665), .ZN(
        n18679) );
  NOR2_X1 U21721 ( .A1(n18667), .A2(n18666), .ZN(n18670) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18668), .B1(
        n18670), .B2(n18831), .ZN(n18827) );
  OAI22_X1 U21723 ( .A1(n18670), .A2(n18818), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18669), .ZN(n18823) );
  AOI222_X1 U21724 ( .A1(n18827), .A2(n18823), .B1(n18827), .B2(n18672), .C1(
        n18823), .C2(n18671), .ZN(n18674) );
  OAI21_X1 U21725 ( .B1(n18675), .B2(n18674), .A(n18673), .ZN(n18678) );
  AND2_X1 U21726 ( .A1(n18679), .A2(n18678), .ZN(n18676) );
  OAI221_X1 U21727 ( .B1(n18679), .B2(n18678), .C1(n18677), .C2(n18676), .A(
        n18681), .ZN(n18683) );
  AOI21_X1 U21728 ( .B1(n18681), .B2(n18680), .A(n18679), .ZN(n18682) );
  AOI222_X1 U21729 ( .A1(n18684), .A2(n18683), .B1(n18684), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18683), .C2(n18682), .ZN(
        n18685) );
  NOR4_X1 U21730 ( .A1(n18687), .A2(n18844), .A3(n18686), .A4(n18685), .ZN(
        n18698) );
  AOI22_X1 U21731 ( .A1(n18826), .A2(n18853), .B1(n18722), .B2(n17449), .ZN(
        n18688) );
  INV_X1 U21732 ( .A(n18688), .ZN(n18694) );
  INV_X1 U21733 ( .A(n18689), .ZN(n18690) );
  OAI211_X1 U21734 ( .C1(n18691), .C2(n18690), .A(n18846), .B(n18698), .ZN(
        n18802) );
  OAI21_X1 U21735 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18851), .A(n18802), 
        .ZN(n18699) );
  NOR2_X1 U21736 ( .A1(n18692), .A2(n18699), .ZN(n18693) );
  MUX2_X1 U21737 ( .A(n18694), .B(n18693), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18696) );
  OAI211_X1 U21738 ( .C1(n18698), .C2(n18697), .A(n18696), .B(n18695), .ZN(
        P3_U2996) );
  NAND2_X1 U21739 ( .A1(n18722), .A2(n17449), .ZN(n18703) );
  NAND4_X1 U21740 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18722), .A4(n18862), .ZN(n18705) );
  OR3_X1 U21741 ( .A1(n9706), .A2(n18700), .A3(n18699), .ZN(n18702) );
  NAND4_X1 U21742 ( .A1(n18704), .A2(n18703), .A3(n18705), .A4(n18702), .ZN(
        P3_U2997) );
  INV_X1 U21743 ( .A(n18705), .ZN(n18707) );
  INV_X1 U21744 ( .A(n18801), .ZN(n18706) );
  NOR4_X1 U21745 ( .A1(n18853), .A2(n18708), .A3(n18707), .A4(n18706), .ZN(
        P3_U2998) );
  AND2_X1 U21746 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18713), .ZN(
        P3_U2999) );
  AND2_X1 U21747 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18713), .ZN(
        P3_U3000) );
  NOR2_X1 U21748 ( .A1(n18709), .A2(n18800), .ZN(P3_U3001) );
  AND2_X1 U21749 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18713), .ZN(
        P3_U3002) );
  AND2_X1 U21750 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18713), .ZN(
        P3_U3003) );
  AND2_X1 U21751 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18713), .ZN(
        P3_U3004) );
  NOR2_X1 U21752 ( .A1(n18710), .A2(n18800), .ZN(P3_U3005) );
  AND2_X1 U21753 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18713), .ZN(
        P3_U3006) );
  AND2_X1 U21754 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18713), .ZN(
        P3_U3007) );
  AND2_X1 U21755 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18713), .ZN(
        P3_U3008) );
  AND2_X1 U21756 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18713), .ZN(
        P3_U3009) );
  AND2_X1 U21757 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18713), .ZN(
        P3_U3010) );
  AND2_X1 U21758 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18713), .ZN(
        P3_U3011) );
  AND2_X1 U21759 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18713), .ZN(
        P3_U3012) );
  AND2_X1 U21760 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18713), .ZN(
        P3_U3013) );
  AND2_X1 U21761 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18713), .ZN(
        P3_U3014) );
  AND2_X1 U21762 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18713), .ZN(
        P3_U3015) );
  AND2_X1 U21763 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18711), .ZN(
        P3_U3016) );
  AND2_X1 U21764 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18711), .ZN(
        P3_U3017) );
  AND2_X1 U21765 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18711), .ZN(
        P3_U3018) );
  AND2_X1 U21766 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18711), .ZN(
        P3_U3019) );
  AND2_X1 U21767 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18711), .ZN(
        P3_U3020) );
  AND2_X1 U21768 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18711), .ZN(P3_U3021) );
  AND2_X1 U21769 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18713), .ZN(P3_U3022) );
  AND2_X1 U21770 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18713), .ZN(P3_U3023) );
  AND2_X1 U21771 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18713), .ZN(P3_U3024) );
  AND2_X1 U21772 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18713), .ZN(P3_U3025) );
  NOR2_X1 U21773 ( .A1(n18712), .A2(n18800), .ZN(P3_U3026) );
  AND2_X1 U21774 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18713), .ZN(P3_U3027) );
  AND2_X1 U21775 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18713), .ZN(P3_U3028) );
  INV_X1 U21776 ( .A(n18719), .ZN(n18718) );
  OAI21_X1 U21777 ( .B1(n18714), .B2(n20773), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18715) );
  AOI22_X1 U21778 ( .A1(n18728), .A2(n18730), .B1(n18841), .B2(n18715), .ZN(
        n18717) );
  NAND3_X1 U21779 ( .A1(NA), .A2(n18728), .A3(n18716), .ZN(n18721) );
  OAI211_X1 U21780 ( .C1(n18851), .C2(n18718), .A(n18717), .B(n18721), .ZN(
        P3_U3029) );
  NAND2_X1 U21781 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n18723) );
  AOI22_X1 U21782 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18723), .B1(HOLD), 
        .B2(n18719), .ZN(n18720) );
  NAND2_X1 U21783 ( .A1(n18722), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18724) );
  OAI211_X1 U21784 ( .C1(n18720), .C2(n18728), .A(n18724), .B(n18848), .ZN(
        P3_U3030) );
  AOI22_X1 U21785 ( .A1(n18722), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18728), 
        .B2(n18721), .ZN(n18729) );
  INV_X1 U21786 ( .A(n18723), .ZN(n18726) );
  OAI22_X1 U21787 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18724), .ZN(n18725) );
  OAI22_X1 U21788 ( .A1(n18726), .A2(n18725), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18727) );
  OAI22_X1 U21789 ( .A1(n18729), .A2(n18730), .B1(n18728), .B2(n18727), .ZN(
        P3_U3031) );
  INV_X1 U21790 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18733) );
  NAND2_X1 U21791 ( .A1(n18788), .A2(n18730), .ZN(n18790) );
  OAI222_X1 U21792 ( .A1(n18839), .A2(n18795), .B1(n18731), .B2(n18788), .C1(
        n18733), .C2(n18791), .ZN(P3_U3032) );
  OAI222_X1 U21793 ( .A1(n18733), .A2(n18795), .B1(n18732), .B2(n18788), .C1(
        n18735), .C2(n18791), .ZN(P3_U3033) );
  OAI222_X1 U21794 ( .A1(n18735), .A2(n18795), .B1(n18734), .B2(n18788), .C1(
        n18737), .C2(n18791), .ZN(P3_U3034) );
  OAI222_X1 U21795 ( .A1(n18737), .A2(n18795), .B1(n18736), .B2(n18788), .C1(
        n18739), .C2(n18791), .ZN(P3_U3035) );
  OAI222_X1 U21796 ( .A1(n18739), .A2(n18795), .B1(n18738), .B2(n18788), .C1(
        n18741), .C2(n18791), .ZN(P3_U3036) );
  OAI222_X1 U21797 ( .A1(n18741), .A2(n18795), .B1(n18740), .B2(n18788), .C1(
        n18743), .C2(n18791), .ZN(P3_U3037) );
  OAI222_X1 U21798 ( .A1(n18743), .A2(n18795), .B1(n18742), .B2(n18788), .C1(
        n18745), .C2(n18791), .ZN(P3_U3038) );
  OAI222_X1 U21799 ( .A1(n18745), .A2(n18795), .B1(n18744), .B2(n18788), .C1(
        n18747), .C2(n18791), .ZN(P3_U3039) );
  OAI222_X1 U21800 ( .A1(n18747), .A2(n18786), .B1(n18746), .B2(n18788), .C1(
        n18749), .C2(n18791), .ZN(P3_U3040) );
  OAI222_X1 U21801 ( .A1(n18749), .A2(n18786), .B1(n18748), .B2(n18788), .C1(
        n18751), .C2(n18791), .ZN(P3_U3041) );
  INV_X1 U21802 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18753) );
  OAI222_X1 U21803 ( .A1(n18751), .A2(n18786), .B1(n18750), .B2(n18788), .C1(
        n18753), .C2(n18791), .ZN(P3_U3042) );
  OAI222_X1 U21804 ( .A1(n18753), .A2(n18786), .B1(n18752), .B2(n18788), .C1(
        n18755), .C2(n18791), .ZN(P3_U3043) );
  INV_X1 U21805 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18757) );
  OAI222_X1 U21806 ( .A1(n18755), .A2(n18786), .B1(n18754), .B2(n18788), .C1(
        n18757), .C2(n18790), .ZN(P3_U3044) );
  OAI222_X1 U21807 ( .A1(n18757), .A2(n18786), .B1(n18756), .B2(n18788), .C1(
        n18758), .C2(n18790), .ZN(P3_U3045) );
  OAI222_X1 U21808 ( .A1(n18790), .A2(n18761), .B1(n18759), .B2(n18788), .C1(
        n18758), .C2(n18786), .ZN(P3_U3046) );
  OAI222_X1 U21809 ( .A1(n18761), .A2(n18786), .B1(n18760), .B2(n18788), .C1(
        n18763), .C2(n18790), .ZN(P3_U3047) );
  OAI222_X1 U21810 ( .A1(n18763), .A2(n18786), .B1(n18762), .B2(n18788), .C1(
        n18764), .C2(n18791), .ZN(P3_U3048) );
  OAI222_X1 U21811 ( .A1(n18790), .A2(n18766), .B1(n18765), .B2(n18788), .C1(
        n18764), .C2(n18786), .ZN(P3_U3049) );
  INV_X1 U21812 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18769) );
  OAI222_X1 U21813 ( .A1(n18791), .A2(n18769), .B1(n18767), .B2(n18788), .C1(
        n18766), .C2(n18786), .ZN(P3_U3050) );
  OAI222_X1 U21814 ( .A1(n18769), .A2(n18786), .B1(n18768), .B2(n18788), .C1(
        n18771), .C2(n18791), .ZN(P3_U3051) );
  OAI222_X1 U21815 ( .A1(n18771), .A2(n18786), .B1(n18770), .B2(n18788), .C1(
        n18772), .C2(n18791), .ZN(P3_U3052) );
  OAI222_X1 U21816 ( .A1(n18790), .A2(n18774), .B1(n18773), .B2(n18788), .C1(
        n18772), .C2(n18786), .ZN(P3_U3053) );
  OAI222_X1 U21817 ( .A1(n18791), .A2(n18776), .B1(n18775), .B2(n18788), .C1(
        n18774), .C2(n18786), .ZN(P3_U3054) );
  OAI222_X1 U21818 ( .A1(n18791), .A2(n18778), .B1(n18777), .B2(n18788), .C1(
        n18776), .C2(n18786), .ZN(P3_U3055) );
  OAI222_X1 U21819 ( .A1(n18790), .A2(n18780), .B1(n18779), .B2(n18788), .C1(
        n18778), .C2(n18786), .ZN(P3_U3056) );
  OAI222_X1 U21820 ( .A1(n18790), .A2(n18782), .B1(n18781), .B2(n18788), .C1(
        n18780), .C2(n18786), .ZN(P3_U3057) );
  OAI222_X1 U21821 ( .A1(n18790), .A2(n18785), .B1(n18783), .B2(n18788), .C1(
        n18782), .C2(n18786), .ZN(P3_U3058) );
  OAI222_X1 U21822 ( .A1(n18785), .A2(n18786), .B1(n18784), .B2(n18788), .C1(
        n18787), .C2(n18791), .ZN(P3_U3059) );
  OAI222_X1 U21823 ( .A1(n18790), .A2(n18794), .B1(n18789), .B2(n18788), .C1(
        n18787), .C2(n18786), .ZN(P3_U3060) );
  OAI222_X1 U21824 ( .A1(n18795), .A2(n18794), .B1(n18793), .B2(n18788), .C1(
        n18792), .C2(n18791), .ZN(P3_U3061) );
  MUX2_X1 U21825 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n18788), .Z(P3_U3274) );
  MUX2_X1 U21826 ( .A(P3_BE_N_REG_2__SCAN_IN), .B(P3_BYTEENABLE_REG_2__SCAN_IN), .S(n18788), .Z(P3_U3275) );
  MUX2_X1 U21827 ( .A(P3_BE_N_REG_1__SCAN_IN), .B(P3_BYTEENABLE_REG_1__SCAN_IN), .S(n18788), .Z(P3_U3276) );
  OAI22_X1 U21828 ( .A1(n18841), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18788), .ZN(n18796) );
  INV_X1 U21829 ( .A(n18796), .ZN(P3_U3277) );
  OAI21_X1 U21830 ( .B1(n18800), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18798), 
        .ZN(n18797) );
  INV_X1 U21831 ( .A(n18797), .ZN(P3_U3280) );
  OAI21_X1 U21832 ( .B1(n18800), .B2(n18799), .A(n18798), .ZN(P3_U3281) );
  OAI221_X1 U21833 ( .B1(n18803), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18803), 
        .C2(n18802), .A(n18801), .ZN(P3_U3282) );
  AOI22_X1 U21834 ( .A1(n18863), .A2(n18805), .B1(n18826), .B2(n18804), .ZN(
        n18806) );
  INV_X1 U21835 ( .A(n18832), .ZN(n18829) );
  AOI22_X1 U21836 ( .A1(n18832), .A2(n18807), .B1(n18806), .B2(n18829), .ZN(
        P3_U3285) );
  AOI22_X1 U21837 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18809), .B2(n18808), .ZN(
        n18819) );
  NOR2_X1 U21838 ( .A1(n18810), .A2(n18828), .ZN(n18820) );
  OAI22_X1 U21839 ( .A1(n18814), .A2(n18813), .B1(n18812), .B2(n18811), .ZN(
        n18815) );
  AOI21_X1 U21840 ( .B1(n18819), .B2(n18820), .A(n18815), .ZN(n18816) );
  AOI22_X1 U21841 ( .A1(n18832), .A2(n18817), .B1(n18816), .B2(n18829), .ZN(
        P3_U3288) );
  INV_X1 U21842 ( .A(n18818), .ZN(n18822) );
  INV_X1 U21843 ( .A(n18819), .ZN(n18821) );
  AOI222_X1 U21844 ( .A1(n18823), .A2(n18863), .B1(n18826), .B2(n18822), .C1(
        n18821), .C2(n18820), .ZN(n18824) );
  AOI22_X1 U21845 ( .A1(n18832), .A2(n18825), .B1(n18824), .B2(n18829), .ZN(
        P3_U3289) );
  AOI222_X1 U21846 ( .A1(n18828), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18863), 
        .B2(n18827), .C1(n18831), .C2(n18826), .ZN(n18830) );
  AOI22_X1 U21847 ( .A1(n18832), .A2(n18831), .B1(n18830), .B2(n18829), .ZN(
        P3_U3290) );
  AOI21_X1 U21848 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18833) );
  OAI22_X1 U21849 ( .A1(n18834), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(n18833), .B2(n18836), .ZN(n18835) );
  AOI21_X1 U21850 ( .B1(n18840), .B2(n18836), .A(n18835), .ZN(P3_U3292) );
  INV_X1 U21851 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18837) );
  AOI22_X1 U21852 ( .A1(n18840), .A2(n18839), .B1(n18838), .B2(n18837), .ZN(
        P3_U3293) );
  INV_X1 U21853 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18842) );
  AOI22_X1 U21854 ( .A1(n18788), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18842), 
        .B2(n18841), .ZN(P3_U3294) );
  MUX2_X1 U21855 ( .A(P3_MORE_REG_SCAN_IN), .B(n18844), .S(n18843), .Z(
        P3_U3295) );
  OAI21_X1 U21856 ( .B1(n18846), .B2(n18845), .A(n18859), .ZN(n18847) );
  AOI21_X1 U21857 ( .B1(n17449), .B2(n18851), .A(n18847), .ZN(n18857) );
  AOI21_X1 U21858 ( .B1(n18850), .B2(n18849), .A(n18848), .ZN(n18852) );
  OAI211_X1 U21859 ( .C1(n18858), .C2(n18852), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18851), .ZN(n18854) );
  AOI21_X1 U21860 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18854), .A(n18853), 
        .ZN(n18856) );
  NAND2_X1 U21861 ( .A1(n18857), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18855) );
  OAI21_X1 U21862 ( .B1(n18857), .B2(n18856), .A(n18855), .ZN(P3_U3296) );
  MUX2_X1 U21863 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n18788), .Z(P3_U3297) );
  INV_X1 U21864 ( .A(n18859), .ZN(n18866) );
  INV_X1 U21865 ( .A(n18858), .ZN(n18861) );
  AOI21_X1 U21866 ( .B1(n18863), .B2(n18862), .A(P3_READREQUEST_REG_SCAN_IN), 
        .ZN(n18860) );
  AOI22_X1 U21867 ( .A1(n18866), .A2(n18861), .B1(n18860), .B2(n18859), .ZN(
        P3_U3298) );
  AOI21_X1 U21868 ( .B1(n18863), .B2(n18862), .A(P3_MEMORYFETCH_REG_SCAN_IN), 
        .ZN(n18865) );
  OAI21_X1 U21869 ( .B1(n18866), .B2(n18865), .A(n18864), .ZN(P3_U3299) );
  INV_X1 U21870 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19835) );
  INV_X1 U21871 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18867) );
  NAND2_X1 U21872 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19852), .ZN(n19843) );
  NAND2_X1 U21873 ( .A1(n19835), .A2(n18871), .ZN(n19840) );
  OAI21_X1 U21874 ( .B1(n19835), .B2(n19843), .A(n19840), .ZN(n19911) );
  OAI21_X1 U21875 ( .B1(n19835), .B2(n18867), .A(n19834), .ZN(P2_U2815) );
  INV_X1 U21876 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18869) );
  OAI22_X1 U21877 ( .A1(n18870), .A2(n18869), .B1(n19969), .B2(n18868), .ZN(
        P2_U2816) );
  OR2_X1 U21878 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n18871), .ZN(n19982) );
  INV_X2 U21879 ( .A(n19982), .ZN(n19985) );
  AOI21_X1 U21880 ( .B1(n19835), .B2(n19852), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18872) );
  AOI22_X1 U21881 ( .A1(n19985), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18872), 
        .B2(n19982), .ZN(P2_U2817) );
  OAI21_X1 U21882 ( .B1(n19837), .B2(BS16), .A(n19911), .ZN(n19909) );
  OAI21_X1 U21883 ( .B1(n19911), .B2(n19914), .A(n19909), .ZN(P2_U2818) );
  NOR2_X1 U21884 ( .A1(n18874), .A2(n18873), .ZN(n19953) );
  OAI21_X1 U21885 ( .B1(n19953), .B2(n18876), .A(n18875), .ZN(P2_U2819) );
  AOI211_X1 U21886 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_9__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18877) );
  AND4_X1 U21887 ( .A1(n18878), .A2(n18877), .A3(n19829), .A4(n19830), .ZN(
        n18886) );
  NOR4_X1 U21888 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_10__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n18885) );
  NOR4_X1 U21889 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18884) );
  NOR4_X1 U21890 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_18__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_20__SCAN_IN), .ZN(n18882) );
  NOR4_X1 U21891 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_14__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n18881) );
  NOR4_X1 U21892 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_27__SCAN_IN), .A3(P2_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18880) );
  NOR4_X1 U21893 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_23__SCAN_IN), .A3(P2_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_25__SCAN_IN), .ZN(n18879) );
  AND4_X1 U21894 ( .A1(n18882), .A2(n18881), .A3(n18880), .A4(n18879), .ZN(
        n18883) );
  NAND4_X1 U21895 ( .A1(n18886), .A2(n18885), .A3(n18884), .A4(n18883), .ZN(
        n18893) );
  NOR2_X1 U21896 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18893), .ZN(n18887) );
  INV_X1 U21897 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U21898 ( .A1(n18887), .A2(n18888), .B1(n18893), .B2(n19907), .ZN(
        P2_U2820) );
  OR3_X1 U21899 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18892) );
  INV_X1 U21900 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U21901 ( .A1(n18887), .A2(n18892), .B1(n18893), .B2(n19905), .ZN(
        P2_U2821) );
  INV_X1 U21902 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19910) );
  NAND2_X1 U21903 ( .A1(n18887), .A2(n19910), .ZN(n18891) );
  INV_X1 U21904 ( .A(n18893), .ZN(n18894) );
  OAI21_X1 U21905 ( .B1(n19853), .B2(n18888), .A(n18894), .ZN(n18889) );
  OAI21_X1 U21906 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18894), .A(n18889), 
        .ZN(n18890) );
  OAI221_X1 U21907 ( .B1(n18891), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18891), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18890), .ZN(P2_U2822) );
  INV_X1 U21908 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19903) );
  OAI221_X1 U21909 ( .B1(n18894), .B2(n19903), .C1(n18893), .C2(n18892), .A(
        n18891), .ZN(P2_U2823) );
  NAND2_X1 U21910 ( .A1(n9716), .A2(n18895), .ZN(n18896) );
  XOR2_X1 U21911 ( .A(n18897), .B(n18896), .Z(n18906) );
  AOI22_X1 U21912 ( .A1(n18898), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n9707), .ZN(n18899) );
  OAI211_X1 U21913 ( .C1(n19880), .C2(n19034), .A(n18899), .B(n9722), .ZN(
        n18900) );
  AOI21_X1 U21914 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19058), .A(n18900), .ZN(
        n18905) );
  INV_X1 U21915 ( .A(n18901), .ZN(n18903) );
  AOI22_X1 U21916 ( .A1(n18903), .A2(n19093), .B1(n18902), .B2(n19019), .ZN(
        n18904) );
  OAI211_X1 U21917 ( .C1(n19825), .C2(n18906), .A(n18905), .B(n18904), .ZN(
        P2_U2836) );
  NOR2_X1 U21918 ( .A1(n19069), .A2(n18907), .ZN(n18909) );
  XOR2_X1 U21919 ( .A(n18909), .B(n18908), .Z(n18917) );
  AOI22_X1 U21920 ( .A1(n18910), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n9707), .ZN(n18911) );
  OAI211_X1 U21921 ( .C1(n12405), .C2(n19034), .A(n18911), .B(n9722), .ZN(
        n18912) );
  AOI21_X1 U21922 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n19058), .A(n18912), .ZN(
        n18916) );
  AOI22_X1 U21923 ( .A1(n18914), .A2(n19093), .B1(n18913), .B2(n19019), .ZN(
        n18915) );
  OAI211_X1 U21924 ( .C1(n19825), .C2(n18917), .A(n18916), .B(n18915), .ZN(
        P2_U2837) );
  NAND2_X1 U21925 ( .A1(n9715), .A2(n18918), .ZN(n18919) );
  XOR2_X1 U21926 ( .A(n18920), .B(n18919), .Z(n18929) );
  OAI21_X1 U21927 ( .B1(n19877), .B2(n19034), .A(n9722), .ZN(n18924) );
  OAI22_X1 U21928 ( .A1(n18922), .A2(n19063), .B1(n18921), .B2(n19079), .ZN(
        n18923) );
  AOI211_X1 U21929 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19058), .A(n18924), .B(
        n18923), .ZN(n18928) );
  AOI22_X1 U21930 ( .A1(n18926), .A2(n19019), .B1(n18925), .B2(n19093), .ZN(
        n18927) );
  OAI211_X1 U21931 ( .C1(n19825), .C2(n18929), .A(n18928), .B(n18927), .ZN(
        P2_U2838) );
  INV_X1 U21932 ( .A(n18930), .ZN(n18932) );
  AOI22_X1 U21933 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n9707), .B1(
        P2_EBX_REG_16__SCAN_IN), .B2(n19058), .ZN(n18931) );
  OAI21_X1 U21934 ( .B1(n18932), .B2(n19063), .A(n18931), .ZN(n18933) );
  AOI211_X1 U21935 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19081), .A(n15077), 
        .B(n18933), .ZN(n18938) );
  NOR2_X1 U21936 ( .A1(n19069), .A2(n18934), .ZN(n18951) );
  XNOR2_X1 U21937 ( .A(n18951), .B(n18935), .ZN(n18936) );
  AOI22_X1 U21938 ( .A1(n19109), .A2(n19019), .B1(n19055), .B2(n18936), .ZN(
        n18937) );
  OAI211_X1 U21939 ( .C1(n18939), .C2(n19075), .A(n18938), .B(n18937), .ZN(
        P2_U2839) );
  OAI21_X1 U21940 ( .B1(n19034), .B2(n18940), .A(n9722), .ZN(n18943) );
  OAI22_X1 U21941 ( .A1(n19091), .A2(n11143), .B1(n18941), .B2(n19079), .ZN(
        n18942) );
  AOI211_X1 U21942 ( .C1(n19086), .C2(n18944), .A(n18943), .B(n18942), .ZN(
        n18945) );
  INV_X1 U21943 ( .A(n18945), .ZN(n18946) );
  AOI21_X1 U21944 ( .B1(n18949), .B2(n18947), .A(n18946), .ZN(n18954) );
  AOI21_X1 U21945 ( .B1(n18949), .B2(n18948), .A(n19825), .ZN(n18950) );
  AOI22_X1 U21946 ( .A1(n18952), .A2(n19093), .B1(n18951), .B2(n18950), .ZN(
        n18953) );
  OAI211_X1 U21947 ( .C1(n19115), .C2(n19083), .A(n18954), .B(n18953), .ZN(
        P2_U2840) );
  INV_X1 U21948 ( .A(n18955), .ZN(n18960) );
  INV_X1 U21949 ( .A(n18962), .ZN(n18956) );
  OAI211_X1 U21950 ( .C1(n19069), .C2(n18957), .A(n18956), .B(n19055), .ZN(
        n18959) );
  AOI22_X1 U21951 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n9707), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19058), .ZN(n18958) );
  OAI211_X1 U21952 ( .C1(n18960), .C2(n19063), .A(n18959), .B(n18958), .ZN(
        n18961) );
  AOI211_X1 U21953 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19081), .A(n15077), 
        .B(n18961), .ZN(n18965) );
  AOI22_X1 U21954 ( .A1(n19019), .A2(n19116), .B1(n18963), .B2(n18962), .ZN(
        n18964) );
  OAI211_X1 U21955 ( .C1(n18966), .C2(n19075), .A(n18965), .B(n18964), .ZN(
        P2_U2841) );
  INV_X1 U21956 ( .A(n18967), .ZN(n18968) );
  AOI22_X1 U21957 ( .A1(n18968), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9707), .ZN(n18969) );
  OAI21_X1 U21958 ( .B1(n19091), .B2(n11128), .A(n18969), .ZN(n18970) );
  AOI211_X1 U21959 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19081), .A(n15077), 
        .B(n18970), .ZN(n18976) );
  NOR2_X1 U21960 ( .A1(n19069), .A2(n18971), .ZN(n18973) );
  XNOR2_X1 U21961 ( .A(n18973), .B(n18972), .ZN(n18974) );
  AOI22_X1 U21962 ( .A1(n19120), .A2(n19019), .B1(n19055), .B2(n18974), .ZN(
        n18975) );
  OAI211_X1 U21963 ( .C1(n18977), .C2(n19075), .A(n18976), .B(n18975), .ZN(
        P2_U2843) );
  OAI21_X1 U21964 ( .B1(n11291), .B2(n19034), .A(n9722), .ZN(n18981) );
  OAI22_X1 U21965 ( .A1(n18979), .A2(n19063), .B1(n18978), .B2(n19079), .ZN(
        n18980) );
  AOI211_X1 U21966 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n19058), .A(n18981), .B(
        n18980), .ZN(n18988) );
  NAND2_X1 U21967 ( .A1(n9716), .A2(n18982), .ZN(n18983) );
  XNOR2_X1 U21968 ( .A(n18984), .B(n18983), .ZN(n18985) );
  AOI22_X1 U21969 ( .A1(n18986), .A2(n19093), .B1(n19055), .B2(n18985), .ZN(
        n18987) );
  OAI211_X1 U21970 ( .C1(n19122), .C2(n19083), .A(n18988), .B(n18987), .ZN(
        P2_U2844) );
  AOI22_X1 U21971 ( .A1(n18989), .A2(n19086), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9707), .ZN(n18990) );
  OAI21_X1 U21972 ( .B1(n19091), .B2(n18991), .A(n18990), .ZN(n18992) );
  AOI211_X1 U21973 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19081), .A(n12404), 
        .B(n18992), .ZN(n18998) );
  NOR2_X1 U21974 ( .A1(n19069), .A2(n18993), .ZN(n18995) );
  XNOR2_X1 U21975 ( .A(n18995), .B(n18994), .ZN(n18996) );
  AOI22_X1 U21976 ( .A1(n19123), .A2(n19019), .B1(n19055), .B2(n18996), .ZN(
        n18997) );
  OAI211_X1 U21977 ( .C1(n18999), .C2(n19075), .A(n18998), .B(n18997), .ZN(
        P2_U2845) );
  OAI21_X1 U21978 ( .B1(n11264), .B2(n19034), .A(n9722), .ZN(n19004) );
  INV_X1 U21979 ( .A(n19000), .ZN(n19002) );
  OAI22_X1 U21980 ( .A1(n19002), .A2(n19063), .B1(n19001), .B2(n19079), .ZN(
        n19003) );
  AOI211_X1 U21981 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19058), .A(n19004), .B(
        n19003), .ZN(n19011) );
  NAND2_X1 U21982 ( .A1(n9715), .A2(n19005), .ZN(n19006) );
  XNOR2_X1 U21983 ( .A(n19007), .B(n19006), .ZN(n19008) );
  AOI22_X1 U21984 ( .A1(n19009), .A2(n19093), .B1(n19055), .B2(n19008), .ZN(
        n19010) );
  OAI211_X1 U21985 ( .C1(n19126), .C2(n19083), .A(n19011), .B(n19010), .ZN(
        P2_U2846) );
  INV_X1 U21986 ( .A(n19012), .ZN(n19014) );
  AOI22_X1 U21987 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n9707), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19058), .ZN(n19013) );
  OAI21_X1 U21988 ( .B1(n19014), .B2(n19063), .A(n19013), .ZN(n19015) );
  AOI211_X1 U21989 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19081), .A(n12404), .B(
        n19015), .ZN(n19022) );
  NOR2_X1 U21990 ( .A1(n19069), .A2(n19016), .ZN(n19018) );
  XNOR2_X1 U21991 ( .A(n19018), .B(n19017), .ZN(n19020) );
  AOI22_X1 U21992 ( .A1(n19055), .A2(n19020), .B1(n19019), .B2(n19127), .ZN(
        n19021) );
  OAI211_X1 U21993 ( .C1(n19075), .C2(n19023), .A(n19022), .B(n19021), .ZN(
        P2_U2847) );
  NAND2_X1 U21994 ( .A1(n9715), .A2(n19024), .ZN(n19026) );
  XOR2_X1 U21995 ( .A(n19026), .B(n19025), .Z(n19033) );
  AOI22_X1 U21996 ( .A1(n19027), .A2(n19086), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19058), .ZN(n19028) );
  OAI211_X1 U21997 ( .C1(n19863), .C2(n19034), .A(n19028), .B(n9722), .ZN(
        n19031) );
  OAI22_X1 U21998 ( .A1(n19083), .A2(n19131), .B1(n19075), .B2(n19029), .ZN(
        n19030) );
  AOI211_X1 U21999 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n9707), .A(
        n19031), .B(n19030), .ZN(n19032) );
  OAI21_X1 U22000 ( .B1(n19033), .B2(n19825), .A(n19032), .ZN(P2_U2848) );
  OAI21_X1 U22001 ( .B1(n19861), .B2(n19034), .A(n9722), .ZN(n19038) );
  OAI22_X1 U22002 ( .A1(n19036), .A2(n19063), .B1(n19091), .B2(n19035), .ZN(
        n19037) );
  AOI211_X1 U22003 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n9707), .A(
        n19038), .B(n19037), .ZN(n19045) );
  NOR2_X1 U22004 ( .A1(n19069), .A2(n19039), .ZN(n19041) );
  XNOR2_X1 U22005 ( .A(n19041), .B(n19040), .ZN(n19043) );
  AOI22_X1 U22006 ( .A1(n19055), .A2(n19043), .B1(n19093), .B2(n19042), .ZN(
        n19044) );
  OAI211_X1 U22007 ( .C1(n19083), .C2(n19133), .A(n19045), .B(n19044), .ZN(
        P2_U2849) );
  AOI22_X1 U22008 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n9707), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19058), .ZN(n19047) );
  OAI21_X1 U22009 ( .B1(n19048), .B2(n19063), .A(n19047), .ZN(n19049) );
  AOI211_X1 U22010 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19081), .A(n12404), .B(
        n19049), .ZN(n19057) );
  NAND2_X1 U22011 ( .A1(n9715), .A2(n19050), .ZN(n19051) );
  XNOR2_X1 U22012 ( .A(n19052), .B(n19051), .ZN(n19054) );
  AOI22_X1 U22013 ( .A1(n19055), .A2(n19054), .B1(n19093), .B2(n19053), .ZN(
        n19056) );
  OAI211_X1 U22014 ( .C1(n19083), .C2(n19141), .A(n19057), .B(n19056), .ZN(
        P2_U2850) );
  INV_X1 U22015 ( .A(n19145), .ZN(n19067) );
  INV_X1 U22016 ( .A(n19143), .ZN(n19060) );
  AOI22_X1 U22017 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n9707), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19058), .ZN(n19059) );
  OAI211_X1 U22018 ( .C1(n19083), .C2(n19060), .A(n19059), .B(n9722), .ZN(
        n19061) );
  AOI21_X1 U22019 ( .B1(n19081), .B2(P2_REIP_REG_4__SCAN_IN), .A(n19061), .ZN(
        n19062) );
  OAI21_X1 U22020 ( .B1(n19064), .B2(n19063), .A(n19062), .ZN(n19065) );
  AOI21_X1 U22021 ( .B1(n19067), .B2(n19066), .A(n19065), .ZN(n19074) );
  INV_X1 U22022 ( .A(n19268), .ZN(n19072) );
  NOR2_X1 U22023 ( .A1(n19069), .A2(n19068), .ZN(n19071) );
  AOI21_X1 U22024 ( .B1(n19072), .B2(n19071), .A(n19825), .ZN(n19070) );
  OAI21_X1 U22025 ( .B1(n19072), .B2(n19071), .A(n19070), .ZN(n19073) );
  OAI211_X1 U22026 ( .C1(n19259), .C2(n19075), .A(n19074), .B(n19073), .ZN(
        P2_U2851) );
  INV_X1 U22027 ( .A(n19076), .ZN(n19100) );
  AOI21_X1 U22028 ( .B1(n19079), .B2(n19078), .A(n19077), .ZN(n19080) );
  AOI21_X1 U22029 ( .B1(n19081), .B2(P2_REIP_REG_0__SCAN_IN), .A(n19080), .ZN(
        n19082) );
  OAI21_X1 U22030 ( .B1(n19084), .B2(n19083), .A(n19082), .ZN(n19085) );
  INV_X1 U22031 ( .A(n19085), .ZN(n19089) );
  NAND2_X1 U22032 ( .A1(n19087), .A2(n19086), .ZN(n19088) );
  OAI211_X1 U22033 ( .C1(n19091), .C2(n19090), .A(n19089), .B(n19088), .ZN(
        n19092) );
  AOI21_X1 U22034 ( .B1(n19094), .B2(n19093), .A(n19092), .ZN(n19095) );
  OAI21_X1 U22035 ( .B1(n19945), .B2(n19096), .A(n19095), .ZN(n19097) );
  INV_X1 U22036 ( .A(n19097), .ZN(n19098) );
  OAI21_X1 U22037 ( .B1(n19100), .B2(n19099), .A(n19098), .ZN(P2_U2855) );
  AOI22_X1 U22038 ( .A1(n19101), .A2(n19158), .B1(n19107), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19103) );
  AOI22_X1 U22039 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19157), .B1(n19106), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19102) );
  NAND2_X1 U22040 ( .A1(n19103), .A2(n19102), .ZN(P2_U2888) );
  AOI22_X1 U22041 ( .A1(n19105), .A2(n19104), .B1(n19157), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19113) );
  AOI22_X1 U22042 ( .A1(n19107), .A2(BUF2_REG_16__SCAN_IN), .B1(n19106), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19112) );
  INV_X1 U22043 ( .A(n19108), .ZN(n19110) );
  AOI22_X1 U22044 ( .A1(n19110), .A2(n19146), .B1(n19158), .B2(n19109), .ZN(
        n19111) );
  NAND3_X1 U22045 ( .A1(n19113), .A2(n19112), .A3(n19111), .ZN(P2_U2903) );
  OAI222_X1 U22046 ( .A1(n19115), .A2(n19142), .B1(n19177), .B2(n19132), .C1(
        n19114), .C2(n19166), .ZN(P2_U2904) );
  INV_X1 U22047 ( .A(n19116), .ZN(n19118) );
  AOI22_X1 U22048 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19157), .B1(n19230), 
        .B2(n19134), .ZN(n19117) );
  OAI21_X1 U22049 ( .B1(n19142), .B2(n19118), .A(n19117), .ZN(P2_U2905) );
  INV_X1 U22050 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19182) );
  OAI222_X1 U22051 ( .A1(n19119), .A2(n19142), .B1(n19182), .B2(n19132), .C1(
        n19166), .C2(n19255), .ZN(P2_U2906) );
  INV_X1 U22052 ( .A(n19120), .ZN(n19121) );
  INV_X1 U22053 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19184) );
  OAI222_X1 U22054 ( .A1(n19121), .A2(n19142), .B1(n19184), .B2(n19132), .C1(
        n19166), .C2(n19252), .ZN(P2_U2907) );
  INV_X1 U22055 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19186) );
  OAI222_X1 U22056 ( .A1(n19122), .A2(n19142), .B1(n19186), .B2(n19132), .C1(
        n19166), .C2(n19250), .ZN(P2_U2908) );
  INV_X1 U22057 ( .A(n19123), .ZN(n19125) );
  AOI22_X1 U22058 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19157), .B1(n19224), 
        .B2(n19134), .ZN(n19124) );
  OAI21_X1 U22059 ( .B1(n19142), .B2(n19125), .A(n19124), .ZN(P2_U2909) );
  INV_X1 U22060 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19192) );
  OAI222_X1 U22061 ( .A1(n19126), .A2(n19142), .B1(n19192), .B2(n19132), .C1(
        n19166), .C2(n19244), .ZN(P2_U2910) );
  INV_X1 U22062 ( .A(n19127), .ZN(n19130) );
  AOI22_X1 U22063 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19157), .B1(n19128), .B2(
        n19134), .ZN(n19129) );
  OAI21_X1 U22064 ( .B1(n19142), .B2(n19130), .A(n19129), .ZN(P2_U2911) );
  OAI222_X1 U22065 ( .A1(n19131), .A2(n19142), .B1(n19196), .B2(n19132), .C1(
        n19166), .C2(n19313), .ZN(P2_U2912) );
  INV_X1 U22066 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19198) );
  OAI222_X1 U22067 ( .A1(n19133), .A2(n19142), .B1(n19198), .B2(n19132), .C1(
        n19166), .C2(n19306), .ZN(P2_U2913) );
  AOI22_X1 U22068 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19157), .B1(n19135), .B2(
        n19134), .ZN(n19140) );
  AOI21_X1 U22069 ( .B1(n19137), .B2(n19929), .A(n19136), .ZN(n19153) );
  XNOR2_X1 U22070 ( .A(n19323), .B(n19923), .ZN(n19152) );
  NOR2_X1 U22071 ( .A1(n19153), .A2(n19152), .ZN(n19151) );
  AOI21_X1 U22072 ( .B1(n19323), .B2(n19923), .A(n19151), .ZN(n19138) );
  NOR2_X1 U22073 ( .A1(n19138), .A2(n19143), .ZN(n19144) );
  OR3_X1 U22074 ( .A1(n19144), .A2(n19145), .A3(n19162), .ZN(n19139) );
  OAI211_X1 U22075 ( .C1(n19142), .C2(n19141), .A(n19140), .B(n19139), .ZN(
        P2_U2914) );
  AOI22_X1 U22076 ( .A1(n19158), .A2(n19143), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19157), .ZN(n19149) );
  XOR2_X1 U22077 ( .A(n19145), .B(n19144), .Z(n19147) );
  NAND2_X1 U22078 ( .A1(n19147), .A2(n19146), .ZN(n19148) );
  OAI211_X1 U22079 ( .C1(n19296), .C2(n19166), .A(n19149), .B(n19148), .ZN(
        P2_U2915) );
  INV_X1 U22080 ( .A(n19923), .ZN(n19150) );
  AOI22_X1 U22081 ( .A1(n19150), .A2(n19158), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19157), .ZN(n19156) );
  AOI21_X1 U22082 ( .B1(n19153), .B2(n19152), .A(n19151), .ZN(n19154) );
  OR2_X1 U22083 ( .A1(n19154), .A2(n19162), .ZN(n19155) );
  OAI211_X1 U22084 ( .C1(n19292), .C2(n19166), .A(n19156), .B(n19155), .ZN(
        P2_U2916) );
  AOI22_X1 U22085 ( .A1(n19941), .A2(n19158), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19157), .ZN(n19165) );
  AOI21_X1 U22086 ( .B1(n19161), .B2(n19160), .A(n19159), .ZN(n19163) );
  OR2_X1 U22087 ( .A1(n19163), .A2(n19162), .ZN(n19164) );
  OAI211_X1 U22088 ( .C1(n19284), .C2(n19166), .A(n19165), .B(n19164), .ZN(
        P2_U2918) );
  NOR2_X1 U22089 ( .A1(n19205), .A2(n19167), .ZN(P2_U2920) );
  INV_X1 U22090 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19170) );
  INV_X1 U22091 ( .A(n19168), .ZN(n19173) );
  AOI22_X1 U22092 ( .A1(n19173), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19212), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19169) );
  OAI21_X1 U22093 ( .B1(n19205), .B2(n19170), .A(n19169), .ZN(P2_U2921) );
  AOI22_X1 U22094 ( .A1(n19173), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n19212), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n19171) );
  OAI21_X1 U22095 ( .B1(n19172), .B2(n19205), .A(n19171), .ZN(P2_U2925) );
  AOI22_X1 U22096 ( .A1(n19173), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n19212), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n19174) );
  OAI21_X1 U22097 ( .B1(n19175), .B2(n19205), .A(n19174), .ZN(P2_U2933) );
  INV_X1 U22098 ( .A(n19203), .ZN(n19214) );
  OAI222_X1 U22099 ( .A1(n19205), .A2(n19178), .B1(n19214), .B2(n19177), .C1(
        n19966), .C2(n19176), .ZN(P2_U2936) );
  AOI22_X1 U22100 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19203), .B1(n19211), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19179) );
  OAI21_X1 U22101 ( .B1(n19180), .B2(n19966), .A(n19179), .ZN(P2_U2937) );
  AOI22_X1 U22102 ( .A1(n19212), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19181) );
  OAI21_X1 U22103 ( .B1(n19182), .B2(n19214), .A(n19181), .ZN(P2_U2938) );
  AOI22_X1 U22104 ( .A1(n19212), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19183) );
  OAI21_X1 U22105 ( .B1(n19184), .B2(n19214), .A(n19183), .ZN(P2_U2939) );
  INV_X1 U22106 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n19185) );
  OAI222_X1 U22107 ( .A1(n19205), .A2(n19187), .B1(n19214), .B2(n19186), .C1(
        n19966), .C2(n19185), .ZN(P2_U2940) );
  INV_X1 U22108 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19189) );
  OAI222_X1 U22109 ( .A1(n19205), .A2(n19190), .B1(n19214), .B2(n19189), .C1(
        n19966), .C2(n19188), .ZN(P2_U2941) );
  AOI22_X1 U22110 ( .A1(n19212), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U22111 ( .B1(n19192), .B2(n19214), .A(n19191), .ZN(P2_U2942) );
  AOI22_X1 U22112 ( .A1(n19212), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19193) );
  OAI21_X1 U22113 ( .B1(n19194), .B2(n19214), .A(n19193), .ZN(P2_U2943) );
  AOI22_X1 U22114 ( .A1(n19212), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19195) );
  OAI21_X1 U22115 ( .B1(n19196), .B2(n19214), .A(n19195), .ZN(P2_U2944) );
  AOI22_X1 U22116 ( .A1(n19212), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19197) );
  OAI21_X1 U22117 ( .B1(n19198), .B2(n19214), .A(n19197), .ZN(P2_U2945) );
  INV_X1 U22118 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19200) );
  AOI22_X1 U22119 ( .A1(n19212), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19199) );
  OAI21_X1 U22120 ( .B1(n19200), .B2(n19214), .A(n19199), .ZN(P2_U2946) );
  INV_X1 U22121 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19202) );
  AOI22_X1 U22122 ( .A1(n19212), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19201) );
  OAI21_X1 U22123 ( .B1(n19202), .B2(n19214), .A(n19201), .ZN(P2_U2947) );
  AOI22_X1 U22124 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n19203), .B1(n19212), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n19204) );
  OAI21_X1 U22125 ( .B1(n19206), .B2(n19205), .A(n19204), .ZN(P2_U2948) );
  AOI22_X1 U22126 ( .A1(n19212), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22127 ( .B1(n19208), .B2(n19214), .A(n19207), .ZN(P2_U2949) );
  AOI22_X1 U22128 ( .A1(n19212), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U22129 ( .B1(n19210), .B2(n19214), .A(n19209), .ZN(P2_U2950) );
  AOI22_X1 U22130 ( .A1(n19212), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U22131 ( .B1(n13554), .B2(n19214), .A(n19213), .ZN(P2_U2951) );
  AOI22_X1 U22132 ( .A1(n19246), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19229), .ZN(n19215) );
  OAI21_X1 U22133 ( .B1(n19234), .B2(n19254), .A(n19215), .ZN(P2_U2952) );
  AOI22_X1 U22134 ( .A1(n19246), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19245), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n19216) );
  OAI21_X1 U22135 ( .B1(n19284), .B2(n19254), .A(n19216), .ZN(P2_U2953) );
  AOI22_X1 U22136 ( .A1(n19246), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19229), .ZN(n19217) );
  OAI21_X1 U22137 ( .B1(n19237), .B2(n19254), .A(n19217), .ZN(P2_U2954) );
  AOI22_X1 U22138 ( .A1(n19246), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n19229), .ZN(n19218) );
  OAI21_X1 U22139 ( .B1(n19292), .B2(n19254), .A(n19218), .ZN(P2_U2955) );
  AOI22_X1 U22140 ( .A1(n19246), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19229), .ZN(n19219) );
  OAI21_X1 U22141 ( .B1(n19296), .B2(n19254), .A(n19219), .ZN(P2_U2956) );
  AOI22_X1 U22142 ( .A1(n19246), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19245), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n19220) );
  OAI21_X1 U22143 ( .B1(n19302), .B2(n19254), .A(n19220), .ZN(P2_U2957) );
  AOI22_X1 U22144 ( .A1(n19246), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19229), .ZN(n19221) );
  OAI21_X1 U22145 ( .B1(n19306), .B2(n19254), .A(n19221), .ZN(P2_U2958) );
  AOI22_X1 U22146 ( .A1(n19246), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19245), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n19222) );
  OAI21_X1 U22147 ( .B1(n19313), .B2(n19254), .A(n19222), .ZN(P2_U2959) );
  AOI22_X1 U22148 ( .A1(n19246), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19245), .ZN(n19223) );
  OAI21_X1 U22149 ( .B1(n19244), .B2(n19254), .A(n19223), .ZN(P2_U2961) );
  AOI22_X1 U22150 ( .A1(n19246), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n19229), .ZN(n19225) );
  NAND2_X1 U22151 ( .A1(n19231), .A2(n19224), .ZN(n19247) );
  NAND2_X1 U22152 ( .A1(n19225), .A2(n19247), .ZN(P2_U2962) );
  AOI22_X1 U22153 ( .A1(n19246), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19245), .ZN(n19226) );
  OAI21_X1 U22154 ( .B1(n19250), .B2(n19254), .A(n19226), .ZN(P2_U2963) );
  AOI22_X1 U22155 ( .A1(n19246), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19245), .ZN(n19227) );
  OAI21_X1 U22156 ( .B1(n19252), .B2(n19254), .A(n19227), .ZN(P2_U2964) );
  AOI22_X1 U22157 ( .A1(n19246), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19229), .ZN(n19228) );
  OAI21_X1 U22158 ( .B1(n19255), .B2(n19254), .A(n19228), .ZN(P2_U2965) );
  AOI22_X1 U22159 ( .A1(n19246), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19229), .ZN(n19232) );
  NAND2_X1 U22160 ( .A1(n19231), .A2(n19230), .ZN(n19256) );
  NAND2_X1 U22161 ( .A1(n19232), .A2(n19256), .ZN(P2_U2966) );
  AOI22_X1 U22162 ( .A1(n19246), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19229), .ZN(n19233) );
  OAI21_X1 U22163 ( .B1(n19234), .B2(n19254), .A(n19233), .ZN(P2_U2967) );
  AOI22_X1 U22164 ( .A1(n19246), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19245), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n19235) );
  OAI21_X1 U22165 ( .B1(n19284), .B2(n19254), .A(n19235), .ZN(P2_U2968) );
  AOI22_X1 U22166 ( .A1(n19246), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19245), .ZN(n19236) );
  OAI21_X1 U22167 ( .B1(n19237), .B2(n19254), .A(n19236), .ZN(P2_U2969) );
  AOI22_X1 U22168 ( .A1(n19246), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19229), .ZN(n19238) );
  OAI21_X1 U22169 ( .B1(n19292), .B2(n19254), .A(n19238), .ZN(P2_U2970) );
  AOI22_X1 U22170 ( .A1(n19246), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19245), .ZN(n19239) );
  OAI21_X1 U22171 ( .B1(n19296), .B2(n19254), .A(n19239), .ZN(P2_U2971) );
  AOI22_X1 U22172 ( .A1(n19246), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19245), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n19240) );
  OAI21_X1 U22173 ( .B1(n19302), .B2(n19254), .A(n19240), .ZN(P2_U2972) );
  AOI22_X1 U22174 ( .A1(n19246), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19245), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n19241) );
  OAI21_X1 U22175 ( .B1(n19306), .B2(n19254), .A(n19241), .ZN(P2_U2973) );
  AOI22_X1 U22176 ( .A1(n19246), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19245), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n19242) );
  OAI21_X1 U22177 ( .B1(n19313), .B2(n19254), .A(n19242), .ZN(P2_U2974) );
  AOI22_X1 U22178 ( .A1(n19246), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n19245), .ZN(n19243) );
  OAI21_X1 U22179 ( .B1(n19244), .B2(n19254), .A(n19243), .ZN(P2_U2976) );
  AOI22_X1 U22180 ( .A1(n19246), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19245), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n19248) );
  NAND2_X1 U22181 ( .A1(n19248), .A2(n19247), .ZN(P2_U2977) );
  AOI22_X1 U22182 ( .A1(n19246), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n19245), .ZN(n19249) );
  OAI21_X1 U22183 ( .B1(n19250), .B2(n19254), .A(n19249), .ZN(P2_U2978) );
  AOI22_X1 U22184 ( .A1(n19246), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19245), .ZN(n19251) );
  OAI21_X1 U22185 ( .B1(n19252), .B2(n19254), .A(n19251), .ZN(P2_U2979) );
  AOI22_X1 U22186 ( .A1(n19246), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19245), .ZN(n19253) );
  OAI21_X1 U22187 ( .B1(n19255), .B2(n19254), .A(n19253), .ZN(P2_U2980) );
  AOI22_X1 U22188 ( .A1(n19246), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19245), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n19257) );
  NAND2_X1 U22189 ( .A1(n19257), .A2(n19256), .ZN(P2_U2981) );
  AOI22_X1 U22190 ( .A1(n19258), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n12404), .ZN(n19267) );
  INV_X1 U22191 ( .A(n19259), .ZN(n19262) );
  AOI222_X1 U22192 ( .A1(n19265), .A2(n19264), .B1(n19263), .B2(n19262), .C1(
        n19261), .C2(n19260), .ZN(n19266) );
  OAI211_X1 U22193 ( .C1(n19269), .C2(n19268), .A(n19267), .B(n19266), .ZN(
        P2_U3010) );
  INV_X1 U22194 ( .A(n19814), .ZN(n19271) );
  NOR2_X2 U22195 ( .A1(n19562), .A2(n19419), .ZN(n19345) );
  INV_X1 U22196 ( .A(n19345), .ZN(n19270) );
  NAND2_X1 U22197 ( .A1(n19271), .A2(n19270), .ZN(n19272) );
  INV_X1 U22198 ( .A(n19934), .ZN(n19913) );
  AOI21_X1 U22199 ( .B1(n19272), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19913), 
        .ZN(n19275) );
  NOR2_X1 U22200 ( .A1(n19273), .A2(n19926), .ZN(n19809) );
  NAND2_X1 U22201 ( .A1(n19382), .A2(n19943), .ZN(n19324) );
  NOR2_X1 U22202 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19324), .ZN(
        n19312) );
  NOR2_X1 U22203 ( .A1(n19809), .A2(n19312), .ZN(n19278) );
  AOI211_X1 U22204 ( .C1(n19276), .C2(n19533), .A(n19312), .B(n19934), .ZN(
        n19274) );
  INV_X1 U22205 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19282) );
  AOI22_X1 U22206 ( .A1(n19715), .A2(n19814), .B1(n19761), .B2(n19312), .ZN(
        n19281) );
  INV_X1 U22207 ( .A(n19275), .ZN(n19279) );
  OAI21_X1 U22208 ( .B1(n19276), .B2(n19312), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19277) );
  AOI22_X1 U22209 ( .A1(n19762), .A2(n19316), .B1(n19345), .B2(n19770), .ZN(
        n19280) );
  OAI211_X1 U22210 ( .C1(n19320), .C2(n19282), .A(n19281), .B(n19280), .ZN(
        P2_U3048) );
  INV_X1 U22211 ( .A(n19779), .ZN(n19689) );
  NOR2_X2 U22212 ( .A1(n19283), .A2(n19310), .ZN(n19774) );
  AOI22_X1 U22213 ( .A1(n19689), .A2(n19814), .B1(n19774), .B2(n19312), .ZN(
        n19286) );
  NOR2_X2 U22214 ( .A1(n19284), .A2(n19357), .ZN(n19775) );
  AOI22_X1 U22215 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19314), .ZN(n19692) );
  AOI22_X1 U22216 ( .A1(n19775), .A2(n19316), .B1(n19345), .B2(n19776), .ZN(
        n19285) );
  OAI211_X1 U22217 ( .C1(n19320), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P2_U3049) );
  INV_X1 U22218 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19290) );
  AOI22_X1 U22219 ( .A1(n19732), .A2(n19814), .B1(n19780), .B2(n19312), .ZN(
        n19289) );
  AOI22_X1 U22220 ( .A1(n19781), .A2(n19316), .B1(n19345), .B2(n19782), .ZN(
        n19288) );
  OAI211_X1 U22221 ( .C1(n19320), .C2(n19290), .A(n19289), .B(n19288), .ZN(
        P2_U3050) );
  INV_X1 U22222 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19295) );
  AOI22_X1 U22223 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19314), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19315), .ZN(n19791) );
  INV_X1 U22224 ( .A(n19791), .ZN(n19736) );
  NOR2_X2 U22225 ( .A1(n19291), .A2(n19310), .ZN(n19786) );
  AOI22_X1 U22226 ( .A1(n19736), .A2(n19814), .B1(n19786), .B2(n19312), .ZN(
        n19294) );
  NOR2_X2 U22227 ( .A1(n19292), .A2(n19357), .ZN(n19787) );
  AOI22_X1 U22228 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19314), .ZN(n19739) );
  AOI22_X1 U22229 ( .A1(n19787), .A2(n19316), .B1(n19345), .B2(n19788), .ZN(
        n19293) );
  OAI211_X1 U22230 ( .C1(n19320), .C2(n19295), .A(n19294), .B(n19293), .ZN(
        P2_U3051) );
  INV_X1 U22231 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19299) );
  AOI22_X1 U22232 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19314), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19315), .ZN(n19797) );
  INV_X1 U22233 ( .A(n19797), .ZN(n19697) );
  NOR2_X2 U22234 ( .A1(n11019), .A2(n19310), .ZN(n19792) );
  AOI22_X1 U22235 ( .A1(n19697), .A2(n19814), .B1(n19792), .B2(n19312), .ZN(
        n19298) );
  NOR2_X2 U22236 ( .A1(n19296), .A2(n19357), .ZN(n19793) );
  AOI22_X1 U22237 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19314), .ZN(n19700) );
  AOI22_X1 U22238 ( .A1(n19793), .A2(n19316), .B1(n19345), .B2(n19794), .ZN(
        n19297) );
  OAI211_X1 U22239 ( .C1(n19320), .C2(n19299), .A(n19298), .B(n19297), .ZN(
        P2_U3052) );
  AOI22_X1 U22240 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19314), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19315), .ZN(n19802) );
  INV_X1 U22241 ( .A(n19802), .ZN(n19701) );
  AOI22_X1 U22242 ( .A1(n19701), .A2(n19814), .B1(n19301), .B2(n19312), .ZN(
        n19304) );
  NOR2_X2 U22243 ( .A1(n19302), .A2(n19357), .ZN(n19798) );
  AOI22_X1 U22244 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19314), .ZN(n19704) );
  AOI22_X1 U22245 ( .A1(n19798), .A2(n19316), .B1(n19345), .B2(n19799), .ZN(
        n19303) );
  OAI211_X1 U22246 ( .C1(n19320), .C2(n13782), .A(n19304), .B(n19303), .ZN(
        P2_U3053) );
  INV_X1 U22247 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19309) );
  AOI22_X1 U22248 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19314), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19315), .ZN(n19808) );
  NOR2_X2 U22249 ( .A1(n19305), .A2(n19310), .ZN(n19803) );
  AOI22_X1 U22250 ( .A1(n19746), .A2(n19814), .B1(n19803), .B2(n19312), .ZN(
        n19308) );
  NOR2_X2 U22251 ( .A1(n19306), .A2(n19357), .ZN(n19804) );
  AOI22_X1 U22252 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19314), .ZN(n19749) );
  INV_X1 U22253 ( .A(n19749), .ZN(n19805) );
  AOI22_X1 U22254 ( .A1(n19804), .A2(n19316), .B1(n19345), .B2(n19805), .ZN(
        n19307) );
  OAI211_X1 U22255 ( .C1(n19320), .C2(n19309), .A(n19308), .B(n19307), .ZN(
        P2_U3054) );
  AOI22_X1 U22256 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19314), .ZN(n19819) );
  INV_X1 U22257 ( .A(n19819), .ZN(n19752) );
  INV_X1 U22258 ( .A(n19310), .ZN(n19311) );
  AND2_X1 U22259 ( .A1(n10547), .A2(n19311), .ZN(n19810) );
  AOI22_X1 U22260 ( .A1(n19752), .A2(n19814), .B1(n19810), .B2(n19312), .ZN(
        n19318) );
  NOR2_X2 U22261 ( .A1(n19313), .A2(n19357), .ZN(n19811) );
  AOI22_X1 U22262 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19315), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19314), .ZN(n19757) );
  AOI22_X1 U22263 ( .A1(n19811), .A2(n19316), .B1(n19345), .B2(n19813), .ZN(
        n19317) );
  OAI211_X1 U22264 ( .C1(n19320), .C2(n19319), .A(n19318), .B(n19317), .ZN(
        P2_U3055) );
  NOR2_X1 U22265 ( .A1(n19562), .A2(n19506), .ZN(n19371) );
  NOR2_X1 U22266 ( .A1(n19679), .A2(n19349), .ZN(n19343) );
  OAI21_X1 U22267 ( .B1(n19321), .B2(n19343), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19322) );
  OAI21_X1 U22268 ( .B1(n19324), .B2(n19913), .A(n19322), .ZN(n19344) );
  AOI22_X1 U22269 ( .A1(n19762), .A2(n19344), .B1(n19761), .B2(n19343), .ZN(
        n19330) );
  AND2_X1 U22270 ( .A1(n19323), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19495) );
  INV_X1 U22271 ( .A(n19495), .ZN(n19446) );
  OAI21_X1 U22272 ( .B1(n19446), .B2(n19562), .A(n19324), .ZN(n19328) );
  INV_X1 U22273 ( .A(n19343), .ZN(n19325) );
  OAI211_X1 U22274 ( .C1(n19326), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19325), 
        .B(n19913), .ZN(n19327) );
  NAND3_X1 U22275 ( .A1(n19328), .A2(n19768), .A3(n19327), .ZN(n19346) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19715), .ZN(n19329) );
  OAI211_X1 U22277 ( .C1(n19729), .C2(n19379), .A(n19330), .B(n19329), .ZN(
        P2_U3056) );
  AOI22_X1 U22278 ( .A1(n19344), .A2(n19775), .B1(n19774), .B2(n19343), .ZN(
        n19332) );
  AOI22_X1 U22279 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19689), .ZN(n19331) );
  OAI211_X1 U22280 ( .C1(n19692), .C2(n19379), .A(n19332), .B(n19331), .ZN(
        P2_U3057) );
  AOI22_X1 U22281 ( .A1(n19781), .A2(n19344), .B1(n19780), .B2(n19343), .ZN(
        n19334) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19732), .ZN(n19333) );
  OAI211_X1 U22283 ( .C1(n19735), .C2(n19379), .A(n19334), .B(n19333), .ZN(
        P2_U3058) );
  AOI22_X1 U22284 ( .A1(n19344), .A2(n19787), .B1(n19786), .B2(n19343), .ZN(
        n19336) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19736), .ZN(n19335) );
  OAI211_X1 U22286 ( .C1(n19739), .C2(n19379), .A(n19336), .B(n19335), .ZN(
        P2_U3059) );
  AOI22_X1 U22287 ( .A1(n19344), .A2(n19793), .B1(n19792), .B2(n19343), .ZN(
        n19338) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19697), .ZN(n19337) );
  OAI211_X1 U22289 ( .C1(n19700), .C2(n19379), .A(n19338), .B(n19337), .ZN(
        P2_U3060) );
  AOI22_X1 U22290 ( .A1(n19344), .A2(n19798), .B1(n19301), .B2(n19343), .ZN(
        n19340) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19701), .ZN(n19339) );
  OAI211_X1 U22292 ( .C1(n19704), .C2(n19379), .A(n19340), .B(n19339), .ZN(
        P2_U3061) );
  AOI22_X1 U22293 ( .A1(n19344), .A2(n19804), .B1(n19803), .B2(n19343), .ZN(
        n19342) );
  AOI22_X1 U22294 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19746), .ZN(n19341) );
  OAI211_X1 U22295 ( .C1(n19749), .C2(n19379), .A(n19342), .B(n19341), .ZN(
        P2_U3062) );
  AOI22_X1 U22296 ( .A1(n19344), .A2(n19811), .B1(n19810), .B2(n19343), .ZN(
        n19348) );
  AOI22_X1 U22297 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19346), .B1(
        n19345), .B2(n19752), .ZN(n19347) );
  OAI211_X1 U22298 ( .C1(n19757), .C2(n19379), .A(n19348), .B(n19347), .ZN(
        P2_U3063) );
  NOR2_X1 U22299 ( .A1(n19593), .A2(n19349), .ZN(n19374) );
  OAI21_X1 U22300 ( .B1(n19352), .B2(n19374), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19351) );
  NOR2_X1 U22301 ( .A1(n19599), .A2(n19349), .ZN(n19353) );
  INV_X1 U22302 ( .A(n19353), .ZN(n19350) );
  NAND2_X1 U22303 ( .A1(n19351), .A2(n19350), .ZN(n19375) );
  AOI22_X1 U22304 ( .A1(n19375), .A2(n19762), .B1(n19761), .B2(n19374), .ZN(
        n19360) );
  AOI21_X1 U22305 ( .B1(n19352), .B2(n19533), .A(n19374), .ZN(n19356) );
  NAND2_X1 U22306 ( .A1(n19410), .A2(n19379), .ZN(n19354) );
  AOI21_X1 U22307 ( .B1(n19354), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19353), 
        .ZN(n19355) );
  MUX2_X1 U22308 ( .A(n19356), .B(n19355), .S(n19934), .Z(n19358) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19376), .B1(
        n19402), .B2(n19770), .ZN(n19359) );
  OAI211_X1 U22310 ( .C1(n19773), .C2(n19379), .A(n19360), .B(n19359), .ZN(
        P2_U3064) );
  AOI22_X1 U22311 ( .A1(n19375), .A2(n19775), .B1(n19774), .B2(n19374), .ZN(
        n19362) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19376), .B1(
        n19402), .B2(n19776), .ZN(n19361) );
  OAI211_X1 U22313 ( .C1(n19779), .C2(n19379), .A(n19362), .B(n19361), .ZN(
        P2_U3065) );
  AOI22_X1 U22314 ( .A1(n19375), .A2(n19781), .B1(n19780), .B2(n19374), .ZN(
        n19364) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19376), .B1(
        n19402), .B2(n19782), .ZN(n19363) );
  OAI211_X1 U22316 ( .C1(n19785), .C2(n19379), .A(n19364), .B(n19363), .ZN(
        P2_U3066) );
  AOI22_X1 U22317 ( .A1(n19375), .A2(n19787), .B1(n19786), .B2(n19374), .ZN(
        n19366) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19376), .B1(
        n19402), .B2(n19788), .ZN(n19365) );
  OAI211_X1 U22319 ( .C1(n19791), .C2(n19379), .A(n19366), .B(n19365), .ZN(
        P2_U3067) );
  AOI22_X1 U22320 ( .A1(n19375), .A2(n19793), .B1(n19792), .B2(n19374), .ZN(
        n19368) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19376), .B1(
        n19402), .B2(n19794), .ZN(n19367) );
  OAI211_X1 U22322 ( .C1(n19797), .C2(n19379), .A(n19368), .B(n19367), .ZN(
        P2_U3068) );
  AOI22_X1 U22323 ( .A1(n19375), .A2(n19798), .B1(n19301), .B2(n19374), .ZN(
        n19370) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19376), .B1(
        n19402), .B2(n19799), .ZN(n19369) );
  OAI211_X1 U22325 ( .C1(n19802), .C2(n19379), .A(n19370), .B(n19369), .ZN(
        P2_U3069) );
  AOI22_X1 U22326 ( .A1(n19375), .A2(n19804), .B1(n19803), .B2(n19374), .ZN(
        n19373) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19376), .B1(
        n19371), .B2(n19746), .ZN(n19372) );
  OAI211_X1 U22328 ( .C1(n19749), .C2(n19410), .A(n19373), .B(n19372), .ZN(
        P2_U3070) );
  AOI22_X1 U22329 ( .A1(n19375), .A2(n19811), .B1(n19810), .B2(n19374), .ZN(
        n19378) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19376), .B1(
        n19402), .B2(n19813), .ZN(n19377) );
  OAI211_X1 U22331 ( .C1(n19819), .C2(n19379), .A(n19378), .B(n19377), .ZN(
        P2_U3071) );
  AND2_X1 U22332 ( .A1(n19380), .A2(n19382), .ZN(n19405) );
  AOI22_X1 U22333 ( .A1(n19715), .A2(n19402), .B1(n19761), .B2(n19405), .ZN(
        n19391) );
  AOI21_X1 U22334 ( .B1(n19381), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19384) );
  INV_X1 U22335 ( .A(n19915), .ZN(n19629) );
  AOI21_X1 U22336 ( .B1(n19495), .B2(n19629), .A(n19913), .ZN(n19385) );
  NAND2_X1 U22337 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19382), .ZN(
        n19388) );
  NAND2_X1 U22338 ( .A1(n19385), .A2(n19388), .ZN(n19383) );
  OAI211_X1 U22339 ( .C1(n19405), .C2(n19384), .A(n19383), .B(n19768), .ZN(
        n19407) );
  INV_X1 U22340 ( .A(n19385), .ZN(n19389) );
  OAI21_X1 U22341 ( .B1(n19386), .B2(n19405), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19387) );
  OAI21_X1 U22342 ( .B1(n19389), .B2(n19388), .A(n19387), .ZN(n19406) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19407), .B1(
        n19762), .B2(n19406), .ZN(n19390) );
  OAI211_X1 U22344 ( .C1(n19729), .C2(n19445), .A(n19391), .B(n19390), .ZN(
        P2_U3072) );
  AOI22_X1 U22345 ( .A1(n19689), .A2(n19402), .B1(n19405), .B2(n19774), .ZN(
        n19393) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19407), .B1(
        n19775), .B2(n19406), .ZN(n19392) );
  OAI211_X1 U22347 ( .C1(n19692), .C2(n19445), .A(n19393), .B(n19392), .ZN(
        P2_U3073) );
  AOI22_X1 U22348 ( .A1(n19732), .A2(n19402), .B1(n19780), .B2(n19405), .ZN(
        n19395) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19407), .B1(
        n19781), .B2(n19406), .ZN(n19394) );
  OAI211_X1 U22350 ( .C1(n19735), .C2(n19445), .A(n19395), .B(n19394), .ZN(
        P2_U3074) );
  AOI22_X1 U22351 ( .A1(n19736), .A2(n19402), .B1(n19405), .B2(n19786), .ZN(
        n19397) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19407), .B1(
        n19787), .B2(n19406), .ZN(n19396) );
  OAI211_X1 U22353 ( .C1(n19739), .C2(n19445), .A(n19397), .B(n19396), .ZN(
        P2_U3075) );
  AOI22_X1 U22354 ( .A1(n19697), .A2(n19402), .B1(n19405), .B2(n19792), .ZN(
        n19399) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19407), .B1(
        n19793), .B2(n19406), .ZN(n19398) );
  OAI211_X1 U22356 ( .C1(n19700), .C2(n19445), .A(n19399), .B(n19398), .ZN(
        P2_U3076) );
  AOI22_X1 U22357 ( .A1(n19701), .A2(n19402), .B1(n19405), .B2(n19301), .ZN(
        n19401) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19407), .B1(
        n19798), .B2(n19406), .ZN(n19400) );
  OAI211_X1 U22359 ( .C1(n19704), .C2(n19445), .A(n19401), .B(n19400), .ZN(
        P2_U3077) );
  AOI22_X1 U22360 ( .A1(n19746), .A2(n19402), .B1(n19405), .B2(n19803), .ZN(
        n19404) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19407), .B1(
        n19804), .B2(n19406), .ZN(n19403) );
  OAI211_X1 U22362 ( .C1(n19749), .C2(n19445), .A(n19404), .B(n19403), .ZN(
        P2_U3078) );
  AOI22_X1 U22363 ( .A1(n19813), .A2(n19437), .B1(n19405), .B2(n19810), .ZN(
        n19409) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19407), .B1(
        n19811), .B2(n19406), .ZN(n19408) );
  OAI211_X1 U22365 ( .C1(n19819), .C2(n19410), .A(n19409), .B(n19408), .ZN(
        P2_U3079) );
  NAND2_X1 U22366 ( .A1(n19926), .A2(n19411), .ZN(n19421) );
  INV_X1 U22367 ( .A(n19412), .ZN(n19415) );
  NAND2_X1 U22368 ( .A1(n19413), .A2(n19943), .ZN(n19452) );
  NOR2_X1 U22369 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19452), .ZN(
        n19440) );
  OAI21_X1 U22370 ( .B1(n10756), .B2(n19440), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19414) );
  OAI21_X1 U22371 ( .B1(n19421), .B2(n19415), .A(n19414), .ZN(n19441) );
  AOI22_X1 U22372 ( .A1(n19441), .A2(n19762), .B1(n19761), .B2(n19440), .ZN(
        n19426) );
  INV_X1 U22373 ( .A(n10756), .ZN(n19417) );
  INV_X1 U22374 ( .A(n19440), .ZN(n19416) );
  OAI211_X1 U22375 ( .C1(n19417), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19416), 
        .B(n19913), .ZN(n19424) );
  INV_X1 U22376 ( .A(n19418), .ZN(n19422) );
  OAI21_X1 U22377 ( .B1(n19437), .B2(n19470), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19420) );
  OAI21_X1 U22378 ( .B1(n19422), .B2(n19421), .A(n19420), .ZN(n19423) );
  NAND3_X1 U22379 ( .A1(n19424), .A2(n19768), .A3(n19423), .ZN(n19442) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19442), .B1(
        n19470), .B2(n19770), .ZN(n19425) );
  OAI211_X1 U22381 ( .C1(n19773), .C2(n19445), .A(n19426), .B(n19425), .ZN(
        P2_U3080) );
  AOI22_X1 U22382 ( .A1(n19441), .A2(n19775), .B1(n19774), .B2(n19440), .ZN(
        n19428) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19442), .B1(
        n19470), .B2(n19776), .ZN(n19427) );
  OAI211_X1 U22384 ( .C1(n19779), .C2(n19445), .A(n19428), .B(n19427), .ZN(
        P2_U3081) );
  AOI22_X1 U22385 ( .A1(n19441), .A2(n19781), .B1(n19780), .B2(n19440), .ZN(
        n19430) );
  AOI22_X1 U22386 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19442), .B1(
        n19437), .B2(n19732), .ZN(n19429) );
  OAI211_X1 U22387 ( .C1(n19735), .C2(n19466), .A(n19430), .B(n19429), .ZN(
        P2_U3082) );
  AOI22_X1 U22388 ( .A1(n19441), .A2(n19787), .B1(n19786), .B2(n19440), .ZN(
        n19432) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19442), .B1(
        n19437), .B2(n19736), .ZN(n19431) );
  OAI211_X1 U22390 ( .C1(n19739), .C2(n19466), .A(n19432), .B(n19431), .ZN(
        P2_U3083) );
  AOI22_X1 U22391 ( .A1(n19441), .A2(n19793), .B1(n19792), .B2(n19440), .ZN(
        n19434) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19442), .B1(
        n19437), .B2(n19697), .ZN(n19433) );
  OAI211_X1 U22393 ( .C1(n19700), .C2(n19466), .A(n19434), .B(n19433), .ZN(
        P2_U3084) );
  AOI22_X1 U22394 ( .A1(n19441), .A2(n19798), .B1(n19301), .B2(n19440), .ZN(
        n19436) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19442), .B1(
        n19470), .B2(n19799), .ZN(n19435) );
  OAI211_X1 U22396 ( .C1(n19802), .C2(n19445), .A(n19436), .B(n19435), .ZN(
        P2_U3085) );
  AOI22_X1 U22397 ( .A1(n19441), .A2(n19804), .B1(n19803), .B2(n19440), .ZN(
        n19439) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19442), .B1(
        n19437), .B2(n19746), .ZN(n19438) );
  OAI211_X1 U22399 ( .C1(n19749), .C2(n19466), .A(n19439), .B(n19438), .ZN(
        P2_U3086) );
  AOI22_X1 U22400 ( .A1(n19441), .A2(n19811), .B1(n19810), .B2(n19440), .ZN(
        n19444) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19442), .B1(
        n19470), .B2(n19813), .ZN(n19443) );
  OAI211_X1 U22402 ( .C1(n19819), .C2(n19445), .A(n19444), .B(n19443), .ZN(
        P2_U3087) );
  NOR2_X1 U22403 ( .A1(n19496), .A2(n19679), .ZN(n19469) );
  AOI22_X1 U22404 ( .A1(n19715), .A2(n19470), .B1(n19761), .B2(n19469), .ZN(
        n19455) );
  OAI21_X1 U22405 ( .B1(n19446), .B2(n19676), .A(n19934), .ZN(n19453) );
  INV_X1 U22406 ( .A(n19452), .ZN(n19450) );
  INV_X1 U22407 ( .A(n19469), .ZN(n19447) );
  OAI211_X1 U22408 ( .C1(n19448), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19447), 
        .B(n19913), .ZN(n19449) );
  OAI211_X1 U22409 ( .C1(n19453), .C2(n19450), .A(n19768), .B(n19449), .ZN(
        n19472) );
  OAI21_X1 U22410 ( .B1(n10749), .B2(n19469), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19451) );
  OAI21_X1 U22411 ( .B1(n19453), .B2(n19452), .A(n19451), .ZN(n19471) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19472), .B1(
        n19762), .B2(n19471), .ZN(n19454) );
  OAI211_X1 U22413 ( .C1(n19729), .C2(n19494), .A(n19455), .B(n19454), .ZN(
        P2_U3088) );
  AOI22_X1 U22414 ( .A1(n19776), .A2(n19486), .B1(n19774), .B2(n19469), .ZN(
        n19457) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19472), .B1(
        n19775), .B2(n19471), .ZN(n19456) );
  OAI211_X1 U22416 ( .C1(n19779), .C2(n19466), .A(n19457), .B(n19456), .ZN(
        P2_U3089) );
  AOI22_X1 U22417 ( .A1(n19782), .A2(n19486), .B1(n19780), .B2(n19469), .ZN(
        n19459) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19472), .B1(
        n19781), .B2(n19471), .ZN(n19458) );
  OAI211_X1 U22419 ( .C1(n19785), .C2(n19466), .A(n19459), .B(n19458), .ZN(
        P2_U3090) );
  AOI22_X1 U22420 ( .A1(n19788), .A2(n19486), .B1(n19469), .B2(n19786), .ZN(
        n19461) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19472), .B1(
        n19787), .B2(n19471), .ZN(n19460) );
  OAI211_X1 U22422 ( .C1(n19791), .C2(n19466), .A(n19461), .B(n19460), .ZN(
        P2_U3091) );
  AOI22_X1 U22423 ( .A1(n19697), .A2(n19470), .B1(n19469), .B2(n19792), .ZN(
        n19463) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19472), .B1(
        n19793), .B2(n19471), .ZN(n19462) );
  OAI211_X1 U22425 ( .C1(n19700), .C2(n19494), .A(n19463), .B(n19462), .ZN(
        P2_U3092) );
  AOI22_X1 U22426 ( .A1(n19799), .A2(n19486), .B1(n19469), .B2(n19301), .ZN(
        n19465) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19472), .B1(
        n19798), .B2(n19471), .ZN(n19464) );
  OAI211_X1 U22428 ( .C1(n19802), .C2(n19466), .A(n19465), .B(n19464), .ZN(
        P2_U3093) );
  AOI22_X1 U22429 ( .A1(n19746), .A2(n19470), .B1(n19803), .B2(n19469), .ZN(
        n19468) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19472), .B1(
        n19804), .B2(n19471), .ZN(n19467) );
  OAI211_X1 U22431 ( .C1(n19749), .C2(n19494), .A(n19468), .B(n19467), .ZN(
        P2_U3094) );
  AOI22_X1 U22432 ( .A1(n19752), .A2(n19470), .B1(n19810), .B2(n19469), .ZN(
        n19474) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19472), .B1(
        n19811), .B2(n19471), .ZN(n19473) );
  OAI211_X1 U22434 ( .C1(n19757), .C2(n19494), .A(n19474), .B(n19473), .ZN(
        P2_U3095) );
  AOI22_X1 U22435 ( .A1(n19490), .A2(n19775), .B1(n19489), .B2(n19774), .ZN(
        n19477) );
  INV_X1 U22436 ( .A(n19475), .ZN(n19491) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19491), .B1(
        n19521), .B2(n19776), .ZN(n19476) );
  OAI211_X1 U22438 ( .C1(n19779), .C2(n19494), .A(n19477), .B(n19476), .ZN(
        P2_U3097) );
  AOI22_X1 U22439 ( .A1(n19490), .A2(n19781), .B1(n19780), .B2(n19489), .ZN(
        n19479) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19491), .B1(
        n19521), .B2(n19782), .ZN(n19478) );
  OAI211_X1 U22441 ( .C1(n19785), .C2(n19494), .A(n19479), .B(n19478), .ZN(
        P2_U3098) );
  AOI22_X1 U22442 ( .A1(n19490), .A2(n19787), .B1(n19489), .B2(n19786), .ZN(
        n19481) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19491), .B1(
        n19521), .B2(n19788), .ZN(n19480) );
  OAI211_X1 U22444 ( .C1(n19791), .C2(n19494), .A(n19481), .B(n19480), .ZN(
        P2_U3099) );
  AOI22_X1 U22445 ( .A1(n19490), .A2(n19793), .B1(n19489), .B2(n19792), .ZN(
        n19483) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19491), .B1(
        n19521), .B2(n19794), .ZN(n19482) );
  OAI211_X1 U22447 ( .C1(n19797), .C2(n19494), .A(n19483), .B(n19482), .ZN(
        P2_U3100) );
  AOI22_X1 U22448 ( .A1(n19490), .A2(n19798), .B1(n19489), .B2(n19301), .ZN(
        n19485) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19491), .B1(
        n19521), .B2(n19799), .ZN(n19484) );
  OAI211_X1 U22450 ( .C1(n19802), .C2(n19494), .A(n19485), .B(n19484), .ZN(
        P2_U3101) );
  INV_X1 U22451 ( .A(n19521), .ZN(n19530) );
  AOI22_X1 U22452 ( .A1(n19490), .A2(n19804), .B1(n19489), .B2(n19803), .ZN(
        n19488) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19491), .B1(
        n19486), .B2(n19746), .ZN(n19487) );
  OAI211_X1 U22454 ( .C1(n19749), .C2(n19530), .A(n19488), .B(n19487), .ZN(
        P2_U3102) );
  AOI22_X1 U22455 ( .A1(n19490), .A2(n19811), .B1(n19489), .B2(n19810), .ZN(
        n19493) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19491), .B1(
        n19521), .B2(n19813), .ZN(n19492) );
  OAI211_X1 U22457 ( .C1(n19819), .C2(n19494), .A(n19493), .B(n19492), .ZN(
        P2_U3103) );
  AND2_X1 U22458 ( .A1(n19495), .A2(n19763), .ZN(n19912) );
  NOR2_X1 U22459 ( .A1(n19943), .A2(n19496), .ZN(n19501) );
  OAI21_X1 U22460 ( .B1(n19912), .B2(n19501), .A(n19768), .ZN(n19500) );
  INV_X1 U22461 ( .A(n19535), .ZN(n19538) );
  AND2_X1 U22462 ( .A1(n19535), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19497) );
  NAND2_X1 U22463 ( .A1(n19498), .A2(n19497), .ZN(n19504) );
  OAI21_X1 U22464 ( .B1(n19538), .B2(n19533), .A(n19504), .ZN(n19499) );
  INV_X1 U22465 ( .A(n19501), .ZN(n19502) );
  OAI21_X1 U22466 ( .B1(n19502), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19973), 
        .ZN(n19503) );
  AOI22_X1 U22467 ( .A1(n19762), .A2(n19526), .B1(n19538), .B2(n19761), .ZN(
        n19508) );
  AOI22_X1 U22468 ( .A1(n19553), .A2(n19770), .B1(n19521), .B2(n19715), .ZN(
        n19507) );
  OAI211_X1 U22469 ( .C1(n19525), .C2(n19509), .A(n19508), .B(n19507), .ZN(
        P2_U3104) );
  AOI22_X1 U22470 ( .A1(n19526), .A2(n19775), .B1(n19538), .B2(n19774), .ZN(
        n19511) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19527), .B1(
        n19553), .B2(n19776), .ZN(n19510) );
  OAI211_X1 U22472 ( .C1(n19779), .C2(n19530), .A(n19511), .B(n19510), .ZN(
        P2_U3105) );
  INV_X1 U22473 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n19514) );
  AOI22_X1 U22474 ( .A1(n19781), .A2(n19526), .B1(n19538), .B2(n19780), .ZN(
        n19513) );
  AOI22_X1 U22475 ( .A1(n19553), .A2(n19782), .B1(n19521), .B2(n19732), .ZN(
        n19512) );
  OAI211_X1 U22476 ( .C1(n19525), .C2(n19514), .A(n19513), .B(n19512), .ZN(
        P2_U3106) );
  AOI22_X1 U22477 ( .A1(n19526), .A2(n19787), .B1(n19538), .B2(n19786), .ZN(
        n19516) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19527), .B1(
        n19553), .B2(n19788), .ZN(n19515) );
  OAI211_X1 U22479 ( .C1(n19791), .C2(n19530), .A(n19516), .B(n19515), .ZN(
        P2_U3107) );
  AOI22_X1 U22480 ( .A1(n19526), .A2(n19793), .B1(n19538), .B2(n19792), .ZN(
        n19518) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19527), .B1(
        n19553), .B2(n19794), .ZN(n19517) );
  OAI211_X1 U22482 ( .C1(n19797), .C2(n19530), .A(n19518), .B(n19517), .ZN(
        P2_U3108) );
  AOI22_X1 U22483 ( .A1(n19526), .A2(n19798), .B1(n19538), .B2(n19301), .ZN(
        n19520) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19527), .B1(
        n19553), .B2(n19799), .ZN(n19519) );
  OAI211_X1 U22485 ( .C1(n19802), .C2(n19530), .A(n19520), .B(n19519), .ZN(
        P2_U3109) );
  AOI22_X1 U22486 ( .A1(n19526), .A2(n19804), .B1(n19538), .B2(n19803), .ZN(
        n19523) );
  AOI22_X1 U22487 ( .A1(n19553), .A2(n19805), .B1(n19521), .B2(n19746), .ZN(
        n19522) );
  OAI211_X1 U22488 ( .C1(n19525), .C2(n19524), .A(n19523), .B(n19522), .ZN(
        P2_U3110) );
  AOI22_X1 U22489 ( .A1(n19526), .A2(n19811), .B1(n19538), .B2(n19810), .ZN(
        n19529) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19527), .B1(
        n19553), .B2(n19813), .ZN(n19528) );
  OAI211_X1 U22491 ( .C1(n19819), .C2(n19530), .A(n19529), .B(n19528), .ZN(
        P2_U3111) );
  NOR2_X2 U22492 ( .A1(n19713), .A2(n19562), .ZN(n19585) );
  NAND2_X1 U22493 ( .A1(n19933), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19624) );
  NOR2_X1 U22494 ( .A1(n19624), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19566) );
  INV_X1 U22495 ( .A(n19566), .ZN(n19569) );
  NOR2_X1 U22496 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19569), .ZN(
        n19556) );
  AOI22_X1 U22497 ( .A1(n19770), .A2(n19585), .B1(n19761), .B2(n19556), .ZN(
        n19542) );
  INV_X1 U22498 ( .A(n19585), .ZN(n19531) );
  NAND2_X1 U22499 ( .A1(n19531), .A2(n19561), .ZN(n19532) );
  AOI21_X1 U22500 ( .B1(n19532), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19913), 
        .ZN(n19537) );
  OAI21_X1 U22501 ( .B1(n10764), .B2(n19973), .A(n19533), .ZN(n19534) );
  AOI21_X1 U22502 ( .B1(n19537), .B2(n19535), .A(n19534), .ZN(n19536) );
  OAI21_X1 U22503 ( .B1(n19556), .B2(n19536), .A(n19768), .ZN(n19558) );
  OAI21_X1 U22504 ( .B1(n19538), .B2(n19556), .A(n19537), .ZN(n19540) );
  OAI21_X1 U22505 ( .B1(n10764), .B2(n19556), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19539) );
  NAND2_X1 U22506 ( .A1(n19540), .A2(n19539), .ZN(n19557) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19558), .B1(
        n19762), .B2(n19557), .ZN(n19541) );
  OAI211_X1 U22508 ( .C1(n19773), .C2(n19561), .A(n19542), .B(n19541), .ZN(
        P2_U3112) );
  AOI22_X1 U22509 ( .A1(n19776), .A2(n19585), .B1(n19556), .B2(n19774), .ZN(
        n19544) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19775), .ZN(n19543) );
  OAI211_X1 U22511 ( .C1(n19779), .C2(n19561), .A(n19544), .B(n19543), .ZN(
        P2_U3113) );
  AOI22_X1 U22512 ( .A1(n19782), .A2(n19585), .B1(n19780), .B2(n19556), .ZN(
        n19546) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19781), .ZN(n19545) );
  OAI211_X1 U22514 ( .C1(n19785), .C2(n19561), .A(n19546), .B(n19545), .ZN(
        P2_U3114) );
  AOI22_X1 U22515 ( .A1(n19788), .A2(n19585), .B1(n19556), .B2(n19786), .ZN(
        n19548) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19787), .ZN(n19547) );
  OAI211_X1 U22517 ( .C1(n19791), .C2(n19561), .A(n19548), .B(n19547), .ZN(
        P2_U3115) );
  AOI22_X1 U22518 ( .A1(n19794), .A2(n19585), .B1(n19556), .B2(n19792), .ZN(
        n19550) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19793), .ZN(n19549) );
  OAI211_X1 U22520 ( .C1(n19797), .C2(n19561), .A(n19550), .B(n19549), .ZN(
        P2_U3116) );
  AOI22_X1 U22521 ( .A1(n19799), .A2(n19585), .B1(n19556), .B2(n19301), .ZN(
        n19552) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19798), .ZN(n19551) );
  OAI211_X1 U22523 ( .C1(n19802), .C2(n19561), .A(n19552), .B(n19551), .ZN(
        P2_U3117) );
  AOI22_X1 U22524 ( .A1(n19746), .A2(n19553), .B1(n19803), .B2(n19556), .ZN(
        n19555) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19804), .ZN(n19554) );
  OAI211_X1 U22526 ( .C1(n19749), .C2(n19531), .A(n19555), .B(n19554), .ZN(
        P2_U3118) );
  AOI22_X1 U22527 ( .A1(n19813), .A2(n19585), .B1(n19810), .B2(n19556), .ZN(
        n19560) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19811), .ZN(n19559) );
  OAI211_X1 U22529 ( .C1(n19819), .C2(n19561), .A(n19560), .B(n19559), .ZN(
        P2_U3119) );
  NOR2_X1 U22530 ( .A1(n19679), .A2(n19624), .ZN(n19590) );
  AOI22_X1 U22531 ( .A1(n19715), .A2(n19585), .B1(n19761), .B2(n19590), .ZN(
        n19572) );
  NAND2_X1 U22532 ( .A1(n19920), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19628) );
  OAI21_X1 U22533 ( .B1(n19628), .B2(n19562), .A(n19934), .ZN(n19570) );
  INV_X1 U22534 ( .A(n19590), .ZN(n19563) );
  OAI211_X1 U22535 ( .C1(n19564), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19563), 
        .B(n19913), .ZN(n19565) );
  OAI211_X1 U22536 ( .C1(n19570), .C2(n19566), .A(n19768), .B(n19565), .ZN(
        n19587) );
  OAI21_X1 U22537 ( .B1(n19567), .B2(n19590), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19568) );
  OAI21_X1 U22538 ( .B1(n19570), .B2(n19569), .A(n19568), .ZN(n19586) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19587), .B1(
        n19762), .B2(n19586), .ZN(n19571) );
  OAI211_X1 U22540 ( .C1(n19729), .C2(n19623), .A(n19572), .B(n19571), .ZN(
        P2_U3120) );
  AOI22_X1 U22541 ( .A1(n19776), .A2(n19614), .B1(n19774), .B2(n19590), .ZN(
        n19574) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19587), .B1(
        n19775), .B2(n19586), .ZN(n19573) );
  OAI211_X1 U22543 ( .C1(n19779), .C2(n19531), .A(n19574), .B(n19573), .ZN(
        P2_U3121) );
  AOI22_X1 U22544 ( .A1(n19732), .A2(n19585), .B1(n19780), .B2(n19590), .ZN(
        n19576) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19587), .B1(
        n19781), .B2(n19586), .ZN(n19575) );
  OAI211_X1 U22546 ( .C1(n19735), .C2(n19623), .A(n19576), .B(n19575), .ZN(
        P2_U3122) );
  AOI22_X1 U22547 ( .A1(n19788), .A2(n19614), .B1(n19786), .B2(n19590), .ZN(
        n19578) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19587), .B1(
        n19787), .B2(n19586), .ZN(n19577) );
  OAI211_X1 U22549 ( .C1(n19791), .C2(n19531), .A(n19578), .B(n19577), .ZN(
        P2_U3123) );
  AOI22_X1 U22550 ( .A1(n19697), .A2(n19585), .B1(n19792), .B2(n19590), .ZN(
        n19580) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19587), .B1(
        n19793), .B2(n19586), .ZN(n19579) );
  OAI211_X1 U22552 ( .C1(n19700), .C2(n19623), .A(n19580), .B(n19579), .ZN(
        P2_U3124) );
  AOI22_X1 U22553 ( .A1(n19701), .A2(n19585), .B1(n19301), .B2(n19590), .ZN(
        n19582) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19587), .B1(
        n19798), .B2(n19586), .ZN(n19581) );
  OAI211_X1 U22555 ( .C1(n19704), .C2(n19623), .A(n19582), .B(n19581), .ZN(
        P2_U3125) );
  AOI22_X1 U22556 ( .A1(n19805), .A2(n19614), .B1(n19803), .B2(n19590), .ZN(
        n19584) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19587), .B1(
        n19804), .B2(n19586), .ZN(n19583) );
  OAI211_X1 U22558 ( .C1(n19808), .C2(n19531), .A(n19584), .B(n19583), .ZN(
        P2_U3126) );
  AOI22_X1 U22559 ( .A1(n19752), .A2(n19585), .B1(n19810), .B2(n19590), .ZN(
        n19589) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19587), .B1(
        n19811), .B2(n19586), .ZN(n19588) );
  OAI211_X1 U22561 ( .C1(n19757), .C2(n19623), .A(n19589), .B(n19588), .ZN(
        P2_U3127) );
  INV_X1 U22562 ( .A(n19597), .ZN(n19592) );
  AOI221_X1 U22563 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19614), .C1(
        P2_STATEBS16_REG_SCAN_IN), .C2(n19619), .A(n19590), .ZN(n19591) );
  MUX2_X1 U22564 ( .A(n19592), .B(n19591), .S(n19973), .Z(n19595) );
  NOR2_X1 U22565 ( .A1(n19593), .A2(n19624), .ZN(n19617) );
  INV_X1 U22566 ( .A(n19617), .ZN(n19594) );
  OAI21_X1 U22567 ( .B1(n19595), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19594), 
        .ZN(n19596) );
  AND2_X1 U22568 ( .A1(n19596), .A2(n19768), .ZN(n19603) );
  INV_X1 U22569 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n19602) );
  OAI21_X1 U22570 ( .B1(n19597), .B2(n19617), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19598) );
  OAI21_X1 U22571 ( .B1(n19624), .B2(n19599), .A(n19598), .ZN(n19618) );
  AOI22_X1 U22572 ( .A1(n19618), .A2(n19762), .B1(n19761), .B2(n19617), .ZN(
        n19601) );
  AOI22_X1 U22573 ( .A1(n19619), .A2(n19770), .B1(n19614), .B2(n19715), .ZN(
        n19600) );
  OAI211_X1 U22574 ( .C1(n19603), .C2(n19602), .A(n19601), .B(n19600), .ZN(
        P2_U3128) );
  AOI22_X1 U22575 ( .A1(n19618), .A2(n19775), .B1(n19774), .B2(n19617), .ZN(
        n19605) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19776), .ZN(n19604) );
  OAI211_X1 U22577 ( .C1(n19779), .C2(n19623), .A(n19605), .B(n19604), .ZN(
        P2_U3129) );
  AOI22_X1 U22578 ( .A1(n19618), .A2(n19781), .B1(n19780), .B2(n19617), .ZN(
        n19607) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19782), .ZN(n19606) );
  OAI211_X1 U22580 ( .C1(n19785), .C2(n19623), .A(n19607), .B(n19606), .ZN(
        P2_U3130) );
  AOI22_X1 U22581 ( .A1(n19618), .A2(n19787), .B1(n19786), .B2(n19617), .ZN(
        n19609) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19788), .ZN(n19608) );
  OAI211_X1 U22583 ( .C1(n19791), .C2(n19623), .A(n19609), .B(n19608), .ZN(
        P2_U3131) );
  AOI22_X1 U22584 ( .A1(n19618), .A2(n19793), .B1(n19792), .B2(n19617), .ZN(
        n19611) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19794), .ZN(n19610) );
  OAI211_X1 U22586 ( .C1(n19797), .C2(n19623), .A(n19611), .B(n19610), .ZN(
        P2_U3132) );
  AOI22_X1 U22587 ( .A1(n19618), .A2(n19798), .B1(n19301), .B2(n19617), .ZN(
        n19613) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19799), .ZN(n19612) );
  OAI211_X1 U22589 ( .C1(n19802), .C2(n19623), .A(n19613), .B(n19612), .ZN(
        P2_U3133) );
  AOI22_X1 U22590 ( .A1(n19618), .A2(n19804), .B1(n19803), .B2(n19617), .ZN(
        n19616) );
  AOI22_X1 U22591 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19620), .B1(
        n19614), .B2(n19746), .ZN(n19615) );
  OAI211_X1 U22592 ( .C1(n19749), .C2(n19653), .A(n19616), .B(n19615), .ZN(
        P2_U3134) );
  AOI22_X1 U22593 ( .A1(n19618), .A2(n19811), .B1(n19810), .B2(n19617), .ZN(
        n19622) );
  AOI22_X1 U22594 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n19813), .ZN(n19621) );
  OAI211_X1 U22595 ( .C1(n19819), .C2(n19623), .A(n19622), .B(n19621), .ZN(
        P2_U3135) );
  OR2_X1 U22596 ( .A1(n19943), .A2(n19624), .ZN(n19631) );
  OR2_X1 U22597 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19631), .ZN(n19627) );
  NOR2_X1 U22598 ( .A1(n19625), .A2(n19624), .ZN(n19648) );
  NOR3_X1 U22599 ( .A1(n19626), .A2(n19648), .A3(n19973), .ZN(n19630) );
  AOI21_X1 U22600 ( .B1(n19973), .B2(n19627), .A(n19630), .ZN(n19649) );
  AOI22_X1 U22601 ( .A1(n19649), .A2(n19762), .B1(n19761), .B2(n19648), .ZN(
        n19635) );
  INV_X1 U22602 ( .A(n19628), .ZN(n19764) );
  NAND2_X1 U22603 ( .A1(n19764), .A2(n19629), .ZN(n19632) );
  AOI21_X1 U22604 ( .B1(n19632), .B2(n19631), .A(n19630), .ZN(n19633) );
  OAI211_X1 U22605 ( .C1(n19648), .C2(n19533), .A(n19633), .B(n19768), .ZN(
        n19650) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19650), .B1(
        n19670), .B2(n19770), .ZN(n19634) );
  OAI211_X1 U22607 ( .C1(n19773), .C2(n19653), .A(n19635), .B(n19634), .ZN(
        P2_U3136) );
  AOI22_X1 U22608 ( .A1(n19649), .A2(n19775), .B1(n19774), .B2(n19648), .ZN(
        n19637) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19650), .B1(
        n19670), .B2(n19776), .ZN(n19636) );
  OAI211_X1 U22610 ( .C1(n19779), .C2(n19653), .A(n19637), .B(n19636), .ZN(
        P2_U3137) );
  AOI22_X1 U22611 ( .A1(n19649), .A2(n19781), .B1(n19780), .B2(n19648), .ZN(
        n19639) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19650), .B1(
        n19670), .B2(n19782), .ZN(n19638) );
  OAI211_X1 U22613 ( .C1(n19785), .C2(n19653), .A(n19639), .B(n19638), .ZN(
        P2_U3138) );
  AOI22_X1 U22614 ( .A1(n19649), .A2(n19787), .B1(n19786), .B2(n19648), .ZN(
        n19641) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19650), .B1(
        n19670), .B2(n19788), .ZN(n19640) );
  OAI211_X1 U22616 ( .C1(n19791), .C2(n19653), .A(n19641), .B(n19640), .ZN(
        P2_U3139) );
  AOI22_X1 U22617 ( .A1(n19649), .A2(n19793), .B1(n19792), .B2(n19648), .ZN(
        n19643) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19650), .B1(
        n19670), .B2(n19794), .ZN(n19642) );
  OAI211_X1 U22619 ( .C1(n19797), .C2(n19653), .A(n19643), .B(n19642), .ZN(
        P2_U3140) );
  AOI22_X1 U22620 ( .A1(n19649), .A2(n19798), .B1(n19301), .B2(n19648), .ZN(
        n19645) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19650), .B1(
        n19670), .B2(n19799), .ZN(n19644) );
  OAI211_X1 U22622 ( .C1(n19802), .C2(n19653), .A(n19645), .B(n19644), .ZN(
        P2_U3141) );
  AOI22_X1 U22623 ( .A1(n19649), .A2(n19804), .B1(n19803), .B2(n19648), .ZN(
        n19647) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19650), .B1(
        n19670), .B2(n19805), .ZN(n19646) );
  OAI211_X1 U22625 ( .C1(n19808), .C2(n19653), .A(n19647), .B(n19646), .ZN(
        P2_U3142) );
  AOI22_X1 U22626 ( .A1(n19649), .A2(n19811), .B1(n19810), .B2(n19648), .ZN(
        n19652) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19650), .B1(
        n19670), .B2(n19813), .ZN(n19651) );
  OAI211_X1 U22628 ( .C1(n19819), .C2(n19653), .A(n19652), .B(n19651), .ZN(
        P2_U3143) );
  AOI22_X1 U22629 ( .A1(n19669), .A2(n19775), .B1(n19668), .B2(n19774), .ZN(
        n19655) );
  AOI22_X1 U22630 ( .A1(n19709), .A2(n19776), .B1(n19670), .B2(n19689), .ZN(
        n19654) );
  OAI211_X1 U22631 ( .C1(n19674), .C2(n9847), .A(n19655), .B(n19654), .ZN(
        P2_U3145) );
  INV_X1 U22632 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n19658) );
  AOI22_X1 U22633 ( .A1(n19669), .A2(n19787), .B1(n19668), .B2(n19786), .ZN(
        n19657) );
  AOI22_X1 U22634 ( .A1(n19709), .A2(n19788), .B1(n19670), .B2(n19736), .ZN(
        n19656) );
  OAI211_X1 U22635 ( .C1(n19674), .C2(n19658), .A(n19657), .B(n19656), .ZN(
        P2_U3147) );
  INV_X1 U22636 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n19661) );
  AOI22_X1 U22637 ( .A1(n19669), .A2(n19793), .B1(n19668), .B2(n19792), .ZN(
        n19660) );
  AOI22_X1 U22638 ( .A1(n19709), .A2(n19794), .B1(n19670), .B2(n19697), .ZN(
        n19659) );
  OAI211_X1 U22639 ( .C1(n19674), .C2(n19661), .A(n19660), .B(n19659), .ZN(
        P2_U3148) );
  INV_X1 U22640 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n19664) );
  AOI22_X1 U22641 ( .A1(n19669), .A2(n19798), .B1(n19668), .B2(n19301), .ZN(
        n19663) );
  AOI22_X1 U22642 ( .A1(n19709), .A2(n19799), .B1(n19670), .B2(n19701), .ZN(
        n19662) );
  OAI211_X1 U22643 ( .C1(n19674), .C2(n19664), .A(n19663), .B(n19662), .ZN(
        P2_U3149) );
  INV_X1 U22644 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n19667) );
  AOI22_X1 U22645 ( .A1(n19669), .A2(n19804), .B1(n19668), .B2(n19803), .ZN(
        n19666) );
  AOI22_X1 U22646 ( .A1(n19670), .A2(n19746), .B1(n19709), .B2(n19805), .ZN(
        n19665) );
  OAI211_X1 U22647 ( .C1(n19674), .C2(n19667), .A(n19666), .B(n19665), .ZN(
        P2_U3150) );
  INV_X1 U22648 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n19673) );
  AOI22_X1 U22649 ( .A1(n19669), .A2(n19811), .B1(n19668), .B2(n19810), .ZN(
        n19672) );
  AOI22_X1 U22650 ( .A1(n19709), .A2(n19813), .B1(n19670), .B2(n19752), .ZN(
        n19671) );
  OAI211_X1 U22651 ( .C1(n19674), .C2(n19673), .A(n19672), .B(n19671), .ZN(
        P2_U3151) );
  INV_X1 U22652 ( .A(n19675), .ZN(n19677) );
  INV_X1 U22653 ( .A(n19676), .ZN(n19682) );
  INV_X1 U22654 ( .A(n19717), .ZN(n19678) );
  NOR2_X1 U22655 ( .A1(n19679), .A2(n19678), .ZN(n19707) );
  NOR3_X1 U22656 ( .A1(n19680), .A2(n19707), .A3(n19973), .ZN(n19683) );
  AOI211_X2 U22657 ( .C1(n19684), .C2(n19973), .A(n19681), .B(n19683), .ZN(
        n19708) );
  AOI22_X1 U22658 ( .A1(n19708), .A2(n19762), .B1(n19761), .B2(n19707), .ZN(
        n19688) );
  NAND2_X1 U22659 ( .A1(n19764), .A2(n19682), .ZN(n19685) );
  AOI21_X1 U22660 ( .B1(n19685), .B2(n19684), .A(n19683), .ZN(n19686) );
  OAI211_X1 U22661 ( .C1(n19707), .C2(n19533), .A(n19686), .B(n19768), .ZN(
        n19710) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19710), .B1(
        n19709), .B2(n19715), .ZN(n19687) );
  OAI211_X1 U22663 ( .C1(n19729), .C2(n19745), .A(n19688), .B(n19687), .ZN(
        P2_U3152) );
  AOI22_X1 U22664 ( .A1(n19708), .A2(n19775), .B1(n19774), .B2(n19707), .ZN(
        n19691) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19710), .B1(
        n19709), .B2(n19689), .ZN(n19690) );
  OAI211_X1 U22666 ( .C1(n19692), .C2(n19745), .A(n19691), .B(n19690), .ZN(
        P2_U3153) );
  AOI22_X1 U22667 ( .A1(n19708), .A2(n19781), .B1(n19780), .B2(n19707), .ZN(
        n19694) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19710), .B1(
        n19709), .B2(n19732), .ZN(n19693) );
  OAI211_X1 U22669 ( .C1(n19735), .C2(n19745), .A(n19694), .B(n19693), .ZN(
        P2_U3154) );
  AOI22_X1 U22670 ( .A1(n19708), .A2(n19787), .B1(n19786), .B2(n19707), .ZN(
        n19696) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19710), .B1(
        n19709), .B2(n19736), .ZN(n19695) );
  OAI211_X1 U22672 ( .C1(n19739), .C2(n19745), .A(n19696), .B(n19695), .ZN(
        P2_U3155) );
  AOI22_X1 U22673 ( .A1(n19708), .A2(n19793), .B1(n19792), .B2(n19707), .ZN(
        n19699) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19710), .B1(
        n19709), .B2(n19697), .ZN(n19698) );
  OAI211_X1 U22675 ( .C1(n19700), .C2(n19745), .A(n19699), .B(n19698), .ZN(
        P2_U3156) );
  AOI22_X1 U22676 ( .A1(n19708), .A2(n19798), .B1(n19301), .B2(n19707), .ZN(
        n19703) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19710), .B1(
        n19709), .B2(n19701), .ZN(n19702) );
  OAI211_X1 U22678 ( .C1(n19704), .C2(n19745), .A(n19703), .B(n19702), .ZN(
        P2_U3157) );
  AOI22_X1 U22679 ( .A1(n19708), .A2(n19804), .B1(n19803), .B2(n19707), .ZN(
        n19706) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19710), .B1(
        n19709), .B2(n19746), .ZN(n19705) );
  OAI211_X1 U22681 ( .C1(n19749), .C2(n19745), .A(n19706), .B(n19705), .ZN(
        P2_U3158) );
  AOI22_X1 U22682 ( .A1(n19708), .A2(n19811), .B1(n19810), .B2(n19707), .ZN(
        n19712) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19710), .B1(
        n19709), .B2(n19752), .ZN(n19711) );
  OAI211_X1 U22684 ( .C1(n19757), .C2(n19745), .A(n19712), .B(n19711), .ZN(
        P2_U3159) );
  INV_X1 U22685 ( .A(n19713), .ZN(n19714) );
  NAND2_X1 U22686 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19717), .ZN(
        n19766) );
  NOR2_X1 U22687 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19766), .ZN(
        n19750) );
  AOI22_X1 U22688 ( .A1(n19715), .A2(n19751), .B1(n19761), .B2(n19750), .ZN(
        n19728) );
  OAI21_X1 U22689 ( .B1(n19751), .B2(n19742), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19716) );
  NAND2_X1 U22690 ( .A1(n19716), .A2(n19934), .ZN(n19726) );
  AND2_X1 U22691 ( .A1(n19718), .A2(n19717), .ZN(n19722) );
  INV_X1 U22692 ( .A(n19750), .ZN(n19719) );
  OAI211_X1 U22693 ( .C1(n19720), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19719), 
        .B(n19913), .ZN(n19721) );
  OAI211_X1 U22694 ( .C1(n19726), .C2(n19722), .A(n19768), .B(n19721), .ZN(
        n19754) );
  INV_X1 U22695 ( .A(n19722), .ZN(n19725) );
  OAI21_X1 U22696 ( .B1(n19723), .B2(n19750), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19724) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19754), .B1(
        n19762), .B2(n19753), .ZN(n19727) );
  OAI211_X1 U22698 ( .C1(n19729), .C2(n19818), .A(n19728), .B(n19727), .ZN(
        P2_U3160) );
  AOI22_X1 U22699 ( .A1(n19742), .A2(n19776), .B1(n19774), .B2(n19750), .ZN(
        n19731) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19754), .B1(
        n19775), .B2(n19753), .ZN(n19730) );
  OAI211_X1 U22701 ( .C1(n19779), .C2(n19745), .A(n19731), .B(n19730), .ZN(
        P2_U3161) );
  AOI22_X1 U22702 ( .A1(n19732), .A2(n19751), .B1(n19780), .B2(n19750), .ZN(
        n19734) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19754), .B1(
        n19781), .B2(n19753), .ZN(n19733) );
  OAI211_X1 U22704 ( .C1(n19735), .C2(n19818), .A(n19734), .B(n19733), .ZN(
        P2_U3162) );
  AOI22_X1 U22705 ( .A1(n19736), .A2(n19751), .B1(n19786), .B2(n19750), .ZN(
        n19738) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19754), .B1(
        n19787), .B2(n19753), .ZN(n19737) );
  OAI211_X1 U22707 ( .C1(n19739), .C2(n19818), .A(n19738), .B(n19737), .ZN(
        P2_U3163) );
  AOI22_X1 U22708 ( .A1(n19794), .A2(n19742), .B1(n19792), .B2(n19750), .ZN(
        n19741) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19754), .B1(
        n19793), .B2(n19753), .ZN(n19740) );
  OAI211_X1 U22710 ( .C1(n19797), .C2(n19745), .A(n19741), .B(n19740), .ZN(
        P2_U3164) );
  AOI22_X1 U22711 ( .A1(n19742), .A2(n19799), .B1(n19301), .B2(n19750), .ZN(
        n19744) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19754), .B1(
        n19798), .B2(n19753), .ZN(n19743) );
  OAI211_X1 U22713 ( .C1(n19802), .C2(n19745), .A(n19744), .B(n19743), .ZN(
        P2_U3165) );
  AOI22_X1 U22714 ( .A1(n19751), .A2(n19746), .B1(n19803), .B2(n19750), .ZN(
        n19748) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19754), .B1(
        n19804), .B2(n19753), .ZN(n19747) );
  OAI211_X1 U22716 ( .C1(n19749), .C2(n19818), .A(n19748), .B(n19747), .ZN(
        P2_U3166) );
  AOI22_X1 U22717 ( .A1(n19752), .A2(n19751), .B1(n19810), .B2(n19750), .ZN(
        n19756) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19754), .B1(
        n19811), .B2(n19753), .ZN(n19755) );
  OAI211_X1 U22719 ( .C1(n19757), .C2(n19818), .A(n19756), .B(n19755), .ZN(
        P2_U3167) );
  NOR3_X1 U22720 ( .A1(n19758), .A2(n19809), .A3(n19973), .ZN(n19765) );
  INV_X1 U22721 ( .A(n19766), .ZN(n19759) );
  AOI21_X1 U22722 ( .B1(n19533), .B2(n19759), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19760) );
  NOR2_X1 U22723 ( .A1(n19765), .A2(n19760), .ZN(n19812) );
  AOI22_X1 U22724 ( .A1(n19812), .A2(n19762), .B1(n19761), .B2(n19809), .ZN(
        n19772) );
  NAND2_X1 U22725 ( .A1(n19764), .A2(n19763), .ZN(n19767) );
  AOI21_X1 U22726 ( .B1(n19767), .B2(n19766), .A(n19765), .ZN(n19769) );
  OAI211_X1 U22727 ( .C1(n19809), .C2(n19533), .A(n19769), .B(n19768), .ZN(
        n19815) );
  AOI22_X1 U22728 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19770), .ZN(n19771) );
  OAI211_X1 U22729 ( .C1(n19773), .C2(n19818), .A(n19772), .B(n19771), .ZN(
        P2_U3168) );
  AOI22_X1 U22730 ( .A1(n19812), .A2(n19775), .B1(n19774), .B2(n19809), .ZN(
        n19778) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19776), .ZN(n19777) );
  OAI211_X1 U22732 ( .C1(n19779), .C2(n19818), .A(n19778), .B(n19777), .ZN(
        P2_U3169) );
  AOI22_X1 U22733 ( .A1(n19812), .A2(n19781), .B1(n19780), .B2(n19809), .ZN(
        n19784) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19782), .ZN(n19783) );
  OAI211_X1 U22735 ( .C1(n19785), .C2(n19818), .A(n19784), .B(n19783), .ZN(
        P2_U3170) );
  AOI22_X1 U22736 ( .A1(n19812), .A2(n19787), .B1(n19786), .B2(n19809), .ZN(
        n19790) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19788), .ZN(n19789) );
  OAI211_X1 U22738 ( .C1(n19791), .C2(n19818), .A(n19790), .B(n19789), .ZN(
        P2_U3171) );
  AOI22_X1 U22739 ( .A1(n19812), .A2(n19793), .B1(n19792), .B2(n19809), .ZN(
        n19796) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19794), .ZN(n19795) );
  OAI211_X1 U22741 ( .C1(n19797), .C2(n19818), .A(n19796), .B(n19795), .ZN(
        P2_U3172) );
  AOI22_X1 U22742 ( .A1(n19812), .A2(n19798), .B1(n19301), .B2(n19809), .ZN(
        n19801) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19799), .ZN(n19800) );
  OAI211_X1 U22744 ( .C1(n19802), .C2(n19818), .A(n19801), .B(n19800), .ZN(
        P2_U3173) );
  AOI22_X1 U22745 ( .A1(n19812), .A2(n19804), .B1(n19803), .B2(n19809), .ZN(
        n19807) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19805), .ZN(n19806) );
  OAI211_X1 U22747 ( .C1(n19808), .C2(n19818), .A(n19807), .B(n19806), .ZN(
        P2_U3174) );
  AOI22_X1 U22748 ( .A1(n19812), .A2(n19811), .B1(n19810), .B2(n19809), .ZN(
        n19817) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n19813), .ZN(n19816) );
  OAI211_X1 U22750 ( .C1(n19819), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        P2_U3175) );
  OAI211_X1 U22751 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19822), .A(n19821), 
        .B(n19820), .ZN(n19827) );
  NOR2_X1 U22752 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19969), .ZN(n19823) );
  OAI211_X1 U22753 ( .C1(n19824), .C2(n19823), .A(n19974), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19826) );
  OAI211_X1 U22754 ( .C1(n19828), .C2(n19827), .A(n19826), .B(n19825), .ZN(
        P2_U3177) );
  AND2_X1 U22755 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19834), .ZN(
        P2_U3179) );
  NOR2_X1 U22756 ( .A1(n19829), .A2(n19911), .ZN(P2_U3180) );
  NOR2_X1 U22757 ( .A1(n19830), .A2(n19911), .ZN(P2_U3181) );
  AND2_X1 U22758 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19834), .ZN(
        P2_U3182) );
  AND2_X1 U22759 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19834), .ZN(
        P2_U3183) );
  AND2_X1 U22760 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19834), .ZN(
        P2_U3184) );
  AND2_X1 U22761 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19834), .ZN(
        P2_U3185) );
  AND2_X1 U22762 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19834), .ZN(
        P2_U3186) );
  AND2_X1 U22763 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19834), .ZN(
        P2_U3187) );
  NOR2_X1 U22764 ( .A1(n19831), .A2(n19911), .ZN(P2_U3188) );
  AND2_X1 U22765 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19834), .ZN(
        P2_U3189) );
  AND2_X1 U22766 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19834), .ZN(
        P2_U3190) );
  AND2_X1 U22767 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19834), .ZN(
        P2_U3191) );
  AND2_X1 U22768 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19834), .ZN(
        P2_U3192) );
  AND2_X1 U22769 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19834), .ZN(
        P2_U3193) );
  AND2_X1 U22770 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19834), .ZN(
        P2_U3194) );
  AND2_X1 U22771 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19834), .ZN(
        P2_U3195) );
  AND2_X1 U22772 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19834), .ZN(
        P2_U3196) );
  AND2_X1 U22773 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19834), .ZN(
        P2_U3197) );
  AND2_X1 U22774 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19834), .ZN(
        P2_U3198) );
  AND2_X1 U22775 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19834), .ZN(
        P2_U3199) );
  AND2_X1 U22776 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19834), .ZN(
        P2_U3200) );
  NOR2_X1 U22777 ( .A1(n19832), .A2(n19911), .ZN(P2_U3201) );
  AND2_X1 U22778 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19834), .ZN(P2_U3202) );
  AND2_X1 U22779 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19834), .ZN(P2_U3203) );
  AND2_X1 U22780 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19834), .ZN(P2_U3204) );
  AND2_X1 U22781 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19834), .ZN(P2_U3205) );
  NOR2_X1 U22782 ( .A1(n19833), .A2(n19911), .ZN(P2_U3206) );
  AND2_X1 U22783 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19834), .ZN(P2_U3207) );
  AND2_X1 U22784 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19834), .ZN(P2_U3208) );
  INV_X1 U22785 ( .A(NA), .ZN(n20778) );
  NOR2_X1 U22786 ( .A1(n20778), .A2(n19840), .ZN(n19851) );
  INV_X1 U22787 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19980) );
  NOR2_X1 U22788 ( .A1(n19835), .A2(n19980), .ZN(n19836) );
  NAND2_X1 U22789 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19974), .ZN(n19846) );
  AOI21_X1 U22790 ( .B1(n19836), .B2(n19846), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19839) );
  AOI211_X1 U22791 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20773), .A(
        n19837), .B(n19985), .ZN(n19838) );
  OR3_X1 U22792 ( .A1(n19851), .A2(n19839), .A3(n19838), .ZN(P2_U3209) );
  AOI21_X1 U22793 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20773), .A(n19852), 
        .ZN(n19844) );
  NOR2_X1 U22794 ( .A1(n19980), .A2(n19844), .ZN(n19841) );
  AOI21_X1 U22795 ( .B1(n19841), .B2(n19840), .A(n19970), .ZN(n19842) );
  OAI211_X1 U22796 ( .C1(n20773), .C2(n19843), .A(n19842), .B(n19846), .ZN(
        P2_U3210) );
  AOI21_X1 U22797 ( .B1(n19974), .B2(n19845), .A(n19844), .ZN(n19850) );
  OAI22_X1 U22798 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19847), .B1(NA), 
        .B2(n19846), .ZN(n19848) );
  OAI211_X1 U22799 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19848), .ZN(n19849) );
  OAI21_X1 U22800 ( .B1(n19851), .B2(n19850), .A(n19849), .ZN(P2_U3211) );
  OAI222_X1 U22801 ( .A1(n19901), .A2(n19855), .B1(n19854), .B2(n19985), .C1(
        n19853), .C2(n19898), .ZN(P2_U3212) );
  OAI222_X1 U22802 ( .A1(n19901), .A2(n11214), .B1(n19856), .B2(n19985), .C1(
        n19855), .C2(n19898), .ZN(P2_U3213) );
  OAI222_X1 U22803 ( .A1(n19901), .A2(n11221), .B1(n19857), .B2(n19985), .C1(
        n11214), .C2(n19898), .ZN(P2_U3214) );
  INV_X1 U22804 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19859) );
  OAI222_X1 U22805 ( .A1(n19901), .A2(n19859), .B1(n19858), .B2(n19985), .C1(
        n11221), .C2(n19898), .ZN(P2_U3215) );
  OAI222_X1 U22806 ( .A1(n19901), .A2(n19861), .B1(n19860), .B2(n19985), .C1(
        n19859), .C2(n19898), .ZN(P2_U3216) );
  OAI222_X1 U22807 ( .A1(n19901), .A2(n19863), .B1(n19862), .B2(n19985), .C1(
        n19861), .C2(n19898), .ZN(P2_U3217) );
  INV_X1 U22808 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19865) );
  OAI222_X1 U22809 ( .A1(n19901), .A2(n19865), .B1(n19864), .B2(n19985), .C1(
        n19863), .C2(n19898), .ZN(P2_U3218) );
  OAI222_X1 U22810 ( .A1(n19901), .A2(n11264), .B1(n19866), .B2(n19985), .C1(
        n19865), .C2(n19898), .ZN(P2_U3219) );
  OAI222_X1 U22811 ( .A1(n19901), .A2(n11267), .B1(n19867), .B2(n19985), .C1(
        n11264), .C2(n19898), .ZN(P2_U3220) );
  OAI222_X1 U22812 ( .A1(n19901), .A2(n11291), .B1(n19868), .B2(n19985), .C1(
        n11267), .C2(n19898), .ZN(P2_U3221) );
  OAI222_X1 U22813 ( .A1(n19901), .A2(n11295), .B1(n19869), .B2(n19985), .C1(
        n11291), .C2(n19898), .ZN(P2_U3222) );
  OAI222_X1 U22814 ( .A1(n19901), .A2(n19871), .B1(n19870), .B2(n19985), .C1(
        n11295), .C2(n19898), .ZN(P2_U3223) );
  INV_X1 U22815 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19873) );
  OAI222_X1 U22816 ( .A1(n19901), .A2(n19873), .B1(n19872), .B2(n19985), .C1(
        n19871), .C2(n19898), .ZN(P2_U3224) );
  OAI222_X1 U22817 ( .A1(n19901), .A2(n18940), .B1(n19874), .B2(n19985), .C1(
        n19873), .C2(n19898), .ZN(P2_U3225) );
  OAI222_X1 U22818 ( .A1(n19901), .A2(n15264), .B1(n19875), .B2(n19985), .C1(
        n18940), .C2(n19898), .ZN(P2_U3226) );
  OAI222_X1 U22819 ( .A1(n19901), .A2(n19877), .B1(n19876), .B2(n19985), .C1(
        n15264), .C2(n19898), .ZN(P2_U3227) );
  OAI222_X1 U22820 ( .A1(n19901), .A2(n12405), .B1(n19878), .B2(n19985), .C1(
        n19877), .C2(n19898), .ZN(P2_U3228) );
  OAI222_X1 U22821 ( .A1(n19901), .A2(n19880), .B1(n19879), .B2(n19985), .C1(
        n12405), .C2(n19898), .ZN(P2_U3229) );
  OAI222_X1 U22822 ( .A1(n19901), .A2(n15116), .B1(n19881), .B2(n19985), .C1(
        n19880), .C2(n19898), .ZN(P2_U3230) );
  OAI222_X1 U22823 ( .A1(n19901), .A2(n19883), .B1(n19882), .B2(n19985), .C1(
        n15116), .C2(n19898), .ZN(P2_U3231) );
  OAI222_X1 U22824 ( .A1(n19901), .A2(n12550), .B1(n19884), .B2(n19985), .C1(
        n19883), .C2(n19898), .ZN(P2_U3232) );
  OAI222_X1 U22825 ( .A1(n19901), .A2(n19886), .B1(n19885), .B2(n19985), .C1(
        n12550), .C2(n19898), .ZN(P2_U3233) );
  OAI222_X1 U22826 ( .A1(n19901), .A2(n12555), .B1(n19887), .B2(n19985), .C1(
        n19886), .C2(n19898), .ZN(P2_U3234) );
  OAI222_X1 U22827 ( .A1(n19901), .A2(n19889), .B1(n19888), .B2(n19985), .C1(
        n12555), .C2(n19898), .ZN(P2_U3235) );
  OAI222_X1 U22828 ( .A1(n19901), .A2(n15066), .B1(n19890), .B2(n19985), .C1(
        n19889), .C2(n19898), .ZN(P2_U3236) );
  OAI222_X1 U22829 ( .A1(n19901), .A2(n19893), .B1(n19891), .B2(n19985), .C1(
        n15066), .C2(n19898), .ZN(P2_U3237) );
  OAI222_X1 U22830 ( .A1(n19898), .A2(n19893), .B1(n19892), .B2(n19985), .C1(
        n19894), .C2(n19901), .ZN(P2_U3238) );
  OAI222_X1 U22831 ( .A1(n19901), .A2(n19896), .B1(n19895), .B2(n19985), .C1(
        n19894), .C2(n19898), .ZN(P2_U3239) );
  OAI222_X1 U22832 ( .A1(n19901), .A2(n14308), .B1(n19897), .B2(n19985), .C1(
        n19896), .C2(n19898), .ZN(P2_U3240) );
  INV_X1 U22833 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19900) );
  OAI222_X1 U22834 ( .A1(n19901), .A2(n19900), .B1(n19899), .B2(n19985), .C1(
        n14308), .C2(n19898), .ZN(P2_U3241) );
  AOI22_X1 U22835 ( .A1(n19985), .A2(n19903), .B1(n19902), .B2(n19982), .ZN(
        P2_U3585) );
  MUX2_X1 U22836 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19985), .Z(P2_U3586) );
  INV_X1 U22837 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19904) );
  AOI22_X1 U22838 ( .A1(n19985), .A2(n19905), .B1(n19904), .B2(n19982), .ZN(
        P2_U3587) );
  INV_X1 U22839 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19906) );
  AOI22_X1 U22840 ( .A1(n19985), .A2(n19907), .B1(n19906), .B2(n19982), .ZN(
        P2_U3588) );
  OAI21_X1 U22841 ( .B1(n19911), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19909), 
        .ZN(n19908) );
  INV_X1 U22842 ( .A(n19908), .ZN(P2_U3591) );
  OAI21_X1 U22843 ( .B1(n19911), .B2(n19910), .A(n19909), .ZN(P2_U3592) );
  NAND2_X1 U22844 ( .A1(n19912), .A2(n19934), .ZN(n19922) );
  OR3_X1 U22845 ( .A1(n19915), .A2(n19914), .A3(n19913), .ZN(n19927) );
  NAND3_X1 U22846 ( .A1(n19917), .A2(n19916), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19918) );
  NAND2_X1 U22847 ( .A1(n19918), .A2(n19935), .ZN(n19928) );
  NAND2_X1 U22848 ( .A1(n19927), .A2(n19928), .ZN(n19919) );
  NAND2_X1 U22849 ( .A1(n19920), .A2(n19919), .ZN(n19921) );
  OAI211_X1 U22850 ( .C1(n19923), .C2(n19533), .A(n19922), .B(n19921), .ZN(
        n19924) );
  INV_X1 U22851 ( .A(n19924), .ZN(n19925) );
  AOI22_X1 U22852 ( .A1(n19951), .A2(n19926), .B1(n19925), .B2(n19948), .ZN(
        P2_U3602) );
  OAI21_X1 U22853 ( .B1(n19929), .B2(n19928), .A(n19927), .ZN(n19930) );
  AOI21_X1 U22854 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19931), .A(n19930), 
        .ZN(n19932) );
  AOI22_X1 U22855 ( .A1(n19951), .A2(n19933), .B1(n19932), .B2(n19948), .ZN(
        P2_U3603) );
  NAND3_X1 U22856 ( .A1(n19937), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19934), 
        .ZN(n19939) );
  INV_X1 U22857 ( .A(n19935), .ZN(n19944) );
  OR3_X1 U22858 ( .A1(n19937), .A2(n19944), .A3(n19936), .ZN(n19938) );
  NAND2_X1 U22859 ( .A1(n19939), .A2(n19938), .ZN(n19940) );
  AOI21_X1 U22860 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19941), .A(n19940), 
        .ZN(n19942) );
  AOI22_X1 U22861 ( .A1(n19951), .A2(n19943), .B1(n19942), .B2(n19948), .ZN(
        P2_U3604) );
  OAI22_X1 U22862 ( .A1(n19945), .A2(n19944), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19533), .ZN(n19946) );
  AOI21_X1 U22863 ( .B1(n19947), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19946), 
        .ZN(n19949) );
  AOI22_X1 U22864 ( .A1(n19951), .A2(n19950), .B1(n19949), .B2(n19948), .ZN(
        P2_U3605) );
  AOI22_X1 U22865 ( .A1(n19985), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19952), 
        .B2(n19982), .ZN(P2_U3608) );
  INV_X1 U22866 ( .A(n19953), .ZN(n19962) );
  INV_X1 U22867 ( .A(n19954), .ZN(n19958) );
  AOI22_X1 U22868 ( .A1(n19958), .A2(n19957), .B1(n19956), .B2(n19955), .ZN(
        n19961) );
  NOR2_X1 U22869 ( .A1(n19962), .A2(n19959), .ZN(n19960) );
  AOI22_X1 U22870 ( .A1(n16349), .A2(n19962), .B1(n19961), .B2(n19960), .ZN(
        P2_U3609) );
  OAI21_X1 U22871 ( .B1(n19963), .B2(n19973), .A(n19533), .ZN(n19964) );
  OAI211_X1 U22872 ( .C1(n19966), .C2(n19974), .A(n19965), .B(n19964), .ZN(
        n19981) );
  AOI21_X1 U22873 ( .B1(n19970), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19967), 
        .ZN(n19972) );
  NOR3_X1 U22874 ( .A1(n19970), .A2(n19969), .A3(n19968), .ZN(n19971) );
  MUX2_X1 U22875 ( .A(n19972), .B(n19971), .S(n11196), .Z(n19978) );
  OAI22_X1 U22876 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19975), .B1(n19974), 
        .B2(n19973), .ZN(n19976) );
  INV_X1 U22877 ( .A(n19976), .ZN(n19977) );
  OAI21_X1 U22878 ( .B1(n19978), .B2(n19977), .A(n19981), .ZN(n19979) );
  OAI21_X1 U22879 ( .B1(n19981), .B2(n19980), .A(n19979), .ZN(P2_U3610) );
  INV_X1 U22880 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19983) );
  AOI22_X1 U22881 ( .A1(n19985), .A2(n19984), .B1(n19983), .B2(n19982), .ZN(
        P2_U3611) );
  NAND2_X1 U22882 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(n19986), .ZN(n19989)
         );
  INV_X1 U22883 ( .A(n19987), .ZN(n19995) );
  NAND3_X1 U22884 ( .A1(n19989), .A2(n19995), .A3(n19988), .ZN(P1_U2801) );
  AOI21_X1 U22885 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20781), .A(n20772), 
        .ZN(n20774) );
  INV_X1 U22886 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19990) );
  NAND2_X1 U22887 ( .A1(n20772), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20860) );
  INV_X2 U22888 ( .A(n20860), .ZN(n20832) );
  AOI21_X1 U22889 ( .B1(n20774), .B2(n19990), .A(n20832), .ZN(P1_U2802) );
  INV_X1 U22890 ( .A(n19991), .ZN(n19993) );
  OAI21_X1 U22891 ( .B1(n19993), .B2(n19992), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19994) );
  OAI21_X1 U22892 ( .B1(n19995), .B2(n20761), .A(n19994), .ZN(P1_U2803) );
  NOR2_X1 U22893 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19997) );
  OAI21_X1 U22894 ( .B1(n19997), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20860), .ZN(
        n19996) );
  OAI21_X1 U22895 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20860), .A(n19996), 
        .ZN(P1_U2804) );
  NOR2_X1 U22896 ( .A1(n20774), .A2(n20832), .ZN(n20851) );
  OAI21_X1 U22897 ( .B1(BS16), .B2(n19997), .A(n20851), .ZN(n20849) );
  OAI21_X1 U22898 ( .B1(n20851), .B2(n20633), .A(n20849), .ZN(P1_U2805) );
  OAI21_X1 U22899 ( .B1(n19999), .B2(n19998), .A(n20158), .ZN(P1_U2806) );
  NOR4_X1 U22900 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20003) );
  NOR4_X1 U22901 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20002) );
  NOR4_X1 U22902 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20001) );
  NOR4_X1 U22903 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20000) );
  NAND4_X1 U22904 ( .A1(n20003), .A2(n20002), .A3(n20001), .A4(n20000), .ZN(
        n20009) );
  NOR4_X1 U22905 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20007) );
  AOI211_X1 U22906 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_16__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20006) );
  NOR4_X1 U22907 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20005) );
  NOR4_X1 U22908 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20004) );
  NAND4_X1 U22909 ( .A1(n20007), .A2(n20006), .A3(n20005), .A4(n20004), .ZN(
        n20008) );
  NOR2_X1 U22910 ( .A1(n20009), .A2(n20008), .ZN(n20856) );
  INV_X1 U22911 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20844) );
  NOR3_X1 U22912 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20011) );
  OAI21_X1 U22913 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20011), .A(n20856), .ZN(
        n20010) );
  OAI21_X1 U22914 ( .B1(n20856), .B2(n20844), .A(n20010), .ZN(P1_U2807) );
  INV_X1 U22915 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20850) );
  AOI21_X1 U22916 ( .B1(n20852), .B2(n20850), .A(n20011), .ZN(n20012) );
  INV_X1 U22917 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20841) );
  INV_X1 U22918 ( .A(n20856), .ZN(n20858) );
  AOI22_X1 U22919 ( .A1(n20856), .A2(n20012), .B1(n20841), .B2(n20858), .ZN(
        P1_U2808) );
  INV_X1 U22920 ( .A(n20013), .ZN(n20018) );
  AOI22_X1 U22921 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n20093), .B1(n20099), .B2(
        n20014), .ZN(n20015) );
  OAI211_X1 U22922 ( .C1(n20064), .C2(n20016), .A(n20015), .B(n20177), .ZN(
        n20017) );
  AOI221_X1 U22923 ( .B1(n20027), .B2(P1_REIP_REG_9__SCAN_IN), .C1(n20018), 
        .C2(n20796), .A(n20017), .ZN(n20023) );
  INV_X1 U22924 ( .A(n20019), .ZN(n20021) );
  AOI22_X1 U22925 ( .A1(n20021), .A2(n20051), .B1(n20102), .B2(n20020), .ZN(
        n20022) );
  NAND2_X1 U22926 ( .A1(n20023), .A2(n20022), .ZN(P1_U2831) );
  OAI22_X1 U22927 ( .A1(n20064), .A2(n20025), .B1(n20024), .B2(n14034), .ZN(
        n20026) );
  AOI211_X1 U22928 ( .C1(n20027), .C2(P1_REIP_REG_8__SCAN_IN), .A(n16000), .B(
        n20026), .ZN(n20028) );
  OAI21_X1 U22929 ( .B1(n20030), .B2(n20029), .A(n20028), .ZN(n20031) );
  AOI21_X1 U22930 ( .B1(n20032), .B2(n20102), .A(n20031), .ZN(n20035) );
  INV_X1 U22931 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20792) );
  NAND2_X1 U22932 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20039) );
  NOR2_X1 U22933 ( .A1(n20792), .A2(n20039), .ZN(n20033) );
  NAND3_X1 U22934 ( .A1(n20033), .A2(n20067), .A3(n20793), .ZN(n20034) );
  OAI211_X1 U22935 ( .C1(n20036), .C2(n20081), .A(n20035), .B(n20034), .ZN(
        P1_U2832) );
  NOR2_X1 U22936 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20039), .ZN(n20037) );
  AOI22_X1 U22937 ( .A1(n20099), .A2(n20038), .B1(n20067), .B2(n20037), .ZN(
        n20046) );
  INV_X1 U22938 ( .A(n20039), .ZN(n20040) );
  AOI21_X1 U22939 ( .B1(n20040), .B2(n20059), .A(n20060), .ZN(n20050) );
  AOI22_X1 U22940 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n20093), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20050), .ZN(n20042) );
  NAND2_X1 U22941 ( .A1(n20092), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n20041) );
  NAND3_X1 U22942 ( .A1(n20042), .A2(n20177), .A3(n20041), .ZN(n20043) );
  AOI21_X1 U22943 ( .B1(n20051), .B2(n20044), .A(n20043), .ZN(n20045) );
  OAI211_X1 U22944 ( .C1(n20047), .C2(n20088), .A(n20046), .B(n20045), .ZN(
        P1_U2833) );
  INV_X1 U22945 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20789) );
  NOR2_X1 U22946 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20789), .ZN(n20048) );
  AOI22_X1 U22947 ( .A1(n20099), .A2(n20049), .B1(n20067), .B2(n20048), .ZN(
        n20057) );
  AOI22_X1 U22948 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n20093), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20050), .ZN(n20055) );
  NAND2_X1 U22949 ( .A1(n20052), .A2(n20051), .ZN(n20054) );
  NAND2_X1 U22950 ( .A1(n20092), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20053) );
  AND4_X1 U22951 ( .A1(n20055), .A2(n20054), .A3(n20177), .A4(n20053), .ZN(
        n20056) );
  OAI211_X1 U22952 ( .C1(n20058), .C2(n20088), .A(n20057), .B(n20056), .ZN(
        P1_U2834) );
  NOR2_X1 U22953 ( .A1(n20060), .A2(n20059), .ZN(n20084) );
  AOI22_X1 U22954 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n20093), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20084), .ZN(n20072) );
  INV_X1 U22955 ( .A(n20061), .ZN(n20062) );
  NAND2_X1 U22956 ( .A1(n20099), .A2(n20062), .ZN(n20063) );
  OAI211_X1 U22957 ( .C1(n20065), .C2(n20064), .A(n20177), .B(n20063), .ZN(
        n20066) );
  AOI21_X1 U22958 ( .B1(n20067), .B2(n20789), .A(n20066), .ZN(n20071) );
  INV_X1 U22959 ( .A(n20068), .ZN(n20069) );
  NAND2_X1 U22960 ( .A1(n20069), .A2(n20104), .ZN(n20070) );
  AND3_X1 U22961 ( .A1(n20072), .A2(n20071), .A3(n20070), .ZN(n20073) );
  OAI21_X1 U22962 ( .B1(n20074), .B2(n20088), .A(n20073), .ZN(P1_U2835) );
  NAND3_X1 U22963 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .ZN(n20075) );
  NOR3_X1 U22964 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20091), .A3(n20075), .ZN(
        n20083) );
  INV_X1 U22965 ( .A(n20076), .ZN(n20078) );
  AOI22_X1 U22966 ( .A1(n20078), .A2(n20077), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20092), .ZN(n20079) );
  OAI211_X1 U22967 ( .C1(n20081), .C2(n20080), .A(n20079), .B(n20177), .ZN(
        n20082) );
  AOI211_X1 U22968 ( .C1(n20093), .C2(P1_EBX_REG_4__SCAN_IN), .A(n20083), .B(
        n20082), .ZN(n20087) );
  AOI22_X1 U22969 ( .A1(n20085), .A2(n20104), .B1(n20084), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20086) );
  OAI211_X1 U22970 ( .C1(n20089), .C2(n20088), .A(n20087), .B(n20086), .ZN(
        P1_U2836) );
  NAND2_X1 U22971 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n20090) );
  NOR3_X1 U22972 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20091), .A3(n20090), .ZN(
        n20098) );
  INV_X1 U22973 ( .A(n13653), .ZN(n20096) );
  AOI22_X1 U22974 ( .A1(n20093), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20092), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20094) );
  OAI21_X1 U22975 ( .B1(n20096), .B2(n20095), .A(n20094), .ZN(n20097) );
  AOI211_X1 U22976 ( .C1(n20100), .C2(n20099), .A(n20098), .B(n20097), .ZN(
        n20107) );
  INV_X1 U22977 ( .A(n20101), .ZN(n20103) );
  AOI22_X1 U22978 ( .A1(n20105), .A2(n20104), .B1(n20103), .B2(n20102), .ZN(
        n20106) );
  OAI211_X1 U22979 ( .C1(n20108), .C2(n13769), .A(n20107), .B(n20106), .ZN(
        P1_U2837) );
  INV_X1 U22980 ( .A(n20109), .ZN(n20110) );
  AOI22_X1 U22981 ( .A1(n20144), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n20110), 
        .B2(P1_EAX_REG_29__SCAN_IN), .ZN(n20111) );
  OAI21_X1 U22982 ( .B1(n20150), .B2(n20133), .A(n20111), .ZN(P1_U2907) );
  AOI22_X1 U22983 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20120), .B1(n20144), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20112) );
  OAI21_X1 U22984 ( .B1(n20113), .B2(n20133), .A(n20112), .ZN(P1_U2921) );
  AOI22_X1 U22985 ( .A1(n9726), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20114) );
  OAI21_X1 U22986 ( .B1(n20115), .B2(n20146), .A(n20114), .ZN(P1_U2922) );
  AOI22_X1 U22987 ( .A1(n9726), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20116) );
  OAI21_X1 U22988 ( .B1(n20117), .B2(n20146), .A(n20116), .ZN(P1_U2923) );
  AOI22_X1 U22989 ( .A1(n9726), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20118) );
  OAI21_X1 U22990 ( .B1(n20119), .B2(n20146), .A(n20118), .ZN(P1_U2924) );
  AOI22_X1 U22991 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n20120), .B1(n9726), .B2(
        P1_LWORD_REG_11__SCAN_IN), .ZN(n20121) );
  OAI21_X1 U22992 ( .B1(n20122), .B2(n20135), .A(n20121), .ZN(P1_U2925) );
  AOI22_X1 U22993 ( .A1(n9726), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20123) );
  OAI21_X1 U22994 ( .B1(n20124), .B2(n20146), .A(n20123), .ZN(P1_U2926) );
  AOI22_X1 U22995 ( .A1(n9726), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20125) );
  OAI21_X1 U22996 ( .B1(n20126), .B2(n20146), .A(n20125), .ZN(P1_U2927) );
  AOI22_X1 U22997 ( .A1(n9726), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20127) );
  OAI21_X1 U22998 ( .B1(n20128), .B2(n20146), .A(n20127), .ZN(P1_U2928) );
  AOI22_X1 U22999 ( .A1(n9726), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20129) );
  OAI21_X1 U23000 ( .B1(n20130), .B2(n20146), .A(n20129), .ZN(P1_U2929) );
  AOI22_X1 U23001 ( .A1(n9726), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20131) );
  OAI21_X1 U23002 ( .B1(n11862), .B2(n20146), .A(n20131), .ZN(P1_U2930) );
  INV_X1 U23003 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n20132) );
  OAI222_X1 U23004 ( .A1(n20135), .A2(n20134), .B1(n20146), .B2(n11786), .C1(
        n20133), .C2(n20132), .ZN(P1_U2931) );
  AOI22_X1 U23005 ( .A1(n9726), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20136) );
  OAI21_X1 U23006 ( .B1(n20137), .B2(n20146), .A(n20136), .ZN(P1_U2932) );
  AOI22_X1 U23007 ( .A1(n9726), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20138) );
  OAI21_X1 U23008 ( .B1(n20139), .B2(n20146), .A(n20138), .ZN(P1_U2933) );
  AOI22_X1 U23009 ( .A1(n9726), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20140) );
  OAI21_X1 U23010 ( .B1(n20141), .B2(n20146), .A(n20140), .ZN(P1_U2934) );
  AOI22_X1 U23011 ( .A1(n9726), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20142) );
  OAI21_X1 U23012 ( .B1(n20143), .B2(n20146), .A(n20142), .ZN(P1_U2935) );
  AOI22_X1 U23013 ( .A1(n9726), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20144), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20145) );
  OAI21_X1 U23014 ( .B1(n20147), .B2(n20146), .A(n20145), .ZN(P1_U2936) );
  AOI21_X1 U23015 ( .B1(n20153), .B2(P1_EAX_REG_29__SCAN_IN), .A(n20148), .ZN(
        n20149) );
  OAI21_X1 U23016 ( .B1(n20151), .B2(n20150), .A(n20149), .ZN(P1_U2950) );
  AOI22_X1 U23017 ( .A1(n20153), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20152), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20155) );
  NAND2_X1 U23018 ( .A1(n20155), .A2(n20154), .ZN(P1_U2963) );
  INV_X1 U23019 ( .A(n20156), .ZN(n20159) );
  OAI22_X1 U23020 ( .A1(n20159), .A2(n20158), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20157), .ZN(n20160) );
  AOI211_X1 U23021 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20165), .A(
        n20161), .B(n20160), .ZN(n20162) );
  OAI21_X1 U23022 ( .B1(n20191), .B2(n20163), .A(n20162), .ZN(P1_U2998) );
  OR2_X1 U23023 ( .A1(n20165), .A2(n20164), .ZN(n20166) );
  AOI22_X1 U23024 ( .A1(n20168), .A2(n20167), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20166), .ZN(n20170) );
  OAI211_X1 U23025 ( .C1(n20171), .C2(n20191), .A(n20170), .B(n20169), .ZN(
        P1_U2999) );
  NOR2_X1 U23026 ( .A1(n20172), .A2(n13589), .ZN(n20174) );
  AOI21_X1 U23027 ( .B1(n20175), .B2(n20174), .A(n20173), .ZN(n20185) );
  INV_X1 U23028 ( .A(n20176), .ZN(n20183) );
  OAI22_X1 U23029 ( .A1(n20179), .A2(n20178), .B1(n20784), .B2(n20177), .ZN(
        n20180) );
  AOI211_X1 U23030 ( .C1(n20183), .C2(n20182), .A(n20181), .B(n20180), .ZN(
        n20184) );
  OAI221_X1 U23031 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20186), .C1(
        n12621), .C2(n20185), .A(n20184), .ZN(P1_U3029) );
  NOR2_X1 U23032 ( .A1(n20188), .A2(n20187), .ZN(P1_U3032) );
  NOR2_X2 U23033 ( .A1(n20191), .A2(n20189), .ZN(n20233) );
  NOR2_X2 U23034 ( .A1(n20191), .A2(n20190), .ZN(n20232) );
  AOI22_X1 U23035 ( .A1(DATAI_16_), .A2(n20233), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20232), .ZN(n20671) );
  AOI22_X1 U23036 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20232), .B1(DATAI_24_), 
        .B2(n20233), .ZN(n20710) );
  INV_X1 U23037 ( .A(n20710), .ZN(n20668) );
  NOR2_X2 U23038 ( .A1(n20235), .A2(n20196), .ZN(n20701) );
  NAND3_X1 U23039 ( .A1(n20549), .A2(n12247), .A3(n20587), .ZN(n20245) );
  NOR2_X1 U23040 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20245), .ZN(
        n20236) );
  AOI22_X1 U23041 ( .A1(n20732), .A2(n20668), .B1(n20701), .B2(n20236), .ZN(
        n20209) );
  INV_X1 U23042 ( .A(n20268), .ZN(n20197) );
  OAI21_X1 U23043 ( .B1(n20197), .B2(n20732), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20198) );
  NAND2_X1 U23044 ( .A1(n20198), .A2(n20636), .ZN(n20207) );
  OR2_X1 U23045 ( .A1(n13653), .A2(n20199), .ZN(n20299) );
  NOR2_X1 U23046 ( .A1(n20299), .A2(n20659), .ZN(n20204) );
  INV_X1 U23047 ( .A(n20519), .ZN(n20200) );
  OR2_X1 U23048 ( .A1(n20455), .A2(n20200), .ZN(n20338) );
  INV_X1 U23049 ( .A(n20236), .ZN(n20201) );
  AOI22_X1 U23050 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20338), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20201), .ZN(n20202) );
  NAND2_X1 U23051 ( .A1(n20205), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20660) );
  NAND2_X1 U23052 ( .A1(n20238), .A2(n20660), .ZN(n20452) );
  INV_X1 U23053 ( .A(n20452), .ZN(n20523) );
  OAI211_X1 U23054 ( .C1(n20207), .C2(n20204), .A(n20202), .B(n20523), .ZN(
        n20240) );
  NAND2_X1 U23055 ( .A1(n20238), .A2(n20203), .ZN(n20597) );
  INV_X1 U23056 ( .A(n20204), .ZN(n20206) );
  NOR2_X1 U23057 ( .A1(n20205), .A2(n20764), .ZN(n20521) );
  INV_X1 U23058 ( .A(n20521), .ZN(n20456) );
  OAI22_X1 U23059 ( .A1(n20207), .A2(n20206), .B1(n20456), .B2(n20338), .ZN(
        n20239) );
  AOI22_X1 U23060 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20240), .B1(
        n20700), .B2(n20239), .ZN(n20208) );
  OAI211_X1 U23061 ( .C1(n20671), .C2(n20268), .A(n20209), .B(n20208), .ZN(
        P1_U3033) );
  AOI22_X1 U23062 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20232), .B1(DATAI_17_), 
        .B2(n20233), .ZN(n20675) );
  AOI22_X1 U23063 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20232), .B1(DATAI_25_), 
        .B2(n20233), .ZN(n20716) );
  INV_X1 U23064 ( .A(n20716), .ZN(n20672) );
  NOR2_X2 U23065 ( .A1(n20235), .A2(n12214), .ZN(n20712) );
  AOI22_X1 U23066 ( .A1(n20732), .A2(n20672), .B1(n20712), .B2(n20236), .ZN(
        n20212) );
  NAND2_X1 U23067 ( .A1(n20238), .A2(n20210), .ZN(n20600) );
  AOI22_X1 U23068 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20240), .B1(
        n20711), .B2(n20239), .ZN(n20211) );
  OAI211_X1 U23069 ( .C1(n20675), .C2(n20268), .A(n20212), .B(n20211), .ZN(
        P1_U3034) );
  AOI22_X1 U23070 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20232), .B1(DATAI_18_), 
        .B2(n20233), .ZN(n20722) );
  NOR2_X2 U23071 ( .A1(n20213), .A2(n20235), .ZN(n20718) );
  AOI22_X1 U23072 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20232), .B1(DATAI_26_), 
        .B2(n20233), .ZN(n20499) );
  INV_X1 U23073 ( .A(n20499), .ZN(n20719) );
  AOI22_X1 U23074 ( .A1(n20236), .A2(n20718), .B1(n20732), .B2(n20719), .ZN(
        n20216) );
  NOR2_X2 U23075 ( .A1(n20342), .A2(n20214), .ZN(n20717) );
  AOI22_X1 U23076 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20240), .B1(
        n20717), .B2(n20239), .ZN(n20215) );
  OAI211_X1 U23077 ( .C1(n20722), .C2(n20268), .A(n20216), .B(n20215), .ZN(
        P1_U3035) );
  AOI22_X1 U23078 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20232), .B1(DATAI_19_), 
        .B2(n20233), .ZN(n20681) );
  AOI22_X1 U23079 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20232), .B1(DATAI_27_), 
        .B2(n20233), .ZN(n20728) );
  INV_X1 U23080 ( .A(n20728), .ZN(n20678) );
  NOR2_X2 U23081 ( .A1(n20235), .A2(n20217), .ZN(n20724) );
  AOI22_X1 U23082 ( .A1(n20732), .A2(n20678), .B1(n20724), .B2(n20236), .ZN(
        n20220) );
  NAND2_X1 U23083 ( .A1(n20238), .A2(n20218), .ZN(n20607) );
  AOI22_X1 U23084 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20240), .B1(
        n20723), .B2(n20239), .ZN(n20219) );
  OAI211_X1 U23085 ( .C1(n20681), .C2(n20268), .A(n20220), .B(n20219), .ZN(
        P1_U3036) );
  AOI22_X1 U23086 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20232), .B1(DATAI_20_), 
        .B2(n20233), .ZN(n20685) );
  AOI22_X1 U23087 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20232), .B1(DATAI_28_), 
        .B2(n20233), .ZN(n20736) );
  INV_X1 U23088 ( .A(n20736), .ZN(n20682) );
  NOR2_X2 U23089 ( .A1(n20235), .A2(n20221), .ZN(n20729) );
  AOI22_X1 U23090 ( .A1(n20732), .A2(n20682), .B1(n20729), .B2(n20236), .ZN(
        n20224) );
  NOR2_X2 U23091 ( .A1(n20342), .A2(n20222), .ZN(n20730) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20240), .B1(
        n20730), .B2(n20239), .ZN(n20223) );
  OAI211_X1 U23093 ( .C1(n20685), .C2(n20268), .A(n20224), .B(n20223), .ZN(
        P1_U3037) );
  AOI22_X1 U23094 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20232), .B1(DATAI_21_), 
        .B2(n20233), .ZN(n20742) );
  AOI22_X1 U23095 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20232), .B1(DATAI_29_), 
        .B2(n20233), .ZN(n20506) );
  INV_X1 U23096 ( .A(n20506), .ZN(n20739) );
  NOR2_X2 U23097 ( .A1(n20235), .A2(n11608), .ZN(n20737) );
  AOI22_X1 U23098 ( .A1(n20732), .A2(n20739), .B1(n20737), .B2(n20236), .ZN(
        n20227) );
  NOR2_X2 U23099 ( .A1(n20342), .A2(n20225), .ZN(n20738) );
  AOI22_X1 U23100 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20240), .B1(
        n20738), .B2(n20239), .ZN(n20226) );
  OAI211_X1 U23101 ( .C1(n20742), .C2(n20268), .A(n20227), .B(n20226), .ZN(
        P1_U3038) );
  AOI22_X1 U23102 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20232), .B1(DATAI_22_), 
        .B2(n20233), .ZN(n20748) );
  AOI22_X1 U23103 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20232), .B1(DATAI_30_), 
        .B2(n20233), .ZN(n20509) );
  INV_X1 U23104 ( .A(n20509), .ZN(n20745) );
  NOR2_X2 U23105 ( .A1(n20235), .A2(n20228), .ZN(n20743) );
  AOI22_X1 U23106 ( .A1(n20732), .A2(n20745), .B1(n20743), .B2(n20236), .ZN(
        n20231) );
  NOR2_X2 U23107 ( .A1(n20342), .A2(n20229), .ZN(n20744) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20240), .B1(
        n20744), .B2(n20239), .ZN(n20230) );
  OAI211_X1 U23109 ( .C1(n20748), .C2(n20268), .A(n20231), .B(n20230), .ZN(
        P1_U3039) );
  AOI22_X1 U23110 ( .A1(DATAI_23_), .A2(n20233), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20232), .ZN(n20759) );
  AOI22_X1 U23111 ( .A1(DATAI_31_), .A2(n20233), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20232), .ZN(n20516) );
  INV_X1 U23112 ( .A(n20516), .ZN(n20753) );
  NOR2_X2 U23113 ( .A1(n20235), .A2(n20234), .ZN(n20752) );
  AOI22_X1 U23114 ( .A1(n20732), .A2(n20753), .B1(n20752), .B2(n20236), .ZN(
        n20242) );
  NAND2_X1 U23115 ( .A1(n20238), .A2(n20237), .ZN(n20625) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20240), .B1(
        n20750), .B2(n20239), .ZN(n20241) );
  OAI211_X1 U23117 ( .C1(n20759), .C2(n20268), .A(n20242), .B(n20241), .ZN(
        P1_U3040) );
  NOR2_X1 U23118 ( .A1(n20628), .A2(n20245), .ZN(n20264) );
  INV_X1 U23119 ( .A(n20299), .ZN(n20244) );
  INV_X1 U23120 ( .A(n20243), .ZN(n20630) );
  AOI21_X1 U23121 ( .B1(n20244), .B2(n20630), .A(n20264), .ZN(n20246) );
  OAI22_X1 U23122 ( .A1(n20246), .A2(n20698), .B1(n20245), .B2(n20764), .ZN(
        n20263) );
  AOI22_X1 U23123 ( .A1(n20701), .A2(n20264), .B1(n20263), .B2(n20700), .ZN(
        n20250) );
  INV_X1 U23124 ( .A(n20245), .ZN(n20248) );
  OAI211_X1 U23125 ( .C1(n20307), .C2(n20633), .A(n20636), .B(n20246), .ZN(
        n20247) );
  OAI211_X1 U23126 ( .C1(n20636), .C2(n20248), .A(n20705), .B(n20247), .ZN(
        n20265) );
  OR2_X1 U23127 ( .A1(n9717), .A2(n20579), .ZN(n20368) );
  INV_X1 U23128 ( .A(n20671), .ZN(n20707) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20265), .B1(
        n20292), .B2(n20707), .ZN(n20249) );
  OAI211_X1 U23130 ( .C1(n20710), .C2(n20268), .A(n20250), .B(n20249), .ZN(
        P1_U3041) );
  AOI22_X1 U23131 ( .A1(n20712), .A2(n20264), .B1(n20263), .B2(n20711), .ZN(
        n20252) );
  INV_X1 U23132 ( .A(n20675), .ZN(n20713) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20265), .B1(
        n20292), .B2(n20713), .ZN(n20251) );
  OAI211_X1 U23134 ( .C1(n20716), .C2(n20268), .A(n20252), .B(n20251), .ZN(
        P1_U3042) );
  AOI22_X1 U23135 ( .A1(n20717), .A2(n20263), .B1(n20718), .B2(n20264), .ZN(
        n20254) );
  INV_X1 U23136 ( .A(n20722), .ZN(n20601) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20265), .B1(
        n20292), .B2(n20601), .ZN(n20253) );
  OAI211_X1 U23138 ( .C1(n20499), .C2(n20268), .A(n20254), .B(n20253), .ZN(
        P1_U3043) );
  AOI22_X1 U23139 ( .A1(n20724), .A2(n20264), .B1(n20263), .B2(n20723), .ZN(
        n20256) );
  INV_X1 U23140 ( .A(n20681), .ZN(n20725) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20265), .B1(
        n20292), .B2(n20725), .ZN(n20255) );
  OAI211_X1 U23142 ( .C1(n20728), .C2(n20268), .A(n20256), .B(n20255), .ZN(
        P1_U3044) );
  AOI22_X1 U23143 ( .A1(n20730), .A2(n20263), .B1(n20729), .B2(n20264), .ZN(
        n20258) );
  INV_X1 U23144 ( .A(n20685), .ZN(n20731) );
  AOI22_X1 U23145 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20265), .B1(
        n20292), .B2(n20731), .ZN(n20257) );
  OAI211_X1 U23146 ( .C1(n20736), .C2(n20268), .A(n20258), .B(n20257), .ZN(
        P1_U3045) );
  AOI22_X1 U23147 ( .A1(n20738), .A2(n20263), .B1(n20737), .B2(n20264), .ZN(
        n20260) );
  INV_X1 U23148 ( .A(n20742), .ZN(n20611) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20265), .B1(
        n20292), .B2(n20611), .ZN(n20259) );
  OAI211_X1 U23150 ( .C1(n20506), .C2(n20268), .A(n20260), .B(n20259), .ZN(
        P1_U3046) );
  AOI22_X1 U23151 ( .A1(n20744), .A2(n20263), .B1(n20743), .B2(n20264), .ZN(
        n20262) );
  INV_X1 U23152 ( .A(n20748), .ZN(n20615) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20265), .B1(
        n20292), .B2(n20615), .ZN(n20261) );
  OAI211_X1 U23154 ( .C1(n20509), .C2(n20268), .A(n20262), .B(n20261), .ZN(
        P1_U3047) );
  AOI22_X1 U23155 ( .A1(n20752), .A2(n20264), .B1(n20263), .B2(n20750), .ZN(
        n20267) );
  INV_X1 U23156 ( .A(n20759), .ZN(n20620) );
  AOI22_X1 U23157 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20265), .B1(
        n20292), .B2(n20620), .ZN(n20266) );
  OAI211_X1 U23158 ( .C1(n20516), .C2(n20268), .A(n20267), .B(n20266), .ZN(
        P1_U3048) );
  INV_X1 U23159 ( .A(n20292), .ZN(n20269) );
  NAND2_X1 U23160 ( .A1(n20269), .A2(n20636), .ZN(n20271) );
  OAI21_X1 U23161 ( .B1(n20271), .B2(n20330), .A(n20582), .ZN(n20272) );
  NOR2_X1 U23162 ( .A1(n20299), .A2(n20392), .ZN(n20275) );
  NAND3_X1 U23163 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20549), .A3(
        n12247), .ZN(n20304) );
  NOR2_X1 U23164 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20304), .ZN(
        n20291) );
  AOI22_X1 U23165 ( .A1(n20292), .A2(n20668), .B1(n20701), .B2(n20291), .ZN(
        n20278) );
  INV_X1 U23166 ( .A(n20272), .ZN(n20276) );
  INV_X1 U23167 ( .A(n20291), .ZN(n20273) );
  NOR2_X1 U23168 ( .A1(n10073), .A2(n20764), .ZN(n20395) );
  AOI211_X1 U23169 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20273), .A(n20395), 
        .B(n20452), .ZN(n20274) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20293), .B1(
        n20330), .B2(n20707), .ZN(n20277) );
  OAI211_X1 U23171 ( .C1(n20296), .C2(n20597), .A(n20278), .B(n20277), .ZN(
        P1_U3049) );
  AOI22_X1 U23172 ( .A1(n20330), .A2(n20713), .B1(n20291), .B2(n20712), .ZN(
        n20280) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20672), .ZN(n20279) );
  OAI211_X1 U23174 ( .C1(n20296), .C2(n20600), .A(n20280), .B(n20279), .ZN(
        P1_U3050) );
  INV_X1 U23175 ( .A(n20717), .ZN(n20604) );
  AOI22_X1 U23176 ( .A1(n20330), .A2(n20601), .B1(n20291), .B2(n20718), .ZN(
        n20282) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20719), .ZN(n20281) );
  OAI211_X1 U23178 ( .C1(n20296), .C2(n20604), .A(n20282), .B(n20281), .ZN(
        P1_U3051) );
  AOI22_X1 U23179 ( .A1(n20330), .A2(n20725), .B1(n20291), .B2(n20724), .ZN(
        n20284) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20678), .ZN(n20283) );
  OAI211_X1 U23181 ( .C1(n20296), .C2(n20607), .A(n20284), .B(n20283), .ZN(
        P1_U3052) );
  INV_X1 U23182 ( .A(n20730), .ZN(n20610) );
  AOI22_X1 U23183 ( .A1(n20292), .A2(n20682), .B1(n20291), .B2(n20729), .ZN(
        n20286) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20293), .B1(
        n20330), .B2(n20731), .ZN(n20285) );
  OAI211_X1 U23185 ( .C1(n20296), .C2(n20610), .A(n20286), .B(n20285), .ZN(
        P1_U3053) );
  INV_X1 U23186 ( .A(n20738), .ZN(n20614) );
  AOI22_X1 U23187 ( .A1(n20330), .A2(n20611), .B1(n20291), .B2(n20737), .ZN(
        n20288) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20739), .ZN(n20287) );
  OAI211_X1 U23189 ( .C1(n20296), .C2(n20614), .A(n20288), .B(n20287), .ZN(
        P1_U3054) );
  INV_X1 U23190 ( .A(n20744), .ZN(n20618) );
  AOI22_X1 U23191 ( .A1(n20330), .A2(n20615), .B1(n20291), .B2(n20743), .ZN(
        n20290) );
  AOI22_X1 U23192 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20293), .B1(
        n20292), .B2(n20745), .ZN(n20289) );
  OAI211_X1 U23193 ( .C1(n20296), .C2(n20618), .A(n20290), .B(n20289), .ZN(
        P1_U3055) );
  AOI22_X1 U23194 ( .A1(n20292), .A2(n20753), .B1(n20291), .B2(n20752), .ZN(
        n20295) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20293), .B1(
        n20330), .B2(n20620), .ZN(n20294) );
  OAI211_X1 U23196 ( .C1(n20296), .C2(n20625), .A(n20295), .B(n20294), .ZN(
        P1_U3056) );
  AOI21_X1 U23197 ( .B1(n20307), .B2(n20636), .A(n20556), .ZN(n20306) );
  AND2_X1 U23198 ( .A1(n20297), .A2(n11833), .ZN(n20696) );
  INV_X1 U23199 ( .A(n20696), .ZN(n20298) );
  OR2_X1 U23200 ( .A1(n20299), .A2(n20298), .ZN(n20301) );
  NOR2_X1 U23201 ( .A1(n20550), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20329) );
  INV_X1 U23202 ( .A(n20329), .ZN(n20300) );
  AND2_X1 U23203 ( .A1(n20301), .A2(n20300), .ZN(n20305) );
  INV_X1 U23204 ( .A(n20305), .ZN(n20302) );
  OAI21_X1 U23205 ( .B1(n20306), .B2(n20302), .A(n20705), .ZN(n20303) );
  AOI22_X1 U23206 ( .A1(n20330), .A2(n20668), .B1(n20701), .B2(n20329), .ZN(
        n20309) );
  OAI22_X1 U23207 ( .A1(n20306), .A2(n20305), .B1(n20764), .B2(n20304), .ZN(
        n20331) );
  AOI22_X1 U23208 ( .A1(n20700), .A2(n20331), .B1(n20360), .B2(n20707), .ZN(
        n20308) );
  OAI211_X1 U23209 ( .C1(n20335), .C2(n20310), .A(n20309), .B(n20308), .ZN(
        P1_U3057) );
  INV_X1 U23210 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n20313) );
  AOI22_X1 U23211 ( .A1(n20330), .A2(n20672), .B1(n20712), .B2(n20329), .ZN(
        n20312) );
  AOI22_X1 U23212 ( .A1(n20711), .A2(n20331), .B1(n20360), .B2(n20713), .ZN(
        n20311) );
  OAI211_X1 U23213 ( .C1(n20335), .C2(n20313), .A(n20312), .B(n20311), .ZN(
        P1_U3058) );
  INV_X1 U23214 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n20316) );
  AOI22_X1 U23215 ( .A1(n20329), .A2(n20718), .B1(n20360), .B2(n20601), .ZN(
        n20315) );
  AOI22_X1 U23216 ( .A1(n20330), .A2(n20719), .B1(n20717), .B2(n20331), .ZN(
        n20314) );
  OAI211_X1 U23217 ( .C1(n20335), .C2(n20316), .A(n20315), .B(n20314), .ZN(
        P1_U3059) );
  INV_X1 U23218 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n20319) );
  AOI22_X1 U23219 ( .A1(n20330), .A2(n20678), .B1(n20724), .B2(n20329), .ZN(
        n20318) );
  AOI22_X1 U23220 ( .A1(n20723), .A2(n20331), .B1(n20360), .B2(n20725), .ZN(
        n20317) );
  OAI211_X1 U23221 ( .C1(n20335), .C2(n20319), .A(n20318), .B(n20317), .ZN(
        P1_U3060) );
  INV_X1 U23222 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n20322) );
  AOI22_X1 U23223 ( .A1(n20330), .A2(n20682), .B1(n20729), .B2(n20329), .ZN(
        n20321) );
  AOI22_X1 U23224 ( .A1(n20730), .A2(n20331), .B1(n20360), .B2(n20731), .ZN(
        n20320) );
  OAI211_X1 U23225 ( .C1(n20335), .C2(n20322), .A(n20321), .B(n20320), .ZN(
        P1_U3061) );
  INV_X1 U23226 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n20325) );
  AOI22_X1 U23227 ( .A1(n20330), .A2(n20739), .B1(n20737), .B2(n20329), .ZN(
        n20324) );
  AOI22_X1 U23228 ( .A1(n20738), .A2(n20331), .B1(n20360), .B2(n20611), .ZN(
        n20323) );
  OAI211_X1 U23229 ( .C1(n20335), .C2(n20325), .A(n20324), .B(n20323), .ZN(
        P1_U3062) );
  INV_X1 U23230 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n20328) );
  AOI22_X1 U23231 ( .A1(n20330), .A2(n20745), .B1(n20743), .B2(n20329), .ZN(
        n20327) );
  AOI22_X1 U23232 ( .A1(n20744), .A2(n20331), .B1(n20360), .B2(n20615), .ZN(
        n20326) );
  OAI211_X1 U23233 ( .C1(n20335), .C2(n20328), .A(n20327), .B(n20326), .ZN(
        P1_U3063) );
  AOI22_X1 U23234 ( .A1(n20330), .A2(n20753), .B1(n20752), .B2(n20329), .ZN(
        n20333) );
  AOI22_X1 U23235 ( .A1(n20750), .A2(n20331), .B1(n20360), .B2(n20620), .ZN(
        n20332) );
  OAI211_X1 U23236 ( .C1(n20335), .C2(n20334), .A(n20333), .B(n20332), .ZN(
        P1_U3064) );
  NAND3_X1 U23237 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20549), .A3(
        n20587), .ZN(n20364) );
  NOR2_X1 U23238 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20364), .ZN(
        n20359) );
  OR2_X1 U23239 ( .A1(n13643), .A2(n20336), .ZN(n20393) );
  INV_X1 U23240 ( .A(n20393), .ZN(n20421) );
  NAND3_X1 U23241 ( .A1(n20421), .A2(n20636), .A3(n20392), .ZN(n20337) );
  OAI21_X1 U23242 ( .B1(n20660), .B2(n20338), .A(n20337), .ZN(n20358) );
  AOI22_X1 U23243 ( .A1(n20701), .A2(n20359), .B1(n20700), .B2(n20358), .ZN(
        n20345) );
  INV_X1 U23244 ( .A(n20360), .ZN(n20339) );
  AOI21_X1 U23245 ( .B1(n20339), .B2(n20388), .A(n20633), .ZN(n20340) );
  AOI21_X1 U23246 ( .B1(n20421), .B2(n20392), .A(n20340), .ZN(n20341) );
  NOR2_X1 U23247 ( .A1(n20341), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20343) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20668), .ZN(n20344) );
  OAI211_X1 U23249 ( .C1(n20671), .C2(n20388), .A(n20345), .B(n20344), .ZN(
        P1_U3065) );
  AOI22_X1 U23250 ( .A1(n20712), .A2(n20359), .B1(n20711), .B2(n20358), .ZN(
        n20347) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20672), .ZN(n20346) );
  OAI211_X1 U23252 ( .C1(n20675), .C2(n20388), .A(n20347), .B(n20346), .ZN(
        P1_U3066) );
  AOI22_X1 U23253 ( .A1(n20717), .A2(n20358), .B1(n20718), .B2(n20359), .ZN(
        n20349) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20719), .ZN(n20348) );
  OAI211_X1 U23255 ( .C1(n20722), .C2(n20388), .A(n20349), .B(n20348), .ZN(
        P1_U3067) );
  AOI22_X1 U23256 ( .A1(n20724), .A2(n20359), .B1(n20723), .B2(n20358), .ZN(
        n20351) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20678), .ZN(n20350) );
  OAI211_X1 U23258 ( .C1(n20681), .C2(n20388), .A(n20351), .B(n20350), .ZN(
        P1_U3068) );
  AOI22_X1 U23259 ( .A1(n20730), .A2(n20358), .B1(n20729), .B2(n20359), .ZN(
        n20353) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20682), .ZN(n20352) );
  OAI211_X1 U23261 ( .C1(n20685), .C2(n20388), .A(n20353), .B(n20352), .ZN(
        P1_U3069) );
  AOI22_X1 U23262 ( .A1(n20738), .A2(n20358), .B1(n20737), .B2(n20359), .ZN(
        n20355) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20739), .ZN(n20354) );
  OAI211_X1 U23264 ( .C1(n20742), .C2(n20388), .A(n20355), .B(n20354), .ZN(
        P1_U3070) );
  AOI22_X1 U23265 ( .A1(n20744), .A2(n20358), .B1(n20743), .B2(n20359), .ZN(
        n20357) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20745), .ZN(n20356) );
  OAI211_X1 U23267 ( .C1(n20748), .C2(n20388), .A(n20357), .B(n20356), .ZN(
        P1_U3071) );
  AOI22_X1 U23268 ( .A1(n20752), .A2(n20359), .B1(n20750), .B2(n20358), .ZN(
        n20363) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20361), .B1(
        n20360), .B2(n20753), .ZN(n20362) );
  OAI211_X1 U23270 ( .C1(n20759), .C2(n20388), .A(n20363), .B(n20362), .ZN(
        P1_U3072) );
  NOR2_X1 U23271 ( .A1(n20628), .A2(n20364), .ZN(n20384) );
  AOI21_X1 U23272 ( .B1(n20421), .B2(n20630), .A(n20384), .ZN(n20365) );
  OAI22_X1 U23273 ( .A1(n20365), .A2(n20698), .B1(n20364), .B2(n20764), .ZN(
        n20383) );
  AOI22_X1 U23274 ( .A1(n20701), .A2(n20384), .B1(n20700), .B2(n20383), .ZN(
        n20370) );
  INV_X1 U23275 ( .A(n20364), .ZN(n20367) );
  OAI21_X1 U23276 ( .B1(n20427), .B2(n20633), .A(n20365), .ZN(n20366) );
  OAI221_X1 U23277 ( .B1(n20636), .B2(n20367), .C1(n20698), .C2(n20366), .A(
        n20705), .ZN(n20385) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20707), .ZN(n20369) );
  OAI211_X1 U23279 ( .C1(n20710), .C2(n20388), .A(n20370), .B(n20369), .ZN(
        P1_U3073) );
  AOI22_X1 U23280 ( .A1(n20712), .A2(n20384), .B1(n20711), .B2(n20383), .ZN(
        n20372) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20713), .ZN(n20371) );
  OAI211_X1 U23282 ( .C1(n20716), .C2(n20388), .A(n20372), .B(n20371), .ZN(
        P1_U3074) );
  AOI22_X1 U23283 ( .A1(n20717), .A2(n20383), .B1(n20718), .B2(n20384), .ZN(
        n20374) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20601), .ZN(n20373) );
  OAI211_X1 U23285 ( .C1(n20499), .C2(n20388), .A(n20374), .B(n20373), .ZN(
        P1_U3075) );
  AOI22_X1 U23286 ( .A1(n20724), .A2(n20384), .B1(n20723), .B2(n20383), .ZN(
        n20376) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20725), .ZN(n20375) );
  OAI211_X1 U23288 ( .C1(n20728), .C2(n20388), .A(n20376), .B(n20375), .ZN(
        P1_U3076) );
  AOI22_X1 U23289 ( .A1(n20730), .A2(n20383), .B1(n20729), .B2(n20384), .ZN(
        n20378) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20731), .ZN(n20377) );
  OAI211_X1 U23291 ( .C1(n20736), .C2(n20388), .A(n20378), .B(n20377), .ZN(
        P1_U3077) );
  AOI22_X1 U23292 ( .A1(n20738), .A2(n20383), .B1(n20737), .B2(n20384), .ZN(
        n20380) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20611), .ZN(n20379) );
  OAI211_X1 U23294 ( .C1(n20506), .C2(n20388), .A(n20380), .B(n20379), .ZN(
        P1_U3078) );
  AOI22_X1 U23295 ( .A1(n20744), .A2(n20383), .B1(n20743), .B2(n20384), .ZN(
        n20382) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20615), .ZN(n20381) );
  OAI211_X1 U23297 ( .C1(n20509), .C2(n20388), .A(n20382), .B(n20381), .ZN(
        P1_U3079) );
  AOI22_X1 U23298 ( .A1(n20752), .A2(n20384), .B1(n20750), .B2(n20383), .ZN(
        n20387) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20620), .ZN(n20386) );
  OAI211_X1 U23300 ( .C1(n20516), .C2(n20388), .A(n20387), .B(n20386), .ZN(
        P1_U3080) );
  INV_X1 U23301 ( .A(n20414), .ZN(n20390) );
  NAND3_X1 U23302 ( .A1(n20390), .A2(n20636), .A3(n20447), .ZN(n20391) );
  NAND2_X1 U23303 ( .A1(n20391), .A2(n20582), .ZN(n20397) );
  NOR2_X1 U23304 ( .A1(n20393), .A2(n20392), .ZN(n20394) );
  INV_X1 U23305 ( .A(n20660), .ZN(n20586) );
  INV_X1 U23306 ( .A(n20425), .ZN(n20422) );
  NOR2_X1 U23307 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20422), .ZN(
        n20413) );
  AOI22_X1 U23308 ( .A1(n20414), .A2(n20668), .B1(n20701), .B2(n20413), .ZN(
        n20400) );
  INV_X1 U23309 ( .A(n20394), .ZN(n20396) );
  AOI21_X1 U23310 ( .B1(n20397), .B2(n20396), .A(n20395), .ZN(n20398) );
  OAI211_X1 U23311 ( .C1(n20413), .C2(n20593), .A(n20666), .B(n20398), .ZN(
        n20416) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20707), .ZN(n20399) );
  OAI211_X1 U23313 ( .C1(n20419), .C2(n20597), .A(n20400), .B(n20399), .ZN(
        P1_U3081) );
  AOI22_X1 U23314 ( .A1(n20415), .A2(n20713), .B1(n20712), .B2(n20413), .ZN(
        n20402) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20416), .B1(
        n20414), .B2(n20672), .ZN(n20401) );
  OAI211_X1 U23316 ( .C1(n20419), .C2(n20600), .A(n20402), .B(n20401), .ZN(
        P1_U3082) );
  AOI22_X1 U23317 ( .A1(n20413), .A2(n20718), .B1(n20414), .B2(n20719), .ZN(
        n20404) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20601), .ZN(n20403) );
  OAI211_X1 U23319 ( .C1(n20419), .C2(n20604), .A(n20404), .B(n20403), .ZN(
        P1_U3083) );
  AOI22_X1 U23320 ( .A1(n20414), .A2(n20678), .B1(n20724), .B2(n20413), .ZN(
        n20406) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20725), .ZN(n20405) );
  OAI211_X1 U23322 ( .C1(n20419), .C2(n20607), .A(n20406), .B(n20405), .ZN(
        P1_U3084) );
  AOI22_X1 U23323 ( .A1(n20415), .A2(n20731), .B1(n20729), .B2(n20413), .ZN(
        n20408) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20416), .B1(
        n20414), .B2(n20682), .ZN(n20407) );
  OAI211_X1 U23325 ( .C1(n20419), .C2(n20610), .A(n20408), .B(n20407), .ZN(
        P1_U3085) );
  AOI22_X1 U23326 ( .A1(n20415), .A2(n20611), .B1(n20737), .B2(n20413), .ZN(
        n20410) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20416), .B1(
        n20414), .B2(n20739), .ZN(n20409) );
  OAI211_X1 U23328 ( .C1(n20419), .C2(n20614), .A(n20410), .B(n20409), .ZN(
        P1_U3086) );
  AOI22_X1 U23329 ( .A1(n20414), .A2(n20745), .B1(n20743), .B2(n20413), .ZN(
        n20412) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20615), .ZN(n20411) );
  OAI211_X1 U23331 ( .C1(n20419), .C2(n20618), .A(n20412), .B(n20411), .ZN(
        P1_U3087) );
  AOI22_X1 U23332 ( .A1(n20414), .A2(n20753), .B1(n20752), .B2(n20413), .ZN(
        n20418) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20620), .ZN(n20417) );
  OAI211_X1 U23334 ( .C1(n20419), .C2(n20625), .A(n20418), .B(n20417), .ZN(
        P1_U3088) );
  INV_X1 U23335 ( .A(n20420), .ZN(n20443) );
  AOI21_X1 U23336 ( .B1(n20421), .B2(n20696), .A(n20443), .ZN(n20423) );
  OAI22_X1 U23337 ( .A1(n20423), .A2(n20698), .B1(n20422), .B2(n20764), .ZN(
        n20442) );
  AOI22_X1 U23338 ( .A1(n20701), .A2(n20443), .B1(n20700), .B2(n20442), .ZN(
        n20429) );
  OAI21_X1 U23339 ( .B1(n20425), .B2(n20424), .A(n20705), .ZN(n20444) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20444), .B1(
        n20483), .B2(n20707), .ZN(n20428) );
  OAI211_X1 U23341 ( .C1(n20710), .C2(n20447), .A(n20429), .B(n20428), .ZN(
        P1_U3089) );
  AOI22_X1 U23342 ( .A1(n20712), .A2(n20443), .B1(n20711), .B2(n20442), .ZN(
        n20431) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20444), .B1(
        n20483), .B2(n20713), .ZN(n20430) );
  OAI211_X1 U23344 ( .C1(n20716), .C2(n20447), .A(n20431), .B(n20430), .ZN(
        P1_U3090) );
  AOI22_X1 U23345 ( .A1(n20443), .A2(n20718), .B1(n20717), .B2(n20442), .ZN(
        n20433) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20444), .B1(
        n20483), .B2(n20601), .ZN(n20432) );
  OAI211_X1 U23347 ( .C1(n20499), .C2(n20447), .A(n20433), .B(n20432), .ZN(
        P1_U3091) );
  AOI22_X1 U23348 ( .A1(n20724), .A2(n20443), .B1(n20723), .B2(n20442), .ZN(
        n20435) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20444), .B1(
        n20483), .B2(n20725), .ZN(n20434) );
  OAI211_X1 U23350 ( .C1(n20728), .C2(n20447), .A(n20435), .B(n20434), .ZN(
        P1_U3092) );
  AOI22_X1 U23351 ( .A1(n20730), .A2(n20442), .B1(n20729), .B2(n20443), .ZN(
        n20437) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20444), .B1(
        n20483), .B2(n20731), .ZN(n20436) );
  OAI211_X1 U23353 ( .C1(n20736), .C2(n20447), .A(n20437), .B(n20436), .ZN(
        P1_U3093) );
  AOI22_X1 U23354 ( .A1(n20738), .A2(n20442), .B1(n20737), .B2(n20443), .ZN(
        n20439) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20444), .B1(
        n20483), .B2(n20611), .ZN(n20438) );
  OAI211_X1 U23356 ( .C1(n20506), .C2(n20447), .A(n20439), .B(n20438), .ZN(
        P1_U3094) );
  AOI22_X1 U23357 ( .A1(n20744), .A2(n20442), .B1(n20743), .B2(n20443), .ZN(
        n20441) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20444), .B1(
        n20483), .B2(n20615), .ZN(n20440) );
  OAI211_X1 U23359 ( .C1(n20509), .C2(n20447), .A(n20441), .B(n20440), .ZN(
        P1_U3095) );
  AOI22_X1 U23360 ( .A1(n20752), .A2(n20443), .B1(n20750), .B2(n20442), .ZN(
        n20446) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20444), .B1(
        n20483), .B2(n20620), .ZN(n20445) );
  OAI211_X1 U23362 ( .C1(n20516), .C2(n20447), .A(n20446), .B(n20445), .ZN(
        P1_U3096) );
  NOR3_X1 U23363 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20549), .ZN(n20492) );
  NAND2_X1 U23364 ( .A1(n20492), .A2(n20628), .ZN(n20458) );
  INV_X1 U23365 ( .A(n20483), .ZN(n20449) );
  AOI21_X1 U23366 ( .B1(n20449), .B2(n20515), .A(n20633), .ZN(n20451) );
  AND2_X1 U23367 ( .A1(n13653), .A2(n13643), .ZN(n20551) );
  INV_X1 U23368 ( .A(n20551), .ZN(n20450) );
  OAI21_X1 U23369 ( .B1(n20450), .B2(n20659), .A(n20458), .ZN(n20454) );
  NOR2_X1 U23370 ( .A1(n20451), .A2(n20454), .ZN(n20453) );
  AOI211_X2 U23371 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20458), .A(n20453), 
        .B(n20452), .ZN(n20487) );
  INV_X1 U23372 ( .A(n20454), .ZN(n20457) );
  AND2_X1 U23373 ( .A1(n20455), .A2(n20519), .ZN(n20585) );
  INV_X1 U23374 ( .A(n20585), .ZN(n20589) );
  OAI22_X1 U23375 ( .A1(n20457), .A2(n20698), .B1(n20456), .B2(n20589), .ZN(
        n20481) );
  INV_X1 U23376 ( .A(n20458), .ZN(n20480) );
  AOI22_X1 U23377 ( .A1(n20481), .A2(n20700), .B1(n20701), .B2(n20480), .ZN(
        n20460) );
  AOI22_X1 U23378 ( .A1(n20483), .A2(n20668), .B1(n20482), .B2(n20707), .ZN(
        n20459) );
  OAI211_X1 U23379 ( .C1(n20487), .C2(n20461), .A(n20460), .B(n20459), .ZN(
        P1_U3097) );
  AOI22_X1 U23380 ( .A1(n20481), .A2(n20711), .B1(n20712), .B2(n20480), .ZN(
        n20463) );
  AOI22_X1 U23381 ( .A1(n20482), .A2(n20713), .B1(n20483), .B2(n20672), .ZN(
        n20462) );
  OAI211_X1 U23382 ( .C1(n20487), .C2(n20464), .A(n20463), .B(n20462), .ZN(
        P1_U3098) );
  INV_X1 U23383 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n20467) );
  AOI22_X1 U23384 ( .A1(n20717), .A2(n20481), .B1(n20718), .B2(n20480), .ZN(
        n20466) );
  AOI22_X1 U23385 ( .A1(n20482), .A2(n20601), .B1(n20483), .B2(n20719), .ZN(
        n20465) );
  OAI211_X1 U23386 ( .C1(n20487), .C2(n20467), .A(n20466), .B(n20465), .ZN(
        P1_U3099) );
  INV_X1 U23387 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20470) );
  AOI22_X1 U23388 ( .A1(n20481), .A2(n20723), .B1(n20724), .B2(n20480), .ZN(
        n20469) );
  AOI22_X1 U23389 ( .A1(n20482), .A2(n20725), .B1(n20483), .B2(n20678), .ZN(
        n20468) );
  OAI211_X1 U23390 ( .C1(n20487), .C2(n20470), .A(n20469), .B(n20468), .ZN(
        P1_U3100) );
  INV_X1 U23391 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n20473) );
  AOI22_X1 U23392 ( .A1(n20730), .A2(n20481), .B1(n20729), .B2(n20480), .ZN(
        n20472) );
  AOI22_X1 U23393 ( .A1(n20483), .A2(n20682), .B1(n20482), .B2(n20731), .ZN(
        n20471) );
  OAI211_X1 U23394 ( .C1(n20487), .C2(n20473), .A(n20472), .B(n20471), .ZN(
        P1_U3101) );
  INV_X1 U23395 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n20476) );
  AOI22_X1 U23396 ( .A1(n20738), .A2(n20481), .B1(n20737), .B2(n20480), .ZN(
        n20475) );
  AOI22_X1 U23397 ( .A1(n20482), .A2(n20611), .B1(n20483), .B2(n20739), .ZN(
        n20474) );
  OAI211_X1 U23398 ( .C1(n20487), .C2(n20476), .A(n20475), .B(n20474), .ZN(
        P1_U3102) );
  INV_X1 U23399 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n20479) );
  AOI22_X1 U23400 ( .A1(n20744), .A2(n20481), .B1(n20743), .B2(n20480), .ZN(
        n20478) );
  AOI22_X1 U23401 ( .A1(n20482), .A2(n20615), .B1(n20483), .B2(n20745), .ZN(
        n20477) );
  OAI211_X1 U23402 ( .C1(n20487), .C2(n20479), .A(n20478), .B(n20477), .ZN(
        P1_U3103) );
  INV_X1 U23403 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n20486) );
  AOI22_X1 U23404 ( .A1(n20481), .A2(n20750), .B1(n20752), .B2(n20480), .ZN(
        n20485) );
  AOI22_X1 U23405 ( .A1(n20483), .A2(n20753), .B1(n20482), .B2(n20620), .ZN(
        n20484) );
  OAI211_X1 U23406 ( .C1(n20487), .C2(n20486), .A(n20485), .B(n20484), .ZN(
        P1_U3104) );
  INV_X1 U23407 ( .A(n20492), .ZN(n20488) );
  NOR2_X1 U23408 ( .A1(n20628), .A2(n20488), .ZN(n20511) );
  AOI21_X1 U23409 ( .B1(n20551), .B2(n20630), .A(n20511), .ZN(n20489) );
  OAI22_X1 U23410 ( .A1(n20489), .A2(n20698), .B1(n20488), .B2(n20764), .ZN(
        n20510) );
  AOI22_X1 U23411 ( .A1(n20701), .A2(n20511), .B1(n20700), .B2(n20510), .ZN(
        n20494) );
  INV_X1 U23412 ( .A(n20553), .ZN(n20490) );
  OAI211_X1 U23413 ( .C1(n20490), .C2(n20633), .A(n20636), .B(n20489), .ZN(
        n20491) );
  OAI211_X1 U23414 ( .C1(n20636), .C2(n20492), .A(n20705), .B(n20491), .ZN(
        n20512) );
  AOI22_X1 U23415 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20707), .ZN(n20493) );
  OAI211_X1 U23416 ( .C1(n20710), .C2(n20515), .A(n20494), .B(n20493), .ZN(
        P1_U3105) );
  AOI22_X1 U23417 ( .A1(n20712), .A2(n20511), .B1(n20711), .B2(n20510), .ZN(
        n20496) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20713), .ZN(n20495) );
  OAI211_X1 U23419 ( .C1(n20716), .C2(n20515), .A(n20496), .B(n20495), .ZN(
        P1_U3106) );
  AOI22_X1 U23420 ( .A1(n20717), .A2(n20510), .B1(n20718), .B2(n20511), .ZN(
        n20498) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20601), .ZN(n20497) );
  OAI211_X1 U23422 ( .C1(n20499), .C2(n20515), .A(n20498), .B(n20497), .ZN(
        P1_U3107) );
  AOI22_X1 U23423 ( .A1(n20724), .A2(n20511), .B1(n20723), .B2(n20510), .ZN(
        n20501) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20725), .ZN(n20500) );
  OAI211_X1 U23425 ( .C1(n20728), .C2(n20515), .A(n20501), .B(n20500), .ZN(
        P1_U3108) );
  AOI22_X1 U23426 ( .A1(n20730), .A2(n20510), .B1(n20729), .B2(n20511), .ZN(
        n20503) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20731), .ZN(n20502) );
  OAI211_X1 U23428 ( .C1(n20736), .C2(n20515), .A(n20503), .B(n20502), .ZN(
        P1_U3109) );
  AOI22_X1 U23429 ( .A1(n20738), .A2(n20510), .B1(n20737), .B2(n20511), .ZN(
        n20505) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20611), .ZN(n20504) );
  OAI211_X1 U23431 ( .C1(n20506), .C2(n20515), .A(n20505), .B(n20504), .ZN(
        P1_U3110) );
  AOI22_X1 U23432 ( .A1(n20744), .A2(n20510), .B1(n20743), .B2(n20511), .ZN(
        n20508) );
  AOI22_X1 U23433 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20615), .ZN(n20507) );
  OAI211_X1 U23434 ( .C1(n20509), .C2(n20515), .A(n20508), .B(n20507), .ZN(
        P1_U3111) );
  AOI22_X1 U23435 ( .A1(n20752), .A2(n20511), .B1(n20750), .B2(n20510), .ZN(
        n20514) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20512), .B1(
        n20543), .B2(n20620), .ZN(n20513) );
  OAI211_X1 U23437 ( .C1(n20516), .C2(n20515), .A(n20514), .B(n20513), .ZN(
        P1_U3112) );
  INV_X1 U23438 ( .A(n20543), .ZN(n20517) );
  NAND2_X1 U23439 ( .A1(n20517), .A2(n20636), .ZN(n20518) );
  OAI21_X1 U23440 ( .B1(n20518), .B2(n20575), .A(n20582), .ZN(n20526) );
  AND2_X1 U23441 ( .A1(n20551), .A2(n20659), .ZN(n20522) );
  OR2_X1 U23442 ( .A1(n20519), .A2(n20549), .ZN(n20661) );
  INV_X1 U23443 ( .A(n20661), .ZN(n20520) );
  NAND3_X1 U23444 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n12247), .ZN(n20552) );
  NOR2_X1 U23445 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20552), .ZN(
        n20542) );
  AOI22_X1 U23446 ( .A1(n20543), .A2(n20668), .B1(n20701), .B2(n20542), .ZN(
        n20529) );
  INV_X1 U23447 ( .A(n20522), .ZN(n20525) );
  NAND2_X1 U23448 ( .A1(n20661), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20665) );
  OAI211_X1 U23449 ( .C1(n20593), .C2(n20542), .A(n20665), .B(n20523), .ZN(
        n20524) );
  AOI21_X1 U23450 ( .B1(n20526), .B2(n20525), .A(n20524), .ZN(n20527) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20544), .B1(
        n20575), .B2(n20707), .ZN(n20528) );
  OAI211_X1 U23452 ( .C1(n20547), .C2(n20597), .A(n20529), .B(n20528), .ZN(
        P1_U3113) );
  AOI22_X1 U23453 ( .A1(n20575), .A2(n20713), .B1(n20712), .B2(n20542), .ZN(
        n20531) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20672), .ZN(n20530) );
  OAI211_X1 U23455 ( .C1(n20547), .C2(n20600), .A(n20531), .B(n20530), .ZN(
        P1_U3114) );
  AOI22_X1 U23456 ( .A1(n20542), .A2(n20718), .B1(n20575), .B2(n20601), .ZN(
        n20533) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20719), .ZN(n20532) );
  OAI211_X1 U23458 ( .C1(n20547), .C2(n20604), .A(n20533), .B(n20532), .ZN(
        P1_U3115) );
  AOI22_X1 U23459 ( .A1(n20543), .A2(n20678), .B1(n20724), .B2(n20542), .ZN(
        n20535) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20544), .B1(
        n20575), .B2(n20725), .ZN(n20534) );
  OAI211_X1 U23461 ( .C1(n20547), .C2(n20607), .A(n20535), .B(n20534), .ZN(
        P1_U3116) );
  AOI22_X1 U23462 ( .A1(n20575), .A2(n20731), .B1(n20729), .B2(n20542), .ZN(
        n20537) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20682), .ZN(n20536) );
  OAI211_X1 U23464 ( .C1(n20547), .C2(n20610), .A(n20537), .B(n20536), .ZN(
        P1_U3117) );
  AOI22_X1 U23465 ( .A1(n20543), .A2(n20739), .B1(n20737), .B2(n20542), .ZN(
        n20539) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20544), .B1(
        n20575), .B2(n20611), .ZN(n20538) );
  OAI211_X1 U23467 ( .C1(n20547), .C2(n20614), .A(n20539), .B(n20538), .ZN(
        P1_U3118) );
  AOI22_X1 U23468 ( .A1(n20543), .A2(n20745), .B1(n20743), .B2(n20542), .ZN(
        n20541) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20544), .B1(
        n20575), .B2(n20615), .ZN(n20540) );
  OAI211_X1 U23470 ( .C1(n20547), .C2(n20618), .A(n20541), .B(n20540), .ZN(
        P1_U3119) );
  AOI22_X1 U23471 ( .A1(n20543), .A2(n20753), .B1(n20752), .B2(n20542), .ZN(
        n20546) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20544), .B1(
        n20575), .B2(n20620), .ZN(n20545) );
  OAI211_X1 U23473 ( .C1(n20547), .C2(n20625), .A(n20546), .B(n20545), .ZN(
        P1_U3120) );
  NOR2_X1 U23474 ( .A1(n20550), .A2(n20549), .ZN(n20574) );
  AOI21_X1 U23475 ( .B1(n20551), .B2(n20696), .A(n20574), .ZN(n20554) );
  OAI22_X1 U23476 ( .A1(n20554), .A2(n20698), .B1(n20552), .B2(n20764), .ZN(
        n20573) );
  AOI22_X1 U23477 ( .A1(n20701), .A2(n20574), .B1(n20573), .B2(n20700), .ZN(
        n20560) );
  INV_X1 U23478 ( .A(n20552), .ZN(n20558) );
  NOR2_X1 U23479 ( .A1(n20553), .A2(n20698), .ZN(n20555) );
  OAI21_X1 U23480 ( .B1(n20556), .B2(n20555), .A(n20554), .ZN(n20557) );
  OAI211_X1 U23481 ( .C1(n20636), .C2(n20558), .A(n20705), .B(n20557), .ZN(
        n20576) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20668), .ZN(n20559) );
  OAI211_X1 U23483 ( .C1(n20671), .C2(n20594), .A(n20560), .B(n20559), .ZN(
        P1_U3121) );
  AOI22_X1 U23484 ( .A1(n20712), .A2(n20574), .B1(n20573), .B2(n20711), .ZN(
        n20562) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20672), .ZN(n20561) );
  OAI211_X1 U23486 ( .C1(n20675), .C2(n20594), .A(n20562), .B(n20561), .ZN(
        P1_U3122) );
  AOI22_X1 U23487 ( .A1(n20717), .A2(n20573), .B1(n20718), .B2(n20574), .ZN(
        n20564) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20719), .ZN(n20563) );
  OAI211_X1 U23489 ( .C1(n20722), .C2(n20594), .A(n20564), .B(n20563), .ZN(
        P1_U3123) );
  AOI22_X1 U23490 ( .A1(n20724), .A2(n20574), .B1(n20573), .B2(n20723), .ZN(
        n20566) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20678), .ZN(n20565) );
  OAI211_X1 U23492 ( .C1(n20681), .C2(n20594), .A(n20566), .B(n20565), .ZN(
        P1_U3124) );
  AOI22_X1 U23493 ( .A1(n20730), .A2(n20573), .B1(n20729), .B2(n20574), .ZN(
        n20568) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20682), .ZN(n20567) );
  OAI211_X1 U23495 ( .C1(n20685), .C2(n20594), .A(n20568), .B(n20567), .ZN(
        P1_U3125) );
  AOI22_X1 U23496 ( .A1(n20738), .A2(n20573), .B1(n20737), .B2(n20574), .ZN(
        n20570) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20739), .ZN(n20569) );
  OAI211_X1 U23498 ( .C1(n20742), .C2(n20594), .A(n20570), .B(n20569), .ZN(
        P1_U3126) );
  AOI22_X1 U23499 ( .A1(n20744), .A2(n20573), .B1(n20743), .B2(n20574), .ZN(
        n20572) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20745), .ZN(n20571) );
  OAI211_X1 U23501 ( .C1(n20748), .C2(n20594), .A(n20572), .B(n20571), .ZN(
        P1_U3127) );
  AOI22_X1 U23502 ( .A1(n20752), .A2(n20574), .B1(n20573), .B2(n20750), .ZN(
        n20578) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20753), .ZN(n20577) );
  OAI211_X1 U23504 ( .C1(n20759), .C2(n20594), .A(n20578), .B(n20577), .ZN(
        P1_U3128) );
  INV_X1 U23505 ( .A(n20653), .ZN(n20581) );
  NAND3_X1 U23506 ( .A1(n20581), .A2(n20636), .A3(n20594), .ZN(n20583) );
  NAND2_X1 U23507 ( .A1(n20583), .A2(n20582), .ZN(n20591) );
  OR2_X1 U23508 ( .A1(n13643), .A2(n20584), .ZN(n20629) );
  NOR2_X1 U23509 ( .A1(n20629), .A2(n20659), .ZN(n20588) );
  NAND3_X1 U23510 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20587), .ZN(n20631) );
  NOR2_X1 U23511 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20631), .ZN(
        n20619) );
  AOI22_X1 U23512 ( .A1(n20653), .A2(n20707), .B1(n20701), .B2(n20619), .ZN(
        n20596) );
  INV_X1 U23513 ( .A(n20588), .ZN(n20590) );
  AOI22_X1 U23514 ( .A1(n20591), .A2(n20590), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20589), .ZN(n20592) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20668), .ZN(n20595) );
  OAI211_X1 U23516 ( .C1(n20626), .C2(n20597), .A(n20596), .B(n20595), .ZN(
        P1_U3129) );
  AOI22_X1 U23517 ( .A1(n20653), .A2(n20713), .B1(n20712), .B2(n20619), .ZN(
        n20599) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20672), .ZN(n20598) );
  OAI211_X1 U23519 ( .C1(n20626), .C2(n20600), .A(n20599), .B(n20598), .ZN(
        P1_U3130) );
  AOI22_X1 U23520 ( .A1(n20619), .A2(n20718), .B1(n20653), .B2(n20601), .ZN(
        n20603) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20719), .ZN(n20602) );
  OAI211_X1 U23522 ( .C1(n20626), .C2(n20604), .A(n20603), .B(n20602), .ZN(
        P1_U3131) );
  AOI22_X1 U23523 ( .A1(n20653), .A2(n20725), .B1(n20724), .B2(n20619), .ZN(
        n20606) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20678), .ZN(n20605) );
  OAI211_X1 U23525 ( .C1(n20626), .C2(n20607), .A(n20606), .B(n20605), .ZN(
        P1_U3132) );
  AOI22_X1 U23526 ( .A1(n20653), .A2(n20731), .B1(n20729), .B2(n20619), .ZN(
        n20609) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20682), .ZN(n20608) );
  OAI211_X1 U23528 ( .C1(n20626), .C2(n20610), .A(n20609), .B(n20608), .ZN(
        P1_U3133) );
  AOI22_X1 U23529 ( .A1(n20653), .A2(n20611), .B1(n20737), .B2(n20619), .ZN(
        n20613) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20739), .ZN(n20612) );
  OAI211_X1 U23531 ( .C1(n20626), .C2(n20614), .A(n20613), .B(n20612), .ZN(
        P1_U3134) );
  AOI22_X1 U23532 ( .A1(n20653), .A2(n20615), .B1(n20743), .B2(n20619), .ZN(
        n20617) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20745), .ZN(n20616) );
  OAI211_X1 U23534 ( .C1(n20626), .C2(n20618), .A(n20617), .B(n20616), .ZN(
        P1_U3135) );
  AOI22_X1 U23535 ( .A1(n20653), .A2(n20620), .B1(n20752), .B2(n20619), .ZN(
        n20624) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20753), .ZN(n20623) );
  OAI211_X1 U23537 ( .C1(n20626), .C2(n20625), .A(n20624), .B(n20623), .ZN(
        P1_U3136) );
  NOR2_X1 U23538 ( .A1(n20628), .A2(n20631), .ZN(n20652) );
  INV_X1 U23539 ( .A(n20629), .ZN(n20697) );
  AOI21_X1 U23540 ( .B1(n20697), .B2(n20630), .A(n20652), .ZN(n20632) );
  OAI22_X1 U23541 ( .A1(n20632), .A2(n20698), .B1(n20631), .B2(n20764), .ZN(
        n20651) );
  AOI22_X1 U23542 ( .A1(n20701), .A2(n20652), .B1(n20700), .B2(n20651), .ZN(
        n20638) );
  INV_X1 U23543 ( .A(n20631), .ZN(n20635) );
  OAI21_X1 U23544 ( .B1(n20704), .B2(n20633), .A(n20632), .ZN(n20634) );
  OAI221_X1 U23545 ( .B1(n20636), .B2(n20635), .C1(n20698), .C2(n20634), .A(
        n20705), .ZN(n20654) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20668), .ZN(n20637) );
  OAI211_X1 U23547 ( .C1(n20671), .C2(n20662), .A(n20638), .B(n20637), .ZN(
        P1_U3137) );
  AOI22_X1 U23548 ( .A1(n20712), .A2(n20652), .B1(n20711), .B2(n20651), .ZN(
        n20640) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20672), .ZN(n20639) );
  OAI211_X1 U23550 ( .C1(n20675), .C2(n20662), .A(n20640), .B(n20639), .ZN(
        P1_U3138) );
  AOI22_X1 U23551 ( .A1(n20717), .A2(n20651), .B1(n20718), .B2(n20652), .ZN(
        n20642) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20719), .ZN(n20641) );
  OAI211_X1 U23553 ( .C1(n20722), .C2(n20662), .A(n20642), .B(n20641), .ZN(
        P1_U3139) );
  AOI22_X1 U23554 ( .A1(n20724), .A2(n20652), .B1(n20723), .B2(n20651), .ZN(
        n20644) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20678), .ZN(n20643) );
  OAI211_X1 U23556 ( .C1(n20681), .C2(n20662), .A(n20644), .B(n20643), .ZN(
        P1_U3140) );
  AOI22_X1 U23557 ( .A1(n20730), .A2(n20651), .B1(n20729), .B2(n20652), .ZN(
        n20646) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20682), .ZN(n20645) );
  OAI211_X1 U23559 ( .C1(n20685), .C2(n20662), .A(n20646), .B(n20645), .ZN(
        P1_U3141) );
  AOI22_X1 U23560 ( .A1(n20738), .A2(n20651), .B1(n20737), .B2(n20652), .ZN(
        n20648) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20739), .ZN(n20647) );
  OAI211_X1 U23562 ( .C1(n20742), .C2(n20662), .A(n20648), .B(n20647), .ZN(
        P1_U3142) );
  AOI22_X1 U23563 ( .A1(n20744), .A2(n20651), .B1(n20743), .B2(n20652), .ZN(
        n20650) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20745), .ZN(n20649) );
  OAI211_X1 U23565 ( .C1(n20748), .C2(n20662), .A(n20650), .B(n20649), .ZN(
        P1_U3143) );
  AOI22_X1 U23566 ( .A1(n20752), .A2(n20652), .B1(n20750), .B2(n20651), .ZN(
        n20656) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20753), .ZN(n20655) );
  OAI211_X1 U23568 ( .C1(n20759), .C2(n20662), .A(n20656), .B(n20655), .ZN(
        P1_U3144) );
  NOR2_X1 U23569 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20702), .ZN(
        n20691) );
  NAND2_X1 U23570 ( .A1(n20697), .A2(n20659), .ZN(n20663) );
  OAI22_X1 U23571 ( .A1(n20663), .A2(n20698), .B1(n20661), .B2(n20660), .ZN(
        n20690) );
  AOI22_X1 U23572 ( .A1(n20701), .A2(n20691), .B1(n20700), .B2(n20690), .ZN(
        n20670) );
  OAI21_X1 U23573 ( .B1(n20754), .B2(n20692), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20664) );
  AOI21_X1 U23574 ( .B1(n20664), .B2(n20663), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20667) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20693), .B1(
        n20692), .B2(n20668), .ZN(n20669) );
  OAI211_X1 U23576 ( .C1(n20671), .C2(n20735), .A(n20670), .B(n20669), .ZN(
        P1_U3145) );
  AOI22_X1 U23577 ( .A1(n20712), .A2(n20691), .B1(n20711), .B2(n20690), .ZN(
        n20674) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20693), .B1(
        n20692), .B2(n20672), .ZN(n20673) );
  OAI211_X1 U23579 ( .C1(n20675), .C2(n20735), .A(n20674), .B(n20673), .ZN(
        P1_U3146) );
  AOI22_X1 U23580 ( .A1(n20717), .A2(n20690), .B1(n20718), .B2(n20691), .ZN(
        n20677) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20693), .B1(
        n20692), .B2(n20719), .ZN(n20676) );
  OAI211_X1 U23582 ( .C1(n20722), .C2(n20735), .A(n20677), .B(n20676), .ZN(
        P1_U3147) );
  AOI22_X1 U23583 ( .A1(n20724), .A2(n20691), .B1(n20723), .B2(n20690), .ZN(
        n20680) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20693), .B1(
        n20692), .B2(n20678), .ZN(n20679) );
  OAI211_X1 U23585 ( .C1(n20681), .C2(n20735), .A(n20680), .B(n20679), .ZN(
        P1_U3148) );
  AOI22_X1 U23586 ( .A1(n20730), .A2(n20690), .B1(n20729), .B2(n20691), .ZN(
        n20684) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20693), .B1(
        n20692), .B2(n20682), .ZN(n20683) );
  OAI211_X1 U23588 ( .C1(n20685), .C2(n20735), .A(n20684), .B(n20683), .ZN(
        P1_U3149) );
  AOI22_X1 U23589 ( .A1(n20738), .A2(n20690), .B1(n20737), .B2(n20691), .ZN(
        n20687) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20693), .B1(
        n20692), .B2(n20739), .ZN(n20686) );
  OAI211_X1 U23591 ( .C1(n20742), .C2(n20735), .A(n20687), .B(n20686), .ZN(
        P1_U3150) );
  AOI22_X1 U23592 ( .A1(n20744), .A2(n20690), .B1(n20743), .B2(n20691), .ZN(
        n20689) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20693), .B1(
        n20692), .B2(n20745), .ZN(n20688) );
  OAI211_X1 U23594 ( .C1(n20748), .C2(n20735), .A(n20689), .B(n20688), .ZN(
        P1_U3151) );
  AOI22_X1 U23595 ( .A1(n20752), .A2(n20691), .B1(n20750), .B2(n20690), .ZN(
        n20695) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20693), .B1(
        n20692), .B2(n20753), .ZN(n20694) );
  OAI211_X1 U23597 ( .C1(n20759), .C2(n20735), .A(n20695), .B(n20694), .ZN(
        P1_U3152) );
  AOI21_X1 U23598 ( .B1(n20697), .B2(n20696), .A(n20751), .ZN(n20699) );
  OAI22_X1 U23599 ( .A1(n20699), .A2(n20698), .B1(n20702), .B2(n20764), .ZN(
        n20749) );
  AOI22_X1 U23600 ( .A1(n20701), .A2(n20751), .B1(n20700), .B2(n20749), .ZN(
        n20709) );
  OAI21_X1 U23601 ( .B1(n20704), .B2(n20703), .A(n20702), .ZN(n20706) );
  NAND2_X1 U23602 ( .A1(n20706), .A2(n20705), .ZN(n20755) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20755), .B1(
        n20732), .B2(n20707), .ZN(n20708) );
  OAI211_X1 U23604 ( .C1(n20710), .C2(n20735), .A(n20709), .B(n20708), .ZN(
        P1_U3153) );
  AOI22_X1 U23605 ( .A1(n20712), .A2(n20751), .B1(n20711), .B2(n20749), .ZN(
        n20715) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20755), .B1(
        n20732), .B2(n20713), .ZN(n20714) );
  OAI211_X1 U23607 ( .C1(n20716), .C2(n20735), .A(n20715), .B(n20714), .ZN(
        P1_U3154) );
  AOI22_X1 U23608 ( .A1(n20751), .A2(n20718), .B1(n20717), .B2(n20749), .ZN(
        n20721) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20755), .B1(
        n20754), .B2(n20719), .ZN(n20720) );
  OAI211_X1 U23610 ( .C1(n20722), .C2(n20758), .A(n20721), .B(n20720), .ZN(
        P1_U3155) );
  AOI22_X1 U23611 ( .A1(n20724), .A2(n20751), .B1(n20723), .B2(n20749), .ZN(
        n20727) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20755), .B1(
        n20732), .B2(n20725), .ZN(n20726) );
  OAI211_X1 U23613 ( .C1(n20728), .C2(n20735), .A(n20727), .B(n20726), .ZN(
        P1_U3156) );
  AOI22_X1 U23614 ( .A1(n20730), .A2(n20749), .B1(n20729), .B2(n20751), .ZN(
        n20734) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20755), .B1(
        n20732), .B2(n20731), .ZN(n20733) );
  OAI211_X1 U23616 ( .C1(n20736), .C2(n20735), .A(n20734), .B(n20733), .ZN(
        P1_U3157) );
  AOI22_X1 U23617 ( .A1(n20738), .A2(n20749), .B1(n20737), .B2(n20751), .ZN(
        n20741) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20755), .B1(
        n20754), .B2(n20739), .ZN(n20740) );
  OAI211_X1 U23619 ( .C1(n20742), .C2(n20758), .A(n20741), .B(n20740), .ZN(
        P1_U3158) );
  AOI22_X1 U23620 ( .A1(n20744), .A2(n20749), .B1(n20743), .B2(n20751), .ZN(
        n20747) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20755), .B1(
        n20754), .B2(n20745), .ZN(n20746) );
  OAI211_X1 U23622 ( .C1(n20748), .C2(n20758), .A(n20747), .B(n20746), .ZN(
        P1_U3159) );
  AOI22_X1 U23623 ( .A1(n20752), .A2(n20751), .B1(n20750), .B2(n20749), .ZN(
        n20757) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20755), .B1(
        n20754), .B2(n20753), .ZN(n20756) );
  OAI211_X1 U23625 ( .C1(n20759), .C2(n20758), .A(n20757), .B(n20756), .ZN(
        P1_U3160) );
  NOR2_X1 U23626 ( .A1(n20761), .A2(n20760), .ZN(n20765) );
  INV_X1 U23627 ( .A(n20762), .ZN(n20763) );
  OAI21_X1 U23628 ( .B1(n20765), .B2(n20764), .A(n20763), .ZN(P1_U3163) );
  AND2_X1 U23629 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20847), .ZN(
        P1_U3164) );
  AND2_X1 U23630 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20847), .ZN(
        P1_U3165) );
  AND2_X1 U23631 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20847), .ZN(
        P1_U3166) );
  AND2_X1 U23632 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20847), .ZN(
        P1_U3167) );
  AND2_X1 U23633 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20847), .ZN(
        P1_U3168) );
  AND2_X1 U23634 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20847), .ZN(
        P1_U3169) );
  AND2_X1 U23635 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20847), .ZN(
        P1_U3170) );
  AND2_X1 U23636 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20847), .ZN(
        P1_U3171) );
  AND2_X1 U23637 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20847), .ZN(
        P1_U3172) );
  AND2_X1 U23638 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20847), .ZN(
        P1_U3173) );
  AND2_X1 U23639 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20847), .ZN(
        P1_U3174) );
  AND2_X1 U23640 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20847), .ZN(
        P1_U3175) );
  AND2_X1 U23641 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20847), .ZN(
        P1_U3176) );
  AND2_X1 U23642 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20847), .ZN(
        P1_U3177) );
  AND2_X1 U23643 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20847), .ZN(
        P1_U3178) );
  NOR2_X1 U23644 ( .A1(n20851), .A2(n20766), .ZN(P1_U3179) );
  AND2_X1 U23645 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20847), .ZN(
        P1_U3180) );
  AND2_X1 U23646 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20847), .ZN(
        P1_U3181) );
  AND2_X1 U23647 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20847), .ZN(
        P1_U3182) );
  AND2_X1 U23648 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20847), .ZN(
        P1_U3183) );
  AND2_X1 U23649 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20847), .ZN(
        P1_U3184) );
  AND2_X1 U23650 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20847), .ZN(
        P1_U3185) );
  AND2_X1 U23651 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20847), .ZN(P1_U3186) );
  AND2_X1 U23652 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20847), .ZN(P1_U3187) );
  AND2_X1 U23653 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20847), .ZN(P1_U3188) );
  AND2_X1 U23654 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20847), .ZN(P1_U3189) );
  AND2_X1 U23655 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20847), .ZN(P1_U3190) );
  AND2_X1 U23656 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20847), .ZN(P1_U3191) );
  AND2_X1 U23657 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20847), .ZN(P1_U3192) );
  AND2_X1 U23658 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20847), .ZN(P1_U3193) );
  NAND2_X1 U23659 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20771), .ZN(n20777) );
  INV_X1 U23660 ( .A(n20777), .ZN(n20770) );
  NOR2_X1 U23661 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20767) );
  OAI21_X1 U23662 ( .B1(n20767), .B2(n20773), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20768) );
  AOI21_X1 U23663 ( .B1(NA), .B2(n20772), .A(n20768), .ZN(n20769) );
  OAI22_X1 U23664 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20770), .B1(n20832), 
        .B2(n20769), .ZN(P1_U3194) );
  NOR3_X1 U23665 ( .A1(NA), .A2(n20772), .A3(n20771), .ZN(n20776) );
  AOI21_X1 U23666 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20781), .A(n20773), .ZN(n20775) );
  AOI222_X1 U23667 ( .A1(n20776), .A2(n20775), .B1(n20776), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .C1(n20775), .C2(n20774), .ZN(n20780)
         );
  OAI211_X1 U23668 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20778), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20777), .ZN(n20779) );
  NAND2_X1 U23669 ( .A1(n20780), .A2(n20779), .ZN(P1_U3196) );
  AND2_X1 U23670 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20832), .ZN(n20838) );
  INV_X1 U23671 ( .A(n20838), .ZN(n20835) );
  INV_X1 U23672 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20782) );
  AND2_X1 U23673 ( .A1(n20832), .A2(n20781), .ZN(n20837) );
  OAI222_X1 U23674 ( .A1(n20835), .A2(n20852), .B1(n20782), .B2(n20832), .C1(
        n20784), .C2(n20830), .ZN(P1_U3197) );
  INV_X1 U23675 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20783) );
  OAI222_X1 U23676 ( .A1(n20835), .A2(n20784), .B1(n20783), .B2(n20832), .C1(
        n13769), .C2(n20830), .ZN(P1_U3198) );
  OAI222_X1 U23677 ( .A1(n20835), .A2(n13769), .B1(n20785), .B2(n20832), .C1(
        n20786), .C2(n20830), .ZN(P1_U3199) );
  INV_X1 U23678 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20787) );
  OAI222_X1 U23679 ( .A1(n20830), .A2(n20789), .B1(n20787), .B2(n20832), .C1(
        n20786), .C2(n20835), .ZN(P1_U3200) );
  AOI22_X1 U23680 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20860), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20837), .ZN(n20788) );
  OAI21_X1 U23681 ( .B1(n20789), .B2(n20835), .A(n20788), .ZN(P1_U3201) );
  AOI22_X1 U23682 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20860), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20838), .ZN(n20790) );
  OAI21_X1 U23683 ( .B1(n20792), .B2(n20830), .A(n20790), .ZN(P1_U3202) );
  INV_X1 U23684 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20791) );
  OAI222_X1 U23685 ( .A1(n20835), .A2(n20792), .B1(n20791), .B2(n20832), .C1(
        n20793), .C2(n20830), .ZN(P1_U3203) );
  INV_X1 U23686 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20794) );
  OAI222_X1 U23687 ( .A1(n20830), .A2(n20796), .B1(n20794), .B2(n20832), .C1(
        n20793), .C2(n20835), .ZN(P1_U3204) );
  INV_X1 U23688 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20795) );
  INV_X1 U23689 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20798) );
  OAI222_X1 U23690 ( .A1(n20835), .A2(n20796), .B1(n20795), .B2(n20832), .C1(
        n20798), .C2(n20830), .ZN(P1_U3205) );
  INV_X1 U23691 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20797) );
  OAI222_X1 U23692 ( .A1(n20835), .A2(n20798), .B1(n20797), .B2(n20832), .C1(
        n20800), .C2(n20830), .ZN(P1_U3206) );
  INV_X1 U23693 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20799) );
  OAI222_X1 U23694 ( .A1(n20835), .A2(n20800), .B1(n20799), .B2(n20832), .C1(
        n20802), .C2(n20830), .ZN(P1_U3207) );
  INV_X1 U23695 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20801) );
  OAI222_X1 U23696 ( .A1(n20835), .A2(n20802), .B1(n20801), .B2(n20832), .C1(
        n20804), .C2(n20830), .ZN(P1_U3208) );
  INV_X1 U23697 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20803) );
  OAI222_X1 U23698 ( .A1(n20835), .A2(n20804), .B1(n20803), .B2(n20832), .C1(
        n20805), .C2(n20830), .ZN(P1_U3209) );
  INV_X1 U23699 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20806) );
  OAI222_X1 U23700 ( .A1(n20830), .A2(n20808), .B1(n20806), .B2(n20832), .C1(
        n20805), .C2(n20835), .ZN(P1_U3210) );
  INV_X1 U23701 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20807) );
  INV_X1 U23702 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20810) );
  OAI222_X1 U23703 ( .A1(n20835), .A2(n20808), .B1(n20807), .B2(n20832), .C1(
        n20810), .C2(n20830), .ZN(P1_U3211) );
  AOI22_X1 U23704 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20860), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20837), .ZN(n20809) );
  OAI21_X1 U23705 ( .B1(n20810), .B2(n20835), .A(n20809), .ZN(P1_U3212) );
  INV_X1 U23706 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20813) );
  AOI22_X1 U23707 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20860), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20838), .ZN(n20811) );
  OAI21_X1 U23708 ( .B1(n20813), .B2(n20830), .A(n20811), .ZN(P1_U3213) );
  INV_X1 U23709 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20812) );
  OAI222_X1 U23710 ( .A1(n20835), .A2(n20813), .B1(n20812), .B2(n20832), .C1(
        n20814), .C2(n20830), .ZN(P1_U3214) );
  INV_X1 U23711 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20815) );
  OAI222_X1 U23712 ( .A1(n20830), .A2(n20817), .B1(n20815), .B2(n20832), .C1(
        n20814), .C2(n20835), .ZN(P1_U3215) );
  INV_X1 U23713 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20816) );
  OAI222_X1 U23714 ( .A1(n20835), .A2(n20817), .B1(n20816), .B2(n20832), .C1(
        n20818), .C2(n20830), .ZN(P1_U3216) );
  INV_X1 U23715 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20819) );
  OAI222_X1 U23716 ( .A1(n20830), .A2(n20821), .B1(n20819), .B2(n20832), .C1(
        n20818), .C2(n20835), .ZN(P1_U3217) );
  AOI22_X1 U23717 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20860), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20837), .ZN(n20820) );
  OAI21_X1 U23718 ( .B1(n20821), .B2(n20835), .A(n20820), .ZN(P1_U3218) );
  AOI22_X1 U23719 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20860), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20838), .ZN(n20822) );
  OAI21_X1 U23720 ( .B1(n20824), .B2(n20830), .A(n20822), .ZN(P1_U3219) );
  INV_X1 U23721 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20823) );
  OAI222_X1 U23722 ( .A1(n20835), .A2(n20824), .B1(n20823), .B2(n20832), .C1(
        n20826), .C2(n20830), .ZN(P1_U3220) );
  INV_X1 U23723 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20825) );
  OAI222_X1 U23724 ( .A1(n20835), .A2(n20826), .B1(n20825), .B2(n20832), .C1(
        n20828), .C2(n20830), .ZN(P1_U3221) );
  AOI22_X1 U23725 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20837), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20860), .ZN(n20827) );
  OAI21_X1 U23726 ( .B1(n20828), .B2(n20835), .A(n20827), .ZN(P1_U3222) );
  INV_X1 U23727 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20834) );
  AOI22_X1 U23728 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20838), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20860), .ZN(n20829) );
  OAI21_X1 U23729 ( .B1(n20834), .B2(n20830), .A(n20829), .ZN(P1_U3223) );
  INV_X1 U23730 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20833) );
  OAI222_X1 U23731 ( .A1(n20835), .A2(n20834), .B1(n20833), .B2(n20832), .C1(
        n20831), .C2(n20830), .ZN(P1_U3224) );
  AOI222_X1 U23732 ( .A1(n20837), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20860), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20838), .ZN(n20836) );
  INV_X1 U23733 ( .A(n20836), .ZN(P1_U3225) );
  AOI222_X1 U23734 ( .A1(n20838), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20860), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20837), .ZN(n20839) );
  INV_X1 U23735 ( .A(n20839), .ZN(P1_U3226) );
  INV_X1 U23736 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U23737 ( .A1(n20832), .A2(n20841), .B1(n20840), .B2(n20860), .ZN(
        P1_U3458) );
  AOI22_X1 U23738 ( .A1(n20832), .A2(n20854), .B1(n20842), .B2(n20860), .ZN(
        P1_U3459) );
  AOI22_X1 U23739 ( .A1(n20832), .A2(n20844), .B1(n20843), .B2(n20860), .ZN(
        P1_U3460) );
  INV_X1 U23740 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20859) );
  INV_X1 U23741 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20845) );
  AOI22_X1 U23742 ( .A1(n20832), .A2(n20859), .B1(n20845), .B2(n20860), .ZN(
        P1_U3461) );
  INV_X1 U23743 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20848) );
  INV_X1 U23744 ( .A(n20849), .ZN(n20846) );
  AOI21_X1 U23745 ( .B1(n20848), .B2(n20847), .A(n20846), .ZN(P1_U3464) );
  OAI21_X1 U23746 ( .B1(n20851), .B2(n20850), .A(n20849), .ZN(P1_U3465) );
  AOI21_X1 U23747 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20853) );
  AOI22_X1 U23748 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20853), .B2(n20852), .ZN(n20855) );
  AOI22_X1 U23749 ( .A1(n20856), .A2(n20855), .B1(n20854), .B2(n20858), .ZN(
        P1_U3481) );
  NOR2_X1 U23750 ( .A1(n20858), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20857) );
  AOI22_X1 U23751 ( .A1(n20859), .A2(n20858), .B1(n13549), .B2(n20857), .ZN(
        P1_U3482) );
  AOI22_X1 U23752 ( .A1(n20832), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20861), 
        .B2(n20860), .ZN(P1_U3483) );
  AOI211_X1 U23753 ( .C1(n9726), .C2(n20864), .A(n20863), .B(n20862), .ZN(
        n20871) );
  INV_X1 U23754 ( .A(n20865), .ZN(n20866) );
  OAI211_X1 U23755 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n11631), .A(n20866), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20868) );
  AOI21_X1 U23756 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20868), .A(n20867), 
        .ZN(n20870) );
  NAND2_X1 U23757 ( .A1(n20871), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20869) );
  OAI21_X1 U23758 ( .B1(n20871), .B2(n20870), .A(n20869), .ZN(P1_U3485) );
  MUX2_X1 U23759 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20832), .Z(P1_U3486) );
  INV_X1 U11520 ( .A(n13129), .ZN(n9737) );
  CLKBUF_X3 U13596 ( .A(n10509), .Z(n13132) );
  XNOR2_X1 U11229 ( .A(n12617), .B(n13544), .ZN(n13587) );
  BUF_X4 U11233 ( .A(n15790), .Z(n9712) );
  NAND2_X1 U14925 ( .A1(n20297), .A2(n11701), .ZN(n11724) );
  CLKBUF_X3 U11458 ( .A(n13273), .Z(n9729) );
  NAND2_X1 U11159 ( .A1(n11676), .A2(n11675), .ZN(n11707) );
  CLKBUF_X1 U11199 ( .A(n11713), .Z(n11714) );
  CLKBUF_X1 U11204 ( .A(n11694), .Z(n11695) );
  NOR2_X2 U11217 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10441) );
  CLKBUF_X1 U11225 ( .A(n14182), .Z(n14186) );
  CLKBUF_X1 U11226 ( .A(n14692), .Z(n14727) );
  AOI21_X1 U11235 ( .B1(n13653), .B2(n20761), .A(n11761), .ZN(n11800) );
  CLKBUF_X1 U11236 ( .A(n11232), .Z(n12564) );
  AND4_X1 U11246 ( .A1(n11603), .A2(n11602), .A3(n11601), .A4(n11600), .ZN(
        n11604) );
  CLKBUF_X1 U11270 ( .A(n13703), .Z(n9715) );
  CLKBUF_X1 U11291 ( .A(n17588), .Z(n9740) );
  CLKBUF_X1 U11522 ( .A(n13934), .Z(n20392) );
  CLKBUF_X1 U11736 ( .A(n16353), .Z(n9710) );
  CLKBUF_X1 U11932 ( .A(n10646), .Z(n14399) );
  CLKBUF_X1 U11991 ( .A(n16534), .Z(n16540) );
endmodule

