

module b17_C_gen_AntiSAT_k_128_2 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9631, n9632, n9633, n9634, n9635, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028;

  CLKBUF_X1 U11075 ( .A(n19111), .Z(n9634) );
  AND2_X1 U11076 ( .A1(n9904), .A2(n10679), .ZN(n9674) );
  INV_X2 U11077 ( .A(n18687), .ZN(n18679) );
  OR2_X1 U11078 ( .A1(n13388), .A2(n13377), .ZN(n13658) );
  OR2_X1 U11079 ( .A1(n13388), .A2(n13383), .ZN(n19351) );
  NAND2_X1 U11080 ( .A1(n10173), .A2(n10449), .ZN(n10602) );
  AOI211_X1 U11081 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n12294), .B(n12293), .ZN(n17401) );
  INV_X1 U11082 ( .A(n17168), .ZN(n17147) );
  CLKBUF_X1 U11083 ( .A(n12309), .Z(n9659) );
  INV_X1 U11084 ( .A(n12308), .ZN(n9657) );
  CLKBUF_X1 U11085 ( .A(n12309), .Z(n9658) );
  AND2_X2 U11086 ( .A1(n12036), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12180) );
  INV_X1 U11087 ( .A(n12307), .ZN(n17169) );
  AND2_X1 U11088 ( .A1(n13136), .A2(n11549), .ZN(n12160) );
  AND2_X1 U11089 ( .A1(n11544), .A2(n11376), .ZN(n11703) );
  AND2_X1 U11090 ( .A1(n11544), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11874) );
  AND2_X1 U11091 ( .A1(n9661), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12103) );
  INV_X2 U11092 ( .A(n12308), .ZN(n9651) );
  BUF_X1 U11094 ( .A(n15623), .Z(n17211) );
  INV_X1 U11095 ( .A(n11440), .ZN(n16348) );
  CLKBUF_X2 U11096 ( .A(n11431), .Z(n12259) );
  AND2_X1 U11097 ( .A1(n10278), .A2(n10277), .ZN(n10743) );
  INV_X1 U11098 ( .A(n10894), .ZN(n11033) );
  AND2_X1 U11099 ( .A1(n13306), .A2(n10277), .ZN(n11064) );
  CLKBUF_X2 U11100 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n16308) );
  INV_X1 U11101 ( .A(n11380), .ZN(n9638) );
  INV_X1 U11102 ( .A(n11430), .ZN(n12923) );
  AND3_X1 U11103 ( .A1(n10469), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10280) );
  NAND2_X1 U11104 ( .A1(n10422), .A2(n10421), .ZN(n10463) );
  BUF_X1 U11105 ( .A(n15623), .Z(n17150) );
  NAND2_X1 U11106 ( .A1(n9704), .A2(n10450), .ZN(n10468) );
  AND2_X1 U11107 ( .A1(n9663), .A2(n11376), .ZN(n11589) );
  OR2_X1 U11108 ( .A1(n13388), .A2(n13387), .ZN(n13881) );
  OR2_X1 U11109 ( .A1(n13023), .A2(n20184), .ZN(n14066) );
  AND3_X1 U11111 ( .A1(n9792), .A2(n9790), .A3(n9789), .ZN(n14251) );
  AND2_X1 U11112 ( .A1(n12037), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12188) );
  INV_X1 U11113 ( .A(n17168), .ZN(n17217) );
  AND2_X1 U11115 ( .A1(n13738), .A2(n13739), .ZN(n10647) );
  NAND2_X1 U11116 ( .A1(n11171), .A2(n11170), .ZN(n11182) );
  INV_X1 U11117 ( .A(n9972), .ZN(n9971) );
  OAI21_X1 U11118 ( .B1(n20812), .B2(n11192), .A(n11187), .ZN(n11189) );
  OR2_X1 U11119 ( .A1(n15391), .A2(n10216), .ZN(n10220) );
  OR2_X1 U11120 ( .A1(n12270), .A2(n18675), .ZN(n9695) );
  INV_X1 U11121 ( .A(n18664), .ZN(n18689) );
  INV_X2 U11122 ( .A(n10265), .ZN(n14293) );
  OR2_X1 U11123 ( .A1(n14520), .A2(n14017), .ZN(n14521) );
  NAND2_X1 U11124 ( .A1(n10825), .A2(n10824), .ZN(n14419) );
  XNOR2_X1 U11125 ( .A(n11182), .B(n20180), .ZN(n13487) );
  INV_X2 U11126 ( .A(n20073), .ZN(n9645) );
  NAND2_X1 U11127 ( .A1(n11414), .A2(n11413), .ZN(n19988) );
  NOR2_X1 U11128 ( .A1(n14989), .A2(n14239), .ZN(n14967) );
  AND2_X1 U11129 ( .A1(n9835), .A2(n9834), .ZN(n11839) );
  INV_X1 U11130 ( .A(n12881), .ZN(n12824) );
  INV_X1 U11132 ( .A(n19269), .ZN(n19267) );
  INV_X1 U11133 ( .A(n12843), .ZN(n13355) );
  INV_X1 U11134 ( .A(n19998), .ZN(n19880) );
  XNOR2_X1 U11135 ( .A(n10463), .B(n10437), .ZN(n10603) );
  AND4_X2 U11136 ( .A1(n13407), .A2(n13406), .A3(n13405), .A4(n13404), .ZN(
        n9707) );
  AOI22_X2 U11137 ( .A1(n19704), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n19576), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13406) );
  AND2_X4 U11139 ( .A1(n9809), .A2(n13424), .ZN(n9942) );
  NOR2_X4 U11140 ( .A1(n16414), .A2(n17903), .ZN(n17815) );
  NOR2_X2 U11141 ( .A1(n12599), .A2(n16083), .ZN(n12597) );
  AND2_X4 U11142 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13134) );
  NAND2_X2 U11143 ( .A1(n11505), .A2(n11506), .ZN(n13358) );
  AND2_X2 U11144 ( .A1(n11465), .A2(n11487), .ZN(n11505) );
  NOR2_X2 U11145 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15740), .ZN(
        n12405) );
  INV_X2 U11146 ( .A(n15763), .ZN(n9939) );
  INV_X1 U11147 ( .A(n11319), .ZN(n9631) );
  AND2_X1 U11148 ( .A1(n13132), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9632) );
  AND2_X1 U11149 ( .A1(n13132), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9633) );
  NAND3_X2 U11150 ( .A1(n9910), .A2(n9967), .A3(n9909), .ZN(n10472) );
  AND2_X2 U11151 ( .A1(n9678), .A2(n9882), .ZN(n12396) );
  NOR2_X2 U11152 ( .A1(n12391), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12392) );
  AND2_X4 U11153 ( .A1(n13811), .A2(n16308), .ZN(n12033) );
  NOR2_X2 U11154 ( .A1(n15036), .A2(n12224), .ZN(n15039) );
  INV_X1 U11155 ( .A(n13176), .ZN(n9635) );
  INV_X1 U11157 ( .A(n9635), .ZN(n9637) );
  INV_X2 U11158 ( .A(n9638), .ZN(n9639) );
  INV_X2 U11159 ( .A(n9638), .ZN(n9640) );
  INV_X2 U11160 ( .A(n9638), .ZN(n9641) );
  INV_X1 U11161 ( .A(n10890), .ZN(n9642) );
  NOR2_X2 U11163 ( .A1(n15085), .A2(n10238), .ZN(n11728) );
  NOR2_X4 U11164 ( .A1(n17629), .A2(n17639), .ZN(n17677) );
  XNOR2_X1 U11166 ( .A(n12535), .B(n18842), .ZN(n17890) );
  NAND2_X2 U11169 ( .A1(n13894), .A2(n13893), .ZN(n14249) );
  OR2_X4 U11170 ( .A1(n16894), .A2(n12272), .ZN(n17181) );
  AND2_X4 U11172 ( .A1(n13307), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13302) );
  XNOR2_X2 U11173 ( .A(n12388), .B(n12387), .ZN(n17819) );
  NAND2_X2 U11174 ( .A1(n17833), .A2(n12385), .ZN(n12388) );
  NAND2_X1 U11175 ( .A1(n9939), .A2(n15762), .ZN(n15282) );
  NOR2_X1 U11176 ( .A1(n15216), .A2(n15327), .ZN(n15346) );
  NAND2_X1 U11177 ( .A1(n15548), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16199) );
  NAND2_X1 U11178 ( .A1(n15548), .A2(n9948), .ZN(n15216) );
  INV_X1 U11179 ( .A(n11236), .ZN(n14884) );
  NAND2_X1 U11180 ( .A1(n13478), .A2(n9683), .ZN(n15085) );
  NAND2_X1 U11181 ( .A1(n13441), .A2(n13440), .ZN(n13496) );
  AND2_X1 U11182 ( .A1(n13289), .A2(n13288), .ZN(n13441) );
  NOR2_X2 U11183 ( .A1(n17802), .A2(n18011), .ZN(n17702) );
  NAND2_X1 U11184 ( .A1(n10619), .A2(n10612), .ZN(n20812) );
  NAND2_X1 U11185 ( .A1(n9785), .A2(n13367), .ZN(n19785) );
  CLKBUF_X1 U11186 ( .A(n13508), .Z(n9656) );
  OAI22_X1 U11187 ( .A1(n13095), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11176), 
        .B2(n11159), .ZN(n10497) );
  OR2_X1 U11188 ( .A1(n18957), .A2(n10106), .ZN(n10105) );
  CLKBUF_X2 U11189 ( .A(n12631), .Z(n19021) );
  NAND2_X1 U11190 ( .A1(n20234), .A2(n10483), .ZN(n13176) );
  OAI22_X1 U11191 ( .A1(n15163), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19986), 
        .B2(n12596), .ZN(n13601) );
  NAND2_X2 U11192 ( .A1(n18689), .A2(n18679), .ZN(n18165) );
  AND2_X1 U11193 ( .A1(n13359), .A2(n11506), .ZN(n15590) );
  NAND2_X1 U11194 ( .A1(n11501), .A2(n11502), .ZN(n11506) );
  AOI21_X1 U11195 ( .B1(n12885), .B2(n10434), .A(n10433), .ZN(n10435) );
  INV_X4 U11196 ( .A(n10056), .ZN(n16860) );
  NOR2_X1 U11197 ( .A1(n13809), .A2(n11484), .ZN(n13133) );
  AND2_X1 U11198 ( .A1(n13132), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11966) );
  AND2_X1 U11199 ( .A1(n12927), .A2(n11459), .ZN(n13132) );
  AND2_X1 U11200 ( .A1(n10404), .A2(n14525), .ZN(n10416) );
  NOR2_X1 U11201 ( .A1(n17609), .A2(n17584), .ZN(n17582) );
  CLKBUF_X1 U11202 ( .A(n11420), .Z(n12260) );
  INV_X1 U11204 ( .A(n12536), .ZN(n17413) );
  INV_X1 U11205 ( .A(n13536), .ZN(n13070) );
  INV_X1 U11206 ( .A(n11420), .ZN(n19305) );
  INV_X1 U11208 ( .A(n13398), .ZN(n9957) );
  NAND2_X1 U11209 ( .A1(n11365), .A2(n11364), .ZN(n11431) );
  INV_X1 U11210 ( .A(n11443), .ZN(n11421) );
  OR2_X1 U11211 ( .A1(n10346), .A2(n10345), .ZN(n13122) );
  INV_X1 U11213 ( .A(n15626), .ZN(n12308) );
  INV_X4 U11214 ( .A(n21028), .ZN(n9646) );
  AND2_X2 U11216 ( .A1(n10278), .A2(n13307), .ZN(n10575) );
  INV_X1 U11217 ( .A(n15668), .ZN(n12309) );
  BUF_X4 U11218 ( .A(n10548), .Z(n9647) );
  OR2_X1 U11219 ( .A1(n12268), .A2(n12271), .ZN(n17080) );
  INV_X1 U11220 ( .A(n11319), .ZN(n9663) );
  OR3_X1 U11222 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n18675), .ZN(n12283) );
  NAND2_X2 U11223 ( .A1(n18866), .A2(n18859), .ZN(n16894) );
  AND2_X1 U11224 ( .A1(n11305), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11380) );
  INV_X2 U11225 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10613) );
  AND4_X1 U11226 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10113) );
  INV_X2 U11227 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11846) );
  NOR2_X1 U11228 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13107) );
  AND2_X1 U11229 ( .A1(n10190), .A2(n11259), .ZN(n14608) );
  OAI21_X1 U11230 ( .B1(n14529), .B2(n15934), .A(n11274), .ZN(n9915) );
  XNOR2_X1 U11231 ( .A(n14305), .B(n11267), .ZN(n14529) );
  INV_X1 U11232 ( .A(n15530), .ZN(n15517) );
  NOR2_X1 U11233 ( .A1(n15216), .A2(n15301), .ZN(n15186) );
  AOI21_X1 U11234 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(n15945) );
  OR2_X1 U11235 ( .A1(n14595), .A2(n14596), .ZN(n14593) );
  OR2_X1 U11236 ( .A1(n15941), .A2(n15940), .ZN(n15943) );
  NAND2_X1 U11237 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  NAND2_X1 U11238 ( .A1(n11250), .A2(n9974), .ZN(n9976) );
  AND2_X1 U11239 ( .A1(n10194), .A2(n10196), .ZN(n14458) );
  NAND2_X1 U11240 ( .A1(n13900), .A2(n13899), .ZN(n14101) );
  NAND2_X1 U11241 ( .A1(n10178), .A2(n14929), .ZN(n9848) );
  INV_X1 U11242 ( .A(n16418), .ZN(n17552) );
  NAND2_X1 U11243 ( .A1(n17553), .A2(n17813), .ZN(n16413) );
  NAND2_X1 U11244 ( .A1(n9881), .A2(n9880), .ZN(n16418) );
  NAND2_X1 U11245 ( .A1(n14103), .A2(n10225), .ZN(n10224) );
  INV_X1 U11246 ( .A(n16403), .ZN(n9881) );
  AND2_X1 U11247 ( .A1(n16403), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17553) );
  AND2_X1 U11248 ( .A1(n9979), .A2(n9709), .ZN(n9977) );
  OR2_X1 U11249 ( .A1(n17564), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10008) );
  AND2_X1 U11250 ( .A1(n14761), .A2(n14757), .ZN(n14739) );
  INV_X1 U11251 ( .A(n9980), .ZN(n9979) );
  AND2_X1 U11252 ( .A1(n10177), .A2(n14079), .ZN(n9974) );
  AND2_X1 U11253 ( .A1(n14716), .A2(n10179), .ZN(n10177) );
  NAND2_X1 U11254 ( .A1(n9837), .A2(n11208), .ZN(n13706) );
  INV_X1 U11255 ( .A(n9975), .ZN(n9972) );
  NAND2_X1 U11256 ( .A1(n9923), .A2(n19081), .ZN(n13898) );
  NAND2_X1 U11257 ( .A1(n9858), .A2(n13728), .ZN(n13637) );
  INV_X2 U11258 ( .A(n11236), .ZN(n9648) );
  INV_X1 U11259 ( .A(n14884), .ZN(n9975) );
  NAND2_X1 U11260 ( .A1(n10071), .A2(n9760), .ZN(n10076) );
  AND2_X1 U11261 ( .A1(n11236), .A2(n11233), .ZN(n13845) );
  INV_X1 U11262 ( .A(n14884), .ZN(n9649) );
  AND2_X1 U11263 ( .A1(n12401), .A2(n17949), .ZN(n9889) );
  AND2_X1 U11264 ( .A1(n13674), .A2(n13673), .ZN(n13893) );
  NOR2_X1 U11265 ( .A1(n13467), .A2(n13470), .ZN(n13468) );
  NAND2_X1 U11266 ( .A1(n9952), .A2(n9956), .ZN(n9810) );
  NAND2_X1 U11267 ( .A1(n12395), .A2(n10010), .ZN(n17648) );
  NAND2_X1 U11268 ( .A1(n11196), .A2(n11195), .ZN(n11197) );
  OAI21_X1 U11269 ( .B1(n11193), .B2(n9914), .A(n10628), .ZN(n13440) );
  OR2_X1 U11270 ( .A1(n11193), .A2(n11192), .ZN(n11196) );
  NOR2_X1 U11271 ( .A1(n15112), .A2(n15110), .ZN(n15104) );
  INV_X1 U11272 ( .A(n17684), .ZN(n12395) );
  NOR2_X1 U11273 ( .A1(n17685), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17684) );
  AND2_X1 U11274 ( .A1(n9927), .A2(n15496), .ZN(n9925) );
  AND2_X1 U11275 ( .A1(n14916), .A2(n14891), .ZN(n14867) );
  NAND2_X1 U11276 ( .A1(n12988), .A2(n11540), .ZN(n13460) );
  INV_X2 U11277 ( .A(n19572), .ZN(n19576) );
  OR2_X1 U11278 ( .A1(n13091), .A2(n13087), .ZN(n14892) );
  AND2_X1 U11279 ( .A1(n11537), .A2(n11539), .ZN(n12987) );
  OAI22_X1 U11280 ( .A1(n13402), .A2(n19380), .B1(n13658), .B2(n13401), .ZN(
        n13403) );
  NOR2_X1 U11281 ( .A1(n20330), .A2(n13625), .ZN(n20708) );
  NOR2_X1 U11282 ( .A1(n20330), .A2(n20214), .ZN(n20702) );
  NOR2_X1 U11283 ( .A1(n20330), .A2(n13540), .ZN(n20695) );
  NOR2_X1 U11284 ( .A1(n20330), .A2(n20185), .ZN(n20665) );
  NOR2_X1 U11285 ( .A1(n20330), .A2(n20206), .ZN(n20689) );
  NOR2_X1 U11286 ( .A1(n20330), .A2(n20199), .ZN(n20683) );
  NOR2_X1 U11287 ( .A1(n20330), .A2(n20193), .ZN(n20677) );
  NAND2_X1 U11288 ( .A1(n13065), .A2(n13064), .ZN(n13091) );
  NOR2_X1 U11289 ( .A1(n20330), .A2(n20228), .ZN(n20718) );
  INV_X1 U11290 ( .A(n17892), .ZN(n17904) );
  AND2_X1 U11291 ( .A1(n10610), .A2(n10172), .ZN(n10171) );
  NAND2_X1 U11292 ( .A1(n10516), .A2(n10515), .ZN(n10610) );
  INV_X2 U11293 ( .A(n13224), .ZN(n9650) );
  AND2_X1 U11294 ( .A1(n15883), .A2(n9753), .ZN(n14434) );
  XNOR2_X1 U11295 ( .A(n11168), .B(n11169), .ZN(n9839) );
  NAND2_X1 U11296 ( .A1(n10227), .A2(n11500), .ZN(n9830) );
  NAND2_X1 U11297 ( .A1(n12568), .A2(n16544), .ZN(n17903) );
  NAND2_X1 U11298 ( .A1(n13047), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11168) );
  NAND2_X1 U11299 ( .A1(n11167), .A2(n9744), .ZN(n11169) );
  AND2_X1 U11300 ( .A1(n10105), .A2(n19111), .ZN(n18934) );
  NAND2_X1 U11301 ( .A1(n10468), .A2(n10460), .ZN(n10595) );
  NAND2_X2 U11302 ( .A1(n13145), .A2(n10484), .ZN(n13095) );
  NAND2_X1 U11303 ( .A1(n11149), .A2(n11148), .ZN(n13126) );
  OAI21_X1 U11304 ( .B1(n20261), .B2(n11192), .A(n11163), .ZN(n13047) );
  NAND2_X1 U11306 ( .A1(n17365), .A2(n17270), .ZN(n17412) );
  AND2_X1 U11307 ( .A1(n10459), .A2(n10458), .ZN(n10460) );
  NAND2_X1 U11308 ( .A1(n11504), .A2(n11503), .ZN(n15594) );
  NAND2_X1 U11309 ( .A1(n15590), .A2(n11528), .ZN(n11504) );
  NAND2_X1 U11310 ( .A1(n11921), .A2(n11521), .ZN(n11526) );
  NOR2_X1 U11311 ( .A1(n13782), .A2(n13781), .ZN(n13925) );
  XNOR2_X1 U11312 ( .A(n12595), .B(n12594), .ZN(n15163) );
  INV_X2 U11313 ( .A(n19148), .ZN(n12991) );
  OR2_X1 U11314 ( .A1(n11502), .A2(n11501), .ZN(n13359) );
  AOI221_X1 U11315 ( .B1(n18051), .B2(n18687), .C1(n18050), .C2(n18687), .A(
        n18089), .ZN(n18068) );
  OR2_X1 U11316 ( .A1(n11520), .A2(n11519), .ZN(n11921) );
  INV_X1 U11317 ( .A(n13447), .ZN(n10027) );
  AOI21_X2 U11318 ( .B1(n15738), .B2(n15737), .A(n18732), .ZN(n18215) );
  NAND4_X1 U11319 ( .A1(n9851), .A2(n9857), .A3(n9855), .A4(n9856), .ZN(n11487) );
  NAND2_X1 U11320 ( .A1(n9808), .A2(n11489), .ZN(n11917) );
  OR2_X1 U11321 ( .A1(n13295), .A2(n13294), .ZN(n13447) );
  NOR2_X2 U11322 ( .A1(n12717), .A2(n19282), .ZN(n12718) );
  NOR2_X2 U11323 ( .A1(n17394), .A2(n12386), .ZN(n17813) );
  NOR2_X1 U11324 ( .A1(n15718), .A2(n9900), .ZN(n12518) );
  OR2_X2 U11325 ( .A1(n17466), .A2(n18724), .ZN(n17533) );
  AND2_X1 U11326 ( .A1(n12513), .A2(n12514), .ZN(n9900) );
  NAND2_X1 U11327 ( .A1(n18898), .A2(n16522), .ZN(n17427) );
  AND4_X1 U11328 ( .A1(n11469), .A2(n11468), .A3(n11467), .A4(n11466), .ZN(
        n11475) );
  NAND2_X1 U11329 ( .A1(n11462), .A2(n11461), .ZN(n9854) );
  AND2_X1 U11330 ( .A1(n12887), .A2(n12886), .ZN(n12132) );
  NAND2_X1 U11331 ( .A1(n9846), .A2(n9845), .ZN(n13326) );
  INV_X1 U11332 ( .A(n10637), .ZN(n10557) );
  NAND2_X1 U11333 ( .A1(n12941), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11457) );
  OR2_X1 U11334 ( .A1(n12933), .A2(n19986), .ZN(n11429) );
  CLKBUF_X1 U11335 ( .A(n11908), .Z(n14959) );
  AND2_X1 U11336 ( .A1(n16348), .A2(n9836), .ZN(n11908) );
  CLKBUF_X1 U11337 ( .A(n12712), .Z(n16328) );
  OR2_X1 U11338 ( .A1(n10417), .A2(n10430), .ZN(n13058) );
  NAND2_X1 U11339 ( .A1(n10384), .A2(n10385), .ZN(n10429) );
  NAND2_X1 U11340 ( .A1(n10428), .A2(n10408), .ZN(n13098) );
  NAND2_X1 U11341 ( .A1(n17278), .A2(n12529), .ZN(n12508) );
  INV_X1 U11342 ( .A(n18884), .ZN(n16544) );
  AND2_X1 U11343 ( .A1(n10434), .A2(n10402), .ZN(n10384) );
  NAND2_X1 U11344 ( .A1(n10362), .A2(n10361), .ZN(n10385) );
  INV_X1 U11345 ( .A(n15867), .ZN(n18688) );
  NAND2_X2 U11346 ( .A1(n11159), .A2(n10504), .ZN(n11143) );
  NOR3_X1 U11347 ( .A1(n12528), .A2(n15735), .A3(n12529), .ZN(n12505) );
  NAND2_X2 U11348 ( .A1(n12078), .A2(n12079), .ZN(n12257) );
  AND2_X2 U11349 ( .A1(n10069), .A2(n19310), .ZN(n12927) );
  AND2_X1 U11350 ( .A1(n11451), .A2(n10230), .ZN(n12925) );
  NAND2_X1 U11351 ( .A1(n13070), .A2(n9714), .ZN(n10362) );
  NAND2_X1 U11352 ( .A1(n20184), .A2(n9660), .ZN(n13565) );
  INV_X1 U11353 ( .A(n18262), .ZN(n12529) );
  NAND2_X1 U11354 ( .A1(n10405), .A2(n13070), .ZN(n10406) );
  INV_X1 U11355 ( .A(n11431), .ZN(n19310) );
  AND2_X1 U11356 ( .A1(n12370), .A2(n12369), .ZN(n17899) );
  AND2_X1 U11357 ( .A1(n12303), .A2(n9883), .ZN(n17408) );
  AOI211_X2 U11358 ( .C1(n17030), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n12478), .B(n12477), .ZN(n18262) );
  NAND2_X1 U11359 ( .A1(n10359), .A2(n20205), .ZN(n13304) );
  AOI211_X2 U11360 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n12282), .B(n12281), .ZN(n17394) );
  NAND2_X1 U11361 ( .A1(n10299), .A2(n10300), .ZN(n13536) );
  INV_X2 U11362 ( .A(U212), .ZN(n16460) );
  AND2_X1 U11363 ( .A1(n19988), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12774) );
  NAND2_X1 U11364 ( .A1(n9825), .A2(n9824), .ZN(n11430) );
  INV_X2 U11365 ( .A(n20184), .ZN(n13581) );
  INV_X1 U11366 ( .A(n11449), .ZN(n11418) );
  AND2_X1 U11367 ( .A1(n9806), .A2(n9805), .ZN(n11449) );
  NAND2_X1 U11368 ( .A1(n9820), .A2(n9819), .ZN(n9825) );
  NAND2_X1 U11369 ( .A1(n9822), .A2(n9821), .ZN(n9824) );
  OR2_X2 U11370 ( .A1(n16472), .A2(n16423), .ZN(n16474) );
  AND2_X1 U11371 ( .A1(n10399), .A2(n10398), .ZN(n10400) );
  NAND2_X1 U11372 ( .A1(n9803), .A2(n9801), .ZN(n19287) );
  NAND2_X1 U11373 ( .A1(n11359), .A2(n11358), .ZN(n11445) );
  AND4_X1 U11374 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10300) );
  AND4_X1 U11375 ( .A1(n10274), .A2(n10273), .A3(n10272), .A4(n10271), .ZN(
        n10287) );
  AND4_X1 U11376 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(
        n10399) );
  OR2_X2 U11377 ( .A1(n10336), .A2(n10335), .ZN(n9908) );
  NAND2_X2 U11378 ( .A1(n19880), .A2(n19869), .ZN(n19922) );
  AND4_X1 U11379 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10358) );
  AND3_X1 U11380 ( .A1(n11357), .A2(n11356), .A3(n11355), .ZN(n11359) );
  NAND2_X2 U11381 ( .A1(n18893), .A2(n18760), .ZN(n18810) );
  NAND2_X2 U11382 ( .A1(n18893), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18822) );
  AND2_X2 U11383 ( .A1(n12036), .A2(n11376), .ZN(n12194) );
  CLKBUF_X3 U11384 ( .A(n10548), .Z(n10949) );
  OR2_X2 U11385 ( .A1(n12271), .A2(n16894), .ZN(n10251) );
  BUF_X4 U11386 ( .A(n10391), .Z(n9652) );
  OR2_X1 U11387 ( .A1(n18841), .A2(n12269), .ZN(n10258) );
  AND2_X2 U11388 ( .A1(n13177), .A2(n10268), .ZN(n11013) );
  OR2_X2 U11389 ( .A1(n12271), .A2(n18675), .ZN(n10260) );
  INV_X2 U11390 ( .A(n20766), .ZN(n9653) );
  AND2_X2 U11391 ( .A1(n10278), .A2(n13177), .ZN(n10548) );
  AND2_X2 U11392 ( .A1(n10280), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9666) );
  AND2_X1 U11393 ( .A1(n10280), .A2(n10613), .ZN(n10330) );
  AND2_X2 U11394 ( .A1(n10280), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10329) );
  INV_X2 U11395 ( .A(n11319), .ZN(n9662) );
  INV_X2 U11396 ( .A(n16513), .ZN(n16515) );
  NAND2_X1 U11397 ( .A1(n13107), .A2(n10279), .ZN(n10890) );
  NAND2_X1 U11398 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18866), .ZN(
        n12268) );
  OR2_X1 U11399 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15726), .ZN(
        n12295) );
  NAND2_X1 U11400 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18841), .ZN(
        n12271) );
  AND2_X1 U11401 ( .A1(n10275), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10277) );
  NAND4_X2 U11402 ( .A1(n18841), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        n18852), .A4(n9988), .ZN(n17172) );
  AND2_X2 U11403 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13136) );
  AND2_X1 U11404 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10279) );
  AND2_X1 U11405 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13305) );
  NOR2_X2 U11406 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13306) );
  INV_X2 U11407 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11376) );
  AND2_X1 U11408 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10269) );
  NOR2_X2 U11409 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13177) );
  AND2_X1 U11410 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11306) );
  NAND2_X2 U11411 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18675) );
  NAND2_X1 U11412 ( .A1(n9850), .A2(n11253), .ZN(n11254) );
  AND2_X2 U11413 ( .A1(n13811), .A2(n11846), .ZN(n9654) );
  AND2_X2 U11414 ( .A1(n13811), .A2(n11846), .ZN(n11371) );
  NOR3_X1 U11415 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n16894), .ZN(n9655) );
  NOR3_X2 U11416 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n16894), .ZN(n12266) );
  NAND2_X2 U11417 ( .A1(n14136), .A2(n15524), .ZN(n14137) );
  XNOR2_X1 U11418 ( .A(n10595), .B(n10594), .ZN(n13508) );
  INV_X1 U11419 ( .A(n10638), .ZN(n10558) );
  NAND2_X1 U11420 ( .A1(n10542), .A2(n10629), .ZN(n10638) );
  AOI211_X2 U11421 ( .C1(n17940), .C2(n17912), .A(n17911), .B(n17910), .ZN(
        n17919) );
  NOR2_X1 U11422 ( .A1(n14329), .A2(n10204), .ZN(n14305) );
  NAND2_X2 U11423 ( .A1(n14135), .A2(n15519), .ZN(n14138) );
  NAND2_X1 U11425 ( .A1(n9785), .A2(n13378), .ZN(n19677) );
  NAND2_X2 U11426 ( .A1(n10570), .A2(n10569), .ZN(n13738) );
  OAI21_X1 U11427 ( .B1(n12990), .B2(n12767), .A(n11532), .ZN(n11536) );
  NAND2_X1 U11428 ( .A1(n14101), .A2(n14100), .ZN(n14104) );
  INV_X4 U11429 ( .A(n17172), .ZN(n17151) );
  OR2_X2 U11430 ( .A1(n14329), .A2(n10205), .ZN(n9697) );
  OAI22_X2 U11431 ( .A1(n14251), .A2(n10078), .B1(n14253), .B2(n15568), .ZN(
        n16223) );
  INV_X1 U11432 ( .A(n10412), .ZN(n9660) );
  NAND2_X4 U11433 ( .A1(n10400), .A2(n10401), .ZN(n10412) );
  OAI21_X2 U11434 ( .B1(n13775), .B2(n9906), .A(n9905), .ZN(n13982) );
  NAND3_X2 U11435 ( .A1(n10647), .A2(n13776), .A3(n13915), .ZN(n13775) );
  NOR2_X4 U11436 ( .A1(n13496), .A2(n9918), .ZN(n13915) );
  AND2_X2 U11437 ( .A1(n13811), .A2(n16308), .ZN(n9661) );
  NAND2_X2 U11438 ( .A1(n12965), .A2(n13581), .ZN(n12752) );
  NOR2_X4 U11439 ( .A1(n10407), .A2(n9903), .ZN(n12965) );
  NOR2_X1 U11440 ( .A1(n14419), .A2(n9921), .ZN(n14406) );
  NAND2_X2 U11441 ( .A1(n10479), .A2(n10478), .ZN(n13145) );
  AOI22_X2 U11442 ( .A1(n16404), .A2(n17892), .B1(n17815), .B2(n18093), .ZN(
        n17802) );
  AND2_X2 U11443 ( .A1(n10280), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9665) );
  AND2_X1 U11444 ( .A1(n13305), .A2(n10266), .ZN(n9667) );
  AND2_X1 U11445 ( .A1(n13305), .A2(n10266), .ZN(n9668) );
  AND2_X1 U11446 ( .A1(n13305), .A2(n10266), .ZN(n10347) );
  OAI21_X2 U11447 ( .B1(n18680), .B2(n18667), .A(n18666), .ZN(n18687) );
  AND2_X4 U11448 ( .A1(n10270), .A2(n13305), .ZN(n11038) );
  AND2_X2 U11449 ( .A1(n10278), .A2(n13307), .ZN(n9669) );
  INV_X4 U11450 ( .A(n10894), .ZN(n9670) );
  AOI21_X1 U11452 ( .B1(n9956), .B2(n9957), .A(n12094), .ZN(n9953) );
  AOI21_X1 U11453 ( .B1(n11848), .B2(n11843), .A(n11844), .ZN(n11871) );
  NAND2_X1 U11454 ( .A1(n17468), .A2(n16544), .ZN(n15716) );
  NOR2_X1 U11455 ( .A1(n10423), .A2(n20728), .ZN(n10795) );
  AND2_X1 U11456 ( .A1(n11087), .A2(n13536), .ZN(n11133) );
  NOR2_X1 U11457 ( .A1(n15061), .A2(n10255), .ZN(n11808) );
  AND2_X1 U11458 ( .A1(n11786), .A2(n9774), .ZN(n10255) );
  INV_X1 U11459 ( .A(n11808), .ZN(n10234) );
  NAND2_X1 U11460 ( .A1(n10221), .A2(n10217), .ZN(n10216) );
  INV_X1 U11461 ( .A(n14205), .ZN(n10217) );
  INV_X1 U11462 ( .A(n15376), .ZN(n10221) );
  INV_X1 U11463 ( .A(n13426), .ZN(n15158) );
  NAND2_X1 U11464 ( .A1(n12921), .A2(n12920), .ZN(n12954) );
  AND2_X1 U11465 ( .A1(n10556), .A2(n10555), .ZN(n10637) );
  AND2_X2 U11466 ( .A1(n13107), .A2(n10276), .ZN(n10391) );
  NOR2_X1 U11467 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10275), .ZN(
        n10276) );
  NAND2_X1 U11468 ( .A1(n16348), .A2(n12774), .ZN(n11460) );
  NAND2_X1 U11469 ( .A1(n13400), .A2(n9957), .ZN(n9956) );
  NOR2_X1 U11470 ( .A1(n14378), .A2(n10203), .ZN(n10202) );
  INV_X1 U11471 ( .A(n14393), .ZN(n10203) );
  NAND2_X1 U11472 ( .A1(n14404), .A2(n9922), .ZN(n9921) );
  INV_X1 U11473 ( .A(n14418), .ZN(n9922) );
  INV_X1 U11474 ( .A(n11133), .ZN(n11130) );
  OR2_X1 U11475 ( .A1(n13068), .A2(n10411), .ZN(n9911) );
  INV_X1 U11476 ( .A(n10586), .ZN(n10498) );
  OAI21_X1 U11477 ( .B1(n9721), .B2(n9968), .A(P1_STATE2_REG_0__SCAN_IN), .ZN(
        n9967) );
  NOR2_X1 U11478 ( .A1(n10298), .A2(n10297), .ZN(n10299) );
  NOR2_X1 U11479 ( .A1(n14140), .A2(n14139), .ZN(n10148) );
  AND2_X1 U11480 ( .A1(n13398), .A2(n12774), .ZN(n9836) );
  AND2_X1 U11481 ( .A1(n9737), .A2(n13839), .ZN(n10244) );
  AND2_X1 U11482 ( .A1(n12928), .A2(n11450), .ZN(n12056) );
  NOR2_X1 U11483 ( .A1(n10094), .A2(n13043), .ZN(n10093) );
  INV_X1 U11484 ( .A(n13608), .ZN(n10094) );
  NAND2_X1 U11485 ( .A1(n11917), .A2(n11522), .ZN(n10087) );
  OR2_X1 U11486 ( .A1(n15280), .A2(n15237), .ZN(n9936) );
  NOR2_X1 U11487 ( .A1(n15237), .A2(n15234), .ZN(n9937) );
  NAND2_X1 U11488 ( .A1(n16178), .A2(n9929), .ZN(n9928) );
  INV_X1 U11489 ( .A(n16177), .ZN(n9929) );
  INV_X1 U11490 ( .A(n13678), .ZN(n13894) );
  AND2_X1 U11491 ( .A1(n13890), .A2(n13889), .ZN(n14247) );
  NAND2_X1 U11492 ( .A1(n10129), .A2(n13338), .ZN(n10133) );
  INV_X1 U11493 ( .A(n12150), .ZN(n10129) );
  NAND2_X1 U11494 ( .A1(n11449), .A2(n19287), .ZN(n11484) );
  MUX2_X1 U11495 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11894), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12909) );
  NAND2_X1 U11496 ( .A1(n11330), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11331) );
  XNOR2_X1 U11497 ( .A(n17413), .B(n12535), .ZN(n12358) );
  NAND2_X1 U11498 ( .A1(n17365), .A2(n18237), .ZN(n12506) );
  AOI21_X1 U11499 ( .B1(n15725), .B2(n15716), .A(n9746), .ZN(n15865) );
  OAI21_X1 U11500 ( .B1(n11172), .B2(n10592), .A(n9912), .ZN(n13244) );
  AOI21_X1 U11501 ( .B1(n10593), .B2(n9914), .A(n9913), .ZN(n9912) );
  INV_X1 U11502 ( .A(n10609), .ZN(n9913) );
  NAND2_X1 U11503 ( .A1(n14614), .A2(n11252), .ZN(n11253) );
  NAND2_X1 U11504 ( .A1(n11147), .A2(n11146), .ZN(n11148) );
  OAI21_X1 U11505 ( .B1(n11147), .B2(n11145), .A(n11144), .ZN(n11149) );
  INV_X1 U11506 ( .A(n15244), .ZN(n10112) );
  NAND2_X1 U11507 ( .A1(n10234), .A2(n10231), .ZN(n9834) );
  NAND2_X1 U11508 ( .A1(n11809), .A2(n10233), .ZN(n9835) );
  NOR2_X1 U11509 ( .A1(n11807), .A2(n10232), .ZN(n10231) );
  NAND2_X1 U11510 ( .A1(n11728), .A2(n11729), .ZN(n11730) );
  AOI21_X1 U11511 ( .B1(n15194), .B2(n9776), .A(n9694), .ZN(n9826) );
  NOR2_X1 U11512 ( .A1(n15194), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9827) );
  NAND2_X1 U11513 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  NOR2_X1 U11514 ( .A1(n13680), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10075) );
  INV_X1 U11515 ( .A(n13680), .ZN(n10070) );
  INV_X1 U11516 ( .A(n19781), .ZN(n19708) );
  INV_X1 U11517 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17214) );
  NAND2_X1 U11518 ( .A1(n10006), .A2(n18843), .ZN(n10004) );
  OR2_X1 U11519 ( .A1(n12407), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12408) );
  AOI21_X1 U11520 ( .B1(n16052), .B2(n19248), .A(n15314), .ZN(n15320) );
  OR2_X1 U11521 ( .A1(n14259), .A2(n9944), .ZN(n9943) );
  AND2_X1 U11522 ( .A1(n15336), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9944) );
  CLKBUF_X1 U11523 ( .A(n10367), .Z(n11063) );
  NAND2_X1 U11524 ( .A1(n10171), .A2(n10517), .ZN(n10630) );
  INV_X1 U11525 ( .A(n9745), .ZN(n10172) );
  INV_X1 U11526 ( .A(n12898), .ZN(n10504) );
  NOR2_X1 U11527 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U11528 ( .A1(n11434), .A2(n11449), .ZN(n11435) );
  NAND2_X1 U11529 ( .A1(n12934), .A2(n19291), .ZN(n11436) );
  NOR2_X1 U11530 ( .A1(n13398), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12079) );
  AND2_X1 U11531 ( .A1(n11420), .A2(n11443), .ZN(n11439) );
  AOI21_X1 U11532 ( .B1(n19291), .B2(n11479), .A(n12922), .ZN(n11399) );
  AND2_X2 U11533 ( .A1(n11439), .A2(n11430), .ZN(n10069) );
  NAND2_X1 U11534 ( .A1(n11430), .A2(n11431), .ZN(n11419) );
  AND2_X1 U11535 ( .A1(n11852), .A2(n11842), .ZN(n11848) );
  OR2_X1 U11536 ( .A1(n11851), .A2(n11850), .ZN(n11852) );
  NOR2_X1 U11537 ( .A1(n12374), .A2(n17408), .ZN(n12376) );
  AOI21_X1 U11538 ( .B1(n17086), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(n9893), .ZN(n9892) );
  OAI21_X1 U11539 ( .B1(n21028), .B2(n17189), .A(n9894), .ZN(n9893) );
  NAND2_X1 U11540 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n9894) );
  AND2_X1 U11541 ( .A1(n11142), .A2(n11140), .ZN(n11280) );
  INV_X1 U11542 ( .A(n14367), .ZN(n10201) );
  AND2_X1 U11543 ( .A1(n10197), .A2(n14508), .ZN(n10196) );
  NOR2_X1 U11544 ( .A1(n13991), .A2(n10198), .ZN(n10197) );
  INV_X1 U11545 ( .A(n14515), .ZN(n10198) );
  NAND2_X1 U11546 ( .A1(n9648), .A2(n14781), .ZN(n10183) );
  NAND2_X1 U11547 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  NAND2_X1 U11548 ( .A1(n9971), .A2(n10191), .ZN(n10186) );
  NAND2_X1 U11549 ( .A1(n10188), .A2(n9971), .ZN(n10187) );
  NAND2_X1 U11550 ( .A1(n9648), .A2(n9778), .ZN(n10188) );
  INV_X1 U11551 ( .A(n9778), .ZN(n10189) );
  OR2_X1 U11552 ( .A1(n10310), .A2(n10309), .ZN(n11222) );
  INV_X1 U11553 ( .A(n10029), .ZN(n10028) );
  INV_X1 U11554 ( .A(n14057), .ZN(n14048) );
  NAND2_X1 U11555 ( .A1(n13530), .A2(n10030), .ZN(n10029) );
  INV_X1 U11556 ( .A(n13446), .ZN(n10030) );
  NAND2_X1 U11557 ( .A1(n13291), .A2(n14293), .ZN(n14057) );
  NAND2_X1 U11558 ( .A1(n9839), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11171) );
  AND3_X1 U11559 ( .A1(n10264), .A2(n10447), .A3(n10446), .ZN(n11164) );
  AND2_X1 U11560 ( .A1(n10454), .A2(n10175), .ZN(n10174) );
  NAND2_X1 U11561 ( .A1(n10449), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10175) );
  INV_X1 U11562 ( .A(n10449), .ZN(n10176) );
  INV_X1 U11563 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20489) );
  AND2_X1 U11564 ( .A1(n9691), .A2(n15070), .ZN(n10160) );
  NOR2_X1 U11565 ( .A1(n10153), .A2(n10155), .ZN(n10151) );
  INV_X1 U11566 ( .A(n14151), .ZN(n10155) );
  NAND2_X1 U11567 ( .A1(n14220), .A2(n14167), .ZN(n14156) );
  NAND2_X1 U11568 ( .A1(n14126), .A2(n12645), .ZN(n14140) );
  NOR2_X1 U11569 ( .A1(n9854), .A2(n11441), .ZN(n9851) );
  NAND2_X1 U11570 ( .A1(n11514), .A2(n11513), .ZN(n11520) );
  NAND2_X1 U11571 ( .A1(n10243), .A2(n16105), .ZN(n10242) );
  INV_X1 U11572 ( .A(n15087), .ZN(n10243) );
  NOR2_X1 U11573 ( .A1(n10242), .A2(n10241), .ZN(n10240) );
  INV_X1 U11574 ( .A(n15080), .ZN(n10241) );
  NOR2_X1 U11575 ( .A1(n12592), .A2(n10124), .ZN(n10123) );
  INV_X1 U11576 ( .A(n15083), .ZN(n10101) );
  AND2_X1 U11577 ( .A1(n14170), .A2(n13426), .ZN(n14186) );
  INV_X1 U11578 ( .A(n16345), .ZN(n12770) );
  NOR2_X1 U11579 ( .A1(n10098), .A2(n10100), .ZN(n10097) );
  INV_X1 U11580 ( .A(n10259), .ZN(n10100) );
  NAND2_X1 U11581 ( .A1(n10099), .A2(n12665), .ZN(n10098) );
  INV_X1 U11582 ( .A(n14982), .ZN(n10099) );
  NOR2_X1 U11583 ( .A1(n15215), .A2(n10219), .ZN(n10218) );
  OR2_X1 U11584 ( .A1(n16084), .A2(n15158), .ZN(n14230) );
  NOR2_X1 U11585 ( .A1(n15483), .A2(n10103), .ZN(n10102) );
  INV_X1 U11586 ( .A(n13841), .ZN(n10103) );
  INV_X1 U11587 ( .A(n13257), .ZN(n10091) );
  NOR2_X1 U11588 ( .A1(n13606), .A2(n10141), .ZN(n10140) );
  INV_X1 U11589 ( .A(n15556), .ZN(n10141) );
  NAND2_X1 U11590 ( .A1(n14104), .A2(n9951), .ZN(n15532) );
  NOR2_X1 U11591 ( .A1(n10224), .A2(n16227), .ZN(n9951) );
  INV_X1 U11592 ( .A(n12257), .ZN(n14968) );
  NOR2_X1 U11593 ( .A1(n14249), .A2(n14248), .ZN(n14252) );
  NAND2_X1 U11594 ( .A1(n13425), .A2(n12094), .ZN(n9782) );
  NAND2_X1 U11595 ( .A1(n13636), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9815) );
  NAND2_X1 U11596 ( .A1(n13637), .A2(n9817), .ZN(n9816) );
  OR2_X1 U11597 ( .A1(n13636), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9817) );
  INV_X1 U11598 ( .A(n11353), .ZN(n9821) );
  NOR2_X1 U11599 ( .A1(n11354), .A2(n11376), .ZN(n9822) );
  INV_X1 U11600 ( .A(n11343), .ZN(n9819) );
  INV_X1 U11601 ( .A(n19961), .ZN(n19536) );
  AND2_X1 U11602 ( .A1(n11889), .A2(n11872), .ZN(n12060) );
  NAND3_X1 U11603 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18859), .ZN(n12269) );
  NAND2_X1 U11604 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10014) );
  NOR2_X1 U11605 ( .A1(n16378), .A2(n10064), .ZN(n10063) );
  NAND2_X1 U11606 ( .A1(n17591), .A2(n10012), .ZN(n10011) );
  INV_X1 U11607 ( .A(n12402), .ZN(n10012) );
  NOR2_X1 U11608 ( .A1(n17824), .A2(n9879), .ZN(n12559) );
  NOR4_X1 U11609 ( .A1(n12514), .A2(n15735), .A3(n12506), .A4(n12508), .ZN(
        n12515) );
  NAND2_X1 U11610 ( .A1(n15716), .A2(n17427), .ZN(n16539) );
  INV_X1 U11611 ( .A(n12516), .ZN(n18680) );
  NOR2_X1 U11612 ( .A1(n9897), .A2(n12427), .ZN(n9896) );
  AND2_X1 U11613 ( .A1(n9659), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9897)
         );
  AND2_X1 U11614 ( .A1(n13796), .A2(n13797), .ZN(n13999) );
  NAND2_X1 U11615 ( .A1(n13036), .A2(n12882), .ZN(n13583) );
  NAND2_X1 U11616 ( .A1(n10015), .A2(n9765), .ZN(n14369) );
  XNOR2_X1 U11617 ( .A(n11081), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13568) );
  OR2_X1 U11618 ( .A1(n11080), .A2(n14291), .ZN(n11081) );
  INV_X1 U11619 ( .A(n10206), .ZN(n10204) );
  OR2_X1 U11620 ( .A1(n14673), .A2(n11052), .ZN(n10926) );
  NAND2_X1 U11621 ( .A1(n14406), .A2(n10202), .ZN(n14381) );
  AND2_X1 U11622 ( .A1(n10864), .A2(n10863), .ZN(n14404) );
  OR2_X1 U11623 ( .A1(n14691), .A2(n11052), .ZN(n10864) );
  NAND2_X1 U11624 ( .A1(n10679), .A2(n9907), .ZN(n9906) );
  OAI21_X1 U11625 ( .B1(n13775), .B2(n13917), .A(n10695), .ZN(n9905) );
  INV_X1 U11626 ( .A(n10695), .ZN(n9907) );
  AND2_X1 U11627 ( .A1(n10647), .A2(n13915), .ZN(n13737) );
  AOI21_X1 U11628 ( .B1(n11209), .B2(n10795), .A(n10646), .ZN(n13591) );
  NAND2_X1 U11629 ( .A1(n13246), .A2(n10609), .ZN(n13289) );
  OR2_X1 U11630 ( .A1(n13126), .A2(n20001), .ZN(n12966) );
  INV_X1 U11631 ( .A(n11254), .ZN(n14632) );
  NAND2_X1 U11632 ( .A1(n9976), .A2(n11249), .ZN(n14653) );
  AOI21_X1 U11633 ( .B1(n11250), .B2(n9648), .A(n9724), .ZN(n9847) );
  NAND2_X1 U11634 ( .A1(n9648), .A2(n9973), .ZN(n9970) );
  OAI21_X1 U11635 ( .B1(n9705), .B2(n15956), .A(n11235), .ZN(n9980) );
  NAND2_X1 U11636 ( .A1(n9722), .A2(n15955), .ZN(n9978) );
  XNOR2_X1 U11637 ( .A(n10497), .B(n10496), .ZN(n10587) );
  AOI21_X1 U11638 ( .B1(n10472), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10473), .ZN(n10482) );
  INV_X1 U11639 ( .A(n10464), .ZN(n9840) );
  INV_X1 U11640 ( .A(n20819), .ZN(n20518) );
  AOI22_X1 U11641 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U11642 ( .A1(n9656), .A2(n13510), .ZN(n20516) );
  NAND2_X1 U11643 ( .A1(n16039), .A2(n13521), .ZN(n20330) );
  NAND2_X1 U11644 ( .A1(n11407), .A2(n11376), .ZN(n11414) );
  NAND2_X1 U11645 ( .A1(n11412), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11413) );
  INV_X1 U11646 ( .A(n14949), .ZN(n10168) );
  INV_X1 U11647 ( .A(n14226), .ZN(n10169) );
  NAND2_X1 U11648 ( .A1(n14951), .A2(n15154), .ZN(n10166) );
  NAND2_X1 U11649 ( .A1(n15104), .A2(n9764), .ZN(n14989) );
  INV_X1 U11650 ( .A(n14986), .ZN(n10126) );
  INV_X1 U11651 ( .A(n12681), .ZN(n12650) );
  NOR2_X1 U11652 ( .A1(n12651), .A2(n10163), .ZN(n10162) );
  NAND2_X1 U11653 ( .A1(n19021), .A2(n16154), .ZN(n10111) );
  AND2_X1 U11654 ( .A1(n14197), .A2(n14220), .ZN(n12681) );
  INV_X1 U11655 ( .A(n18946), .ZN(n10107) );
  AOI21_X1 U11656 ( .B1(n18965), .B2(n18966), .A(n12631), .ZN(n18957) );
  OR2_X1 U11657 ( .A1(n18957), .A2(n18958), .ZN(n10108) );
  NAND2_X1 U11658 ( .A1(n12648), .A2(n14163), .ZN(n14167) );
  INV_X1 U11659 ( .A(n14176), .ZN(n12648) );
  NAND2_X1 U11660 ( .A1(n9696), .A2(n15154), .ZN(n14220) );
  AND2_X1 U11661 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12620) );
  NAND2_X1 U11662 ( .A1(n11488), .A2(n16308), .ZN(n9808) );
  INV_X1 U11663 ( .A(n11919), .ZN(n9798) );
  INV_X1 U11664 ( .A(n11526), .ZN(n11918) );
  NAND2_X1 U11665 ( .A1(n11526), .A2(n11524), .ZN(n9800) );
  NAND2_X1 U11666 ( .A1(n10234), .A2(n11806), .ZN(n15047) );
  NAND2_X1 U11667 ( .A1(n15104), .A2(n10127), .ZN(n14987) );
  AND2_X1 U11668 ( .A1(n14206), .A2(n12259), .ZN(n12078) );
  OAI22_X1 U11669 ( .A1(n15125), .A2(n9832), .B1(n11730), .B2(n15073), .ZN(
        n15072) );
  NAND2_X1 U11670 ( .A1(n11747), .A2(n9833), .ZN(n9832) );
  INV_X1 U11671 ( .A(n15128), .ZN(n9833) );
  INV_X1 U11672 ( .A(n16109), .ZN(n9831) );
  AND2_X1 U11673 ( .A1(n15039), .A2(n9752), .ZN(n13952) );
  INV_X1 U11674 ( .A(n13964), .ZN(n10142) );
  AND2_X1 U11675 ( .A1(n15039), .A2(n10144), .ZN(n13819) );
  NAND2_X1 U11676 ( .A1(n15039), .A2(n13544), .ZN(n13745) );
  NOR2_X1 U11677 ( .A1(n10133), .A2(n12155), .ZN(n10131) );
  AND2_X1 U11678 ( .A1(n11539), .A2(n11538), .ZN(n11540) );
  NAND2_X1 U11679 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  NOR2_X1 U11680 ( .A1(n10121), .A2(n15246), .ZN(n10119) );
  INV_X1 U11681 ( .A(n12589), .ZN(n10120) );
  CLKBUF_X1 U11682 ( .A(n12602), .Z(n12603) );
  NAND2_X1 U11683 ( .A1(n13934), .A2(n13933), .ZN(n13932) );
  AND3_X1 U11684 ( .A1(n11965), .A2(n11964), .A3(n11963), .ZN(n13627) );
  AND2_X1 U11685 ( .A1(n9949), .A2(n15354), .ZN(n9948) );
  NAND2_X1 U11686 ( .A1(n9814), .A2(n9812), .ZN(n15391) );
  NAND2_X1 U11687 ( .A1(n15390), .A2(n9813), .ZN(n9812) );
  INV_X1 U11688 ( .A(n15405), .ZN(n9813) );
  NOR2_X1 U11689 ( .A1(n14195), .A2(n15293), .ZN(n10222) );
  AND2_X1 U11690 ( .A1(n9934), .A2(n9932), .ZN(n9931) );
  NAND2_X1 U11691 ( .A1(n9937), .A2(n15233), .ZN(n9932) );
  AND2_X1 U11692 ( .A1(n9936), .A2(n15472), .ZN(n9934) );
  INV_X1 U11693 ( .A(n9937), .ZN(n9933) );
  AOI21_X1 U11694 ( .B1(n14178), .B2(n19253), .A(n15761), .ZN(n10080) );
  NAND2_X1 U11695 ( .A1(n15039), .A2(n10143), .ZN(n13963) );
  NOR2_X1 U11696 ( .A1(n15035), .A2(n13474), .ZN(n13934) );
  NAND2_X1 U11697 ( .A1(n14104), .A2(n10223), .ZN(n15572) );
  INV_X1 U11698 ( .A(n10224), .ZN(n10223) );
  NAND2_X1 U11699 ( .A1(n9863), .A2(n9861), .ZN(n9790) );
  NAND2_X1 U11700 ( .A1(n9781), .A2(n19234), .ZN(n10073) );
  INV_X1 U11701 ( .A(n9810), .ZN(n9783) );
  AOI21_X1 U11702 ( .B1(n12867), .B2(n11528), .A(n11510), .ZN(n12903) );
  XNOR2_X1 U11703 ( .A(n15594), .B(n11511), .ZN(n12904) );
  NAND2_X1 U11704 ( .A1(n12904), .A2(n12903), .ZN(n9828) );
  OR2_X1 U11705 ( .A1(n19412), .A2(n19275), .ZN(n19511) );
  AND2_X1 U11706 ( .A1(n19412), .A2(n19275), .ZN(n19567) );
  INV_X1 U11707 ( .A(n19567), .ZN(n19580) );
  AND2_X1 U11708 ( .A1(n19412), .A2(n19953), .ZN(n19932) );
  INV_X1 U11709 ( .A(n19713), .ZN(n19635) );
  OR2_X1 U11710 ( .A1(n19412), .A2(n19953), .ZN(n19706) );
  NAND2_X1 U11711 ( .A1(n9785), .A2(n9784), .ZN(n13654) );
  INV_X1 U11712 ( .A(n13383), .ZN(n9784) );
  NOR2_X1 U11713 ( .A1(n19566), .A2(n19961), .ZN(n19713) );
  AND2_X1 U11714 ( .A1(n15861), .A2(n19986), .ZN(n19781) );
  NOR2_X1 U11715 ( .A1(n18678), .A2(n16539), .ZN(n18710) );
  AOI21_X1 U11716 ( .B1(n10056), .B2(n16595), .A(n16588), .ZN(n10050) );
  AND2_X1 U11717 ( .A1(n16603), .A2(n10056), .ZN(n16594) );
  OR2_X1 U11718 ( .A1(n16594), .A2(n16595), .ZN(n10051) );
  NAND2_X1 U11719 ( .A1(n10056), .A2(n17588), .ZN(n10055) );
  NAND2_X1 U11720 ( .A1(n16627), .A2(n10056), .ZN(n10054) );
  NAND2_X1 U11722 ( .A1(n10054), .A2(n10052), .ZN(n16603) );
  NOR2_X1 U11723 ( .A1(n10053), .A2(n17568), .ZN(n10052) );
  INV_X1 U11724 ( .A(n10055), .ZN(n10053) );
  OR2_X1 U11725 ( .A1(n16629), .A2(n17604), .ZN(n16627) );
  AND2_X1 U11726 ( .A1(n10061), .A2(n12574), .ZN(n10059) );
  NOR2_X1 U11727 ( .A1(n10002), .A2(n9998), .ZN(n9997) );
  INV_X1 U11728 ( .A(n12437), .ZN(n10002) );
  OAI21_X1 U11729 ( .B1(n17190), .B2(n17235), .A(n9999), .ZN(n9998) );
  NOR3_X1 U11730 ( .A1(n9770), .A2(n9993), .A3(n9990), .ZN(n9989) );
  NAND2_X1 U11731 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .ZN(n9993) );
  INV_X1 U11732 ( .A(n9991), .ZN(n9990) );
  CLKBUF_X1 U11733 ( .A(n12295), .Z(n17215) );
  AOI21_X1 U11734 ( .B1(n17192), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n9888), .ZN(n12299) );
  AND3_X1 U11735 ( .A1(n9887), .A2(n9886), .A3(P3_INSTQUEUE_REG_0__3__SCAN_IN), 
        .ZN(n9888) );
  NAND2_X1 U11736 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9885) );
  NOR2_X1 U11737 ( .A1(n12320), .A2(n12319), .ZN(n12321) );
  OAI21_X1 U11738 ( .B1(n15865), .B2(n15864), .A(n18723), .ZN(n15866) );
  AND2_X1 U11739 ( .A1(n17536), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17534) );
  NAND2_X1 U11740 ( .A1(n12400), .A2(n10262), .ZN(n12401) );
  NAND2_X1 U11741 ( .A1(n17694), .A2(n17951), .ZN(n12400) );
  NOR2_X1 U11742 ( .A1(n17826), .A2(n17825), .ZN(n17824) );
  AND2_X1 U11743 ( .A1(n13028), .A2(n13064), .ZN(n20103) );
  NAND2_X1 U11744 ( .A1(n20103), .A2(n20224), .ZN(n14523) );
  INV_X1 U11745 ( .A(n11078), .ZN(n11079) );
  INV_X1 U11746 ( .A(n15963), .ZN(n15950) );
  NAND2_X1 U11747 ( .A1(n14786), .A2(n9778), .ZN(n10021) );
  NOR2_X1 U11748 ( .A1(n14095), .A2(n10020), .ZN(n10019) );
  INV_X1 U11749 ( .A(n14074), .ZN(n10020) );
  NAND2_X1 U11750 ( .A1(n11263), .A2(n9971), .ZN(n11264) );
  NAND2_X1 U11751 ( .A1(n11261), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9843) );
  XNOR2_X1 U11752 ( .A(n14072), .B(n10022), .ZN(n14288) );
  INV_X1 U11753 ( .A(n14073), .ZN(n10022) );
  XNOR2_X1 U11754 ( .A(n11272), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14785) );
  INV_X1 U11755 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20588) );
  INV_X1 U11756 ( .A(n20434), .ZN(n20455) );
  AND2_X1 U11757 ( .A1(n16052), .A2(n19076), .ZN(n16053) );
  INV_X1 U11758 ( .A(n19076), .ZN(n19107) );
  OR2_X1 U11759 ( .A1(n16061), .A2(n12991), .ZN(n12022) );
  INV_X1 U11760 ( .A(n19145), .ZN(n19127) );
  NOR2_X1 U11761 ( .A1(n12027), .A2(n12026), .ZN(n12046) );
  INV_X1 U11762 ( .A(n15131), .ZN(n16127) );
  AND2_X1 U11763 ( .A1(n12064), .A2(n12063), .ZN(n19169) );
  OAI21_X1 U11764 ( .B1(n12020), .B2(n10259), .A(n14958), .ZN(n16061) );
  NOR2_X1 U11765 ( .A1(n16181), .A2(n14178), .ZN(n16166) );
  NAND2_X1 U11766 ( .A1(n16166), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16165) );
  AND2_X1 U11767 ( .A1(n19231), .A2(n19952), .ZN(n16239) );
  INV_X1 U11768 ( .A(n16240), .ZN(n19224) );
  XNOR2_X1 U11769 ( .A(n14965), .B(n14964), .ZN(n16098) );
  AND2_X1 U11770 ( .A1(n15058), .A2(n9768), .ZN(n14965) );
  INV_X1 U11771 ( .A(n15306), .ZN(n10215) );
  XNOR2_X1 U11772 ( .A(n10209), .B(n15161), .ZN(n15310) );
  NAND2_X1 U11773 ( .A1(n10210), .A2(n9713), .ZN(n10209) );
  OR2_X1 U11774 ( .A1(n16057), .A2(n16290), .ZN(n15318) );
  AND2_X1 U11775 ( .A1(n9947), .A2(n14258), .ZN(n15185) );
  NAND2_X1 U11776 ( .A1(n15346), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9947) );
  AND2_X1 U11777 ( .A1(n14985), .A2(n14984), .ZN(n15325) );
  NOR2_X1 U11778 ( .A1(n15757), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9787) );
  AND2_X1 U11779 ( .A1(n9926), .A2(n9927), .ZN(n15499) );
  NAND2_X1 U11780 ( .A1(n16170), .A2(n19250), .ZN(n9788) );
  INV_X1 U11781 ( .A(n19255), .ZN(n16273) );
  INV_X1 U11782 ( .A(n15579), .ZN(n15787) );
  AND2_X1 U11783 ( .A1(n12954), .A2(n12946), .ZN(n19248) );
  INV_X1 U11784 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19959) );
  NOR2_X1 U11785 ( .A1(n19634), .A2(n19512), .ZN(n19430) );
  INV_X1 U11786 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18735) );
  NAND2_X1 U11787 ( .A1(n18723), .A2(n18711), .ZN(n17466) );
  NOR2_X1 U11788 ( .A1(n18710), .A2(n17466), .ZN(n18899) );
  INV_X1 U11789 ( .A(n16572), .ZN(n10034) );
  NOR2_X1 U11790 ( .A1(n16573), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10036) );
  INV_X1 U11791 ( .A(n16889), .ZN(n16874) );
  INV_X1 U11792 ( .A(n17365), .ZN(n18268) );
  NAND2_X1 U11793 ( .A1(n17364), .A2(n9982), .ZN(n17360) );
  AND2_X1 U11794 ( .A1(n17273), .A2(n9775), .ZN(n9982) );
  NOR2_X1 U11795 ( .A1(n15866), .A2(n9986), .ZN(n9985) );
  INV_X1 U11796 ( .A(n12535), .ZN(n17418) );
  NOR2_X1 U11797 ( .A1(n17412), .A2(n18688), .ZN(n17420) );
  CLKBUF_X1 U11798 ( .A(n17530), .Z(n17522) );
  NOR2_X2 U11799 ( .A1(n17394), .A2(n17903), .ZN(n17814) );
  NOR2_X2 U11800 ( .A1(n16544), .A2(n16523), .ZN(n17892) );
  AOI22_X1 U11801 ( .A1(n12412), .A2(n12411), .B1(n12410), .B2(n12409), .ZN(
        n16398) );
  NAND2_X1 U11802 ( .A1(n9872), .A2(n16417), .ZN(n9871) );
  NAND2_X1 U11803 ( .A1(n17546), .A2(n9873), .ZN(n9872) );
  OAI21_X1 U11804 ( .B1(n16420), .B2(n18221), .A(n9868), .ZN(n9867) );
  AOI21_X1 U11805 ( .B1(n17977), .B2(n17544), .A(n17543), .ZN(n9868) );
  NAND2_X1 U11806 ( .A1(n16415), .A2(n18215), .ZN(n18221) );
  INV_X1 U11807 ( .A(n16879), .ZN(n18736) );
  NAND2_X1 U11808 ( .A1(n13306), .A2(n13307), .ZN(n10893) );
  AOI22_X1 U11809 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U11810 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11715) );
  OAI22_X1 U11811 ( .A1(n13654), .A2(n13656), .B1(n19351), .B2(n13655), .ZN(
        n13657) );
  INV_X1 U11812 ( .A(n9956), .ZN(n9955) );
  OAI21_X1 U11813 ( .B1(n13379), .B2(n19469), .A(n9793), .ZN(n13380) );
  NAND2_X1 U11814 ( .A1(n9794), .A2(n9940), .ZN(n9793) );
  OAI21_X1 U11815 ( .B1(n12927), .B2(n12924), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11470) );
  INV_X1 U11816 ( .A(n10630), .ZN(n10542) );
  OR2_X1 U11817 ( .A1(n10554), .A2(n10553), .ZN(n11220) );
  OR2_X1 U11818 ( .A1(n10527), .A2(n10526), .ZN(n11200) );
  OAI21_X1 U11819 ( .B1(n13171), .B2(P1_EBX_REG_1__SCAN_IN), .A(n14293), .ZN(
        n10017) );
  AND2_X1 U11820 ( .A1(n13581), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U11821 ( .A1(n10426), .A2(n13304), .ZN(n9968) );
  OR2_X1 U11822 ( .A1(n10514), .A2(n10513), .ZN(n11186) );
  INV_X1 U11823 ( .A(n13902), .ZN(n10157) );
  AOI22_X1 U11824 ( .A1(n12036), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n10149), .ZN(n11779) );
  AOI22_X1 U11825 ( .A1(n12036), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n10149), .ZN(n11774) );
  NAND2_X1 U11826 ( .A1(n11908), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n9855) );
  AOI22_X1 U11827 ( .A1(n10149), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U11828 ( .A1(n12036), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__2__SCAN_IN), .B2(n10149), .ZN(n11755) );
  AOI22_X1 U11829 ( .A1(n10149), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U11830 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11737) );
  OAI22_X1 U11831 ( .A1(n13654), .A2(n13873), .B1(n19351), .B2(n13872), .ZN(
        n13876) );
  NAND2_X1 U11832 ( .A1(n9795), .A2(n9716), .ZN(n13875) );
  NAND2_X1 U11833 ( .A1(n11908), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11467) );
  OR2_X1 U11834 ( .A1(n12129), .A2(n12128), .ZN(n12844) );
  NAND2_X1 U11835 ( .A1(n9785), .A2(n13382), .ZN(n13866) );
  NOR2_X1 U11836 ( .A1(n17401), .A2(n12357), .ZN(n12383) );
  NOR2_X1 U11837 ( .A1(n10207), .A2(n14306), .ZN(n10206) );
  NAND2_X1 U11838 ( .A1(n10208), .A2(n14317), .ZN(n10207) );
  INV_X1 U11839 ( .A(n14330), .ZN(n10208) );
  INV_X1 U11840 ( .A(n14076), .ZN(n10179) );
  INV_X1 U11841 ( .A(n10632), .ZN(n11052) );
  OR2_X1 U11842 ( .A1(n13179), .A2(n16039), .ZN(n11049) );
  AND2_X1 U11843 ( .A1(n10639), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10563) );
  INV_X1 U11844 ( .A(n14614), .ZN(n14628) );
  AND2_X1 U11845 ( .A1(n14881), .A2(n9725), .ZN(n10178) );
  NAND2_X1 U11846 ( .A1(n9975), .A2(n14888), .ZN(n10180) );
  INV_X1 U11847 ( .A(n14450), .ZN(n10023) );
  NOR2_X1 U11848 ( .A1(n14499), .A2(n10025), .ZN(n10024) );
  INV_X1 U11849 ( .A(n14463), .ZN(n10025) );
  OR2_X1 U11850 ( .A1(n10594), .A2(n20192), .ZN(n11167) );
  INV_X1 U11851 ( .A(n10409), .ZN(n10588) );
  OR2_X1 U11852 ( .A1(n10494), .A2(n10493), .ZN(n10495) );
  INV_X1 U11853 ( .A(n10495), .ZN(n11176) );
  NAND2_X1 U11854 ( .A1(n10463), .A2(n10462), .ZN(n10464) );
  NAND2_X1 U11855 ( .A1(n13076), .A2(n10265), .ZN(n13097) );
  NAND2_X1 U11856 ( .A1(n11133), .A2(n11225), .ZN(n11144) );
  AND2_X1 U11857 ( .A1(n11143), .A2(n11282), .ZN(n11145) );
  NAND2_X1 U11858 ( .A1(n11139), .A2(n11138), .ZN(n11147) );
  OR3_X1 U11859 ( .A1(n13129), .A2(n13128), .A3(n13127), .ZN(n13325) );
  INV_X1 U11860 ( .A(n20261), .ZN(n13510) );
  AOI21_X1 U11861 ( .B1(n11871), .B2(n11870), .A(n11869), .ZN(n11889) );
  INV_X1 U11862 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10161) );
  OR2_X1 U11863 ( .A1(n14148), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14197) );
  NAND2_X1 U11864 ( .A1(n14156), .A2(n14157), .ZN(n14159) );
  AND2_X1 U11865 ( .A1(n14117), .A2(n19138), .ZN(n14123) );
  AND2_X1 U11866 ( .A1(n14108), .A2(n12644), .ZN(n14117) );
  OR2_X1 U11867 ( .A1(n12091), .A2(n12090), .ZN(n12641) );
  NOR2_X1 U11868 ( .A1(n13429), .A2(n13428), .ZN(n13427) );
  INV_X1 U11869 ( .A(n15048), .ZN(n10232) );
  AND2_X1 U11870 ( .A1(n10235), .A2(n15048), .ZN(n10233) );
  INV_X1 U11871 ( .A(n15053), .ZN(n10235) );
  AOI22_X1 U11872 ( .A1(n10149), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11812) );
  NOR2_X1 U11873 ( .A1(n12671), .A2(n10128), .ZN(n10127) );
  INV_X1 U11874 ( .A(n15103), .ZN(n10128) );
  INV_X1 U11875 ( .A(n11542), .ZN(n11804) );
  AND2_X1 U11876 ( .A1(n13544), .A2(n13747), .ZN(n10144) );
  NAND2_X1 U11877 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10121) );
  NOR2_X1 U11878 ( .A1(n10117), .A2(n10116), .ZN(n10115) );
  INV_X1 U11879 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10116) );
  NAND2_X1 U11880 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10117) );
  INV_X1 U11881 ( .A(n13042), .ZN(n10092) );
  OR2_X1 U11882 ( .A1(n12143), .A2(n12142), .ZN(n12846) );
  NOR2_X1 U11883 ( .A1(n15193), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14224) );
  NAND2_X1 U11884 ( .A1(n10089), .A2(n15000), .ZN(n10088) );
  INV_X1 U11885 ( .A(n9773), .ZN(n10089) );
  AND2_X1 U11886 ( .A1(n14256), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9949) );
  AND2_X1 U11887 ( .A1(n12686), .A2(n15416), .ZN(n10147) );
  NAND2_X1 U11888 ( .A1(n9964), .A2(n15404), .ZN(n9963) );
  INV_X1 U11889 ( .A(n14194), .ZN(n9964) );
  AND2_X1 U11890 ( .A1(n15444), .A2(n12686), .ZN(n15415) );
  AND2_X1 U11891 ( .A1(n15442), .A2(n15441), .ZN(n15444) );
  AND2_X1 U11892 ( .A1(n10144), .A2(n13820), .ZN(n10143) );
  AND2_X1 U11893 ( .A1(n14252), .A2(n13426), .ZN(n14254) );
  INV_X1 U11894 ( .A(n15574), .ZN(n10225) );
  AND2_X1 U11895 ( .A1(n13901), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9861) );
  NAND2_X1 U11896 ( .A1(n13681), .A2(n15158), .ZN(n9923) );
  NOR2_X1 U11897 ( .A1(n11884), .A2(n11883), .ZN(n13354) );
  OR2_X1 U11898 ( .A1(n12114), .A2(n12113), .ZN(n12848) );
  NOR2_X1 U11899 ( .A1(n13153), .A2(n12133), .ZN(n12149) );
  NAND2_X1 U11900 ( .A1(n9796), .A2(n12047), .ZN(n12941) );
  NAND2_X1 U11901 ( .A1(n12056), .A2(n9700), .ZN(n9796) );
  INV_X1 U11902 ( .A(n19287), .ZN(n12922) );
  NAND2_X1 U11903 ( .A1(n12867), .A2(n13374), .ZN(n13383) );
  AND2_X1 U11904 ( .A1(n11395), .A2(n11376), .ZN(n9802) );
  AND2_X1 U11905 ( .A1(n11391), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9804) );
  NAND2_X1 U11906 ( .A1(n11390), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9806) );
  NAND2_X1 U11907 ( .A1(n11385), .A2(n11376), .ZN(n9805) );
  NAND3_X1 U11908 ( .A1(n19938), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19781), 
        .ZN(n19268) );
  AND2_X1 U11909 ( .A1(n10001), .A2(n10000), .ZN(n9999) );
  NAND2_X1 U11910 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10001) );
  NAND2_X1 U11911 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10000) );
  NAND2_X1 U11912 ( .A1(n18852), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12270) );
  NAND2_X1 U11913 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12272) );
  INV_X1 U11914 ( .A(n18675), .ZN(n9887) );
  INV_X1 U11915 ( .A(n12272), .ZN(n9886) );
  NAND2_X1 U11916 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12317) );
  OR2_X1 U11917 ( .A1(n12296), .A2(n17063), .ZN(n10254) );
  INV_X1 U11918 ( .A(n10007), .ZN(n10006) );
  OAI21_X1 U11919 ( .B1(n10010), .B2(n18843), .A(n12406), .ZN(n10007) );
  NOR2_X1 U11920 ( .A1(n17631), .A2(n18005), .ZN(n17639) );
  OAI21_X1 U11921 ( .B1(n17791), .B2(n12394), .A(n10010), .ZN(n12398) );
  NAND2_X1 U11922 ( .A1(n17855), .A2(n12378), .ZN(n12381) );
  XNOR2_X1 U11923 ( .A(n12376), .B(n17405), .ZN(n12377) );
  INV_X1 U11924 ( .A(n9899), .ZN(n18666) );
  OAI21_X1 U11925 ( .B1(n12525), .B2(n12524), .A(n12523), .ZN(n16517) );
  NAND2_X1 U11926 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9890) );
  NAND2_X1 U11927 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n9895) );
  NAND2_X1 U11928 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9891) );
  NAND2_X1 U11929 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n9898) );
  OAI211_X1 U11930 ( .C1(n10251), .C2(n17033), .A(n12458), .B(n12457), .ZN(
        n12514) );
  NOR2_X1 U11931 ( .A1(n10770), .A2(n14467), .ZN(n10756) );
  OR2_X1 U11932 ( .A1(n13583), .A2(n13563), .ZN(n13796) );
  INV_X1 U11933 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20074) );
  AND2_X1 U11934 ( .A1(n13796), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13566) );
  NAND2_X1 U11935 ( .A1(n14434), .A2(n14420), .ZN(n14422) );
  AND2_X1 U11936 ( .A1(n14066), .A2(n14293), .ZN(n14058) );
  AND2_X1 U11937 ( .A1(n20728), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11077) );
  NAND2_X1 U11938 ( .A1(n10206), .A2(n11267), .ZN(n10205) );
  AOI21_X1 U11939 ( .B1(n13120), .B2(n15820), .A(n12966), .ZN(n20104) );
  AND2_X2 U11940 ( .A1(n20192), .A2(n13581), .ZN(n13034) );
  AND2_X1 U11941 ( .A1(n11027), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11028) );
  NAND2_X1 U11942 ( .A1(n10985), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11026) );
  NAND2_X1 U11943 ( .A1(n14628), .A2(n14616), .ZN(n14642) );
  OR2_X1 U11944 ( .A1(n10947), .A2(n10946), .ZN(n10984) );
  NAND2_X1 U11945 ( .A1(n9747), .A2(n9920), .ZN(n9919) );
  INV_X1 U11946 ( .A(n9921), .ZN(n9920) );
  AND2_X1 U11947 ( .A1(n10884), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10885) );
  NAND2_X1 U11948 ( .A1(n10845), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10883) );
  NAND2_X1 U11949 ( .A1(n11250), .A2(n10177), .ZN(n14688) );
  NOR2_X1 U11950 ( .A1(n10804), .A2(n14714), .ZN(n10805) );
  NAND2_X1 U11951 ( .A1(n10756), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10804) );
  AND2_X1 U11952 ( .A1(n10803), .A2(n10196), .ZN(n10195) );
  AND2_X1 U11953 ( .A1(n10738), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10786) );
  AND2_X1 U11954 ( .A1(n10734), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10738) );
  NOR2_X1 U11955 ( .A1(n10706), .A2(n15912), .ZN(n10710) );
  NAND2_X1 U11956 ( .A1(n9674), .A2(n10695), .ZN(n13990) );
  NAND2_X1 U11957 ( .A1(n10680), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10706) );
  NOR2_X1 U11958 ( .A1(n10664), .A2(n10663), .ZN(n10680) );
  INV_X1 U11959 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10663) );
  NAND2_X1 U11960 ( .A1(n10658), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10664) );
  AND2_X1 U11961 ( .A1(n10563), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10658) );
  NAND2_X1 U11962 ( .A1(n11226), .A2(n10795), .ZN(n10570) );
  AND2_X1 U11963 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n10631), .ZN(
        n10639) );
  INV_X1 U11964 ( .A(n13591), .ZN(n9916) );
  INV_X1 U11965 ( .A(n13496), .ZN(n9917) );
  NOR2_X1 U11966 ( .A1(n10621), .A2(n20074), .ZN(n10631) );
  NOR2_X1 U11967 ( .A1(n13588), .A2(n10562), .ZN(n10614) );
  INV_X1 U11968 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10562) );
  INV_X1 U11969 ( .A(n13243), .ZN(n10607) );
  NAND2_X1 U11970 ( .A1(n10188), .A2(n9738), .ZN(n10181) );
  NAND2_X1 U11971 ( .A1(n11268), .A2(n10183), .ZN(n10182) );
  NAND2_X1 U11972 ( .A1(n14358), .A2(n14064), .ZN(n14336) );
  INV_X1 U11973 ( .A(n11250), .ZN(n11251) );
  NAND2_X1 U11974 ( .A1(n11250), .A2(n14716), .ZN(n14715) );
  NAND2_X1 U11975 ( .A1(n15883), .A2(n10024), .ZN(n14502) );
  INV_X1 U11976 ( .A(n14722), .ZN(n14883) );
  NAND2_X1 U11977 ( .A1(n15883), .A2(n14463), .ZN(n14500) );
  INV_X1 U11978 ( .A(n13759), .ZN(n10026) );
  NAND2_X1 U11979 ( .A1(n10027), .A2(n9701), .ZN(n16027) );
  AND2_X1 U11980 ( .A1(n13529), .A2(n13528), .ZN(n13530) );
  NOR2_X1 U11981 ( .A1(n13447), .A2(n10029), .ZN(n16026) );
  NOR2_X1 U11982 ( .A1(n13447), .A2(n13446), .ZN(n13531) );
  INV_X1 U11983 ( .A(n13171), .ZN(n13291) );
  OAI21_X1 U11984 ( .B1(n11130), .B2(n20189), .A(n10453), .ZN(n10601) );
  OR2_X1 U11985 ( .A1(n10457), .A2(n10456), .ZN(n10458) );
  OR2_X1 U11986 ( .A1(n20408), .A2(n20623), .ZN(n20383) );
  INV_X1 U11987 ( .A(n9908), .ZN(n20213) );
  NAND2_X1 U11988 ( .A1(n9656), .A2(n20261), .ZN(n20623) );
  AND3_X2 U11989 ( .A1(n10358), .A2(n10357), .A3(n10356), .ZN(n13522) );
  NAND2_X1 U11990 ( .A1(n15960), .A2(n13519), .ZN(n20221) );
  AND2_X1 U11991 ( .A1(n15823), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15822) );
  INV_X1 U11992 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15823) );
  OR2_X1 U11993 ( .A1(n14227), .A2(n14226), .ZN(n14950) );
  NAND2_X1 U11994 ( .A1(n12650), .A2(n14196), .ZN(n14202) );
  NAND2_X1 U11995 ( .A1(n14156), .A2(n10151), .ZN(n14146) );
  NAND2_X1 U11996 ( .A1(n16160), .A2(n10107), .ZN(n10106) );
  NAND2_X1 U11997 ( .A1(n10148), .A2(n9741), .ZN(n14176) );
  INV_X1 U11998 ( .A(n10148), .ZN(n14142) );
  NAND2_X1 U11999 ( .A1(n14133), .A2(n14220), .ZN(n14126) );
  AND2_X1 U12000 ( .A1(n13676), .A2(n10156), .ZN(n14108) );
  AND2_X1 U12001 ( .A1(n9679), .A2(n13598), .ZN(n10156) );
  AND2_X1 U12002 ( .A1(n13427), .A2(n13638), .ZN(n13676) );
  NAND2_X1 U12003 ( .A1(n13676), .A2(n13675), .ZN(n13903) );
  AND3_X1 U12004 ( .A1(n11980), .A2(n11979), .A3(n11978), .ZN(n15083) );
  OR2_X1 U12005 ( .A1(n11599), .A2(n11598), .ZN(n12220) );
  AND2_X1 U12006 ( .A1(n13459), .A2(n9762), .ZN(n10236) );
  OR2_X1 U12007 ( .A1(n15125), .A2(n15128), .ZN(n15126) );
  NAND2_X1 U12008 ( .A1(n10240), .A2(n10239), .ZN(n10238) );
  INV_X1 U12009 ( .A(n16102), .ZN(n10239) );
  OR2_X1 U12010 ( .A1(n11652), .A2(n11651), .ZN(n13839) );
  INV_X1 U12011 ( .A(n16264), .ZN(n10138) );
  AOI21_X1 U12012 ( .B1(n10130), .B2(n10134), .A(n12168), .ZN(n12994) );
  NOR2_X1 U12013 ( .A1(n10133), .A2(n10132), .ZN(n10130) );
  NAND2_X1 U12014 ( .A1(n13456), .A2(n13689), .ZN(n10132) );
  AND2_X1 U12015 ( .A1(n12170), .A2(n12169), .ZN(n12993) );
  INV_X1 U12016 ( .A(n12075), .ZN(n19269) );
  AND2_X1 U12017 ( .A1(n9684), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10122) );
  CLKBUF_X1 U12018 ( .A(n14952), .Z(n14953) );
  NAND2_X1 U12019 ( .A1(n12597), .A2(n10123), .ZN(n14955) );
  CLKBUF_X1 U12020 ( .A(n12599), .Z(n12601) );
  NOR3_X1 U12021 ( .A1(n15412), .A2(n15411), .A3(n9773), .ZN(n15011) );
  NAND2_X1 U12022 ( .A1(n15247), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15477) );
  CLKBUF_X1 U12023 ( .A(n12611), .Z(n12626) );
  NOR2_X1 U12024 ( .A1(n12612), .A2(n10117), .ZN(n12610) );
  CLKBUF_X1 U12025 ( .A(n12612), .Z(n12622) );
  AND3_X1 U12026 ( .A1(n11946), .A2(n11945), .A3(n11944), .ZN(n13257) );
  NAND2_X1 U12027 ( .A1(n10092), .A2(n10093), .ZN(n13609) );
  NOR2_X1 U12028 ( .A1(n15564), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10078) );
  NAND2_X1 U12029 ( .A1(n16223), .A2(n16222), .ZN(n16221) );
  AND3_X1 U12030 ( .A1(n11938), .A2(n11937), .A3(n11936), .ZN(n13043) );
  NAND2_X1 U12031 ( .A1(n13017), .A2(n13018), .ZN(n13042) );
  AND3_X1 U12032 ( .A1(n11930), .A2(n11929), .A3(n11928), .ZN(n12962) );
  NOR2_X1 U12033 ( .A1(n19105), .A2(n12962), .ZN(n13017) );
  OAI21_X1 U12034 ( .B1(n11919), .B2(n10086), .A(n10085), .ZN(n19104) );
  NAND2_X1 U12035 ( .A1(n11524), .A2(n11921), .ZN(n10086) );
  AND2_X1 U12036 ( .A1(n12714), .A2(n12713), .ZN(n12919) );
  INV_X1 U12037 ( .A(n14957), .ZN(n10095) );
  NAND2_X1 U12038 ( .A1(n15152), .A2(n10211), .ZN(n10210) );
  NOR2_X1 U12039 ( .A1(n15174), .A2(n10212), .ZN(n10211) );
  INV_X1 U12040 ( .A(n15151), .ZN(n10212) );
  NAND2_X1 U12041 ( .A1(n15152), .A2(n15151), .ZN(n15171) );
  INV_X1 U12042 ( .A(n10098), .ZN(n10096) );
  AND2_X1 U12043 ( .A1(n10218), .A2(n15223), .ZN(n9966) );
  AND3_X1 U12044 ( .A1(n12011), .A2(n12010), .A3(n12009), .ZN(n15057) );
  NOR2_X1 U12045 ( .A1(n9672), .A2(n15057), .ZN(n15058) );
  NAND2_X1 U12046 ( .A1(n15444), .A2(n10145), .ZN(n15112) );
  AND2_X1 U12047 ( .A1(n9761), .A2(n10146), .ZN(n10145) );
  INV_X1 U12048 ( .A(n15003), .ZN(n10146) );
  AND2_X1 U12049 ( .A1(n15548), .A2(n9949), .ZN(n15379) );
  AND2_X1 U12050 ( .A1(n15444), .A2(n10147), .ZN(n15418) );
  OR2_X1 U12051 ( .A1(n9965), .A2(n9959), .ZN(n9958) );
  AND2_X1 U12052 ( .A1(n10222), .A2(n15404), .ZN(n9965) );
  INV_X1 U12053 ( .A(n9963), .ZN(n9959) );
  NAND2_X1 U12054 ( .A1(n15548), .A2(n14256), .ZN(n15389) );
  OR2_X1 U12055 ( .A1(n12683), .A2(n12685), .ZN(n15412) );
  NOR2_X1 U12056 ( .A1(n15412), .A2(n15411), .ZN(n15413) );
  NAND2_X1 U12057 ( .A1(n9935), .A2(n9936), .ZN(n15272) );
  NAND2_X1 U12058 ( .A1(n15282), .A2(n9937), .ZN(n9935) );
  AND2_X1 U12059 ( .A1(n15489), .A2(n15143), .ZN(n15442) );
  AND3_X1 U12060 ( .A1(n11976), .A2(n11975), .A3(n11974), .ZN(n15483) );
  NAND2_X1 U12061 ( .A1(n15764), .A2(n10102), .ZN(n15486) );
  AND2_X1 U12062 ( .A1(n12237), .A2(n12236), .ZN(n15488) );
  NOR2_X1 U12063 ( .A1(n15487), .A2(n15488), .ZN(n15489) );
  NAND2_X1 U12064 ( .A1(n15764), .A2(n13841), .ZN(n15484) );
  AND2_X1 U12065 ( .A1(n15766), .A2(n13628), .ZN(n15764) );
  OR2_X1 U12066 ( .A1(n18979), .A2(n14168), .ZN(n15281) );
  NAND2_X1 U12067 ( .A1(n15548), .A2(n15285), .ZN(n16181) );
  NAND2_X1 U12068 ( .A1(n9749), .A2(n9928), .ZN(n9927) );
  AND3_X1 U12069 ( .A1(n11958), .A2(n11957), .A3(n11956), .ZN(n13474) );
  NAND2_X1 U12070 ( .A1(n10139), .A2(n10137), .ZN(n15036) );
  AND2_X1 U12071 ( .A1(n9685), .A2(n13298), .ZN(n10137) );
  NAND2_X1 U12072 ( .A1(n10083), .A2(n10082), .ZN(n15035) );
  INV_X1 U12073 ( .A(n15032), .ZN(n10082) );
  INV_X1 U12074 ( .A(n15033), .ZN(n10083) );
  NAND2_X1 U12075 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9865) );
  NOR2_X1 U12076 ( .A1(n13042), .A2(n10090), .ZN(n16209) );
  NAND2_X1 U12077 ( .A1(n9676), .A2(n16207), .ZN(n10090) );
  NAND2_X1 U12078 ( .A1(n16209), .A2(n13465), .ZN(n15033) );
  NAND2_X1 U12079 ( .A1(n10139), .A2(n10140), .ZN(n16265) );
  NOR2_X1 U12080 ( .A1(n13605), .A2(n13606), .ZN(n15557) );
  OAI22_X1 U12081 ( .A1(n12994), .A2(n12993), .B1(n15158), .B2(n12232), .ZN(
        n13033) );
  NAND2_X1 U12082 ( .A1(n13033), .A2(n13032), .ZN(n13605) );
  INV_X1 U12083 ( .A(n10133), .ZN(n10135) );
  NAND2_X1 U12084 ( .A1(n10071), .A2(n15158), .ZN(n9858) );
  INV_X1 U12085 ( .A(n11505), .ZN(n13366) );
  OAI21_X1 U12086 ( .B1(n12257), .B2(n18922), .A(n12102), .ZN(n12887) );
  AND2_X1 U12087 ( .A1(n19986), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11528) );
  NAND2_X1 U12088 ( .A1(n12909), .A2(n11896), .ZN(n16327) );
  AND2_X1 U12089 ( .A1(n19566), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19500) );
  NOR2_X1 U12090 ( .A1(n11344), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9820) );
  NOR2_X2 U12091 ( .A1(n19267), .A2(n19268), .ZN(n19314) );
  NOR2_X1 U12092 ( .A1(n19566), .A2(n19536), .ZN(n19738) );
  INV_X1 U12093 ( .A(n19511), .ZN(n19777) );
  NAND2_X1 U12094 ( .A1(n12705), .A2(n12062), .ZN(n16322) );
  XNOR2_X1 U12095 ( .A(n18884), .B(n18237), .ZN(n18887) );
  INV_X1 U12096 ( .A(n16517), .ZN(n18711) );
  AND2_X1 U12097 ( .A1(n10046), .A2(n10048), .ZN(n16576) );
  AOI21_X1 U12098 ( .B1(n10050), .B2(n16860), .A(n16860), .ZN(n10048) );
  OR2_X1 U12099 ( .A1(n16594), .A2(n10049), .ZN(n10046) );
  INV_X1 U12100 ( .A(n10050), .ZN(n10049) );
  AND2_X1 U12101 ( .A1(n16647), .A2(n10056), .ZN(n16635) );
  NOR2_X1 U12102 ( .A1(n17612), .A2(n16635), .ZN(n16634) );
  OR2_X1 U12103 ( .A1(n16649), .A2(n17628), .ZN(n16647) );
  OR2_X1 U12104 ( .A1(n16673), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n16676) );
  NOR2_X1 U12105 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16721), .ZN(n16710) );
  INV_X1 U12106 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9988) );
  NOR2_X1 U12107 ( .A1(n17470), .A2(n9992), .ZN(n9991) );
  OAI211_X1 U12108 ( .C1(n10251), .C2(n17003), .A(n12489), .B(n12488), .ZN(
        n17278) );
  CLKBUF_X1 U12109 ( .A(n12283), .Z(n16984) );
  CLKBUF_X1 U12110 ( .A(n15623), .Z(n17187) );
  INV_X1 U12111 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17189) );
  OR3_X2 U12112 ( .A1(n12331), .A2(n12332), .A3(n10013), .ZN(n12536) );
  AOI211_X1 U12113 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n12446), .B(n12445), .ZN(n12447) );
  NOR3_X1 U12114 ( .A1(n17427), .A2(n18882), .A3(n17466), .ZN(n17446) );
  NAND2_X1 U12115 ( .A1(n16562), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16561) );
  NOR2_X1 U12116 ( .A1(n17567), .A2(n17566), .ZN(n17536) );
  NOR2_X1 U12117 ( .A1(n9681), .A2(n9748), .ZN(n10067) );
  NOR2_X1 U12118 ( .A1(n17681), .A2(n9681), .ZN(n17622) );
  AND2_X1 U12119 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n9756), .ZN(
        n10068) );
  NOR2_X1 U12120 ( .A1(n17681), .A2(n17680), .ZN(n17669) );
  INV_X1 U12121 ( .A(n17702), .ZN(n17687) );
  INV_X1 U12122 ( .A(n17754), .ZN(n17710) );
  NOR2_X1 U12123 ( .A1(n17753), .A2(n16556), .ZN(n17711) );
  NAND2_X1 U12124 ( .A1(n12564), .A2(n17803), .ZN(n16404) );
  NAND2_X1 U12125 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17807) );
  AND2_X1 U12126 ( .A1(n10043), .A2(n10042), .ZN(n17839) );
  NOR2_X1 U12127 ( .A1(n10045), .A2(n17846), .ZN(n10043) );
  NOR2_X1 U12128 ( .A1(n17886), .A2(n17805), .ZN(n17838) );
  NOR2_X1 U12129 ( .A1(n18717), .A2(n18732), .ZN(n12568) );
  NAND2_X1 U12130 ( .A1(n17552), .A2(n16416), .ZN(n15740) );
  NOR2_X1 U12131 ( .A1(n9875), .A2(n9874), .ZN(n9873) );
  NAND2_X1 U12132 ( .A1(n16415), .A2(n16414), .ZN(n9874) );
  INV_X1 U12133 ( .A(n16413), .ZN(n9875) );
  NOR2_X1 U12134 ( .A1(n10010), .A2(n9777), .ZN(n10032) );
  NOR2_X1 U12135 ( .A1(n16414), .A2(n18713), .ZN(n17940) );
  INV_X1 U12136 ( .A(n17648), .ZN(n17629) );
  INV_X1 U12137 ( .A(n16404), .ZN(n18090) );
  INV_X1 U12138 ( .A(n17777), .ZN(n17790) );
  NAND2_X1 U12139 ( .A1(n12558), .A2(n17831), .ZN(n17825) );
  NAND2_X1 U12140 ( .A1(n17819), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17818) );
  XNOR2_X1 U12141 ( .A(n12381), .B(n12380), .ZN(n17849) );
  INV_X1 U12142 ( .A(n12379), .ZN(n12380) );
  AND2_X1 U12143 ( .A1(n18167), .A2(n18884), .ZN(n18706) );
  NAND2_X1 U12144 ( .A1(n18887), .A2(n15714), .ZN(n18190) );
  XNOR2_X1 U12145 ( .A(n12358), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17879) );
  NAND2_X1 U12146 ( .A1(n17898), .A2(n17890), .ZN(n17889) );
  AOI21_X1 U12147 ( .B1(n12503), .B2(n12502), .A(n16539), .ZN(n12516) );
  NOR2_X1 U12148 ( .A1(n15728), .A2(n15719), .ZN(n16415) );
  OAI211_X1 U12149 ( .C1(n17133), .C2(n17025), .A(n12500), .B(n12499), .ZN(
        n15735) );
  INV_X1 U12150 ( .A(n15725), .ZN(n18678) );
  INV_X1 U12151 ( .A(n18190), .ZN(n18707) );
  NAND2_X1 U12152 ( .A1(n12516), .A2(n9994), .ZN(n15725) );
  INV_X1 U12153 ( .A(n15715), .ZN(n9994) );
  NAND3_X1 U12154 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15726) );
  INV_X1 U12155 ( .A(n17428), .ZN(n18237) );
  INV_X1 U12156 ( .A(n12528), .ZN(n18244) );
  AOI21_X1 U12157 ( .B1(n18706), .B2(n18708), .A(n9902), .ZN(n18717) );
  AND2_X1 U12158 ( .A1(n16415), .A2(n18712), .ZN(n9902) );
  NOR2_X1 U12159 ( .A1(n13581), .A2(n16039), .ZN(n12898) );
  AND2_X1 U12160 ( .A1(n13583), .A2(n13571), .ZN(n20077) );
  AND2_X1 U12161 ( .A1(n13583), .A2(n13577), .ZN(n20053) );
  INV_X1 U12162 ( .A(n20077), .ZN(n20038) );
  NOR2_X2 U12163 ( .A1(n13568), .A2(n13567), .ZN(n20049) );
  INV_X1 U12164 ( .A(n13566), .ZN(n13567) );
  INV_X1 U12165 ( .A(n20049), .ZN(n20087) );
  INV_X1 U12166 ( .A(n20053), .ZN(n20084) );
  INV_X1 U12167 ( .A(n14523), .ZN(n20098) );
  INV_X1 U12168 ( .A(n20103), .ZN(n14485) );
  AND2_X1 U12169 ( .A1(n14603), .A2(n13165), .ZN(n14563) );
  OR2_X1 U12170 ( .A1(n11299), .A2(n13519), .ZN(n14573) );
  INV_X1 U12171 ( .A(n14573), .ZN(n14588) );
  OR2_X1 U12172 ( .A1(n14507), .A2(n14516), .ZN(n14752) );
  OR2_X1 U12173 ( .A1(n13129), .A2(n11286), .ZN(n11287) );
  OR2_X1 U12174 ( .A1(n14569), .A2(n13165), .ZN(n14602) );
  INV_X2 U12175 ( .A(n14563), .ZN(n14605) );
  NOR2_X1 U12176 ( .A1(n20104), .A2(n20130), .ZN(n15855) );
  BUF_X1 U12177 ( .A(n15855), .Z(n20129) );
  BUF_X1 U12178 ( .A(n20120), .Z(n20130) );
  NAND2_X1 U12179 ( .A1(n14406), .A2(n14393), .ZN(n14379) );
  NOR2_X1 U12180 ( .A1(n14419), .A2(n14418), .ZN(n14405) );
  AND2_X1 U12181 ( .A1(n14595), .A2(n14509), .ZN(n15896) );
  AND3_X1 U12182 ( .A1(n14943), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n16039), 
        .ZN(n15960) );
  NAND2_X1 U12183 ( .A1(n11270), .A2(n9971), .ZN(n10190) );
  NAND2_X1 U12184 ( .A1(n11253), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14630) );
  NAND2_X1 U12185 ( .A1(n9978), .A2(n9979), .ZN(n13973) );
  NAND2_X1 U12186 ( .A1(n11229), .A2(n15956), .ZN(n13847) );
  INV_X1 U12187 ( .A(n20164), .ZN(n16033) );
  NOR2_X1 U12188 ( .A1(n14012), .A2(n14912), .ZN(n15998) );
  OR2_X1 U12189 ( .A1(n13091), .A2(n15795), .ZN(n14890) );
  OR2_X1 U12190 ( .A1(n20812), .A2(n13507), .ZN(n20819) );
  OAI21_X1 U12191 ( .B1(n13331), .B2(n16045), .A(n20330), .ZN(n20823) );
  OR2_X1 U12192 ( .A1(n13126), .A2(n13115), .ZN(n20801) );
  NOR2_X1 U12193 ( .A1(n10386), .A2(n10412), .ZN(n9845) );
  INV_X1 U12194 ( .A(n10429), .ZN(n9846) );
  OR2_X1 U12195 ( .A1(n20302), .A2(n20548), .ZN(n20233) );
  INV_X1 U12196 ( .A(n20262), .ZN(n20285) );
  OAI21_X1 U12197 ( .B1(n20269), .B2(n20268), .A(n20267), .ZN(n20286) );
  INV_X1 U12198 ( .A(n20301), .ZN(n20319) );
  OAI21_X1 U12199 ( .B1(n20346), .B2(n20331), .A(n20631), .ZN(n20349) );
  INV_X1 U12200 ( .A(n20383), .ZN(n20426) );
  OAI211_X1 U12201 ( .C1(n20453), .C2(n13115), .A(n20491), .B(n20438), .ZN(
        n20456) );
  NOR2_X2 U12202 ( .A1(n20819), .A2(n20594), .ZN(n20511) );
  INV_X1 U12203 ( .A(n20621), .ZN(n20581) );
  OAI211_X1 U12204 ( .C1(n20654), .C2(n20632), .A(n20631), .B(n20630), .ZN(
        n20657) );
  INV_X1 U12205 ( .A(n20724), .ZN(n20710) );
  OR2_X1 U12206 ( .A1(n20624), .A2(n20516), .ZN(n20724) );
  INV_X2 U12207 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20728) );
  NAND2_X1 U12208 ( .A1(n14227), .A2(n14206), .ZN(n10164) );
  NAND2_X1 U12209 ( .A1(n10167), .A2(n14206), .ZN(n10165) );
  OR2_X1 U12210 ( .A1(n14240), .A2(n14967), .ZN(n16070) );
  NOR2_X1 U12211 ( .A1(n19021), .A2(n16090), .ZN(n16072) );
  NAND2_X1 U12212 ( .A1(n12650), .A2(n10162), .ZN(n14207) );
  NAND2_X1 U12213 ( .A1(n18933), .A2(n10112), .ZN(n10110) );
  NOR2_X1 U12214 ( .A1(n18933), .A2(n19021), .ZN(n12679) );
  NOR2_X1 U12215 ( .A1(n12679), .A2(n15244), .ZN(n12678) );
  NAND2_X1 U12216 ( .A1(n10105), .A2(n10104), .ZN(n18945) );
  NAND2_X1 U12217 ( .A1(n19021), .A2(n10107), .ZN(n10104) );
  INV_X1 U12218 ( .A(n10108), .ZN(n18956) );
  INV_X1 U12219 ( .A(n19093), .ZN(n19095) );
  NAND2_X1 U12220 ( .A1(n14973), .A2(n12663), .ZN(n19096) );
  INV_X1 U12221 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12621) );
  XNOR2_X1 U12222 ( .A(n11920), .B(n11917), .ZN(n9807) );
  AND2_X1 U12223 ( .A1(n18906), .A2(n12668), .ZN(n19076) );
  XNOR2_X1 U12224 ( .A(n14958), .B(n14957), .ZN(n15177) );
  NOR2_X1 U12225 ( .A1(n15054), .A2(n15053), .ZN(n15052) );
  NAND2_X1 U12226 ( .A1(n15047), .A2(n11809), .ZN(n15054) );
  OR2_X1 U12227 ( .A1(n11620), .A2(n11619), .ZN(n19121) );
  NOR2_X1 U12228 ( .A1(n19132), .A2(n19133), .ZN(n11577) );
  NOR2_X1 U12229 ( .A1(n11588), .A2(n11587), .ZN(n13470) );
  CLKBUF_X1 U12230 ( .A(n13468), .Z(n13469) );
  NAND3_X1 U12231 ( .A1(n11527), .A2(n9799), .A3(n9797), .ZN(n12990) );
  OAI21_X1 U12232 ( .B1(n11526), .B2(n11525), .A(n9800), .ZN(n9799) );
  NAND2_X1 U12233 ( .A1(n12989), .A2(n12988), .ZN(n19566) );
  OR2_X1 U12234 ( .A1(n12986), .A2(n12987), .ZN(n12989) );
  INV_X1 U12235 ( .A(n19953), .ZN(n19275) );
  XNOR2_X1 U12236 ( .A(n14972), .B(n14971), .ZN(n19149) );
  AND2_X1 U12237 ( .A1(n14987), .A2(n12672), .ZN(n15343) );
  OR2_X1 U12238 ( .A1(n19169), .A2(n12888), .ZN(n13822) );
  INV_X1 U12239 ( .A(n16119), .ZN(n19150) );
  INV_X1 U12240 ( .A(n16120), .ZN(n19173) );
  BUF_X1 U12241 ( .A(n19198), .Z(n19211) );
  NOR2_X1 U12242 ( .A1(n12824), .A2(n12716), .ZN(n12731) );
  INV_X1 U12243 ( .A(n12784), .ZN(n12878) );
  INV_X1 U12244 ( .A(n16165), .ZN(n15759) );
  AND2_X1 U12245 ( .A1(n13630), .A2(n13629), .ZN(n18990) );
  INV_X1 U12246 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15296) );
  INV_X1 U12247 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16235) );
  INV_X1 U12248 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19068) );
  INV_X1 U12249 ( .A(n10072), .ZN(n19219) );
  INV_X1 U12250 ( .A(n15590), .ZN(n13374) );
  INV_X1 U12251 ( .A(n16239), .ZN(n19223) );
  OR2_X1 U12252 ( .A1(n15391), .A2(n14205), .ZN(n15378) );
  NAND2_X1 U12253 ( .A1(n9962), .A2(n14194), .ZN(n15406) );
  INV_X1 U12254 ( .A(n9938), .ZN(n15276) );
  OAI21_X1 U12255 ( .B1(n9939), .B2(n9933), .A(n9931), .ZN(n9938) );
  AOI21_X1 U12256 ( .B1(n16165), .B2(n10081), .A(n10079), .ZN(n15786) );
  NAND2_X1 U12257 ( .A1(n16292), .A2(n15760), .ZN(n10081) );
  INV_X1 U12258 ( .A(n10080), .ZN(n10079) );
  NAND2_X1 U12259 ( .A1(n14138), .A2(n14137), .ZN(n15295) );
  NAND2_X1 U12260 ( .A1(n14104), .A2(n14103), .ZN(n15573) );
  NAND2_X1 U12261 ( .A1(n15565), .A2(n15564), .ZN(n15563) );
  INV_X1 U12262 ( .A(n14251), .ZN(n15565) );
  NAND2_X1 U12263 ( .A1(n9860), .A2(n9859), .ZN(n14250) );
  AND3_X1 U12264 ( .A1(n10074), .A2(n10073), .A3(n10072), .ZN(n13892) );
  INV_X1 U12265 ( .A(n10076), .ZN(n16294) );
  NOR2_X1 U12266 ( .A1(n10071), .A2(n9760), .ZN(n16293) );
  INV_X1 U12267 ( .A(n16290), .ZN(n19262) );
  OR2_X1 U12268 ( .A1(n19245), .A2(n19253), .ZN(n15579) );
  AND2_X1 U12269 ( .A1(n12954), .A2(n19971), .ZN(n19255) );
  INV_X1 U12270 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19966) );
  OR2_X1 U12271 ( .A1(n15594), .A2(n12840), .ZN(n19961) );
  INV_X1 U12272 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15593) );
  XNOR2_X1 U12273 ( .A(n12904), .B(n12903), .ZN(n19953) );
  NAND2_X1 U12274 ( .A1(n16327), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15860) );
  XNOR2_X1 U12275 ( .A(n12958), .B(n12959), .ZN(n19412) );
  NOR2_X1 U12276 ( .A1(n19580), .A2(n19512), .ZN(n19367) );
  OAI21_X1 U12277 ( .B1(n19417), .B2(n19433), .A(n19416), .ZN(n19435) );
  NOR2_X1 U12278 ( .A1(n19512), .A2(n19706), .ZN(n19486) );
  OAI21_X1 U12279 ( .B1(n19612), .B2(n19628), .A(n19781), .ZN(n19631) );
  NOR2_X2 U12280 ( .A1(n19635), .A2(n19580), .ZN(n19630) );
  INV_X1 U12281 ( .A(n19663), .ZN(n19666) );
  NOR2_X2 U12282 ( .A1(n19635), .A2(n19634), .ZN(n19699) );
  INV_X1 U12283 ( .A(n19830), .ZN(n19761) );
  OAI21_X1 U12284 ( .B1(n13654), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n9924), 
        .ZN(n19741) );
  NOR2_X1 U12285 ( .A1(n19769), .A2(n19938), .ZN(n9924) );
  OAI21_X1 U12286 ( .B1(n19746), .B2(n19745), .A(n19744), .ZN(n19771) );
  AND2_X1 U12287 ( .A1(n19713), .A2(n19712), .ZN(n19770) );
  INV_X1 U12288 ( .A(n19749), .ZN(n19794) );
  INV_X1 U12289 ( .A(n19688), .ZN(n19806) );
  INV_X1 U12290 ( .A(n19724), .ZN(n19813) );
  AND2_X1 U12291 ( .A1(n19291), .A2(n19301), .ZN(n19811) );
  AND2_X1 U12292 ( .A1(n15154), .A2(n19301), .ZN(n19823) );
  INV_X1 U12293 ( .A(n19768), .ZN(n19834) );
  INV_X1 U12294 ( .A(n19829), .ZN(n19841) );
  AND2_X1 U12295 ( .A1(n19738), .A2(n19777), .ZN(n19843) );
  INV_X1 U12296 ( .A(n19605), .ZN(n19842) );
  INV_X1 U12297 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19979) );
  INV_X1 U12298 ( .A(n18887), .ZN(n18898) );
  NOR2_X1 U12299 ( .A1(n16577), .A2(n16576), .ZN(n16575) );
  AND2_X1 U12300 ( .A1(n10051), .A2(n10056), .ZN(n16587) );
  NAND2_X1 U12301 ( .A1(n16594), .A2(n10056), .ZN(n10047) );
  NAND2_X1 U12302 ( .A1(n10054), .A2(n10055), .ZN(n16605) );
  AND2_X1 U12303 ( .A1(n16627), .A2(n10056), .ZN(n16616) );
  NOR2_X1 U12304 ( .A1(n18725), .A2(n16542), .ZN(n16864) );
  AOI21_X1 U12305 ( .B1(n10056), .B2(n17659), .A(n16715), .ZN(n16698) );
  NAND2_X1 U12306 ( .A1(n10062), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10057) );
  NAND2_X1 U12307 ( .A1(n16562), .A2(n10059), .ZN(n10058) );
  OR2_X1 U12308 ( .A1(n16562), .A2(n12574), .ZN(n10060) );
  NOR2_X1 U12309 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16773), .ZN(n16756) );
  NOR2_X1 U12310 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16820), .ZN(n16803) );
  NOR2_X1 U12311 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16844), .ZN(n16825) );
  INV_X1 U12312 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16873) );
  INV_X1 U12313 ( .A(n16864), .ZN(n16892) );
  NOR4_X2 U12314 ( .A1(n18210), .A2(n18899), .A3(n18736), .A4(n16541), .ZN(
        n16899) );
  NOR2_X1 U12315 ( .A1(n16641), .A2(n16976), .ZN(n16982) );
  INV_X1 U12316 ( .A(n12435), .ZN(n9995) );
  INV_X1 U12317 ( .A(n12438), .ZN(n10003) );
  INV_X1 U12318 ( .A(n12436), .ZN(n9996) );
  INV_X1 U12319 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17235) );
  NOR4_X2 U12320 ( .A1(n18884), .A2(n18237), .A3(n15863), .A4(n18732), .ZN(
        n17269) );
  NAND2_X1 U12321 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(P3_EAX_REG_29__SCAN_IN), 
        .ZN(n9987) );
  NOR3_X1 U12322 ( .A1(n17296), .A2(n17492), .A3(n17494), .ZN(n17284) );
  NOR2_X1 U12323 ( .A1(n17296), .A2(n17492), .ZN(n17292) );
  NOR2_X1 U12324 ( .A1(n17488), .A2(n17306), .ZN(n17301) );
  OR2_X1 U12325 ( .A1(n17486), .A2(n17305), .ZN(n17306) );
  AND2_X1 U12326 ( .A1(n17357), .A2(n9692), .ZN(n17311) );
  NAND2_X1 U12327 ( .A1(n17357), .A2(n9989), .ZN(n17312) );
  NOR3_X1 U12328 ( .A1(n17476), .A2(n17474), .A3(n17345), .ZN(n17332) );
  NOR2_X1 U12329 ( .A1(n17472), .A2(n17343), .ZN(n17337) );
  NOR2_X1 U12330 ( .A1(n17412), .A2(n18262), .ZN(n17349) );
  NOR2_X1 U12331 ( .A1(n17529), .A2(n17360), .ZN(n17357) );
  NAND2_X1 U12332 ( .A1(n17357), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n17356) );
  NOR2_X1 U12333 ( .A1(n17271), .A2(n17272), .ZN(n9984) );
  NOR2_X1 U12334 ( .A1(n12306), .A2(n9884), .ZN(n9883) );
  AND2_X1 U12335 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17411), .ZN(n17416) );
  INV_X1 U12336 ( .A(n17420), .ZN(n17417) );
  INV_X1 U12337 ( .A(n15866), .ZN(n17270) );
  CLKBUF_X1 U12338 ( .A(n17443), .Z(n17462) );
  NOR2_X1 U12339 ( .A1(n18884), .A2(n17522), .ZN(n17523) );
  OAI211_X1 U12340 ( .C1(n18884), .C2(n18885), .A(n17468), .B(n17467), .ZN(
        n17530) );
  CLKBUF_X1 U12341 ( .A(n17523), .Z(n17531) );
  NAND2_X1 U12342 ( .A1(n16562), .A2(n10061), .ZN(n16361) );
  OAI21_X1 U12343 ( .B1(n17553), .B2(n10010), .A(n16418), .ZN(n17548) );
  NAND2_X1 U12344 ( .A1(n17633), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17619) );
  NOR2_X1 U12345 ( .A1(n17687), .A2(n17967), .ZN(n17633) );
  NAND2_X1 U12346 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17838), .ZN(n17738) );
  INV_X1 U12347 ( .A(n17738), .ZN(n17756) );
  NAND3_X1 U12348 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(n10040), .ZN(n17820) );
  NOR2_X1 U12349 ( .A1(n16873), .A2(n10041), .ZN(n10040) );
  NAND2_X1 U12350 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U12351 ( .A1(n10044), .A2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17847) );
  NOR2_X1 U12352 ( .A1(n16873), .A2(n10045), .ZN(n10044) );
  AOI21_X2 U12353 ( .B1(n18735), .B2(n15708), .A(n12568), .ZN(n17886) );
  INV_X1 U12354 ( .A(n17894), .ZN(n17884) );
  NAND2_X1 U12355 ( .A1(n17682), .A2(n17738), .ZN(n17894) );
  INV_X1 U12356 ( .A(n17886), .ZN(n17900) );
  NOR2_X1 U12357 ( .A1(n18210), .A2(n16416), .ZN(n9870) );
  INV_X1 U12358 ( .A(n10008), .ZN(n17563) );
  INV_X1 U12359 ( .A(n17591), .ZN(n17595) );
  NOR2_X1 U12360 ( .A1(n18011), .A2(n18090), .ZN(n18034) );
  INV_X1 U12361 ( .A(n18215), .ZN(n18126) );
  NOR2_X1 U12362 ( .A1(n18165), .A2(n18707), .ZN(n18167) );
  INV_X1 U12363 ( .A(n18706), .ZN(n18187) );
  NAND2_X1 U12364 ( .A1(n12516), .A2(n15715), .ZN(n18664) );
  INV_X1 U12365 ( .A(n18209), .ZN(n18223) );
  INV_X1 U12366 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18469) );
  INV_X1 U12367 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18701) );
  NOR2_X1 U12368 ( .A1(n18236), .A2(n15724), .ZN(n18867) );
  INV_X1 U12369 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18719) );
  INV_X1 U12370 ( .A(n18867), .ZN(n18864) );
  NAND2_X1 U12371 ( .A1(n18758), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18894) );
  CLKBUF_X1 U12372 ( .A(n16503), .Z(n16509) );
  INV_X1 U12373 ( .A(n14288), .ZN(n14475) );
  AND2_X1 U12374 ( .A1(n9842), .A2(n9841), .ZN(P1_U2968) );
  NAND2_X1 U12375 ( .A1(n9675), .A2(n20007), .ZN(n9841) );
  OAI21_X1 U12376 ( .B1(n14785), .B2(n20007), .A(n9981), .ZN(P1_U2969) );
  INV_X1 U12377 ( .A(n9915), .ZN(n9981) );
  AOI21_X1 U12378 ( .B1(n14288), .B2(n16032), .A(n10018), .ZN(n14096) );
  NAND2_X1 U12379 ( .A1(n10021), .A2(n10019), .ZN(n10018) );
  AND2_X1 U12380 ( .A1(n12022), .A2(n12021), .ZN(n12023) );
  NAND2_X1 U12381 ( .A1(n14268), .A2(n19127), .ZN(n12024) );
  AND2_X1 U12382 ( .A1(n12263), .A2(n12262), .ZN(n12264) );
  AND2_X1 U12383 ( .A1(n15201), .A2(n15200), .ZN(n15202) );
  NAND2_X1 U12384 ( .A1(n15307), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10213) );
  OR2_X1 U12385 ( .A1(n16098), .A2(n16277), .ZN(n10214) );
  NAND2_X1 U12386 ( .A1(n15320), .A2(n15319), .ZN(n15321) );
  AND2_X1 U12387 ( .A1(n15318), .A2(n15317), .ZN(n15319) );
  AOI21_X1 U12388 ( .B1(n9946), .B2(n9945), .A(n9943), .ZN(n14260) );
  NOR2_X1 U12389 ( .A1(n15186), .A2(n16292), .ZN(n9945) );
  INV_X1 U12390 ( .A(n15185), .ZN(n9946) );
  NAND2_X1 U12391 ( .A1(n9788), .A2(n9786), .ZN(n15505) );
  NOR3_X1 U12392 ( .A1(n9787), .A2(n15503), .A3(n15504), .ZN(n9786) );
  NOR3_X1 U12393 ( .A1(n10036), .A2(n10035), .A3(n10034), .ZN(n10033) );
  OR2_X1 U12394 ( .A1(n16570), .A2(n16569), .ZN(n10035) );
  INV_X1 U12395 ( .A(n9985), .ZN(n17422) );
  AOI21_X1 U12396 ( .B1(n16398), .B2(n17814), .A(n12580), .ZN(n12581) );
  OAI21_X1 U12397 ( .B1(n16402), .B2(n17904), .A(n12579), .ZN(n12580) );
  AOI21_X1 U12398 ( .B1(n16399), .B2(n17815), .A(n12578), .ZN(n12579) );
  INV_X1 U12399 ( .A(n9867), .ZN(n9866) );
  NAND2_X1 U12400 ( .A1(n9871), .A2(n9870), .ZN(n9869) );
  NAND2_X1 U12401 ( .A1(n13478), .A2(n10244), .ZN(n13838) );
  NAND2_X1 U12402 ( .A1(n13306), .A2(n13177), .ZN(n10894) );
  OR3_X1 U12403 ( .A1(n15412), .A2(n10088), .A3(n9763), .ZN(n9672) );
  NAND2_X2 U12404 ( .A1(n13134), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11319) );
  AND2_X1 U12405 ( .A1(n9830), .A2(n10226), .ZN(n12959) );
  INV_X1 U12406 ( .A(n10396), .ZN(n10877) );
  OR2_X1 U12407 ( .A1(n12606), .A2(n12589), .ZN(n9673) );
  AND2_X1 U12408 ( .A1(n10194), .A2(n10200), .ZN(n13989) );
  AND2_X2 U12409 ( .A1(n11266), .A2(n11265), .ZN(n9675) );
  AND2_X1 U12410 ( .A1(n10093), .A2(n10091), .ZN(n9676) );
  AND4_X1 U12411 ( .A1(n13420), .A2(n13419), .A3(n13418), .A4(n13417), .ZN(
        n9677) );
  AND2_X1 U12412 ( .A1(n17791), .A2(n16406), .ZN(n9678) );
  OR2_X1 U12413 ( .A1(n12867), .A2(n15590), .ZN(n13377) );
  AOI21_X1 U12414 ( .B1(n11251), .B2(n10257), .A(n9971), .ZN(n9969) );
  INV_X1 U12415 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17846) );
  AND2_X1 U12416 ( .A1(n9702), .A2(n14105), .ZN(n9679) );
  INV_X1 U12418 ( .A(n12115), .ZN(n12146) );
  NAND2_X1 U12419 ( .A1(n13478), .A2(n11610), .ZN(n13477) );
  INV_X1 U12420 ( .A(n13278), .ZN(n10134) );
  NAND2_X1 U12421 ( .A1(n10237), .A2(n10240), .ZN(n15079) );
  OR3_X1 U12422 ( .A1(n12606), .A2(n12589), .A3(n10121), .ZN(n9680) );
  AND2_X1 U12423 ( .A1(n13478), .A2(n9737), .ZN(n13837) );
  NAND2_X1 U12424 ( .A1(n15444), .A2(n9761), .ZN(n15002) );
  NAND2_X1 U12425 ( .A1(n10068), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9681) );
  AND2_X1 U12426 ( .A1(n10102), .A2(n10101), .ZN(n9682) );
  AND2_X1 U12427 ( .A1(n9639), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12181) );
  AND2_X1 U12428 ( .A1(n10244), .A2(n9831), .ZN(n9683) );
  AND2_X1 U12429 ( .A1(n10123), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9684) );
  AND2_X1 U12430 ( .A1(n10140), .A2(n10138), .ZN(n9685) );
  AND2_X1 U12431 ( .A1(n19121), .A2(n12229), .ZN(n9686) );
  AND2_X1 U12432 ( .A1(n9686), .A2(n11610), .ZN(n9687) );
  AND2_X1 U12433 ( .A1(n10024), .A2(n10023), .ZN(n9688) );
  AND2_X1 U12434 ( .A1(n9682), .A2(n15261), .ZN(n9689) );
  AND2_X1 U12435 ( .A1(n10236), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9690) );
  INV_X1 U12436 ( .A(n20173), .ZN(n16032) );
  INV_X1 U12437 ( .A(n17813), .ZN(n10010) );
  AND2_X1 U12438 ( .A1(n10162), .A2(n10161), .ZN(n9691) );
  AND2_X1 U12439 ( .A1(n9989), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n9692) );
  AND2_X2 U12440 ( .A1(n12033), .A2(n11376), .ZN(n11578) );
  INV_X4 U12441 ( .A(n12283), .ZN(n17186) );
  NAND2_X2 U12442 ( .A1(n13398), .A2(n19988), .ZN(n10230) );
  OR3_X1 U12443 ( .A1(n17296), .A2(n17492), .A3(n9987), .ZN(n9693) );
  INV_X2 U12444 ( .A(n12295), .ZN(n17195) );
  NAND2_X1 U12446 ( .A1(n15224), .A2(n14232), .ZN(n9694) );
  NAND2_X1 U12447 ( .A1(n14355), .A2(n14354), .ZN(n14344) );
  AND2_X1 U12448 ( .A1(n13676), .A2(n9679), .ZN(n9696) );
  NAND2_X1 U12449 ( .A1(n10114), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12613) );
  NOR2_X1 U12450 ( .A1(n11839), .A2(n11840), .ZN(n12027) );
  INV_X1 U12451 ( .A(n17624), .ZN(n17682) );
  NOR2_X1 U12452 ( .A1(n12616), .A2(n19068), .ZN(n12617) );
  NOR2_X1 U12453 ( .A1(n12618), .A2(n19230), .ZN(n12619) );
  AND2_X1 U12454 ( .A1(n17357), .A2(n9991), .ZN(n9698) );
  OR2_X1 U12455 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n14222), .ZN(n9699) );
  AND3_X1 U12456 ( .A1(n11493), .A2(n11492), .A3(n11491), .ZN(n11920) );
  AND2_X1 U12457 ( .A1(n12259), .A2(n11439), .ZN(n9700) );
  AND2_X1 U12458 ( .A1(n10194), .A2(n10197), .ZN(n14507) );
  AND2_X1 U12459 ( .A1(n13754), .A2(n10028), .ZN(n9701) );
  AND2_X1 U12460 ( .A1(n10157), .A2(n13675), .ZN(n9702) );
  AND2_X1 U12461 ( .A1(n12650), .A2(n9691), .ZN(n9703) );
  NOR2_X1 U12462 ( .A1(n10455), .A2(n10324), .ZN(n9704) );
  AND2_X1 U12463 ( .A1(n13845), .A2(n13755), .ZN(n9705) );
  NAND2_X1 U12464 ( .A1(n14929), .A2(n11237), .ZN(n14722) );
  NAND2_X1 U12465 ( .A1(n14156), .A2(n10152), .ZN(n9706) );
  NAND2_X1 U12466 ( .A1(n10220), .A2(n15375), .ZN(n15213) );
  INV_X1 U12467 ( .A(n15375), .ZN(n10219) );
  AND2_X1 U12468 ( .A1(n9811), .A2(n15405), .ZN(n9708) );
  NOR2_X1 U12469 ( .A1(n15060), .A2(n15062), .ZN(n15061) );
  OR2_X1 U12470 ( .A1(n9649), .A2(n13971), .ZN(n9709) );
  OR2_X1 U12471 ( .A1(n15594), .A2(n11512), .ZN(n9710) );
  OR3_X1 U12472 ( .A1(n15412), .A2(n10088), .A3(n15411), .ZN(n9711) );
  AND3_X1 U12473 ( .A1(n9843), .A2(n11264), .A3(n9844), .ZN(n9712) );
  INV_X1 U12474 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13812) );
  AND2_X1 U12475 ( .A1(n15172), .A2(n15170), .ZN(n9713) );
  AND2_X1 U12476 ( .A1(n13122), .A2(n9908), .ZN(n9714) );
  INV_X1 U12477 ( .A(n10170), .ZN(n13076) );
  AND2_X1 U12478 ( .A1(n9781), .A2(n10070), .ZN(n9715) );
  OR2_X1 U12479 ( .A1(n19469), .A2(n13874), .ZN(n9716) );
  AND2_X1 U12480 ( .A1(n9911), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9717) );
  AND4_X1 U12481 ( .A1(n9895), .A2(n9892), .A3(n9891), .A4(n9890), .ZN(n9718)
         );
  OR2_X1 U12482 ( .A1(n13895), .A2(n14247), .ZN(n9719) );
  NAND2_X1 U12483 ( .A1(n15104), .A2(n15103), .ZN(n12670) );
  AND4_X1 U12484 ( .A1(n10215), .A2(n15309), .A3(n10214), .A4(n10213), .ZN(
        n9720) );
  NAND3_X1 U12485 ( .A1(n13097), .A2(n10414), .A3(n10413), .ZN(n9721) );
  OR2_X1 U12486 ( .A1(n14329), .A2(n10207), .ZN(n14304) );
  OR2_X1 U12487 ( .A1(n11917), .A2(n11522), .ZN(n11524) );
  AND2_X1 U12488 ( .A1(n9849), .A2(n15957), .ZN(n9722) );
  OR2_X1 U12489 ( .A1(n11353), .A2(n11354), .ZN(n9723) );
  NAND2_X1 U12490 ( .A1(n9970), .A2(n11249), .ZN(n9724) );
  INV_X1 U12491 ( .A(n9781), .ZN(n10077) );
  NAND2_X1 U12492 ( .A1(n9782), .A2(n13678), .ZN(n9781) );
  INV_X1 U12493 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19017) );
  INV_X1 U12494 ( .A(n17773), .ZN(n18093) );
  OAI21_X1 U12495 ( .B1(n17819), .B2(n9877), .A(n9876), .ZN(n17773) );
  AND2_X1 U12496 ( .A1(n11237), .A2(n10180), .ZN(n9725) );
  OR2_X1 U12497 ( .A1(n11343), .A2(n11344), .ZN(n9726) );
  NOR2_X1 U12498 ( .A1(n17590), .A2(n10032), .ZN(n9727) );
  AND2_X1 U12499 ( .A1(n11255), .A2(n11254), .ZN(n11268) );
  AND2_X1 U12500 ( .A1(n9963), .A2(n15524), .ZN(n9728) );
  AND2_X1 U12501 ( .A1(n10429), .A2(n12898), .ZN(n9729) );
  AND2_X1 U12502 ( .A1(n9963), .A2(n15519), .ZN(n9730) );
  OR2_X1 U12503 ( .A1(n12307), .A2(n15625), .ZN(n9731) );
  AND2_X1 U12504 ( .A1(n9701), .A2(n10026), .ZN(n9732) );
  NAND2_X1 U12505 ( .A1(n15066), .A2(n11772), .ZN(n11786) );
  AND2_X1 U12506 ( .A1(n10166), .A2(n10165), .ZN(n9733) );
  INV_X1 U12507 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19230) );
  XNOR2_X1 U12508 ( .A(n10587), .B(n10586), .ZN(n11172) );
  INV_X1 U12509 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10469) );
  INV_X1 U12510 ( .A(n13605), .ZN(n10139) );
  NAND2_X1 U12511 ( .A1(n10076), .A2(n9715), .ZN(n10072) );
  INV_X1 U12512 ( .A(n10795), .ZN(n9914) );
  OR2_X1 U12513 ( .A1(n12259), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10263) );
  NAND2_X1 U12514 ( .A1(n9917), .A2(n10636), .ZN(n13494) );
  NOR2_X1 U12515 ( .A1(n13932), .A2(n13627), .ZN(n13628) );
  NOR2_X1 U12516 ( .A1(n15085), .A2(n15087), .ZN(n15086) );
  NOR2_X1 U12517 ( .A1(n12606), .A2(n10118), .ZN(n12604) );
  NOR2_X1 U12518 ( .A1(n12609), .A2(n16176), .ZN(n12607) );
  NOR2_X1 U12519 ( .A1(n12611), .A2(n15296), .ZN(n12608) );
  NOR3_X1 U12520 ( .A1(n17820), .A2(n17807), .A3(n12569), .ZN(n12570) );
  INV_X1 U12521 ( .A(n9983), .ZN(n17364) );
  NAND2_X1 U12522 ( .A1(n9985), .A2(n9984), .ZN(n9983) );
  NAND2_X1 U12523 ( .A1(n13478), .A2(n9687), .ZN(n9734) );
  AND2_X1 U12524 ( .A1(n15883), .A2(n9688), .ZN(n9735) );
  NAND2_X1 U12525 ( .A1(n9816), .A2(n9815), .ZN(n19221) );
  NAND2_X1 U12526 ( .A1(n11218), .A2(n11217), .ZN(n15955) );
  NAND2_X1 U12527 ( .A1(n9838), .A2(n11198), .ZN(n13492) );
  AND2_X1 U12528 ( .A1(n15764), .A2(n9682), .ZN(n9736) );
  AND2_X1 U12529 ( .A1(n9828), .A2(n9710), .ZN(n12958) );
  NOR2_X1 U12530 ( .A1(n10429), .A2(n10386), .ZN(n12753) );
  NOR3_X1 U12531 ( .A1(n12606), .A2(n12589), .A3(n15269), .ZN(n12605) );
  NAND2_X1 U12532 ( .A1(n15065), .A2(n15067), .ZN(n15066) );
  AND2_X1 U12533 ( .A1(n9687), .A2(n13961), .ZN(n9737) );
  AND2_X1 U12534 ( .A1(n9971), .A2(n10189), .ZN(n9738) );
  INV_X1 U12535 ( .A(n10015), .ZN(n14410) );
  NOR2_X1 U12536 ( .A1(n14422), .A2(n14408), .ZN(n10015) );
  INV_X1 U12537 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19986) );
  AND2_X1 U12538 ( .A1(n10047), .A2(n10050), .ZN(n9739) );
  AND2_X1 U12539 ( .A1(n11577), .A2(n12208), .ZN(n9740) );
  OR2_X1 U12540 ( .A1(n15154), .A2(n12647), .ZN(n9741) );
  NOR2_X1 U12541 ( .A1(n16616), .A2(n17588), .ZN(n9742) );
  AND2_X1 U12542 ( .A1(n15126), .A2(n11730), .ZN(n9743) );
  AND2_X1 U12543 ( .A1(n11166), .A2(n10192), .ZN(n9744) );
  AND2_X1 U12544 ( .A1(n10529), .A2(n10528), .ZN(n9745) );
  OR2_X1 U12545 ( .A1(n16517), .A2(n18751), .ZN(n9746) );
  INV_X1 U12546 ( .A(n15085), .ZN(n10237) );
  INV_X1 U12547 ( .A(n10153), .ZN(n10152) );
  OR2_X1 U12548 ( .A1(n14152), .A2(n10154), .ZN(n10153) );
  AND2_X1 U12549 ( .A1(n10202), .A2(n10201), .ZN(n9747) );
  NAND2_X1 U12550 ( .A1(n13676), .A2(n9702), .ZN(n10159) );
  NAND2_X1 U12551 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U12552 ( .A1(n16178), .A2(n15291), .ZN(n9749) );
  AND2_X1 U12553 ( .A1(n10139), .A2(n9685), .ZN(n9750) );
  AND2_X1 U12554 ( .A1(n10151), .A2(n10150), .ZN(n9751) );
  INV_X1 U12555 ( .A(n12531), .ZN(n12517) );
  NAND2_X1 U12556 ( .A1(n17365), .A2(n12514), .ZN(n12531) );
  AND2_X1 U12557 ( .A1(n10143), .A2(n10142), .ZN(n9752) );
  AND2_X1 U12558 ( .A1(n9688), .A2(n14432), .ZN(n9753) );
  AND2_X1 U12559 ( .A1(n9928), .A2(n14145), .ZN(n9754) );
  AND2_X1 U12560 ( .A1(n16154), .A2(n10112), .ZN(n9755) );
  AND2_X1 U12561 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9756) );
  NAND2_X1 U12562 ( .A1(n19139), .A2(n12208), .ZN(n13256) );
  INV_X1 U12563 ( .A(n19227), .ZN(n16251) );
  NAND2_X1 U12564 ( .A1(n13460), .A2(n13459), .ZN(n12961) );
  NOR2_X1 U12565 ( .A1(n18093), .A2(n12392), .ZN(n17812) );
  AND2_X1 U12566 ( .A1(n12954), .A2(n19975), .ZN(n19250) );
  NOR2_X1 U12567 ( .A1(n13925), .A2(n13783), .ZN(n9757) );
  NAND2_X1 U12568 ( .A1(n13460), .A2(n10236), .ZN(n13015) );
  NAND2_X1 U12569 ( .A1(n12756), .A2(n12755), .ZN(n19231) );
  NAND2_X1 U12570 ( .A1(n19139), .A2(n9740), .ZN(n13467) );
  NAND2_X1 U12571 ( .A1(n12597), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12590) );
  NAND2_X1 U12572 ( .A1(n10410), .A2(n10588), .ZN(n13066) );
  NOR2_X1 U12573 ( .A1(n12602), .A2(n16140), .ZN(n12600) );
  AND2_X1 U12574 ( .A1(n10066), .A2(n10068), .ZN(n9758) );
  AND2_X1 U12575 ( .A1(n10092), .A2(n9676), .ZN(n9759) );
  INV_X1 U12576 ( .A(n12752), .ZN(n11283) );
  XNOR2_X1 U12577 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13677), .ZN(
        n9760) );
  OR2_X1 U12578 ( .A1(n11868), .A2(n11867), .ZN(n13679) );
  NOR2_X1 U12579 ( .A1(n13042), .A2(n13043), .ZN(n13041) );
  AND2_X1 U12580 ( .A1(n10147), .A2(n15013), .ZN(n9761) );
  INV_X1 U12581 ( .A(n14105), .ZN(n10158) );
  NOR2_X1 U12582 ( .A1(n13278), .A2(n12150), .ZN(n13337) );
  INV_X1 U12583 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n16039) );
  INV_X1 U12584 ( .A(n14196), .ZN(n10163) );
  INV_X1 U12585 ( .A(n14157), .ZN(n10154) );
  NAND2_X1 U12586 ( .A1(n17711), .A2(n10256), .ZN(n17681) );
  AND2_X1 U12587 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9762) );
  OR2_X1 U12588 ( .A1(n12966), .A2(n15808), .ZN(n20007) );
  OR2_X1 U12589 ( .A1(n15411), .A2(n15068), .ZN(n9763) );
  AND2_X1 U12590 ( .A1(n10127), .A2(n10126), .ZN(n9764) );
  AND2_X1 U12591 ( .A1(n14382), .A2(n14396), .ZN(n9765) );
  AND2_X1 U12592 ( .A1(n10110), .A2(n9634), .ZN(n9766) );
  AND2_X1 U12593 ( .A1(n13460), .A2(n9690), .ZN(n19139) );
  NAND2_X1 U12594 ( .A1(n10131), .A2(n10134), .ZN(n10136) );
  INV_X1 U12595 ( .A(n10062), .ZN(n10061) );
  NAND2_X1 U12596 ( .A1(n10063), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10062) );
  AND2_X1 U12597 ( .A1(n10134), .A2(n10135), .ZN(n9767) );
  AND2_X1 U12598 ( .A1(n10097), .A2(n10095), .ZN(n9768) );
  AND2_X1 U12599 ( .A1(n10108), .A2(n9634), .ZN(n9769) );
  NOR2_X1 U12600 ( .A1(n12268), .A2(n12270), .ZN(n15626) );
  INV_X1 U12601 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n9879) );
  OR4_X1 U12602 ( .A1(n17482), .A2(n17480), .A3(n17478), .A4(n17472), .ZN(
        n9770) );
  AND2_X1 U12603 ( .A1(n12597), .A2(n9684), .ZN(n9771) );
  AND2_X1 U12604 ( .A1(n16562), .A2(n10063), .ZN(n9772) );
  AND4_X1 U12605 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        n9773) );
  AND2_X1 U12606 ( .A1(n11785), .A2(n11804), .ZN(n9774) );
  INV_X1 U12607 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17887) );
  AND2_X1 U12608 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n9775) );
  INV_X1 U12609 ( .A(n13991), .ZN(n10200) );
  INV_X1 U12610 ( .A(n19919), .ZN(n19998) );
  NOR2_X2 U12611 ( .A1(n18904), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19919) );
  INV_X1 U12612 ( .A(n19066), .ZN(n15785) );
  INV_X1 U12613 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n9986) );
  NOR2_X1 U12614 ( .A1(n17887), .A2(n16873), .ZN(n10042) );
  INV_X1 U12615 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U12616 ( .A1(n15327), .A2(n15197), .ZN(n9776) );
  INV_X1 U12617 ( .A(n10257), .ZN(n9973) );
  AND2_X1 U12618 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9777) );
  INV_X1 U12619 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10045) );
  INV_X1 U12620 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n9992) );
  INV_X1 U12621 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10065) );
  INV_X1 U12622 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10064) );
  AND2_X1 U12623 ( .A1(n11256), .A2(n14093), .ZN(n9778) );
  INV_X1 U12624 ( .A(n14781), .ZN(n10191) );
  INV_X1 U12625 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9880) );
  INV_X1 U12626 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10150) );
  INV_X1 U12627 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n9878) );
  INV_X1 U12628 ( .A(n20709), .ZN(n9779) );
  INV_X1 U12629 ( .A(n9779), .ZN(n9780) );
  OAI22_X2 U12630 ( .A1(n16425), .A2(n20222), .B1(n20933), .B2(n20221), .ZN(
        n20651) );
  NAND2_X2 U12631 ( .A1(n18906), .A2(n12656), .ZN(n19099) );
  AND2_X1 U12632 ( .A1(n16323), .A2(n12693), .ZN(n18906) );
  OAI22_X2 U12633 ( .A1(n20195), .A2(n20222), .B1(n20194), .B2(n20221), .ZN(
        n20679) );
  OAI22_X2 U12634 ( .A1(n20215), .A2(n20222), .B1(n14567), .B2(n20221), .ZN(
        n20703) );
  NAND2_X1 U12635 ( .A1(n15960), .A2(n14535), .ZN(n20222) );
  NOR2_X1 U12636 ( .A1(n18881), .A2(n17446), .ZN(n17443) );
  AOI22_X2 U12637 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19313), .ZN(n19816) );
  NOR2_X2 U12638 ( .A1(n19269), .A2(n19268), .ZN(n19313) );
  NOR3_X2 U12639 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18726), .A3(
        n18446), .ZN(n18420) );
  NOR2_X2 U12640 ( .A1(n20225), .A2(n13522), .ZN(n20707) );
  NAND3_X1 U12641 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16039), .A3(n13521), 
        .ZN(n20225) );
  NOR2_X2 U12642 ( .A1(n19305), .A2(n19309), .ZN(n19831) );
  NAND2_X1 U12643 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19781), .ZN(n19309) );
  XNOR2_X2 U12644 ( .A(n9783), .B(n9942), .ZN(n10071) );
  NOR2_X2 U12645 ( .A1(n13355), .A2(n13361), .ZN(n9785) );
  AND2_X2 U12646 ( .A1(n11379), .A2(n11378), .ZN(n11443) );
  NAND2_X2 U12647 ( .A1(n11332), .A2(n11331), .ZN(n11420) );
  NAND2_X1 U12648 ( .A1(n9791), .A2(n13901), .ZN(n9789) );
  INV_X1 U12649 ( .A(n9791), .ZN(n9863) );
  NAND2_X1 U12650 ( .A1(n9864), .A2(n13895), .ZN(n9791) );
  NAND2_X1 U12651 ( .A1(n9862), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9792) );
  OAI21_X2 U12652 ( .B1(n9864), .B2(n13901), .A(n9719), .ZN(n9862) );
  NAND2_X2 U12653 ( .A1(n16221), .A2(n14255), .ZN(n15548) );
  AND2_X2 U12654 ( .A1(n9940), .A2(n13378), .ZN(n13649) );
  AND2_X1 U12655 ( .A1(n13378), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U12656 ( .A1(n13649), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n9795) );
  NAND3_X1 U12657 ( .A1(n9798), .A2(n11918), .A3(n11524), .ZN(n9797) );
  NAND2_X2 U12658 ( .A1(n13358), .A2(n11487), .ZN(n11919) );
  NAND4_X1 U12659 ( .A1(n13891), .A2(n10073), .A3(n10074), .A4(n10072), .ZN(
        n9864) );
  OR2_X2 U12660 ( .A1(n16199), .A2(n9865), .ZN(n15530) );
  NAND4_X1 U12661 ( .A1(n11398), .A2(n9802), .A3(n11397), .A4(n11396), .ZN(
        n9801) );
  NAND4_X1 U12662 ( .A1(n11393), .A2(n9804), .A3(n11394), .A4(n11392), .ZN(
        n9803) );
  NAND2_X1 U12663 ( .A1(n15532), .A2(n14128), .ZN(n9950) );
  XNOR2_X2 U12664 ( .A(n14102), .B(n13909), .ZN(n14100) );
  XNOR2_X2 U12665 ( .A(n11919), .B(n9807), .ZN(n12843) );
  NAND2_X1 U12666 ( .A1(n9707), .A2(n9677), .ZN(n9809) );
  NAND2_X1 U12667 ( .A1(n9810), .A2(n9942), .ZN(n13425) );
  NAND3_X1 U12668 ( .A1(n9961), .A2(n9960), .A3(n9958), .ZN(n9811) );
  NAND4_X1 U12669 ( .A1(n9961), .A2(n15390), .A3(n9960), .A4(n9958), .ZN(n9814) );
  NAND2_X1 U12670 ( .A1(n9818), .A2(n13644), .ZN(n13897) );
  NAND2_X1 U12671 ( .A1(n19221), .A2(n19222), .ZN(n9818) );
  NOR2_X2 U12672 ( .A1(n11419), .A2(n9823), .ZN(n11424) );
  NAND2_X1 U12673 ( .A1(n11418), .A2(n19287), .ZN(n9823) );
  OAI21_X2 U12674 ( .B1(n14229), .B2(n9827), .A(n9826), .ZN(n15152) );
  NAND4_X1 U12675 ( .A1(n9830), .A2(n9828), .A3(n9710), .A4(n10226), .ZN(n9829) );
  NAND2_X1 U12676 ( .A1(n9829), .A2(n9830), .ZN(n12986) );
  NOR2_X2 U12677 ( .A1(n15072), .A2(n11751), .ZN(n11771) );
  XNOR2_X1 U12678 ( .A(n11786), .B(n9774), .ZN(n15060) );
  NAND2_X1 U12679 ( .A1(n13492), .A2(n13493), .ZN(n9837) );
  NAND2_X1 U12680 ( .A1(n13451), .A2(n13450), .ZN(n9838) );
  XNOR2_X1 U12681 ( .A(n9839), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13557) );
  NAND2_X2 U12682 ( .A1(n9840), .A2(n20291), .ZN(n10483) );
  NAND4_X1 U12683 ( .A1(n9844), .A2(n9843), .A3(n9675), .A4(n11264), .ZN(n9842) );
  INV_X1 U12684 ( .A(n11260), .ZN(n9844) );
  OAI21_X2 U12685 ( .B1(n12752), .B2(n20192), .A(n13326), .ZN(n13068) );
  NAND2_X2 U12686 ( .A1(n9976), .A2(n9847), .ZN(n14614) );
  NAND2_X2 U12687 ( .A1(n9848), .A2(n11248), .ZN(n11250) );
  NAND2_X1 U12688 ( .A1(n15955), .A2(n15957), .ZN(n11229) );
  INV_X1 U12689 ( .A(n9705), .ZN(n9849) );
  NAND3_X1 U12690 ( .A1(n11253), .A2(n9850), .A3(n14086), .ZN(n11270) );
  NOR2_X2 U12691 ( .A1(n14640), .A2(n14643), .ZN(n9850) );
  NAND2_X1 U12692 ( .A1(n9857), .A2(n11442), .ZN(n11464) );
  NAND2_X1 U12693 ( .A1(n9852), .A2(n9856), .ZN(n11463) );
  NOR2_X1 U12694 ( .A1(n9853), .A2(n9854), .ZN(n9852) );
  INV_X1 U12695 ( .A(n9855), .ZN(n9853) );
  NAND2_X1 U12696 ( .A1(n11903), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9856) );
  NAND2_X1 U12697 ( .A1(n11488), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9857) );
  NAND2_X1 U12698 ( .A1(n9863), .A2(n13901), .ZN(n9859) );
  INV_X1 U12699 ( .A(n9862), .ZN(n9860) );
  NAND3_X1 U12700 ( .A1(n9869), .A2(n16419), .A3(n9866), .ZN(P3_U2834) );
  AOI21_X1 U12701 ( .B1(n12390), .B2(n9879), .A(n9878), .ZN(n9876) );
  INV_X1 U12702 ( .A(n12390), .ZN(n9877) );
  NAND2_X1 U12703 ( .A1(n17818), .A2(n12390), .ZN(n12391) );
  AND2_X2 U12704 ( .A1(n9727), .A2(n10008), .ZN(n16403) );
  NAND2_X1 U12705 ( .A1(n9882), .A2(n17791), .ZN(n17706) );
  OAI21_X1 U12706 ( .B1(n17812), .B2(n17813), .A(n9882), .ZN(n18132) );
  NAND2_X1 U12707 ( .A1(n17773), .A2(n10009), .ZN(n9882) );
  NAND3_X1 U12708 ( .A1(n12304), .A2(n12305), .A3(n9885), .ZN(n9884) );
  NAND2_X2 U12709 ( .A1(n9887), .A2(n9886), .ZN(n17168) );
  NAND2_X1 U12710 ( .A1(n17648), .A2(n12401), .ZN(n17596) );
  NAND2_X1 U12711 ( .A1(n9889), .A2(n17648), .ZN(n17591) );
  NAND4_X1 U12712 ( .A1(n9898), .A2(n12428), .A3(n9896), .A4(n9718), .ZN(
        n12429) );
  OAI21_X1 U12713 ( .B1(n16539), .B2(n9901), .A(n12518), .ZN(n9899) );
  NAND2_X1 U12714 ( .A1(n16544), .A2(n12531), .ZN(n9901) );
  INV_X2 U12715 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18859) );
  NOR2_X1 U12716 ( .A1(n11151), .A2(n9903), .ZN(n13059) );
  NOR2_X1 U12717 ( .A1(n13077), .A2(n9903), .ZN(n13084) );
  NAND2_X2 U12718 ( .A1(n10416), .A2(n10406), .ZN(n9903) );
  INV_X1 U12719 ( .A(n13775), .ZN(n9904) );
  NAND2_X1 U12720 ( .A1(n13982), .A2(n13981), .ZN(n13980) );
  NOR2_X1 U12721 ( .A1(n13536), .A2(n9908), .ZN(n11284) );
  NAND2_X1 U12722 ( .A1(n10415), .A2(n9908), .ZN(n10360) );
  NAND2_X2 U12723 ( .A1(n13522), .A2(n9908), .ZN(n10415) );
  NAND2_X1 U12724 ( .A1(n20192), .A2(n9908), .ZN(n11090) );
  NAND2_X1 U12725 ( .A1(n13070), .A2(n9908), .ZN(n10170) );
  AND2_X1 U12726 ( .A1(n10412), .A2(n9908), .ZN(n11225) );
  NOR2_X1 U12727 ( .A1(n13304), .A2(n9908), .ZN(n10408) );
  AND2_X1 U12728 ( .A1(n13080), .A2(n9908), .ZN(n10192) );
  NAND2_X1 U12729 ( .A1(n13068), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9910) );
  AOI21_X1 U12730 ( .B1(n10411), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9729), 
        .ZN(n9909) );
  NAND2_X1 U12731 ( .A1(n10472), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10422) );
  NAND2_X1 U12732 ( .A1(n10636), .A2(n9916), .ZN(n9918) );
  NOR2_X2 U12733 ( .A1(n14419), .A2(n9919), .ZN(n14355) );
  XNOR2_X2 U12734 ( .A(n13678), .B(n13893), .ZN(n13681) );
  NAND2_X2 U12735 ( .A1(n9941), .A2(n9942), .ZN(n13678) );
  NAND2_X1 U12736 ( .A1(n9926), .A2(n9925), .ZN(n15232) );
  NAND3_X1 U12737 ( .A1(n14138), .A2(n9754), .A3(n14137), .ZN(n9926) );
  NAND3_X1 U12738 ( .A1(n14138), .A2(n14137), .A3(n14145), .ZN(n9930) );
  NAND2_X1 U12739 ( .A1(n9930), .A2(n15291), .ZN(n16180) );
  AOI21_X2 U12740 ( .B1(n15282), .B2(n15236), .A(n15235), .ZN(n15474) );
  NAND2_X2 U12741 ( .A1(n9940), .A2(n13382), .ZN(n19572) );
  NAND2_X2 U12742 ( .A1(n9940), .A2(n13367), .ZN(n19640) );
  INV_X2 U12743 ( .A(n13384), .ZN(n9940) );
  AND2_X2 U12744 ( .A1(n9954), .A2(n9953), .ZN(n9941) );
  NAND2_X2 U12745 ( .A1(n9950), .A2(n14132), .ZN(n15521) );
  NAND2_X1 U12746 ( .A1(n13399), .A2(n13398), .ZN(n9952) );
  OR2_X1 U12747 ( .A1(n13399), .A2(n9955), .ZN(n9954) );
  NAND2_X1 U12748 ( .A1(n14136), .A2(n9728), .ZN(n9960) );
  NAND2_X1 U12749 ( .A1(n14135), .A2(n9730), .ZN(n9961) );
  NAND3_X1 U12750 ( .A1(n14138), .A2(n14137), .A3(n10222), .ZN(n9962) );
  AOI21_X2 U12751 ( .B1(n10220), .B2(n9966), .A(n9694), .ZN(n15191) );
  NOR2_X2 U12752 ( .A1(n10613), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10278) );
  AOI21_X2 U12753 ( .B1(n10472), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10461), .ZN(n10193) );
  NAND2_X2 U12754 ( .A1(n9978), .A2(n9977), .ZN(n14929) );
  AND2_X2 U12755 ( .A1(n10412), .A2(n13023), .ZN(n10265) );
  OR2_X2 U12756 ( .A1(n10373), .A2(n10372), .ZN(n13023) );
  INV_X1 U12757 ( .A(n17284), .ZN(n17287) );
  INV_X2 U12758 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18841) );
  NAND4_X1 U12759 ( .A1(n10003), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(
        n17365) );
  NAND2_X1 U12760 ( .A1(n12405), .A2(n10006), .ZN(n10005) );
  NAND3_X1 U12761 ( .A1(n10005), .A2(n12408), .A3(n10004), .ZN(n12410) );
  NAND2_X1 U12762 ( .A1(n12405), .A2(n10010), .ZN(n10031) );
  NOR2_X1 U12763 ( .A1(n12392), .A2(n10010), .ZN(n10009) );
  NOR2_X2 U12764 ( .A1(n17677), .A2(n10011), .ZN(n12404) );
  NAND3_X1 U12765 ( .A1(n12333), .A2(n10014), .A3(n9731), .ZN(n10013) );
  INV_X2 U12766 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18852) );
  NOR2_X2 U12767 ( .A1(n14369), .A2(n14056), .ZN(n14358) );
  NAND2_X1 U12768 ( .A1(n13170), .A2(n10016), .ZN(n13173) );
  INV_X1 U12769 ( .A(n10017), .ZN(n10016) );
  NAND2_X1 U12770 ( .A1(n10027), .A2(n9732), .ZN(n13782) );
  NAND2_X1 U12771 ( .A1(n15843), .A2(n10031), .ZN(n15844) );
  NOR2_X2 U12773 ( .A1(n16413), .A2(n15846), .ZN(n12407) );
  AND2_X2 U12774 ( .A1(n12322), .A2(n12321), .ZN(n12535) );
  NAND2_X1 U12775 ( .A1(n10037), .A2(n10033), .ZN(P3_U2641) );
  NAND2_X1 U12776 ( .A1(n10038), .A2(n18736), .ZN(n10037) );
  XNOR2_X1 U12777 ( .A(n10039), .B(n16567), .ZN(n10038) );
  NOR2_X1 U12778 ( .A1(n16575), .A2(n16860), .ZN(n10039) );
  INV_X1 U12779 ( .A(n10051), .ZN(n16593) );
  NAND3_X4 U12780 ( .A1(n10060), .A2(n10058), .A3(n10057), .ZN(n10056) );
  INV_X1 U12781 ( .A(n17681), .ZN(n10066) );
  NAND2_X1 U12782 ( .A1(n10066), .A2(n10067), .ZN(n17609) );
  NOR2_X1 U12783 ( .A1(n11432), .A2(n10069), .ZN(n12052) );
  OAI21_X1 U12784 ( .B1(n11400), .B2(n10069), .A(n11399), .ZN(n11417) );
  OAI21_X1 U12785 ( .B1(n16294), .B2(n13680), .A(n10077), .ZN(n19217) );
  NAND2_X1 U12786 ( .A1(n11918), .A2(n10087), .ZN(n10084) );
  NAND2_X1 U12787 ( .A1(n10084), .A2(n11921), .ZN(n10085) );
  AND2_X1 U12788 ( .A1(n15058), .A2(n10096), .ZN(n12020) );
  NAND2_X1 U12789 ( .A1(n15058), .A2(n10097), .ZN(n14958) );
  NAND2_X1 U12790 ( .A1(n15058), .A2(n12665), .ZN(n14983) );
  NAND2_X1 U12791 ( .A1(n15764), .A2(n9689), .ZN(n12683) );
  NAND2_X1 U12792 ( .A1(n10109), .A2(n10111), .ZN(n15777) );
  NAND2_X1 U12793 ( .A1(n18933), .A2(n9755), .ZN(n10109) );
  NAND2_X1 U12794 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10113), .ZN(
        n12616) );
  NAND3_X1 U12795 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12618) );
  INV_X1 U12796 ( .A(n12612), .ZN(n10114) );
  NAND2_X1 U12797 ( .A1(n10114), .A2(n10115), .ZN(n12611) );
  NAND2_X1 U12798 ( .A1(n12597), .A2(n10122), .ZN(n14952) );
  INV_X1 U12799 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10125) );
  AND3_X4 U12800 ( .A1(n11846), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        n13812), .ZN(n11829) );
  INV_X1 U12801 ( .A(n10136), .ZN(n13688) );
  NOR2_X2 U12802 ( .A1(n11543), .A2(n11376), .ZN(n11621) );
  INV_X1 U12803 ( .A(n11543), .ZN(n10149) );
  NAND2_X1 U12804 ( .A1(n14156), .A2(n9751), .ZN(n14148) );
  INV_X1 U12805 ( .A(n10159), .ZN(n14106) );
  NAND2_X1 U12806 ( .A1(n12650), .A2(n10160), .ZN(n14222) );
  NAND2_X1 U12807 ( .A1(n9733), .A2(n10164), .ZN(n15159) );
  NOR3_X1 U12808 ( .A1(n14227), .A2(n14949), .A3(n14226), .ZN(n15156) );
  NAND3_X1 U12809 ( .A1(n10169), .A2(n10168), .A3(n15153), .ZN(n10167) );
  OAI21_X2 U12810 ( .B1(n10595), .B2(n10594), .A(n10468), .ZN(n10586) );
  NAND2_X1 U12811 ( .A1(n10517), .A2(n10610), .ZN(n10619) );
  NAND3_X1 U12812 ( .A1(n11158), .A2(n11209), .A3(n11225), .ZN(n11215) );
  NAND2_X2 U12813 ( .A1(n11158), .A2(n11161), .ZN(n11236) );
  NAND2_X1 U12814 ( .A1(n10603), .A2(n16039), .ZN(n10173) );
  OAI21_X1 U12815 ( .B1(n9664), .B2(n10176), .A(n10174), .ZN(n10459) );
  NAND2_X1 U12816 ( .A1(n11270), .A2(n10185), .ZN(n10184) );
  NAND3_X1 U12817 ( .A1(n10184), .A2(n10182), .A3(n10181), .ZN(n11262) );
  XNOR2_X2 U12818 ( .A(n10193), .B(n9717), .ZN(n20291) );
  NAND2_X1 U12819 ( .A1(n13980), .A2(n13990), .ZN(n10199) );
  NAND2_X1 U12820 ( .A1(n10199), .A2(n10195), .ZN(n14430) );
  CLKBUF_X1 U12821 ( .A(n10199), .Z(n10194) );
  NOR2_X1 U12822 ( .A1(n14329), .A2(n14330), .ZN(n14316) );
  OAI21_X1 U12823 ( .B1(n15310), .B2(n16273), .A(n9720), .ZN(P2_U3015) );
  NAND3_X1 U12824 ( .A1(n10220), .A2(n14225), .A3(n10218), .ZN(n14229) );
  NAND2_X1 U12825 ( .A1(n11499), .A2(n10228), .ZN(n10226) );
  NAND2_X1 U12826 ( .A1(n11499), .A2(n11498), .ZN(n10227) );
  NOR2_X1 U12827 ( .A1(n11500), .A2(n10229), .ZN(n10228) );
  INV_X1 U12828 ( .A(n11498), .ZN(n10229) );
  NOR2_X1 U12829 ( .A1(n10230), .A2(n19986), .ZN(n11477) );
  NAND2_X1 U12830 ( .A1(n11855), .A2(n10230), .ZN(n12634) );
  NOR2_X1 U12831 ( .A1(n10230), .A2(n12655), .ZN(n12656) );
  NOR2_X1 U12832 ( .A1(n10230), .A2(n12667), .ZN(n12668) );
  NOR2_X1 U12833 ( .A1(n11484), .A2(n10230), .ZN(n11459) );
  NOR2_X1 U12834 ( .A1(n16328), .A2(n10230), .ZN(n19971) );
  MUX2_X1 U12835 ( .A(n12848), .B(n12710), .S(n10230), .Z(n12758) );
  MUX2_X1 U12836 ( .A(n13354), .B(n12058), .S(n10230), .Z(n12633) );
  MUX2_X1 U12837 ( .A(n11873), .B(n13679), .S(n12757), .Z(n12639) );
  INV_X1 U12838 ( .A(n10230), .ZN(n12757) );
  NAND2_X1 U12839 ( .A1(n12704), .A2(n10230), .ZN(n11886) );
  NOR2_X4 U12840 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13811) );
  NOR2_X1 U12841 ( .A1(n15085), .A2(n10242), .ZN(n15078) );
  AND2_X1 U12842 ( .A1(n13565), .A2(n14293), .ZN(n12885) );
  NOR2_X2 U12843 ( .A1(n16059), .A2(n16060), .ZN(n16058) );
  OAI211_X1 U12844 ( .C1(n16290), .C2(n16070), .A(n14244), .B(n14243), .ZN(
        n14245) );
  NAND2_X1 U12845 ( .A1(n10409), .A2(n10418), .ZN(n10402) );
  NAND2_X1 U12846 ( .A1(n11426), .A2(n12774), .ZN(n11427) );
  OR2_X2 U12847 ( .A1(n13390), .A2(n13377), .ZN(n19411) );
  INV_X1 U12848 ( .A(n14430), .ZN(n10825) );
  INV_X1 U12849 ( .A(n13244), .ZN(n10608) );
  NAND2_X1 U12850 ( .A1(n11325), .A2(n11376), .ZN(n11332) );
  NAND2_X1 U12851 ( .A1(n11333), .A2(n19305), .ZN(n11542) );
  AND3_X1 U12852 ( .A1(n14206), .A2(n19305), .A3(n9957), .ZN(n11480) );
  NAND2_X1 U12853 ( .A1(n11424), .A2(n11422), .ZN(n11440) );
  NAND2_X1 U12854 ( .A1(n14275), .A2(n10246), .ZN(n11302) );
  AOI22_X1 U12855 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11062), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10340) );
  NOR2_X1 U12856 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10267), .ZN(
        n10268) );
  NOR2_X1 U12857 ( .A1(n20486), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10245) );
  AND2_X1 U12858 ( .A1(n14603), .A2(n20224), .ZN(n10246) );
  INV_X1 U12859 ( .A(n11966), .ZN(n11922) );
  INV_X1 U12860 ( .A(n11922), .ZN(n11962) );
  NOR2_X1 U12861 ( .A1(n16894), .A2(n12270), .ZN(n15623) );
  AND4_X1 U12862 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n10247) );
  OR2_X1 U12863 ( .A1(n15163), .A2(n16236), .ZN(n10248) );
  OR2_X1 U12864 ( .A1(n17663), .A2(n16860), .ZN(n10249) );
  AND2_X1 U12865 ( .A1(n14497), .A2(n14496), .ZN(n10250) );
  INV_X1 U12866 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12751) );
  INV_X1 U12867 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n13115) );
  INV_X1 U12868 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12587) );
  NOR2_X1 U12869 ( .A1(n12587), .A2(n16235), .ZN(n10252) );
  OR2_X1 U12870 ( .A1(n17080), .A2(n17226), .ZN(n10253) );
  AND2_X1 U12871 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10256) );
  AND3_X1 U12872 ( .A1(n14687), .A2(n15835), .A3(n14697), .ZN(n10257) );
  INV_X1 U12873 ( .A(n14615), .ZN(n11252) );
  INV_X1 U12874 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20182) );
  NAND3_X1 U12875 ( .A1(n12019), .A2(n12018), .A3(n12017), .ZN(n10259) );
  INV_X1 U12876 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16213) );
  INV_X1 U12877 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15862) );
  INV_X1 U12878 ( .A(n12108), .ZN(n12179) );
  NOR2_X1 U12879 ( .A1(n18742), .A2(n17886), .ZN(n17624) );
  AND2_X1 U12880 ( .A1(n19287), .A2(n13398), .ZN(n10261) );
  OR3_X1 U12881 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17630), .ZN(n10262) );
  AND4_X1 U12882 ( .A1(n10441), .A2(n10440), .A3(n10439), .A4(n10438), .ZN(
        n10264) );
  INV_X1 U12883 ( .A(n10604), .ZN(n11022) );
  AND2_X1 U12884 ( .A1(n13572), .A2(n13078), .ZN(n10414) );
  NAND2_X1 U12885 ( .A1(n13034), .A2(n10430), .ZN(n10431) );
  OR2_X1 U12886 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11119), .ZN(
        n11117) );
  INV_X1 U12887 ( .A(n10743), .ZN(n10744) );
  OR3_X1 U12888 ( .A1(n11095), .A2(n11143), .A3(n20192), .ZN(n11136) );
  INV_X1 U12889 ( .A(n10415), .ZN(n10405) );
  NAND2_X1 U12890 ( .A1(n10360), .A2(n10359), .ZN(n10361) );
  INV_X1 U12891 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11304) );
  INV_X1 U12892 ( .A(n15223), .ZN(n14223) );
  OR2_X1 U12893 ( .A1(n13671), .A2(n13670), .ZN(n13674) );
  INV_X1 U12894 ( .A(n19988), .ZN(n11415) );
  INV_X1 U12895 ( .A(n10883), .ZN(n10884) );
  INV_X1 U12896 ( .A(n10843), .ZN(n10844) );
  OR2_X1 U12897 ( .A1(n10320), .A2(n10319), .ZN(n11173) );
  NAND2_X1 U12898 ( .A1(n13070), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11159) );
  OR2_X1 U12899 ( .A1(n10539), .A2(n10538), .ZN(n11210) );
  NAND2_X1 U12900 ( .A1(n10436), .A2(n10435), .ZN(n10462) );
  AND2_X1 U12901 ( .A1(n13398), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11333) );
  NOR2_X1 U12902 ( .A1(n14224), .A2(n14223), .ZN(n14225) );
  AND2_X1 U12903 ( .A1(n11846), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11844) );
  NOR2_X1 U12904 ( .A1(n16544), .A2(n15690), .ZN(n12502) );
  AOI21_X1 U12905 ( .B1(n11129), .B2(n11128), .A(n11127), .ZN(n11142) );
  AND2_X1 U12906 ( .A1(n14023), .A2(n14022), .ZN(n15880) );
  AOI22_X1 U12907 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10398) );
  NOR2_X1 U12908 ( .A1(n10984), .A2(n14647), .ZN(n10985) );
  OR2_X1 U12909 ( .A1(n10945), .A2(n14667), .ZN(n10947) );
  AND2_X1 U12910 ( .A1(n10844), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10845) );
  AND2_X1 U12911 ( .A1(n10710), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10734) );
  INV_X1 U12912 ( .A(n13497), .ZN(n10636) );
  NAND2_X1 U12913 ( .A1(n10405), .A2(n10419), .ZN(n13179) );
  NAND2_X1 U12914 ( .A1(n20813), .A2(n16039), .ZN(n10516) );
  AND4_X1 U12915 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12171), .ZN(
        n12207) );
  NAND2_X1 U12916 ( .A1(n11444), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11364) );
  AND3_X1 U12917 ( .A1(n11994), .A2(n11993), .A3(n11992), .ZN(n15411) );
  INV_X1 U12918 ( .A(n14247), .ZN(n14248) );
  INV_X1 U12919 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17063) );
  INV_X1 U12920 ( .A(n17181), .ZN(n12323) );
  INV_X1 U12921 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U12922 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12365) );
  NAND2_X1 U12923 ( .A1(n10786), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10770) );
  AND2_X1 U12924 ( .A1(n14034), .A2(n14033), .ZN(n14432) );
  AND4_X1 U12925 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10401) );
  OR2_X1 U12926 ( .A1(n14635), .A2(n11052), .ZN(n11006) );
  NAND2_X1 U12927 ( .A1(n10885), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10945) );
  OR2_X1 U12928 ( .A1(n14595), .A2(n14459), .ZN(n14497) );
  INV_X1 U12929 ( .A(n11022), .ZN(n10922) );
  NAND2_X1 U12930 ( .A1(n10614), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10621) );
  AND2_X1 U12931 ( .A1(n14020), .A2(n14019), .ZN(n14510) );
  INV_X1 U12932 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11119) );
  AND4_X1 U12933 ( .A1(n10284), .A2(n10283), .A3(n10282), .A4(n10281), .ZN(
        n10285) );
  INV_X1 U12934 ( .A(n20589), .ZN(n20662) );
  NOR2_X1 U12935 ( .A1(n19021), .A2(n15019), .ZN(n14996) );
  INV_X1 U12936 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13827) );
  OR2_X1 U12937 ( .A1(n11555), .A2(n11554), .ZN(n12208) );
  NAND2_X1 U12938 ( .A1(n11536), .A2(n11535), .ZN(n11539) );
  NAND2_X1 U12939 ( .A1(n11311), .A2(n11376), .ZN(n11318) );
  NOR2_X1 U12940 ( .A1(n12167), .A2(n12166), .ZN(n13888) );
  AOI21_X1 U12941 ( .B1(n16187), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15329), .ZN(n15200) );
  OR2_X1 U12942 ( .A1(n15316), .A2(n15315), .ZN(n15317) );
  INV_X1 U12943 ( .A(n15293), .ZN(n14145) );
  AND2_X1 U12944 ( .A1(n12234), .A2(n12233), .ZN(n13964) );
  AND3_X1 U12945 ( .A1(n11954), .A2(n11953), .A3(n11952), .ZN(n15032) );
  AND2_X1 U12946 ( .A1(n15532), .A2(n15531), .ZN(n15551) );
  NAND2_X1 U12947 ( .A1(n11494), .A2(n19979), .ZN(n11531) );
  INV_X1 U12948 ( .A(n13866), .ZN(n19704) );
  AND2_X1 U12949 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11495), .ZN(
        n11529) );
  NOR2_X1 U12950 ( .A1(n17813), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17675) );
  NOR2_X1 U12951 ( .A1(n17773), .A2(n18053), .ZN(n17730) );
  INV_X1 U12952 ( .A(n12392), .ZN(n17791) );
  OAI211_X1 U12953 ( .C1(n17190), .C2(n17257), .A(n12468), .B(n12467), .ZN(
        n12528) );
  NAND2_X1 U12954 ( .A1(n11028), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11080) );
  OR2_X1 U12955 ( .A1(n14417), .A2(n14284), .ZN(n14351) );
  NAND2_X1 U12956 ( .A1(n10805), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10843) );
  INV_X1 U12957 ( .A(n15910), .ZN(n14439) );
  NAND2_X1 U12958 ( .A1(n10503), .A2(n10502), .ZN(n20325) );
  INV_X1 U12959 ( .A(n20051), .ZN(n20075) );
  OR2_X1 U12960 ( .A1(n14710), .A2(n11052), .ZN(n10823) );
  AND3_X1 U12961 ( .A1(n10709), .A2(n10708), .A3(n10707), .ZN(n13991) );
  INV_X1 U12962 ( .A(n14431), .ZN(n10824) );
  INV_X1 U12963 ( .A(n11052), .ZN(n13559) );
  INV_X1 U12964 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15912) );
  INV_X1 U12965 ( .A(n20168), .ZN(n14916) );
  AND2_X1 U12966 ( .A1(n13596), .A2(n13595), .ZN(n16024) );
  OR2_X1 U12967 ( .A1(n13091), .A2(n13088), .ZN(n20168) );
  OR2_X1 U12968 ( .A1(n13091), .A2(n13074), .ZN(n20173) );
  OAI21_X1 U12969 ( .B1(n15828), .B2(n20726), .A(n20801), .ZN(n13521) );
  INV_X1 U12970 ( .A(n13325), .ZN(n15798) );
  INV_X1 U12971 ( .A(n13507), .ZN(n13509) );
  OR2_X1 U12972 ( .A1(n20408), .A2(n20594), .ZN(n20376) );
  INV_X1 U12973 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20519) );
  NOR2_X1 U12974 ( .A1(n20488), .A2(n20330), .ZN(n20631) );
  AOI21_X1 U12975 ( .B1(n20588), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20330), 
        .ZN(n20670) );
  OR2_X1 U12976 ( .A1(n13322), .A2(n13321), .ZN(n15814) );
  NAND2_X1 U12977 ( .A1(n11891), .A2(n11890), .ZN(n12705) );
  NOR2_X1 U12978 ( .A1(n19021), .A2(n14956), .ZN(n14980) );
  OR2_X1 U12979 ( .A1(n19169), .A2(n12065), .ZN(n15131) );
  AND3_X1 U12980 ( .A1(n11989), .A2(n11988), .A3(n11987), .ZN(n12685) );
  AND2_X1 U12981 ( .A1(n15281), .A2(n14169), .ZN(n15762) );
  OR2_X1 U12982 ( .A1(n19043), .A2(n14130), .ZN(n16203) );
  INV_X1 U12983 ( .A(n19248), .ZN(n16277) );
  NOR2_X1 U12984 ( .A1(n12738), .A2(n12055), .ZN(n16320) );
  NAND2_X1 U12985 ( .A1(n15860), .A2(n15859), .ZN(n15861) );
  NAND2_X1 U12986 ( .A1(n19566), .A2(n19536), .ZN(n19512) );
  INV_X1 U12987 ( .A(n19932), .ZN(n19634) );
  INV_X1 U12988 ( .A(n13398), .ZN(n19282) );
  AOI21_X1 U12989 ( .B1(n16725), .B2(n16861), .A(n16860), .ZN(n16715) );
  NOR2_X1 U12990 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16746), .ZN(n16733) );
  INV_X1 U12991 ( .A(n16905), .ZN(n16891) );
  NAND2_X1 U12992 ( .A1(n18899), .A2(n17428), .ZN(n16542) );
  NOR3_X1 U12993 ( .A1(n12531), .A2(n12519), .A3(n18668), .ZN(n15714) );
  INV_X1 U12994 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17123) );
  INV_X1 U12995 ( .A(n17412), .ZN(n17384) );
  INV_X1 U12996 ( .A(n12570), .ZN(n17753) );
  NOR2_X1 U12997 ( .A1(n17729), .A2(n18048), .ZN(n18035) );
  NOR2_X1 U12998 ( .A1(n18126), .A2(n17979), .ZN(n18027) );
  NOR2_X1 U12999 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17765), .ZN(
        n17750) );
  INV_X1 U13000 ( .A(n17940), .ZN(n18092) );
  INV_X1 U13001 ( .A(n12389), .ZN(n12387) );
  AOI211_X1 U13002 ( .C1(n15734), .C2(n18712), .A(n15733), .B(n15732), .ZN(
        n15738) );
  NOR2_X1 U13003 ( .A1(n12368), .A2(n12367), .ZN(n12369) );
  INV_X1 U13004 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18693) );
  OR2_X1 U13005 ( .A1(n18574), .A2(n18518), .ZN(n18519) );
  INV_X1 U13006 ( .A(n12501), .ZN(n17468) );
  OR2_X1 U13007 ( .A1(n12827), .A2(n20001), .ZN(n12882) );
  OR2_X1 U13008 ( .A1(n20809), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12894) );
  NOR2_X1 U13009 ( .A1(n15908), .A2(n14282), .ZN(n15875) );
  OR2_X1 U13010 ( .A1(n20042), .A2(n20041), .ZN(n15910) );
  INV_X1 U13011 ( .A(n15914), .ZN(n20055) );
  AND2_X1 U13012 ( .A1(n13583), .A2(n13582), .ZN(n20042) );
  INV_X1 U13013 ( .A(n14568), .ZN(n14589) );
  INV_X1 U13014 ( .A(n14603), .ZN(n14569) );
  INV_X2 U13015 ( .A(n13194), .ZN(n20161) );
  AOI21_X1 U13016 ( .B1(n14461), .B2(n14593), .A(n14460), .ZN(n14737) );
  AND2_X1 U13017 ( .A1(n20007), .A2(n11153), .ZN(n15948) );
  INV_X1 U13018 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13588) );
  INV_X1 U13019 ( .A(n20007), .ZN(n15959) );
  AND2_X1 U13020 ( .A1(n14806), .A2(n14086), .ZN(n14786) );
  NOR2_X1 U13021 ( .A1(n14880), .A2(n14697), .ZN(n15836) );
  NOR3_X1 U13022 ( .A1(n15972), .A2(n16000), .A3(n14907), .ZN(n15991) );
  OR2_X1 U13023 ( .A1(n13350), .A2(n13349), .ZN(n14913) );
  INV_X1 U13024 ( .A(n14890), .ZN(n13349) );
  INV_X1 U13025 ( .A(n20233), .ZN(n20257) );
  NAND2_X1 U13026 ( .A1(n20812), .A2(n13509), .ZN(n20302) );
  NOR2_X2 U13027 ( .A1(n20302), .A2(n20623), .ZN(n20318) );
  NOR2_X2 U13028 ( .A1(n20302), .A2(n20516), .ZN(n20348) );
  INV_X1 U13029 ( .A(n20376), .ZN(n20399) );
  NAND2_X1 U13030 ( .A1(n13507), .A2(n20323), .ZN(n20408) );
  INV_X1 U13031 ( .A(n20548), .ZN(n20430) );
  INV_X1 U13032 ( .A(n20495), .ZN(n20512) );
  NOR2_X2 U13033 ( .A1(n20819), .A2(n20623), .ZN(n20544) );
  INV_X1 U13034 ( .A(n20558), .ZN(n20582) );
  OR2_X1 U13035 ( .A1(n9656), .A2(n13510), .ZN(n20548) );
  INV_X1 U13036 ( .A(n20248), .ZN(n20696) );
  INV_X1 U13037 ( .A(n20713), .ZN(n20720) );
  OR2_X1 U13038 ( .A1(n13073), .A2(n15853), .ZN(n15820) );
  INV_X1 U13039 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20739) );
  NOR2_X1 U13041 ( .A1(n19851), .A2(n9634), .ZN(n19009) );
  OR2_X1 U13042 ( .A1(n18906), .A2(n12659), .ZN(n19067) );
  INV_X1 U13043 ( .A(n19067), .ZN(n19102) );
  NOR2_X1 U13044 ( .A1(n16322), .A2(n12770), .ZN(n12693) );
  NOR2_X1 U13045 ( .A1(n11576), .A2(n11575), .ZN(n19133) );
  OAI211_X1 U13046 ( .C1(n15167), .C2(n16251), .A(n10248), .B(n15166), .ZN(
        n15168) );
  AND2_X1 U13047 ( .A1(n19231), .A2(n12854), .ZN(n19216) );
  AND2_X1 U13048 ( .A1(n12919), .A2(n12763), .ZN(n19227) );
  NOR2_X1 U13049 ( .A1(n15567), .A2(n16281), .ZN(n15540) );
  AND2_X1 U13050 ( .A1(n15041), .A2(n15040), .ZN(n19156) );
  AND2_X1 U13051 ( .A1(n12954), .A2(n16320), .ZN(n19245) );
  AND2_X1 U13052 ( .A1(n12954), .A2(n12940), .ZN(n19253) );
  OAI21_X1 U13053 ( .B1(n19278), .B2(n19311), .A(n19781), .ZN(n19315) );
  INV_X1 U13054 ( .A(n19345), .ZN(n19337) );
  AND2_X1 U13055 ( .A1(n19468), .A2(n19932), .ZN(n19395) );
  NOR2_X1 U13056 ( .A1(n19413), .A2(n19706), .ZN(n19460) );
  AND2_X1 U13057 ( .A1(n19566), .A2(n19961), .ZN(n19468) );
  INV_X1 U13058 ( .A(n19489), .ZN(n19532) );
  NOR2_X1 U13059 ( .A1(n19512), .A2(n19511), .ZN(n19561) );
  INV_X1 U13060 ( .A(n19588), .ZN(n19601) );
  AND2_X1 U13061 ( .A1(n19645), .A2(n19643), .ZN(n19665) );
  NOR2_X1 U13062 ( .A1(n19670), .A2(n19706), .ZN(n19734) );
  INV_X1 U13063 ( .A(n19822), .ZN(n19757) );
  AND2_X1 U13064 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11900), .ZN(n16345) );
  INV_X1 U13065 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18904) );
  INV_X1 U13066 ( .A(n12424), .ZN(n18708) );
  INV_X1 U13067 ( .A(n16904), .ZN(n16896) );
  NOR2_X1 U13068 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16676), .ZN(n16665) );
  NAND2_X1 U13069 ( .A1(n16698), .A2(n10249), .ZN(n16684) );
  NOR2_X1 U13070 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16796), .ZN(n16778) );
  INV_X1 U13071 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18727) );
  NOR2_X2 U13072 ( .A1(n18833), .A2(n16899), .ZN(n16889) );
  NOR2_X1 U13073 ( .A1(n17011), .A2(n17015), .ZN(n16983) );
  NOR2_X1 U13074 ( .A1(n17059), .A2(n17058), .ZN(n17057) );
  INV_X1 U13075 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17240) );
  AOI21_X1 U13076 ( .B1(n15714), .B2(n18708), .A(n15691), .ZN(n15863) );
  NAND2_X1 U13077 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17301), .ZN(n17296) );
  INV_X1 U13078 ( .A(n17337), .ZN(n17345) );
  INV_X2 U13079 ( .A(n17080), .ZN(n17210) );
  OAI211_X1 U13080 ( .C1(n17190), .C2(n17214), .A(n12448), .B(n12447), .ZN(
        n17428) );
  NOR2_X1 U13081 ( .A1(n18210), .A2(n18215), .ZN(n18084) );
  NAND2_X1 U13082 ( .A1(n18735), .A2(n18235), .ZN(n18518) );
  INV_X1 U13083 ( .A(n18846), .ZN(n18860) );
  INV_X1 U13084 ( .A(n18374), .ZN(n18376) );
  INV_X1 U13085 ( .A(n18563), .ZN(n18569) );
  INV_X1 U13086 ( .A(n18519), .ZN(n18548) );
  OR3_X1 U13087 ( .A1(n13126), .A2(n12752), .A3(n20001), .ZN(n13036) );
  NAND2_X1 U13088 ( .A1(n13568), .A2(n13566), .ZN(n15914) );
  OR2_X1 U13089 ( .A1(n11299), .A2(n14535), .ZN(n14568) );
  OR2_X1 U13090 ( .A1(n10250), .A2(n14498), .ZN(n15935) );
  AND2_X2 U13091 ( .A1(n11287), .A2(n13064), .ZN(n14603) );
  INV_X1 U13092 ( .A(n20104), .ZN(n20132) );
  NOR2_X1 U13093 ( .A1(n13036), .A2(n13035), .ZN(n13224) );
  AND2_X1 U13094 ( .A1(n15943), .A2(n15942), .ZN(n15993) );
  OR2_X1 U13095 ( .A1(n15948), .A2(n13261), .ZN(n15963) );
  OR3_X1 U13096 ( .A1(n15966), .A2(n14075), .A3(n14889), .ZN(n14880) );
  OR2_X1 U13097 ( .A1(n13091), .A2(n13069), .ZN(n20164) );
  OR2_X1 U13098 ( .A1(n20302), .A2(n20594), .ZN(n20262) );
  AOI22_X1 U13099 ( .A1(n20264), .A2(n20268), .B1(n20488), .B2(n10245), .ZN(
        n20289) );
  NAND2_X1 U13100 ( .A1(n20324), .A2(n20430), .ZN(n20375) );
  AOI22_X1 U13101 ( .A1(n20381), .A2(n20378), .B1(n10245), .B2(n20552), .ZN(
        n20403) );
  OR2_X1 U13102 ( .A1(n20408), .A2(n20516), .ZN(n20434) );
  NAND2_X1 U13103 ( .A1(n20518), .A2(n20430), .ZN(n20482) );
  AOI22_X1 U13104 ( .A1(n20494), .A2(n20490), .B1(n20488), .B2(n20487), .ZN(
        n20515) );
  NAND2_X1 U13105 ( .A1(n20518), .A2(n20517), .ZN(n20558) );
  AOI22_X1 U13106 ( .A1(n20556), .A2(n20553), .B1(n20552), .B2(n20551), .ZN(
        n20587) );
  OR2_X1 U13107 ( .A1(n20624), .A2(n20548), .ZN(n20621) );
  OR2_X1 U13108 ( .A1(n20624), .A2(n20623), .ZN(n20713) );
  INV_X1 U13109 ( .A(n20794), .ZN(n20730) );
  OR2_X1 U13110 ( .A1(n12660), .A2(n12942), .ZN(n12715) );
  INV_X1 U13111 ( .A(n19096), .ZN(n19082) );
  AND2_X2 U13112 ( .A1(n11901), .A2(n16345), .ZN(n19148) );
  OR2_X1 U13113 ( .A1(n19169), .A2(n11479), .ZN(n16120) );
  INV_X1 U13114 ( .A(n19169), .ZN(n15130) );
  NOR2_X1 U13115 ( .A1(n19173), .A2(n19150), .ZN(n19179) );
  NOR2_X1 U13116 ( .A1(n19180), .A2(n19212), .ZN(n19198) );
  INV_X1 U13117 ( .A(n19180), .ZN(n19214) );
  OR2_X1 U13118 ( .A1(n12715), .A2(n13398), .ZN(n12881) );
  INV_X1 U13119 ( .A(n19216), .ZN(n16236) );
  INV_X1 U13120 ( .A(n19250), .ZN(n16292) );
  NAND2_X1 U13121 ( .A1(n19567), .A2(n19468), .ZN(n19345) );
  INV_X1 U13122 ( .A(n19367), .ZN(n19375) );
  INV_X1 U13123 ( .A(n19395), .ZN(n19405) );
  INV_X1 U13124 ( .A(n19430), .ZN(n19438) );
  INV_X1 U13125 ( .A(n19460), .ZN(n19467) );
  INV_X1 U13126 ( .A(n19486), .ZN(n19499) );
  AND2_X1 U13127 ( .A1(n19507), .A2(n19506), .ZN(n19526) );
  INV_X1 U13128 ( .A(n19561), .ZN(n19557) );
  AND2_X1 U13129 ( .A1(n19575), .A2(n19574), .ZN(n19588) );
  NAND2_X1 U13130 ( .A1(n19738), .A2(n19567), .ZN(n19604) );
  INV_X1 U13131 ( .A(n19630), .ZN(n19625) );
  NAND2_X1 U13132 ( .A1(n19738), .A2(n19932), .ZN(n19663) );
  INV_X1 U13133 ( .A(n19734), .ZN(n19729) );
  INV_X1 U13134 ( .A(n19825), .ZN(n19764) );
  NAND2_X1 U13135 ( .A1(n19777), .A2(n19713), .ZN(n19829) );
  INV_X1 U13136 ( .A(n19931), .ZN(n19928) );
  OR2_X1 U13137 ( .A1(n16892), .A2(n16645), .ZN(n16663) );
  NOR2_X1 U13138 ( .A1(n16623), .A2(n16966), .ZN(n16971) );
  AND2_X1 U13139 ( .A1(n17269), .A2(n17365), .ZN(n17266) );
  INV_X2 U13140 ( .A(n17266), .ZN(n17256) );
  INV_X1 U13141 ( .A(n17266), .ZN(n17260) );
  INV_X1 U13142 ( .A(n17349), .ZN(n17322) );
  NOR2_X1 U13143 ( .A1(n17517), .A2(n17383), .ZN(n17388) );
  INV_X1 U13144 ( .A(n17419), .ZN(n17414) );
  INV_X1 U13145 ( .A(n17446), .ZN(n17465) );
  INV_X1 U13146 ( .A(n17815), .ZN(n17744) );
  INV_X1 U13147 ( .A(n17814), .ZN(n17789) );
  INV_X1 U13148 ( .A(n18133), .ZN(n18111) );
  INV_X1 U13149 ( .A(n18084), .ZN(n18205) );
  INV_X1 U13150 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18698) );
  INV_X1 U13151 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18833) );
  INV_X1 U13152 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18758) );
  OAI21_X1 U13153 ( .B1(n12027), .B2(n12024), .A(n12023), .ZN(P2_U2858) );
  INV_X1 U13154 ( .A(n12581), .ZN(P3_U2799) );
  AND2_X4 U13155 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13307) );
  AOI22_X1 U13156 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10274) );
  INV_X2 U13157 ( .A(n10893), .ZN(n10865) );
  NOR2_X1 U13158 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13159 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10273) );
  INV_X1 U13160 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U13161 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10272) );
  AND2_X2 U13162 ( .A1(n13177), .A2(n10269), .ZN(n10367) );
  NOR2_X1 U13163 ( .A1(n10613), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10270) );
  AOI22_X1 U13164 ( .A1(n10367), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10271) );
  AND2_X4 U13165 ( .A1(n13302), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10397) );
  AND2_X4 U13166 ( .A1(n13302), .A2(n10613), .ZN(n10396) );
  INV_X1 U13167 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13168 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9652), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10284) );
  INV_X2 U13169 ( .A(n10890), .ZN(n10543) );
  AOI22_X1 U13170 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U13171 ( .A1(n10330), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10282) );
  NAND2_X1 U13172 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10281) );
  AND3_X4 U13173 ( .A1(n10287), .A2(n10286), .A3(n10285), .ZN(n20184) );
  AOI22_X1 U13174 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9647), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10291) );
  INV_X2 U13175 ( .A(n10893), .ZN(n11062) );
  AOI22_X1 U13176 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13177 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13178 ( .A1(n10367), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13179 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10391), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U13180 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10294) );
  NAND2_X1 U13181 ( .A1(n10330), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10293) );
  NAND2_X1 U13182 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10292) );
  NAND4_X1 U13183 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10298) );
  AOI22_X1 U13184 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10296) );
  INV_X1 U13185 ( .A(n10296), .ZN(n10297) );
  INV_X1 U13186 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10323) );
  INV_X1 U13187 ( .A(n10397), .ZN(n10900) );
  AOI22_X1 U13188 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10396), .B1(
        n10397), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13189 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11032), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13190 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13191 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10301) );
  NAND4_X1 U13192 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10310) );
  AOI22_X1 U13193 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n9644), .B1(
        n11062), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13194 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13195 ( .A1(n10949), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13196 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10305) );
  NAND4_X1 U13197 ( .A1(n10308), .A2(n10307), .A3(n10306), .A4(n10305), .ZN(
        n10309) );
  OR2_X1 U13198 ( .A1(n11159), .A2(n11222), .ZN(n10322) );
  AOI22_X1 U13199 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13200 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10313) );
  INV_X2 U13201 ( .A(n10744), .ZN(n10913) );
  AOI22_X1 U13202 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13204 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10311) );
  NAND4_X1 U13205 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10320) );
  AOI22_X1 U13206 ( .A1(n10949), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U13207 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13208 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13209 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10315) );
  NAND4_X1 U13210 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10319) );
  NAND2_X1 U13211 ( .A1(n12898), .A2(n11173), .ZN(n10321) );
  OAI211_X1 U13212 ( .C1(n11130), .C2(n10323), .A(n10322), .B(n10321), .ZN(
        n10455) );
  INV_X1 U13213 ( .A(n11159), .ZN(n10466) );
  NAND2_X1 U13214 ( .A1(n10466), .A2(n11222), .ZN(n10456) );
  INV_X1 U13215 ( .A(n10456), .ZN(n10324) );
  AOI22_X1 U13216 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13217 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13218 ( .A1(n10548), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13219 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10325) );
  NAND4_X1 U13220 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10336) );
  AOI22_X1 U13221 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13222 ( .A1(n10330), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13223 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13224 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10391), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10331) );
  NAND4_X1 U13225 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10335) );
  AOI22_X1 U13226 ( .A1(n10548), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U13227 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13228 ( .A1(n10367), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10337) );
  NAND4_X1 U13229 ( .A1(n10340), .A2(n10339), .A3(n10338), .A4(n10337), .ZN(
        n10346) );
  AOI22_X1 U13230 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13231 ( .A1(n11056), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13232 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13233 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10341) );
  NAND4_X1 U13234 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10345) );
  AOI22_X1 U13235 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10548), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13236 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13237 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13238 ( .A1(n10367), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13239 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13240 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10391), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13241 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U13242 ( .A1(n10330), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10353) );
  NAND2_X1 U13243 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10352) );
  AND4_X1 U13244 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n10356) );
  AOI22_X1 U13246 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13247 ( .A1(n11056), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13248 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13249 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U13250 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n10373) );
  AOI22_X1 U13251 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13252 ( .A1(n10367), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13253 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13254 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10368) );
  NAND4_X1 U13255 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        n10372) );
  NAND2_X1 U13256 ( .A1(n10415), .A2(n13023), .ZN(n10434) );
  AOI22_X1 U13257 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13258 ( .A1(n10330), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10329), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13259 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U13260 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10374) );
  NAND4_X1 U13261 ( .A1(n10377), .A2(n10376), .A3(n10375), .A4(n10374), .ZN(
        n10383) );
  AOI22_X1 U13262 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11062), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13263 ( .A1(n10548), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13264 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13265 ( .A1(n11013), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10378) );
  NAND4_X1 U13266 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10382) );
  OR2_X2 U13267 ( .A1(n10383), .A2(n10382), .ZN(n14525) );
  INV_X2 U13268 ( .A(n13522), .ZN(n10423) );
  NAND2_X1 U13269 ( .A1(n14525), .A2(n13536), .ZN(n10418) );
  NAND2_X1 U13270 ( .A1(n13076), .A2(n20184), .ZN(n10386) );
  AOI22_X1 U13271 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13272 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13273 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13274 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13275 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U13276 ( .A1(n10391), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U13277 ( .A1(n10330), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10393) );
  NAND2_X1 U13278 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10392) );
  INV_X2 U13279 ( .A(n10412), .ZN(n20192) );
  INV_X1 U13280 ( .A(n10402), .ZN(n10403) );
  AND2_X2 U13281 ( .A1(n10359), .A2(n13023), .ZN(n13080) );
  NAND2_X1 U13282 ( .A1(n10403), .A2(n13080), .ZN(n10407) );
  NAND2_X1 U13283 ( .A1(n20213), .A2(n10423), .ZN(n10404) );
  XNOR2_X1 U13284 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12829) );
  INV_X1 U13285 ( .A(n13023), .ZN(n20205) );
  INV_X1 U13286 ( .A(n13098), .ZN(n10410) );
  OAI21_X1 U13287 ( .B1(n12752), .B2(n12829), .A(n13066), .ZN(n10411) );
  NAND2_X1 U13288 ( .A1(n20184), .A2(n10412), .ZN(n13572) );
  NAND2_X1 U13289 ( .A1(n13581), .A2(n13122), .ZN(n13078) );
  NAND2_X1 U13290 ( .A1(n13034), .A2(n13536), .ZN(n10413) );
  NAND2_X1 U13291 ( .A1(n10415), .A2(n13070), .ZN(n10417) );
  INV_X1 U13292 ( .A(n10416), .ZN(n10430) );
  INV_X1 U13293 ( .A(n10418), .ZN(n10419) );
  NAND2_X1 U13294 ( .A1(n13058), .A2(n13179), .ZN(n10426) );
  INV_X1 U13295 ( .A(n15822), .ZN(n15818) );
  NAND2_X1 U13296 ( .A1(n15823), .A2(n13115), .ZN(n20809) );
  INV_X1 U13297 ( .A(n12894), .ZN(n10477) );
  MUX2_X1 U13298 ( .A(n15818), .B(n10477), .S(n20588), .Z(n10420) );
  INV_X1 U13299 ( .A(n10420), .ZN(n10421) );
  OR2_X1 U13300 ( .A1(n13304), .A2(n10423), .ZN(n13085) );
  OR2_X1 U13301 ( .A1(n20809), .A2(n16039), .ZN(n20004) );
  INV_X1 U13302 ( .A(n20004), .ZN(n10424) );
  NAND2_X1 U13303 ( .A1(n13085), .A2(n10424), .ZN(n10425) );
  NOR2_X1 U13304 ( .A1(n9721), .A2(n10425), .ZN(n10436) );
  INV_X1 U13305 ( .A(n10426), .ZN(n10427) );
  NAND2_X1 U13306 ( .A1(n10427), .A2(n10412), .ZN(n10432) );
  INV_X1 U13307 ( .A(n13565), .ZN(n10428) );
  NAND2_X1 U13308 ( .A1(n10429), .A2(n10428), .ZN(n13082) );
  NAND3_X1 U13309 ( .A1(n10432), .A2(n13082), .A3(n10431), .ZN(n10433) );
  INV_X1 U13310 ( .A(n10462), .ZN(n10437) );
  AOI22_X1 U13311 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13312 ( .A1(n10949), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11062), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13313 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13314 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13315 ( .A1(n10743), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13316 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10444) );
  NAND2_X1 U13317 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10443) );
  NAND2_X1 U13318 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10442) );
  AND4_X1 U13319 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10447) );
  AOI22_X1 U13320 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10446) );
  XNOR2_X1 U13321 ( .A(n11164), .B(n11222), .ZN(n10448) );
  NAND2_X1 U13322 ( .A1(n10448), .A2(n10466), .ZN(n10449) );
  INV_X1 U13323 ( .A(n10602), .ZN(n10450) );
  INV_X1 U13324 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20189) );
  INV_X1 U13325 ( .A(n11222), .ZN(n11231) );
  INV_X1 U13326 ( .A(n11164), .ZN(n11174) );
  NAND2_X1 U13327 ( .A1(n20184), .A2(n11174), .ZN(n10451) );
  OAI211_X1 U13328 ( .C1(n11231), .C2(n13536), .A(n10451), .B(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n10452) );
  INV_X1 U13329 ( .A(n10452), .ZN(n10453) );
  AND2_X1 U13330 ( .A1(n10601), .A2(n10455), .ZN(n10454) );
  INV_X1 U13331 ( .A(n10455), .ZN(n10457) );
  NAND2_X1 U13332 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10475) );
  OAI21_X1 U13333 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10475), .ZN(n20486) );
  OR2_X1 U13334 ( .A1(n15822), .A2(n20489), .ZN(n10470) );
  OAI21_X1 U13335 ( .B1(n12894), .B2(n20486), .A(n10470), .ZN(n10461) );
  INV_X1 U13336 ( .A(n20291), .ZN(n10465) );
  NAND2_X1 U13337 ( .A1(n10465), .A2(n10464), .ZN(n20234) );
  NAND2_X1 U13338 ( .A1(n10466), .A2(n11173), .ZN(n10467) );
  NAND2_X1 U13339 ( .A1(n10470), .A2(n10469), .ZN(n10471) );
  NAND2_X1 U13340 ( .A1(n9717), .A2(n10471), .ZN(n10481) );
  NAND2_X1 U13341 ( .A1(n10483), .A2(n10481), .ZN(n10479) );
  NOR2_X1 U13342 ( .A1(n15822), .A2(n11119), .ZN(n10473) );
  INV_X1 U13343 ( .A(n10475), .ZN(n10474) );
  NAND2_X1 U13344 ( .A1(n10474), .A2(n11119), .ZN(n20520) );
  NAND2_X1 U13345 ( .A1(n10475), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10476) );
  NAND2_X1 U13346 ( .A1(n20520), .A2(n10476), .ZN(n13516) );
  NAND2_X1 U13347 ( .A1(n10477), .A2(n13516), .ZN(n10480) );
  NAND2_X1 U13348 ( .A1(n10482), .A2(n10480), .ZN(n10478) );
  NAND4_X1 U13349 ( .A1(n10483), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(
        n10484) );
  INV_X1 U13350 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20203) );
  AOI22_X1 U13351 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13352 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10329), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13353 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13354 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9652), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10485) );
  NAND4_X1 U13355 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10494) );
  AOI22_X1 U13356 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13357 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13358 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13359 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10489) );
  NAND4_X1 U13360 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10493) );
  AOI22_X1 U13361 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12898), .B2(n10495), .ZN(n10496) );
  NAND2_X1 U13362 ( .A1(n10498), .A2(n10587), .ZN(n10611) );
  INV_X1 U13363 ( .A(n10611), .ZN(n10517) );
  NAND2_X1 U13364 ( .A1(n10472), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10503) );
  NAND3_X1 U13365 ( .A1(n20519), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20409) );
  INV_X1 U13366 ( .A(n20409), .ZN(n10499) );
  NAND2_X1 U13367 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10499), .ZN(
        n20404) );
  NAND2_X1 U13368 ( .A1(n20519), .A2(n20404), .ZN(n10500) );
  NOR3_X1 U13369 ( .A1(n20519), .A2(n11119), .A3(n20489), .ZN(n20672) );
  NAND2_X1 U13370 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20672), .ZN(
        n20660) );
  NAND2_X1 U13371 ( .A1(n10500), .A2(n20660), .ZN(n20431) );
  OAI22_X1 U13372 ( .A1(n12894), .A2(n20431), .B1(n15822), .B2(n20519), .ZN(
        n10501) );
  INV_X1 U13373 ( .A(n10501), .ZN(n10502) );
  XNOR2_X2 U13374 ( .A(n13145), .B(n20325), .ZN(n20813) );
  INV_X1 U13375 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20211) );
  AOI22_X1 U13376 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13377 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13378 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13379 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9652), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10505) );
  NAND4_X1 U13380 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10514) );
  AOI22_X1 U13381 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13382 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13383 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13384 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10509) );
  NAND4_X1 U13385 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10513) );
  AOI22_X1 U13386 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11133), .B1(
        n11143), .B2(n11186), .ZN(n10515) );
  NAND2_X1 U13387 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10529) );
  AOI22_X1 U13388 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13389 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13390 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13391 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10518) );
  NAND4_X1 U13392 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10527) );
  AOI22_X1 U13393 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13394 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13395 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13396 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10522) );
  NAND4_X1 U13397 ( .A1(n10525), .A2(n10524), .A3(n10523), .A4(n10522), .ZN(
        n10526) );
  NAND2_X1 U13398 ( .A1(n11143), .A2(n11200), .ZN(n10528) );
  NAND2_X1 U13399 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10541) );
  INV_X1 U13400 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20218) );
  AOI22_X1 U13401 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13402 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13403 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13404 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n9652), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10530) );
  NAND4_X1 U13405 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10539) );
  AOI22_X1 U13406 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13407 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13408 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13409 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10534) );
  NAND4_X1 U13410 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10538) );
  NAND2_X1 U13411 ( .A1(n11143), .A2(n11210), .ZN(n10540) );
  NAND2_X1 U13412 ( .A1(n10541), .A2(n10540), .ZN(n10629) );
  NAND2_X1 U13413 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10556) );
  AOI22_X1 U13414 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13415 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13416 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13417 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10544) );
  NAND4_X1 U13418 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n10554) );
  AOI22_X1 U13419 ( .A1(n10949), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13420 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13421 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10865), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13422 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10549) );
  NAND4_X1 U13423 ( .A1(n10552), .A2(n10551), .A3(n10550), .A4(n10549), .ZN(
        n10553) );
  NAND2_X1 U13424 ( .A1(n11143), .A2(n11220), .ZN(n10555) );
  NAND2_X2 U13425 ( .A1(n10558), .A2(n10557), .ZN(n11158) );
  INV_X1 U13426 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10560) );
  NAND2_X1 U13427 ( .A1(n11143), .A2(n11222), .ZN(n10559) );
  OAI21_X1 U13428 ( .B1(n11130), .B2(n10560), .A(n10559), .ZN(n10561) );
  XNOR2_X2 U13429 ( .A(n11158), .B(n10561), .ZN(n11226) );
  NOR2_X2 U13430 ( .A1(n14525), .A2(n20728), .ZN(n10604) );
  INV_X1 U13431 ( .A(n10658), .ZN(n10565) );
  INV_X1 U13432 ( .A(n10563), .ZN(n10643) );
  INV_X1 U13433 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20037) );
  NAND2_X1 U13434 ( .A1(n10643), .A2(n20037), .ZN(n10564) );
  NAND2_X1 U13435 ( .A1(n10565), .A2(n10564), .ZN(n20034) );
  NOR2_X1 U13436 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10632) );
  NAND2_X1 U13437 ( .A1(n20034), .A2(n13559), .ZN(n10567) );
  NAND2_X1 U13438 ( .A1(n11077), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10566) );
  NAND2_X1 U13439 ( .A1(n10567), .A2(n10566), .ZN(n10568) );
  AOI21_X1 U13440 ( .B1(n10922), .B2(P1_EAX_REG_7__SCAN_IN), .A(n10568), .ZN(
        n10569) );
  AOI22_X1 U13441 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13442 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13443 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13444 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10571) );
  NAND4_X1 U13445 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n10581) );
  AOI22_X1 U13446 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13447 ( .A1(n10949), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13448 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13449 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9667), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10576) );
  NAND4_X1 U13450 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n10580) );
  NOR2_X1 U13451 ( .A1(n10581), .A2(n10580), .ZN(n10585) );
  XOR2_X1 U13452 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10658), .Z(n20023) );
  INV_X1 U13453 ( .A(n20023), .ZN(n10582) );
  AOI22_X1 U13454 ( .A1(n11077), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13559), .B2(n10582), .ZN(n10584) );
  NAND2_X1 U13455 ( .A1(n10922), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10583) );
  OAI211_X1 U13456 ( .C1(n9914), .C2(n10585), .A(n10584), .B(n10583), .ZN(
        n13739) );
  NAND2_X1 U13457 ( .A1(n10588), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10626) );
  NAND2_X1 U13458 ( .A1(n10604), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10591) );
  INV_X1 U13459 ( .A(n10614), .ZN(n10589) );
  OAI21_X1 U13460 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n10589), .ZN(n13769) );
  OAI21_X1 U13461 ( .B1(n13769), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20728), 
        .ZN(n10590) );
  OAI211_X1 U13462 ( .C1(n10626), .C2(n10267), .A(n10591), .B(n10590), .ZN(
        n10592) );
  INV_X1 U13463 ( .A(n10592), .ZN(n10593) );
  NAND2_X1 U13464 ( .A1(n11077), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10609) );
  NAND2_X1 U13465 ( .A1(n13508), .A2(n10795), .ZN(n10600) );
  NAND2_X1 U13466 ( .A1(n20728), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10597) );
  NAND2_X1 U13467 ( .A1(n10922), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n10596) );
  OAI211_X1 U13468 ( .C1(n10626), .C2(n10469), .A(n10597), .B(n10596), .ZN(
        n10598) );
  INV_X1 U13469 ( .A(n10598), .ZN(n10599) );
  NAND2_X1 U13470 ( .A1(n10600), .A2(n10599), .ZN(n13167) );
  XNOR2_X2 U13471 ( .A(n10602), .B(n10601), .ZN(n20261) );
  AOI21_X1 U13472 ( .B1(n20261), .B2(n13522), .A(n20728), .ZN(n13030) );
  NAND2_X1 U13473 ( .A1(n9664), .A2(n10795), .ZN(n10606) );
  AOI22_X1 U13474 ( .A1(n10604), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20728), .ZN(n10605) );
  OAI211_X1 U13475 ( .C1(n10626), .C2(n10275), .A(n10606), .B(n10605), .ZN(
        n13029) );
  MUX2_X1 U13476 ( .A(n10632), .B(n13030), .S(n13029), .Z(n13166) );
  NAND2_X1 U13477 ( .A1(n13167), .A2(n13166), .ZN(n13243) );
  NAND2_X1 U13478 ( .A1(n10608), .A2(n10607), .ZN(n13246) );
  INV_X1 U13479 ( .A(n10610), .ZN(n20323) );
  NAND2_X1 U13480 ( .A1(n10611), .A2(n20323), .ZN(n10612) );
  OAI21_X1 U13481 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10614), .A(
        n10621), .ZN(n13789) );
  AOI22_X1 U13482 ( .A1(n10632), .A2(n13789), .B1(n11077), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U13483 ( .A1(n10922), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10615) );
  OAI211_X1 U13484 ( .C1(n10626), .C2(n10613), .A(n10616), .B(n10615), .ZN(
        n10617) );
  INV_X1 U13485 ( .A(n10617), .ZN(n10618) );
  OAI21_X1 U13486 ( .B1(n20812), .B2(n9914), .A(n10618), .ZN(n13288) );
  NAND2_X1 U13487 ( .A1(n10619), .A2(n9745), .ZN(n10620) );
  NAND2_X1 U13488 ( .A1(n10630), .A2(n10620), .ZN(n11193) );
  INV_X1 U13489 ( .A(n10621), .ZN(n10623) );
  INV_X1 U13490 ( .A(n10631), .ZN(n10622) );
  OAI21_X1 U13491 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10623), .A(
        n10622), .ZN(n20086) );
  INV_X1 U13492 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11134) );
  NAND2_X1 U13493 ( .A1(n10922), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10625) );
  INV_X1 U13494 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20974) );
  OAI21_X1 U13495 ( .B1(n20974), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20728), .ZN(n10624) );
  OAI211_X1 U13496 ( .C1(n10626), .C2(n11134), .A(n10625), .B(n10624), .ZN(
        n10627) );
  OAI21_X1 U13497 ( .B1(n11052), .B2(n20086), .A(n10627), .ZN(n10628) );
  XNOR2_X1 U13498 ( .A(n10630), .B(n10629), .ZN(n11199) );
  INV_X1 U13499 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n10634) );
  XNOR2_X1 U13500 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B(n10631), .ZN(
        n20068) );
  AOI22_X1 U13501 ( .A1(n10632), .A2(n20068), .B1(n11077), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10633) );
  OAI21_X1 U13502 ( .B1(n11022), .B2(n10634), .A(n10633), .ZN(n10635) );
  AOI21_X1 U13503 ( .B1(n11199), .B2(n10795), .A(n10635), .ZN(n13497) );
  NAND2_X1 U13504 ( .A1(n10638), .A2(n10637), .ZN(n11209) );
  INV_X1 U13505 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10645) );
  INV_X1 U13506 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10641) );
  INV_X1 U13507 ( .A(n10639), .ZN(n10640) );
  NAND2_X1 U13508 ( .A1(n10641), .A2(n10640), .ZN(n10642) );
  NAND2_X1 U13509 ( .A1(n10643), .A2(n10642), .ZN(n20047) );
  AOI22_X1 U13510 ( .A1(n20047), .A2(n13559), .B1(n11077), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10644) );
  OAI21_X1 U13511 ( .B1(n11022), .B2(n10645), .A(n10644), .ZN(n10646) );
  AOI22_X1 U13512 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13513 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10329), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13514 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13515 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10648) );
  NAND4_X1 U13516 ( .A1(n10651), .A2(n10650), .A3(n10649), .A4(n10648), .ZN(
        n10657) );
  AOI22_X1 U13517 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9647), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13518 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13519 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10865), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13520 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9667), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10652) );
  NAND4_X1 U13521 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(
        n10656) );
  NOR2_X1 U13522 ( .A1(n10657), .A2(n10656), .ZN(n10662) );
  INV_X1 U13523 ( .A(n10664), .ZN(n10659) );
  XNOR2_X1 U13524 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10659), .ZN(
        n13975) );
  AOI22_X1 U13525 ( .A1(n13559), .A2(n13975), .B1(n11077), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10661) );
  NAND2_X1 U13526 ( .A1(n10922), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10660) );
  OAI211_X1 U13527 ( .C1(n9914), .C2(n10662), .A(n10661), .B(n10660), .ZN(
        n13776) );
  XOR2_X1 U13528 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n10680), .Z(
        n15949) );
  INV_X1 U13529 ( .A(n15949), .ZN(n15923) );
  AOI22_X1 U13530 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13531 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10865), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13532 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13533 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9668), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10665) );
  NAND4_X1 U13534 ( .A1(n10668), .A2(n10667), .A3(n10666), .A4(n10665), .ZN(
        n10674) );
  AOI22_X1 U13535 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13536 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10329), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13537 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U13538 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10669) );
  NAND4_X1 U13539 ( .A1(n10672), .A2(n10671), .A3(n10670), .A4(n10669), .ZN(
        n10673) );
  OAI21_X1 U13540 ( .B1(n10674), .B2(n10673), .A(n10795), .ZN(n10677) );
  NAND2_X1 U13541 ( .A1(n10922), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n10676) );
  NAND2_X1 U13542 ( .A1(n11077), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10675) );
  NAND3_X1 U13543 ( .A1(n10677), .A2(n10676), .A3(n10675), .ZN(n10678) );
  AOI21_X1 U13544 ( .B1(n15923), .B2(n13559), .A(n10678), .ZN(n13917) );
  INV_X1 U13545 ( .A(n13917), .ZN(n10679) );
  XNOR2_X1 U13546 ( .A(n10706), .B(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15918) );
  INV_X1 U13547 ( .A(n11077), .ZN(n10681) );
  NOR2_X1 U13548 ( .A1(n10681), .A2(n15912), .ZN(n10682) );
  AOI21_X1 U13549 ( .B1(n10922), .B2(P1_EAX_REG_11__SCAN_IN), .A(n10682), .ZN(
        n10683) );
  OAI21_X1 U13550 ( .B1(n15918), .B2(n11052), .A(n10683), .ZN(n10695) );
  AOI22_X1 U13551 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13552 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13553 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13554 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10684) );
  NAND4_X1 U13555 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10693) );
  AOI22_X1 U13556 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13557 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11062), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13558 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13559 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10688) );
  NAND4_X1 U13560 ( .A1(n10691), .A2(n10690), .A3(n10689), .A4(n10688), .ZN(
        n10692) );
  OR2_X1 U13561 ( .A1(n10693), .A2(n10692), .ZN(n10694) );
  AND2_X1 U13562 ( .A1(n10795), .A2(n10694), .ZN(n13981) );
  AOI22_X1 U13563 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13564 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13565 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11062), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13566 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10696) );
  NAND4_X1 U13567 ( .A1(n10699), .A2(n10698), .A3(n10697), .A4(n10696), .ZN(
        n10705) );
  AOI22_X1 U13568 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13569 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13570 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13571 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10700) );
  NAND4_X1 U13572 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n10704) );
  OAI21_X1 U13573 ( .B1(n10705), .B2(n10704), .A(n10795), .ZN(n10709) );
  NAND2_X1 U13574 ( .A1(n10922), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10708) );
  XNOR2_X1 U13575 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10710), .ZN(
        n14766) );
  AOI22_X1 U13576 ( .A1(n13559), .A2(n14766), .B1(n11077), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10707) );
  XOR2_X1 U13577 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10734), .Z(
        n14753) );
  AOI22_X1 U13578 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13579 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13580 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13581 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10711) );
  NAND4_X1 U13582 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n10720) );
  AOI22_X1 U13583 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9647), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13584 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13585 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11062), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13586 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9668), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10715) );
  NAND4_X1 U13587 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10719) );
  OR2_X1 U13588 ( .A1(n10720), .A2(n10719), .ZN(n10721) );
  AOI22_X1 U13589 ( .A1(n10795), .A2(n10721), .B1(n11077), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10723) );
  NAND2_X1 U13590 ( .A1(n10604), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10722) );
  OAI211_X1 U13591 ( .C1(n14753), .C2(n11052), .A(n10723), .B(n10722), .ZN(
        n14515) );
  AOI22_X1 U13592 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13593 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10329), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13594 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13595 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10865), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10724) );
  NAND4_X1 U13596 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n10733) );
  AOI22_X1 U13597 ( .A1(n10949), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13598 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13599 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13600 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9668), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10728) );
  NAND4_X1 U13601 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10732) );
  NOR2_X1 U13602 ( .A1(n10733), .A2(n10732), .ZN(n10737) );
  XNOR2_X1 U13603 ( .A(n10738), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15890) );
  NAND2_X1 U13604 ( .A1(n15890), .A2(n13559), .ZN(n10736) );
  AOI22_X1 U13605 ( .A1(n10604), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n11077), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10735) );
  OAI211_X1 U13606 ( .C1(n10737), .C2(n9914), .A(n10736), .B(n10735), .ZN(
        n14508) );
  INV_X1 U13607 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14467) );
  XNOR2_X1 U13608 ( .A(n10804), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14719) );
  AOI22_X1 U13609 ( .A1(n10604), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20728), .ZN(n10755) );
  AOI22_X1 U13610 ( .A1(n10949), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13611 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13612 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10740) );
  NAND2_X1 U13613 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10739) );
  NAND4_X1 U13614 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n10753) );
  INV_X1 U13615 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13616 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10865), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13617 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10747) );
  AOI21_X1 U13618 ( .B1(n10913), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n13559), .ZN(n10746) );
  NAND2_X1 U13619 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10745) );
  AND4_X1 U13620 ( .A1(n10748), .A2(n10747), .A3(n10746), .A4(n10745), .ZN(
        n10750) );
  AOI22_X1 U13621 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9669), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10749) );
  OAI211_X1 U13622 ( .C1(n10877), .C2(n10751), .A(n10750), .B(n10749), .ZN(
        n10752) );
  NAND2_X1 U13623 ( .A1(n11049), .A2(n11052), .ZN(n10878) );
  OAI21_X1 U13624 ( .B1(n10753), .B2(n10752), .A(n10878), .ZN(n10754) );
  AOI22_X1 U13625 ( .A1(n14719), .A2(n13559), .B1(n10755), .B2(n10754), .ZN(
        n14449) );
  XOR2_X1 U13626 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10756), .Z(
        n15870) );
  INV_X1 U13627 ( .A(n15870), .ZN(n15933) );
  AOI22_X1 U13628 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13629 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10329), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13630 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13631 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10865), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10757) );
  NAND4_X1 U13632 ( .A1(n10760), .A2(n10759), .A3(n10758), .A4(n10757), .ZN(
        n10766) );
  AOI22_X1 U13633 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13634 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13635 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13636 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10761) );
  NAND4_X1 U13637 ( .A1(n10764), .A2(n10763), .A3(n10762), .A4(n10761), .ZN(
        n10765) );
  NOR2_X1 U13638 ( .A1(n10766), .A2(n10765), .ZN(n10768) );
  AOI22_X1 U13639 ( .A1(n10604), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n11077), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10767) );
  OAI21_X1 U13640 ( .B1(n11049), .B2(n10768), .A(n10767), .ZN(n10769) );
  AOI21_X1 U13641 ( .B1(n15933), .B2(n13559), .A(n10769), .ZN(n14496) );
  XNOR2_X1 U13642 ( .A(n10770), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14733) );
  NAND2_X1 U13643 ( .A1(n14733), .A2(n13559), .ZN(n10785) );
  AOI22_X1 U13644 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13645 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13646 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13647 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10771) );
  NAND4_X1 U13648 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n10780) );
  AOI22_X1 U13649 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13650 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13651 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13652 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9667), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10775) );
  NAND4_X1 U13653 ( .A1(n10778), .A2(n10777), .A3(n10776), .A4(n10775), .ZN(
        n10779) );
  NOR2_X1 U13654 ( .A1(n10780), .A2(n10779), .ZN(n10783) );
  AOI21_X1 U13655 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14467), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10781) );
  AOI21_X1 U13656 ( .B1(n10922), .B2(P1_EAX_REG_16__SCAN_IN), .A(n10781), .ZN(
        n10782) );
  OAI21_X1 U13657 ( .B1(n11049), .B2(n10783), .A(n10782), .ZN(n10784) );
  NAND2_X1 U13658 ( .A1(n10785), .A2(n10784), .ZN(n14461) );
  XOR2_X1 U13659 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n10786), .Z(
        n15944) );
  INV_X1 U13660 ( .A(n15944), .ZN(n10802) );
  AOI22_X1 U13661 ( .A1(n10949), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13662 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9643), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13663 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13664 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10787) );
  NAND4_X1 U13665 ( .A1(n10790), .A2(n10789), .A3(n10788), .A4(n10787), .ZN(
        n10797) );
  AOI22_X1 U13666 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13667 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n9665), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13668 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13669 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10791) );
  NAND4_X1 U13670 ( .A1(n10794), .A2(n10793), .A3(n10792), .A4(n10791), .ZN(
        n10796) );
  OAI21_X1 U13671 ( .B1(n10797), .B2(n10796), .A(n10795), .ZN(n10800) );
  NAND2_X1 U13672 ( .A1(n10604), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U13673 ( .A1(n11077), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10798) );
  NAND3_X1 U13674 ( .A1(n10800), .A2(n10799), .A3(n10798), .ZN(n10801) );
  AOI21_X1 U13675 ( .B1(n10802), .B2(n13559), .A(n10801), .ZN(n14596) );
  OR2_X1 U13676 ( .A1(n14461), .A2(n14596), .ZN(n14459) );
  NOR2_X1 U13677 ( .A1(n14496), .A2(n14459), .ZN(n14448) );
  AND2_X1 U13678 ( .A1(n14449), .A2(n14448), .ZN(n10803) );
  INV_X1 U13679 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14714) );
  INV_X1 U13680 ( .A(n10805), .ZN(n10807) );
  INV_X1 U13681 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10806) );
  NAND2_X1 U13682 ( .A1(n10807), .A2(n10806), .ZN(n10808) );
  NAND2_X1 U13683 ( .A1(n10843), .A2(n10808), .ZN(n14710) );
  AOI22_X1 U13684 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13685 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U13686 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13687 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10809) );
  NAND4_X1 U13688 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(
        n10818) );
  AOI22_X1 U13689 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U13690 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13691 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13692 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9667), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10813) );
  NAND4_X1 U13693 ( .A1(n10816), .A2(n10815), .A3(n10814), .A4(n10813), .ZN(
        n10817) );
  NOR2_X1 U13694 ( .A1(n10818), .A2(n10817), .ZN(n10821) );
  OAI21_X1 U13695 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20974), .A(
        n20728), .ZN(n10820) );
  NAND2_X1 U13696 ( .A1(n10604), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n10819) );
  OAI211_X1 U13697 ( .C1(n11049), .C2(n10821), .A(n10820), .B(n10819), .ZN(
        n10822) );
  NAND2_X1 U13698 ( .A1(n10823), .A2(n10822), .ZN(n14431) );
  XNOR2_X1 U13699 ( .A(n10843), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14699) );
  NAND2_X1 U13700 ( .A1(n14699), .A2(n13559), .ZN(n10842) );
  AOI22_X1 U13701 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10865), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13702 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10367), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13703 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10827) );
  NAND2_X1 U13704 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10826) );
  NAND4_X1 U13705 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10838) );
  INV_X1 U13706 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13707 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13708 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10832) );
  AOI21_X1 U13709 ( .B1(n10913), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n13559), .ZN(n10831) );
  NAND2_X1 U13710 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10830) );
  AND4_X1 U13711 ( .A1(n10833), .A2(n10832), .A3(n10831), .A4(n10830), .ZN(
        n10835) );
  AOI22_X1 U13712 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10575), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10834) );
  OAI211_X1 U13713 ( .C1(n10877), .C2(n10836), .A(n10835), .B(n10834), .ZN(
        n10837) );
  OAI21_X1 U13714 ( .B1(n10838), .B2(n10837), .A(n10878), .ZN(n10840) );
  AOI22_X1 U13715 ( .A1(n10604), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20728), .ZN(n10839) );
  NAND2_X1 U13716 ( .A1(n10840), .A2(n10839), .ZN(n10841) );
  NAND2_X1 U13717 ( .A1(n10842), .A2(n10841), .ZN(n14418) );
  INV_X1 U13718 ( .A(n10845), .ZN(n10847) );
  INV_X1 U13719 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10846) );
  NAND2_X1 U13720 ( .A1(n10847), .A2(n10846), .ZN(n10848) );
  NAND2_X1 U13721 ( .A1(n10883), .A2(n10848), .ZN(n14691) );
  AOI22_X1 U13722 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13723 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10329), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U13724 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13725 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10849) );
  NAND4_X1 U13726 ( .A1(n10852), .A2(n10851), .A3(n10850), .A4(n10849), .ZN(
        n10858) );
  AOI22_X1 U13727 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13728 ( .A1(n10865), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13729 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13730 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10853) );
  NAND4_X1 U13731 ( .A1(n10856), .A2(n10855), .A3(n10854), .A4(n10853), .ZN(
        n10857) );
  NOR2_X1 U13732 ( .A1(n10858), .A2(n10857), .ZN(n10862) );
  NAND2_X1 U13733 ( .A1(n20728), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10859) );
  NAND2_X1 U13734 ( .A1(n11052), .A2(n10859), .ZN(n10860) );
  AOI21_X1 U13735 ( .B1(n10922), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10860), .ZN(
        n10861) );
  OAI21_X1 U13736 ( .B1(n11049), .B2(n10862), .A(n10861), .ZN(n10863) );
  XNOR2_X1 U13737 ( .A(n10883), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14681) );
  AOI22_X1 U13738 ( .A1(n10604), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20728), .ZN(n10882) );
  AOI22_X1 U13739 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10865), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13740 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13741 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10867) );
  NAND2_X1 U13742 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10866) );
  NAND4_X1 U13743 ( .A1(n10869), .A2(n10868), .A3(n10867), .A4(n10866), .ZN(
        n10880) );
  INV_X1 U13744 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13745 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13746 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10872) );
  AOI21_X1 U13747 ( .B1(n10913), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n13559), .ZN(n10871) );
  NAND2_X1 U13748 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10870) );
  AND4_X1 U13749 ( .A1(n10873), .A2(n10872), .A3(n10871), .A4(n10870), .ZN(
        n10875) );
  AOI22_X1 U13750 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9669), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10874) );
  OAI211_X1 U13751 ( .C1(n10877), .C2(n10876), .A(n10875), .B(n10874), .ZN(
        n10879) );
  OAI21_X1 U13752 ( .B1(n10880), .B2(n10879), .A(n10878), .ZN(n10881) );
  AOI22_X1 U13753 ( .A1(n14681), .A2(n13559), .B1(n10882), .B2(n10881), .ZN(
        n14393) );
  INV_X1 U13754 ( .A(n10885), .ZN(n10887) );
  INV_X1 U13755 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10886) );
  NAND2_X1 U13756 ( .A1(n10887), .A2(n10886), .ZN(n10888) );
  NAND2_X1 U13757 ( .A1(n10945), .A2(n10888), .ZN(n14673) );
  INV_X1 U13758 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10901) );
  INV_X1 U13759 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10891) );
  INV_X1 U13760 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10889) );
  OAI22_X1 U13761 ( .A1(n10744), .A2(n10891), .B1(n10890), .B2(n10889), .ZN(
        n10897) );
  INV_X1 U13762 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10895) );
  INV_X1 U13763 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10892) );
  OAI22_X1 U13764 ( .A1(n10895), .A2(n10894), .B1(n10893), .B2(n10892), .ZN(
        n10896) );
  AOI211_X1 U13765 ( .C1(n10396), .C2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n10897), .B(n10896), .ZN(n10899) );
  AOI22_X1 U13766 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10898) );
  OAI211_X1 U13767 ( .C1(n10901), .C2(n10900), .A(n10899), .B(n10898), .ZN(
        n10907) );
  AOI22_X1 U13768 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11032), .B1(
        n10329), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U13769 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9652), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13770 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13771 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10902) );
  NAND4_X1 U13772 ( .A1(n10905), .A2(n10904), .A3(n10903), .A4(n10902), .ZN(
        n10906) );
  NOR2_X1 U13773 ( .A1(n10907), .A2(n10906), .ZN(n10927) );
  AOI22_X1 U13774 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13775 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13776 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13777 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9667), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10909) );
  NAND4_X1 U13778 ( .A1(n10912), .A2(n10911), .A3(n10910), .A4(n10909), .ZN(
        n10919) );
  AOI22_X1 U13779 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13780 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13781 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13782 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10914) );
  NAND4_X1 U13783 ( .A1(n10917), .A2(n10916), .A3(n10915), .A4(n10914), .ZN(
        n10918) );
  NOR2_X1 U13784 ( .A1(n10919), .A2(n10918), .ZN(n10928) );
  XNOR2_X1 U13785 ( .A(n10927), .B(n10928), .ZN(n10924) );
  NAND2_X1 U13786 ( .A1(n20728), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10920) );
  NAND2_X1 U13787 ( .A1(n11052), .A2(n10920), .ZN(n10921) );
  AOI21_X1 U13788 ( .B1(n10922), .B2(P1_EAX_REG_23__SCAN_IN), .A(n10921), .ZN(
        n10923) );
  OAI21_X1 U13789 ( .B1(n10924), .B2(n11049), .A(n10923), .ZN(n10925) );
  NAND2_X1 U13790 ( .A1(n10926), .A2(n10925), .ZN(n14378) );
  XNOR2_X1 U13791 ( .A(n10945), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14665) );
  NAND2_X1 U13792 ( .A1(n14665), .A2(n13559), .ZN(n10944) );
  NOR2_X1 U13793 ( .A1(n10928), .A2(n10927), .ZN(n10961) );
  AOI22_X1 U13794 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13795 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13796 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U13797 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9652), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10929) );
  NAND4_X1 U13798 ( .A1(n10932), .A2(n10931), .A3(n10930), .A4(n10929), .ZN(
        n10938) );
  AOI22_X1 U13799 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13800 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U13801 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13802 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10933) );
  NAND4_X1 U13803 ( .A1(n10936), .A2(n10935), .A3(n10934), .A4(n10933), .ZN(
        n10937) );
  OR2_X1 U13804 ( .A1(n10938), .A2(n10937), .ZN(n10960) );
  XNOR2_X1 U13805 ( .A(n10961), .B(n10960), .ZN(n10942) );
  NAND2_X1 U13806 ( .A1(n20728), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10939) );
  NAND2_X1 U13807 ( .A1(n11052), .A2(n10939), .ZN(n10940) );
  AOI21_X1 U13808 ( .B1(n10604), .B2(P1_EAX_REG_24__SCAN_IN), .A(n10940), .ZN(
        n10941) );
  OAI21_X1 U13809 ( .B1(n10942), .B2(n11049), .A(n10941), .ZN(n10943) );
  NAND2_X1 U13810 ( .A1(n10944), .A2(n10943), .ZN(n14367) );
  INV_X1 U13811 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14667) );
  INV_X1 U13812 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10946) );
  NAND2_X1 U13813 ( .A1(n10947), .A2(n10946), .ZN(n10948) );
  NAND2_X1 U13814 ( .A1(n10984), .A2(n10948), .ZN(n14658) );
  INV_X1 U13815 ( .A(n14658), .ZN(n14360) );
  AOI22_X1 U13816 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U13817 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U13818 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9668), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U13819 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10950) );
  NAND4_X1 U13820 ( .A1(n10953), .A2(n10952), .A3(n10951), .A4(n10950), .ZN(
        n10959) );
  AOI22_X1 U13821 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9669), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13822 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13823 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U13824 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10954) );
  NAND4_X1 U13825 ( .A1(n10957), .A2(n10956), .A3(n10955), .A4(n10954), .ZN(
        n10958) );
  NOR2_X1 U13826 ( .A1(n10959), .A2(n10958), .ZN(n10967) );
  NAND2_X1 U13827 ( .A1(n10961), .A2(n10960), .ZN(n10966) );
  XOR2_X1 U13828 ( .A(n10967), .B(n10966), .Z(n10964) );
  INV_X1 U13829 ( .A(n11049), .ZN(n11073) );
  INV_X1 U13830 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14548) );
  NAND2_X1 U13831 ( .A1(n20728), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10962) );
  OAI211_X1 U13832 ( .C1(n11022), .C2(n14548), .A(n11052), .B(n10962), .ZN(
        n10963) );
  AOI21_X1 U13833 ( .B1(n10964), .B2(n11073), .A(n10963), .ZN(n10965) );
  AOI21_X1 U13834 ( .B1(n14360), .B2(n13559), .A(n10965), .ZN(n14354) );
  XNOR2_X1 U13835 ( .A(n10984), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14645) );
  NAND2_X1 U13836 ( .A1(n14645), .A2(n13559), .ZN(n10983) );
  NOR2_X1 U13837 ( .A1(n10967), .A2(n10966), .ZN(n11000) );
  AOI22_X1 U13838 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U13839 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U13840 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U13841 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9652), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10968) );
  NAND4_X1 U13842 ( .A1(n10971), .A2(n10970), .A3(n10969), .A4(n10968), .ZN(
        n10977) );
  AOI22_X1 U13843 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U13844 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13845 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U13846 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10972) );
  NAND4_X1 U13847 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n10976) );
  OR2_X1 U13848 ( .A1(n10977), .A2(n10976), .ZN(n10999) );
  XNOR2_X1 U13849 ( .A(n11000), .B(n10999), .ZN(n10981) );
  NAND2_X1 U13850 ( .A1(n20728), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10978) );
  NAND2_X1 U13851 ( .A1(n11052), .A2(n10978), .ZN(n10979) );
  AOI21_X1 U13852 ( .B1(n10604), .B2(P1_EAX_REG_26__SCAN_IN), .A(n10979), .ZN(
        n10980) );
  OAI21_X1 U13853 ( .B1(n10981), .B2(n11049), .A(n10980), .ZN(n10982) );
  NAND2_X1 U13854 ( .A1(n10983), .A2(n10982), .ZN(n14345) );
  OR2_X2 U13855 ( .A1(n14344), .A2(n14345), .ZN(n14329) );
  INV_X1 U13856 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14647) );
  INV_X1 U13857 ( .A(n10985), .ZN(n10987) );
  INV_X1 U13858 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10986) );
  NAND2_X1 U13859 ( .A1(n10987), .A2(n10986), .ZN(n10988) );
  NAND2_X1 U13860 ( .A1(n11026), .A2(n10988), .ZN(n14635) );
  AOI22_X1 U13861 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U13862 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9647), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U13863 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U13864 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10989) );
  NAND4_X1 U13865 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n10998) );
  AOI22_X1 U13866 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9670), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U13867 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U13868 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13869 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10993) );
  NAND4_X1 U13870 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n10997) );
  NOR2_X1 U13871 ( .A1(n10998), .A2(n10997), .ZN(n11008) );
  NAND2_X1 U13872 ( .A1(n11000), .A2(n10999), .ZN(n11007) );
  XNOR2_X1 U13873 ( .A(n11008), .B(n11007), .ZN(n11004) );
  NAND2_X1 U13874 ( .A1(n20728), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11001) );
  NAND2_X1 U13875 ( .A1(n11052), .A2(n11001), .ZN(n11002) );
  AOI21_X1 U13876 ( .B1(n10604), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11002), .ZN(
        n11003) );
  OAI21_X1 U13877 ( .B1(n11004), .B2(n11049), .A(n11003), .ZN(n11005) );
  NAND2_X1 U13878 ( .A1(n11006), .A2(n11005), .ZN(n14330) );
  XNOR2_X1 U13879 ( .A(n11026), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14622) );
  NOR2_X1 U13880 ( .A1(n11008), .A2(n11007), .ZN(n11046) );
  AOI22_X1 U13881 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U13882 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U13883 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U13884 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9652), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11009) );
  NAND4_X1 U13885 ( .A1(n11012), .A2(n11011), .A3(n11010), .A4(n11009), .ZN(
        n11019) );
  AOI22_X1 U13886 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9647), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U13887 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U13888 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11013), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U13889 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11014) );
  NAND4_X1 U13890 ( .A1(n11017), .A2(n11016), .A3(n11015), .A4(n11014), .ZN(
        n11018) );
  OR2_X1 U13891 ( .A1(n11019), .A2(n11018), .ZN(n11045) );
  INV_X1 U13892 ( .A(n11045), .ZN(n11020) );
  XNOR2_X1 U13893 ( .A(n11046), .B(n11020), .ZN(n11024) );
  INV_X1 U13894 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14537) );
  NAND2_X1 U13895 ( .A1(n20728), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11021) );
  OAI211_X1 U13896 ( .C1(n11022), .C2(n14537), .A(n11052), .B(n11021), .ZN(
        n11023) );
  AOI21_X1 U13897 ( .B1(n11024), .B2(n11073), .A(n11023), .ZN(n11025) );
  AOI21_X1 U13898 ( .B1(n14622), .B2(n13559), .A(n11025), .ZN(n14317) );
  INV_X1 U13899 ( .A(n11026), .ZN(n11027) );
  INV_X1 U13900 ( .A(n11028), .ZN(n11030) );
  INV_X1 U13901 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11029) );
  NAND2_X1 U13902 ( .A1(n11030), .A2(n11029), .ZN(n11031) );
  NAND2_X1 U13903 ( .A1(n11080), .A2(n11031), .ZN(n14610) );
  AOI22_X1 U13904 ( .A1(n10397), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U13905 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U13906 ( .A1(n10908), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U13907 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10347), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11034) );
  NAND4_X1 U13908 ( .A1(n11037), .A2(n11036), .A3(n11035), .A4(n11034), .ZN(
        n11044) );
  AOI22_X1 U13909 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U13910 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U13911 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11062), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U13912 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11038), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11039) );
  NAND4_X1 U13913 ( .A1(n11042), .A2(n11041), .A3(n11040), .A4(n11039), .ZN(
        n11043) );
  NOR2_X1 U13914 ( .A1(n11044), .A2(n11043), .ZN(n11055) );
  NAND2_X1 U13915 ( .A1(n11046), .A2(n11045), .ZN(n11054) );
  XNOR2_X1 U13916 ( .A(n11055), .B(n11054), .ZN(n11050) );
  AOI21_X1 U13917 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20728), .A(
        n13559), .ZN(n11048) );
  NAND2_X1 U13918 ( .A1(n10604), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11047) );
  OAI211_X1 U13919 ( .C1(n11050), .C2(n11049), .A(n11048), .B(n11047), .ZN(
        n11051) );
  OAI21_X1 U13920 ( .B1(n14610), .B2(n11052), .A(n11051), .ZN(n14306) );
  XNOR2_X1 U13921 ( .A(n11080), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14298) );
  INV_X1 U13922 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14291) );
  AOI21_X1 U13923 ( .B1(n14291), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11053) );
  AOI21_X1 U13924 ( .B1(n10604), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11053), .ZN(
        n11076) );
  NOR2_X1 U13925 ( .A1(n11055), .A2(n11054), .ZN(n11072) );
  AOI22_X1 U13926 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10397), .B1(
        n10396), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U13927 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U13928 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n9652), .B1(
        n10543), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U13929 ( .A1(n11038), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11058) );
  NAND4_X1 U13930 ( .A1(n11061), .A2(n11060), .A3(n11059), .A4(n11058), .ZN(
        n11070) );
  AOI22_X1 U13931 ( .A1(n10575), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10949), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U13932 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10913), .B1(
        n9670), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U13933 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10908), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U13934 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9643), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11065) );
  NAND4_X1 U13935 ( .A1(n11068), .A2(n11067), .A3(n11066), .A4(n11065), .ZN(
        n11069) );
  NOR2_X1 U13936 ( .A1(n11070), .A2(n11069), .ZN(n11071) );
  XNOR2_X1 U13937 ( .A(n11072), .B(n11071), .ZN(n11074) );
  NAND2_X1 U13938 ( .A1(n11074), .A2(n11073), .ZN(n11075) );
  AOI22_X1 U13939 ( .A1(n14298), .A2(n13559), .B1(n11076), .B2(n11075), .ZN(
        n11267) );
  AOI22_X1 U13940 ( .A1(n10604), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n11077), .ZN(n11078) );
  XNOR2_X2 U13941 ( .A(n9697), .B(n11079), .ZN(n14275) );
  NOR2_X1 U13942 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20671) );
  AND2_X1 U13943 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20671), .ZN(n14943) );
  NAND2_X1 U13944 ( .A1(n14275), .A2(n15960), .ZN(n11266) );
  NAND2_X1 U13945 ( .A1(n20489), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11106) );
  NAND2_X1 U13946 ( .A1(n10469), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11082) );
  NAND2_X1 U13947 ( .A1(n11106), .A2(n11082), .ZN(n11105) );
  NAND2_X1 U13948 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20588), .ZN(
        n11104) );
  XNOR2_X1 U13949 ( .A(n11105), .B(n11104), .ZN(n11277) );
  NAND2_X1 U13950 ( .A1(n11133), .A2(n11277), .ZN(n11084) );
  NAND2_X1 U13951 ( .A1(n11143), .A2(n10412), .ZN(n11083) );
  NAND2_X1 U13952 ( .A1(n20213), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11094) );
  AND3_X1 U13953 ( .A1(n11084), .A2(n11083), .A3(n11094), .ZN(n11099) );
  OAI21_X1 U13954 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20588), .A(
        n11104), .ZN(n11085) );
  INV_X1 U13955 ( .A(n11085), .ZN(n11089) );
  NAND2_X1 U13956 ( .A1(n11143), .A2(n11089), .ZN(n11086) );
  NAND2_X1 U13957 ( .A1(n11144), .A2(n11086), .ZN(n11093) );
  INV_X1 U13958 ( .A(n11087), .ZN(n11088) );
  AOI21_X1 U13959 ( .B1(n10170), .B2(n11089), .A(n11088), .ZN(n11091) );
  NAND2_X1 U13960 ( .A1(n13565), .A2(n11090), .ZN(n11114) );
  OR2_X1 U13961 ( .A1(n11091), .A2(n11114), .ZN(n11092) );
  NAND2_X1 U13962 ( .A1(n11093), .A2(n11092), .ZN(n11098) );
  NAND2_X1 U13963 ( .A1(n11099), .A2(n11098), .ZN(n11097) );
  INV_X1 U13964 ( .A(n11094), .ZN(n11095) );
  NAND2_X1 U13965 ( .A1(n11136), .A2(n11277), .ZN(n11096) );
  NAND2_X1 U13966 ( .A1(n11097), .A2(n11096), .ZN(n11103) );
  INV_X1 U13967 ( .A(n11098), .ZN(n11101) );
  INV_X1 U13968 ( .A(n11099), .ZN(n11100) );
  NAND2_X1 U13969 ( .A1(n11101), .A2(n11100), .ZN(n11102) );
  NAND2_X1 U13970 ( .A1(n11103), .A2(n11102), .ZN(n11112) );
  OR2_X1 U13971 ( .A1(n11105), .A2(n11104), .ZN(n11107) );
  NAND2_X1 U13972 ( .A1(n11107), .A2(n11106), .ZN(n11118) );
  MUX2_X1 U13973 ( .A(n11119), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11108) );
  XNOR2_X1 U13974 ( .A(n11118), .B(n11108), .ZN(n11279) );
  INV_X1 U13975 ( .A(n11279), .ZN(n11113) );
  NAND2_X1 U13976 ( .A1(n11143), .A2(n11113), .ZN(n11110) );
  INV_X1 U13977 ( .A(n11114), .ZN(n11109) );
  OAI211_X1 U13978 ( .C1(n11113), .C2(n11130), .A(n11110), .B(n11109), .ZN(
        n11111) );
  NAND2_X1 U13979 ( .A1(n11112), .A2(n11111), .ZN(n11116) );
  NAND3_X1 U13980 ( .A1(n11143), .A2(n11114), .A3(n11113), .ZN(n11115) );
  NAND2_X1 U13981 ( .A1(n11116), .A2(n11115), .ZN(n11123) );
  NAND2_X1 U13982 ( .A1(n11118), .A2(n11117), .ZN(n11121) );
  NAND2_X1 U13983 ( .A1(n11119), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11120) );
  NAND2_X1 U13984 ( .A1(n11121), .A2(n11120), .ZN(n11129) );
  MUX2_X1 U13985 ( .A(n20519), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11128) );
  XNOR2_X1 U13986 ( .A(n11129), .B(n11128), .ZN(n11278) );
  NAND2_X1 U13987 ( .A1(n11130), .A2(n11278), .ZN(n11122) );
  NAND2_X1 U13988 ( .A1(n11123), .A2(n11122), .ZN(n11126) );
  INV_X1 U13989 ( .A(n11144), .ZN(n11124) );
  NAND2_X1 U13990 ( .A1(n11124), .A2(n11278), .ZN(n11125) );
  NAND2_X1 U13991 ( .A1(n11126), .A2(n11125), .ZN(n11132) );
  NOR2_X1 U13992 ( .A1(n10613), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11127) );
  NOR2_X1 U13993 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20182), .ZN(
        n11140) );
  NAND2_X1 U13994 ( .A1(n11130), .A2(n11280), .ZN(n11131) );
  NAND2_X1 U13995 ( .A1(n11132), .A2(n11131), .ZN(n11139) );
  NAND2_X1 U13996 ( .A1(n11133), .A2(n11280), .ZN(n11135) );
  OAI22_X1 U13997 ( .A1(n11136), .A2(n11135), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n11134), .ZN(n11137) );
  INV_X1 U13998 ( .A(n11137), .ZN(n11138) );
  NAND2_X1 U13999 ( .A1(n20182), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11141) );
  AOI21_X1 U14000 ( .B1(n11142), .B2(n11141), .A(n11140), .ZN(n11282) );
  INV_X1 U14001 ( .A(n11282), .ZN(n11146) );
  NAND2_X1 U14002 ( .A1(n15822), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20001) );
  NAND2_X1 U14003 ( .A1(n10415), .A2(n20184), .ZN(n11150) );
  NAND2_X1 U14004 ( .A1(n11150), .A2(n13080), .ZN(n11151) );
  NAND2_X1 U14005 ( .A1(n13059), .A2(n13076), .ZN(n15808) );
  INV_X1 U14006 ( .A(n20671), .ZN(n20664) );
  NAND2_X1 U14007 ( .A1(n12894), .A2(n20664), .ZN(n11152) );
  NAND2_X1 U14008 ( .A1(n11152), .A2(n16039), .ZN(n11153) );
  NAND2_X1 U14009 ( .A1(n16039), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11155) );
  NAND2_X1 U14010 ( .A1(n20974), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11154) );
  AND2_X1 U14011 ( .A1(n11155), .A2(n11154), .ZN(n13261) );
  INV_X1 U14012 ( .A(n15948), .ZN(n14772) );
  INV_X1 U14013 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11156) );
  NOR2_X1 U14014 ( .A1(n12894), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16031) );
  INV_X2 U14015 ( .A(n16031), .ZN(n20073) );
  NAND2_X1 U14016 ( .A1(n9645), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14074) );
  OAI21_X1 U14017 ( .B1(n14772), .B2(n11156), .A(n14074), .ZN(n11157) );
  AOI21_X1 U14018 ( .B1(n13568), .B2(n15950), .A(n11157), .ZN(n11265) );
  NAND2_X1 U14019 ( .A1(n11225), .A2(n11222), .ZN(n11160) );
  NOR2_X1 U14020 ( .A1(n11160), .A2(n11159), .ZN(n11161) );
  INV_X1 U14021 ( .A(n11225), .ZN(n11192) );
  NAND2_X1 U14022 ( .A1(n13034), .A2(n11164), .ZN(n11162) );
  NAND2_X1 U14023 ( .A1(n20184), .A2(n13023), .ZN(n11177) );
  AND2_X1 U14024 ( .A1(n11162), .A2(n11177), .ZN(n11163) );
  XNOR2_X1 U14025 ( .A(n11164), .B(n11173), .ZN(n11165) );
  NAND2_X1 U14026 ( .A1(n11165), .A2(n13034), .ZN(n11166) );
  INV_X1 U14027 ( .A(n11168), .ZN(n13048) );
  NAND2_X1 U14028 ( .A1(n13048), .A2(n11169), .ZN(n11170) );
  INV_X1 U14029 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20180) );
  NAND2_X1 U14030 ( .A1(n13507), .A2(n11225), .ZN(n11181) );
  NAND2_X1 U14031 ( .A1(n11174), .A2(n11173), .ZN(n11175) );
  NAND2_X1 U14032 ( .A1(n11175), .A2(n11176), .ZN(n11185) );
  OAI21_X1 U14033 ( .B1(n11176), .B2(n11175), .A(n11185), .ZN(n11179) );
  INV_X1 U14034 ( .A(n11177), .ZN(n11178) );
  AOI21_X1 U14035 ( .B1(n11179), .B2(n13034), .A(n11178), .ZN(n11180) );
  NAND2_X1 U14036 ( .A1(n11181), .A2(n11180), .ZN(n13486) );
  NAND2_X1 U14037 ( .A1(n13487), .A2(n13486), .ZN(n11184) );
  NAND2_X1 U14038 ( .A1(n11182), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11183) );
  NAND2_X1 U14039 ( .A1(n11184), .A2(n11183), .ZN(n13348) );
  NAND2_X1 U14040 ( .A1(n11185), .A2(n11186), .ZN(n11202) );
  OAI211_X1 U14041 ( .C1(n11186), .C2(n11185), .A(n11202), .B(n13034), .ZN(
        n11187) );
  INV_X1 U14042 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11188) );
  XNOR2_X1 U14043 ( .A(n11189), .B(n11188), .ZN(n13347) );
  NAND2_X1 U14044 ( .A1(n13348), .A2(n13347), .ZN(n11191) );
  NAND2_X1 U14045 ( .A1(n11189), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11190) );
  NAND2_X1 U14046 ( .A1(n11191), .A2(n11190), .ZN(n13451) );
  XNOR2_X1 U14047 ( .A(n11202), .B(n11200), .ZN(n11194) );
  NAND2_X1 U14048 ( .A1(n11194), .A2(n13034), .ZN(n11195) );
  INV_X1 U14049 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13442) );
  XNOR2_X1 U14050 ( .A(n11197), .B(n13442), .ZN(n13450) );
  NAND2_X1 U14051 ( .A1(n11197), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11198) );
  NAND2_X1 U14052 ( .A1(n11199), .A2(n11225), .ZN(n11205) );
  INV_X1 U14053 ( .A(n11200), .ZN(n11201) );
  OR2_X1 U14054 ( .A1(n11202), .A2(n11201), .ZN(n11212) );
  XNOR2_X1 U14055 ( .A(n11212), .B(n11210), .ZN(n11203) );
  NAND2_X1 U14056 ( .A1(n11203), .A2(n13034), .ZN(n11204) );
  NAND2_X1 U14057 ( .A1(n11205), .A2(n11204), .ZN(n11207) );
  INV_X1 U14058 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11206) );
  XNOR2_X1 U14059 ( .A(n11207), .B(n11206), .ZN(n13493) );
  NAND2_X1 U14060 ( .A1(n11207), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11208) );
  INV_X1 U14061 ( .A(n11210), .ZN(n11211) );
  OR2_X1 U14062 ( .A1(n11212), .A2(n11211), .ZN(n11219) );
  XNOR2_X1 U14063 ( .A(n11219), .B(n11220), .ZN(n11213) );
  NAND2_X1 U14064 ( .A1(n11213), .A2(n13034), .ZN(n11214) );
  NAND2_X1 U14065 ( .A1(n11215), .A2(n11214), .ZN(n11216) );
  INV_X1 U14066 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13592) );
  XNOR2_X1 U14067 ( .A(n11216), .B(n13592), .ZN(n13707) );
  NAND2_X1 U14068 ( .A1(n13706), .A2(n13707), .ZN(n11218) );
  NAND2_X1 U14069 ( .A1(n11216), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11217) );
  INV_X1 U14070 ( .A(n11219), .ZN(n11221) );
  NAND2_X1 U14071 ( .A1(n11221), .A2(n11220), .ZN(n11232) );
  XNOR2_X1 U14072 ( .A(n11232), .B(n11222), .ZN(n11223) );
  AND2_X1 U14073 ( .A1(n11223), .A2(n13034), .ZN(n11224) );
  AOI21_X1 U14074 ( .B1(n11226), .B2(n11225), .A(n11224), .ZN(n11227) );
  INV_X1 U14075 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13854) );
  NAND2_X1 U14076 ( .A1(n11227), .A2(n13854), .ZN(n15957) );
  INV_X1 U14077 ( .A(n11227), .ZN(n11228) );
  NAND2_X1 U14078 ( .A1(n11228), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15956) );
  INV_X1 U14079 ( .A(n13034), .ZN(n11230) );
  OR3_X1 U14080 ( .A1(n11232), .A2(n11231), .A3(n11230), .ZN(n11233) );
  INV_X1 U14081 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13755) );
  INV_X1 U14082 ( .A(n13845), .ZN(n11234) );
  NAND2_X1 U14083 ( .A1(n11234), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11235) );
  INV_X1 U14084 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13971) );
  NAND2_X1 U14085 ( .A1(n9649), .A2(n13971), .ZN(n11237) );
  NAND2_X1 U14086 ( .A1(n14884), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14741) );
  INV_X1 U14087 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U14088 ( .A1(n11236), .A2(n14907), .ZN(n11238) );
  NAND2_X1 U14089 ( .A1(n14741), .A2(n11238), .ZN(n14750) );
  INV_X1 U14090 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13993) );
  NAND2_X1 U14091 ( .A1(n11236), .A2(n13993), .ZN(n14760) );
  NAND2_X1 U14092 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U14093 ( .A1(n11236), .A2(n11239), .ZN(n14748) );
  NAND2_X1 U14094 ( .A1(n14760), .A2(n14748), .ZN(n11240) );
  NOR2_X1 U14095 ( .A1(n14750), .A2(n11240), .ZN(n14740) );
  NAND2_X1 U14096 ( .A1(n9649), .A2(n16000), .ZN(n11241) );
  NAND2_X1 U14097 ( .A1(n14740), .A2(n11241), .ZN(n14723) );
  NAND2_X1 U14098 ( .A1(n9972), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11242) );
  NAND2_X1 U14099 ( .A1(n14741), .A2(n11242), .ZN(n14724) );
  INV_X1 U14100 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15996) );
  NOR2_X1 U14101 ( .A1(n11236), .A2(n15996), .ZN(n14728) );
  NOR2_X1 U14102 ( .A1(n14724), .A2(n14728), .ZN(n11245) );
  XNOR2_X1 U14103 ( .A(n11236), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14732) );
  NAND2_X1 U14104 ( .A1(n11236), .A2(n15996), .ZN(n14730) );
  NAND2_X1 U14105 ( .A1(n14732), .A2(n14730), .ZN(n11243) );
  AOI21_X1 U14106 ( .B1(n14723), .B2(n11245), .A(n11243), .ZN(n14881) );
  NAND2_X1 U14107 ( .A1(n9648), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14761) );
  INV_X1 U14108 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14919) );
  INV_X1 U14109 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14930) );
  NAND2_X1 U14110 ( .A1(n14919), .A2(n14930), .ZN(n11244) );
  NAND2_X1 U14111 ( .A1(n9648), .A2(n11244), .ZN(n14757) );
  NAND2_X1 U14112 ( .A1(n11245), .A2(n14739), .ZN(n14882) );
  NOR2_X1 U14113 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11246) );
  NOR2_X1 U14114 ( .A1(n9649), .A2(n11246), .ZN(n11247) );
  NOR2_X1 U14115 ( .A1(n14882), .A2(n11247), .ZN(n11248) );
  XNOR2_X1 U14116 ( .A(n9649), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14716) );
  NAND2_X1 U14117 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14076) );
  NAND2_X1 U14118 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14862) );
  NAND2_X1 U14119 ( .A1(n9648), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11249) );
  NOR2_X1 U14120 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14687) );
  INV_X1 U14121 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15835) );
  INV_X1 U14122 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14697) );
  NAND2_X1 U14123 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14082) );
  INV_X1 U14124 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14830) );
  NOR2_X1 U14125 ( .A1(n14082), .A2(n14830), .ZN(n14615) );
  NOR2_X1 U14126 ( .A1(n14653), .A2(n9648), .ZN(n14640) );
  AND2_X1 U14127 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14086) );
  INV_X1 U14128 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14837) );
  INV_X1 U14129 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14835) );
  AND3_X1 U14130 ( .A1(n14837), .A2(n14835), .A3(n14830), .ZN(n14616) );
  INV_X1 U14131 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14065) );
  INV_X1 U14132 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14812) );
  NAND2_X1 U14133 ( .A1(n14065), .A2(n14812), .ZN(n14802) );
  NOR2_X1 U14134 ( .A1(n14642), .A2(n14802), .ZN(n11255) );
  INV_X1 U14135 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14091) );
  INV_X1 U14136 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14606) );
  NAND2_X1 U14137 ( .A1(n14091), .A2(n14606), .ZN(n14781) );
  AND2_X1 U14138 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11256) );
  INV_X1 U14139 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14093) );
  INV_X1 U14140 ( .A(n11256), .ZN(n11257) );
  OAI21_X1 U14141 ( .B1(n11270), .B2(n11257), .A(n9971), .ZN(n11258) );
  NAND2_X1 U14142 ( .A1(n11262), .A2(n11258), .ZN(n11261) );
  INV_X1 U14143 ( .A(n11268), .ZN(n11259) );
  NOR4_X1 U14144 ( .A1(n11259), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n9971), .A4(n14781), .ZN(n11260) );
  INV_X1 U14145 ( .A(n11262), .ZN(n11263) );
  INV_X1 U14146 ( .A(n15960), .ZN(n15934) );
  NAND2_X1 U14147 ( .A1(n9971), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11271) );
  NAND3_X1 U14148 ( .A1(n11268), .A2(n14884), .A3(n14606), .ZN(n11269) );
  OAI21_X1 U14149 ( .B1(n11271), .B2(n11270), .A(n11269), .ZN(n11272) );
  NAND2_X1 U14150 ( .A1(n9645), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14777) );
  OAI21_X1 U14151 ( .B1(n14772), .B2(n14291), .A(n14777), .ZN(n11273) );
  AOI21_X1 U14152 ( .B1(n15950), .B2(n14298), .A(n11273), .ZN(n11274) );
  INV_X1 U14153 ( .A(n13179), .ZN(n15793) );
  INV_X1 U14154 ( .A(n13080), .ZN(n11275) );
  NOR2_X1 U14155 ( .A1(n13565), .A2(n11275), .ZN(n11276) );
  NAND2_X1 U14156 ( .A1(n15793), .A2(n11276), .ZN(n13102) );
  NOR4_X1 U14157 ( .A1(n11280), .A2(n11279), .A3(n11278), .A4(n11277), .ZN(
        n11281) );
  NOR2_X1 U14158 ( .A1(n11282), .A2(n11281), .ZN(n12837) );
  NAND2_X1 U14159 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20738) );
  NAND2_X1 U14160 ( .A1(n12837), .A2(n20738), .ZN(n13050) );
  OAI22_X1 U14161 ( .A1(n13126), .A2(n13102), .B1(n13050), .B2(n13326), .ZN(
        n13129) );
  NAND3_X1 U14162 ( .A1(n11283), .A2(n20738), .A3(n10412), .ZN(n11285) );
  INV_X1 U14163 ( .A(n13304), .ZN(n13111) );
  INV_X1 U14164 ( .A(n14525), .ZN(n20224) );
  NAND4_X1 U14165 ( .A1(n13111), .A2(n20224), .A3(n11284), .A4(n10423), .ZN(
        n13026) );
  OAI22_X1 U14166 ( .A1(n13126), .A2(n11285), .B1(n13565), .B2(n13026), .ZN(
        n11286) );
  INV_X1 U14167 ( .A(n20001), .ZN(n13064) );
  OR2_X1 U14168 ( .A1(n14569), .A2(n10409), .ZN(n11299) );
  NOR4_X1 U14169 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11291) );
  NOR4_X1 U14170 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n11290) );
  NOR4_X1 U14171 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11289) );
  NOR4_X1 U14172 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11288) );
  AND4_X1 U14173 ( .A1(n11291), .A2(n11290), .A3(n11289), .A4(n11288), .ZN(
        n11296) );
  NOR4_X1 U14174 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n11294) );
  NOR4_X1 U14175 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n11293) );
  NOR4_X1 U14176 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n11292) );
  INV_X1 U14177 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20749) );
  AND4_X1 U14178 ( .A1(n11294), .A2(n11293), .A3(n11292), .A4(n20749), .ZN(
        n11295) );
  NAND2_X1 U14179 ( .A1(n11296), .A2(n11295), .ZN(n11297) );
  AND2_X2 U14180 ( .A1(n11297), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14535)
         );
  AOI22_X1 U14181 ( .A1(n14589), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14569), .ZN(n11298) );
  INV_X1 U14182 ( .A(n11298), .ZN(n11301) );
  INV_X1 U14183 ( .A(n14535), .ZN(n13519) );
  INV_X1 U14184 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20223) );
  NOR2_X1 U14185 ( .A1(n14573), .A2(n20223), .ZN(n11300) );
  NOR2_X1 U14186 ( .A1(n11301), .A2(n11300), .ZN(n11303) );
  NAND2_X1 U14187 ( .A1(n11303), .A2(n11302), .ZN(P1_U2873) );
  AOI22_X1 U14188 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9663), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11310) );
  AND2_X4 U14189 ( .A1(n13136), .A2(n11304), .ZN(n11544) );
  AND2_X4 U14190 ( .A1(n13134), .A2(n11846), .ZN(n11716) );
  AOI22_X1 U14191 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14192 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11308) );
  AND2_X4 U14193 ( .A1(n11306), .A2(n13812), .ZN(n12037) );
  AOI22_X1 U14194 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11307) );
  NAND4_X1 U14195 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11311) );
  AOI22_X1 U14196 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11544), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14197 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14198 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9641), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14199 ( .A1(n11829), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11312) );
  NAND4_X1 U14200 ( .A1(n11315), .A2(n11314), .A3(n11313), .A4(n11312), .ZN(
        n11316) );
  NAND2_X1 U14201 ( .A1(n11316), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11317) );
  NAND2_X4 U14202 ( .A1(n11318), .A2(n11317), .ZN(n13398) );
  AOI22_X1 U14203 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9631), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14204 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11320) );
  AND2_X1 U14205 ( .A1(n11321), .A2(n11320), .ZN(n11324) );
  AOI22_X1 U14206 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14207 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11322) );
  NAND3_X1 U14208 ( .A1(n11324), .A2(n11323), .A3(n11322), .ZN(n11325) );
  AOI22_X1 U14209 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14210 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14211 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9631), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14212 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11326) );
  NAND4_X1 U14213 ( .A1(n11329), .A2(n11328), .A3(n11327), .A4(n11326), .ZN(
        n11330) );
  INV_X1 U14214 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11334) );
  NOR2_X1 U14215 ( .A1(n11542), .A2(n11334), .ZN(n11500) );
  NAND2_X1 U14216 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11338) );
  NAND2_X1 U14217 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11337) );
  NAND2_X1 U14218 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11336) );
  NAND2_X1 U14219 ( .A1(n11829), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11335) );
  NAND4_X1 U14220 ( .A1(n11338), .A2(n11337), .A3(n11336), .A4(n11335), .ZN(
        n11344) );
  NAND2_X1 U14221 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U14222 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11341) );
  NAND2_X1 U14223 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11340) );
  NAND2_X1 U14224 ( .A1(n11716), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11339) );
  NAND4_X1 U14225 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n11343) );
  NAND2_X1 U14226 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11348) );
  NAND2_X1 U14227 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11347) );
  NAND2_X1 U14228 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U14229 ( .A1(n11829), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11345) );
  NAND4_X1 U14230 ( .A1(n11348), .A2(n11347), .A3(n11346), .A4(n11345), .ZN(
        n11354) );
  NAND2_X1 U14231 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11352) );
  NAND2_X1 U14232 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11351) );
  NAND2_X1 U14233 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11350) );
  NAND2_X1 U14234 ( .A1(n11716), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11349) );
  NAND4_X1 U14235 ( .A1(n11352), .A2(n11351), .A3(n11350), .A4(n11349), .ZN(
        n11353) );
  AOI22_X1 U14236 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9640), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14237 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11716), .B1(
        n11544), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14238 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14239 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11358) );
  NAND2_X1 U14240 ( .A1(n11445), .A2(n11376), .ZN(n11365) );
  AOI22_X1 U14241 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14242 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14243 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14244 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11360) );
  NAND4_X1 U14245 ( .A1(n11363), .A2(n11362), .A3(n11361), .A4(n11360), .ZN(
        n11444) );
  NAND2_X1 U14246 ( .A1(n12923), .A2(n11431), .ZN(n11481) );
  AOI22_X1 U14247 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14248 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14249 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9663), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14250 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11366) );
  NAND4_X1 U14251 ( .A1(n11369), .A2(n11368), .A3(n11367), .A4(n11366), .ZN(
        n11370) );
  NAND2_X1 U14252 ( .A1(n11370), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11379) );
  AOI22_X1 U14253 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14254 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14255 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14256 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11372) );
  NAND4_X1 U14257 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n11377) );
  NAND2_X1 U14258 ( .A1(n11377), .A2(n11376), .ZN(n11378) );
  AND2_X1 U14259 ( .A1(n11421), .A2(n11420), .ZN(n11423) );
  NOR2_X1 U14260 ( .A1(n11481), .A2(n11423), .ZN(n11400) );
  AOI22_X1 U14261 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11544), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14262 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14263 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14264 ( .A1(n11829), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11381) );
  NAND4_X1 U14265 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .ZN(
        n11385) );
  AOI22_X1 U14266 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11544), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14267 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14268 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14269 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11386) );
  NAND4_X1 U14270 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n11390) );
  INV_X1 U14271 ( .A(n11449), .ZN(n19291) );
  NAND2_X2 U14272 ( .A1(n19305), .A2(n11421), .ZN(n11479) );
  AOI22_X1 U14273 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9663), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14274 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14275 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14276 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14277 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14278 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9662), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14279 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14280 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11397) );
  NOR2_X1 U14281 ( .A1(n11418), .A2(n19287), .ZN(n11402) );
  INV_X1 U14282 ( .A(n11419), .ZN(n11401) );
  AND3_X2 U14283 ( .A1(n11402), .A2(n11401), .A3(n11423), .ZN(n11438) );
  INV_X1 U14284 ( .A(n11438), .ZN(n11416) );
  AOI22_X1 U14285 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14286 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14287 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14288 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11403) );
  NAND4_X1 U14289 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11407) );
  AOI22_X1 U14290 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9663), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14291 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14292 ( .A1(n11371), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14293 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11408) );
  NAND4_X1 U14294 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(
        n11412) );
  NAND3_X1 U14295 ( .A1(n11417), .A2(n11416), .A3(n11415), .ZN(n12933) );
  NAND2_X1 U14296 ( .A1(n11479), .A2(n9957), .ZN(n12924) );
  OR2_X1 U14297 ( .A1(n11470), .A2(n19988), .ZN(n11428) );
  NOR2_X1 U14298 ( .A1(n11421), .A2(n12260), .ZN(n11422) );
  NAND2_X1 U14299 ( .A1(n11424), .A2(n11423), .ZN(n12712) );
  NAND2_X1 U14300 ( .A1(n12712), .A2(n10261), .ZN(n11425) );
  NAND2_X1 U14301 ( .A1(n11440), .A2(n11425), .ZN(n11898) );
  INV_X1 U14302 ( .A(n11898), .ZN(n11426) );
  AND3_X2 U14303 ( .A1(n11429), .A2(n11428), .A3(n11427), .ZN(n11476) );
  NAND2_X1 U14304 ( .A1(n11479), .A2(n12923), .ZN(n12048) );
  AND2_X1 U14305 ( .A1(n12048), .A2(n12259), .ZN(n11433) );
  NOR2_X1 U14306 ( .A1(n11479), .A2(n12923), .ZN(n11432) );
  NAND2_X1 U14307 ( .A1(n11433), .A2(n12052), .ZN(n12934) );
  INV_X1 U14308 ( .A(n12927), .ZN(n11434) );
  NAND2_X1 U14309 ( .A1(n11436), .A2(n11435), .ZN(n11472) );
  NAND2_X1 U14310 ( .A1(n11472), .A2(n11477), .ZN(n11437) );
  NAND2_X2 U14311 ( .A1(n11476), .A2(n11437), .ZN(n11488) );
  NOR2_X1 U14312 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19981) );
  INV_X1 U14313 ( .A(n19981), .ZN(n11468) );
  NAND2_X2 U14314 ( .A1(n11438), .A2(n11415), .ZN(n12047) );
  INV_X1 U14315 ( .A(n11484), .ZN(n12928) );
  NOR2_X1 U14316 ( .A1(n13398), .A2(n19988), .ZN(n11450) );
  OAI211_X1 U14317 ( .C1(n19959), .C2(n11468), .A(n11457), .B(n11460), .ZN(
        n11441) );
  INV_X1 U14318 ( .A(n11441), .ZN(n11442) );
  CLKBUF_X3 U14319 ( .A(n11443), .Z(n14206) );
  NAND4_X1 U14320 ( .A1(n9723), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(n11444), .ZN(n11447) );
  NAND4_X1 U14321 ( .A1(n9726), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11376), 
        .A4(n11445), .ZN(n11446) );
  NAND2_X1 U14322 ( .A1(n11447), .A2(n11446), .ZN(n11448) );
  NAND4_X1 U14323 ( .A1(n11480), .A2(n11449), .A3(n19287), .A4(n11448), .ZN(
        n11455) );
  INV_X1 U14324 ( .A(n11450), .ZN(n11451) );
  INV_X1 U14325 ( .A(n12774), .ZN(n11452) );
  NOR2_X1 U14326 ( .A1(n11452), .A2(n13398), .ZN(n11453) );
  NAND2_X1 U14327 ( .A1(n16348), .A2(n11453), .ZN(n11454) );
  OAI21_X1 U14328 ( .B1(n11455), .B2(n12925), .A(n11454), .ZN(n11456) );
  INV_X1 U14329 ( .A(n11456), .ZN(n11458) );
  NAND2_X2 U14330 ( .A1(n11458), .A2(n11457), .ZN(n11903) );
  NAND2_X1 U14331 ( .A1(n9632), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11462) );
  NAND2_X1 U14332 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11461) );
  NAND2_X1 U14333 ( .A1(n11464), .A2(n11463), .ZN(n11465) );
  NAND2_X1 U14334 ( .A1(n9633), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11469) );
  NAND2_X1 U14335 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U14336 ( .A1(n11903), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11474) );
  INV_X1 U14337 ( .A(n11470), .ZN(n11471) );
  NAND2_X1 U14338 ( .A1(n11472), .A2(n11471), .ZN(n11473) );
  NAND4_X1 U14339 ( .A1(n11476), .A2(n11475), .A3(n11474), .A4(n11473), .ZN(
        n11501) );
  AND2_X1 U14340 ( .A1(n11477), .A2(n12928), .ZN(n11478) );
  OAI22_X1 U14341 ( .A1(n11488), .A2(n11478), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11966), .ZN(n11486) );
  INV_X1 U14342 ( .A(n11479), .ZN(n12116) );
  MUX2_X1 U14343 ( .A(n11480), .B(n12116), .S(n19291), .Z(n11483) );
  NOR2_X1 U14344 ( .A1(n12925), .A2(n11481), .ZN(n11482) );
  NAND2_X1 U14345 ( .A1(n11483), .A2(n11482), .ZN(n13809) );
  AOI22_X1 U14346 ( .A1(n13133), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19981), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11485) );
  NAND2_X1 U14347 ( .A1(n11486), .A2(n11485), .ZN(n11502) );
  AOI21_X1 U14348 ( .B1(n19986), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11489) );
  AND2_X1 U14349 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11490) );
  AOI21_X1 U14350 ( .B1(n11908), .B2(P2_REIP_REG_2__SCAN_IN), .A(n11490), .ZN(
        n11493) );
  NAND2_X1 U14351 ( .A1(n11903), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11492) );
  NAND2_X1 U14352 ( .A1(n11966), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11491) );
  NAND2_X1 U14353 ( .A1(n12843), .A2(n11528), .ZN(n11499) );
  NAND2_X1 U14354 ( .A1(n12260), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11494) );
  NOR2_X2 U14355 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19938) );
  NAND2_X1 U14356 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19636) );
  INV_X1 U14357 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19950) );
  NAND2_X1 U14358 ( .A1(n19636), .A2(n19950), .ZN(n11497) );
  NAND2_X1 U14359 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19779) );
  INV_X1 U14360 ( .A(n19779), .ZN(n11495) );
  INV_X1 U14361 ( .A(n11529), .ZN(n11496) );
  AND2_X1 U14362 ( .A1(n11497), .A2(n11496), .ZN(n19406) );
  AOI22_X1 U14363 ( .A1(n11531), .A2(n16308), .B1(n19938), .B2(n19406), .ZN(
        n11498) );
  AOI22_X1 U14364 ( .A1(n11531), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19938), .B2(n19966), .ZN(n11503) );
  NAND2_X1 U14365 ( .A1(n11804), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11511) );
  INV_X1 U14366 ( .A(n11506), .ZN(n11507) );
  XNOR2_X2 U14367 ( .A(n13366), .B(n11507), .ZN(n12867) );
  NAND2_X1 U14368 ( .A1(n11531), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11509) );
  NAND2_X1 U14369 ( .A1(n19966), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14370 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19959), .ZN(
        n19570) );
  NAND2_X1 U14371 ( .A1(n11508), .A2(n19570), .ZN(n19407) );
  NAND2_X1 U14372 ( .A1(n19938), .A2(n19407), .ZN(n19608) );
  NAND2_X1 U14373 ( .A1(n11509), .A2(n19608), .ZN(n11510) );
  INV_X1 U14374 ( .A(n11511), .ZN(n11512) );
  NAND2_X1 U14375 ( .A1(n11488), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11514) );
  NAND2_X1 U14376 ( .A1(n19981), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11513) );
  NAND2_X1 U14377 ( .A1(n11966), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U14378 ( .A1(n11903), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11517) );
  NAND2_X1 U14379 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14380 ( .A1(n11908), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11515) );
  NAND4_X1 U14381 ( .A1(n11518), .A2(n11517), .A3(n11516), .A4(n11515), .ZN(
        n11519) );
  NAND2_X1 U14382 ( .A1(n11520), .A2(n11519), .ZN(n11521) );
  INV_X1 U14383 ( .A(n11920), .ZN(n11522) );
  NAND2_X1 U14384 ( .A1(n11917), .A2(n11522), .ZN(n11523) );
  NAND3_X1 U14385 ( .A1(n11919), .A2(n11526), .A3(n11523), .ZN(n11527) );
  INV_X1 U14386 ( .A(n11523), .ZN(n11525) );
  INV_X1 U14387 ( .A(n11528), .ZN(n12767) );
  NAND2_X1 U14388 ( .A1(n11529), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19786) );
  OAI211_X1 U14389 ( .C1(n11529), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19786), .B(n19938), .ZN(n19674) );
  INV_X1 U14390 ( .A(n19674), .ZN(n11530) );
  AOI21_X1 U14391 ( .B1(n11531), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11530), .ZN(n11532) );
  INV_X1 U14392 ( .A(n11536), .ZN(n11533) );
  NAND2_X1 U14393 ( .A1(n11804), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11534) );
  NAND2_X1 U14394 ( .A1(n11533), .A2(n11534), .ZN(n11537) );
  INV_X1 U14395 ( .A(n11534), .ZN(n11535) );
  NAND2_X1 U14396 ( .A1(n12986), .A2(n12987), .ZN(n12988) );
  NAND2_X1 U14397 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12260), .ZN(
        n11538) );
  INV_X1 U14398 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11541) );
  NOR2_X1 U14399 ( .A1(n11542), .A2(n11541), .ZN(n13459) );
  INV_X1 U14400 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U14401 ( .A1(n12103), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11578), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11548) );
  INV_X1 U14402 ( .A(n11371), .ZN(n11543) );
  AND2_X1 U14403 ( .A1(n11716), .A2(n11376), .ZN(n11556) );
  AOI22_X1 U14404 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14405 ( .A1(n11589), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11546) );
  AND2_X1 U14406 ( .A1(n11716), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11622) );
  AOI22_X1 U14407 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11874), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11545) );
  NAND4_X1 U14408 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n11555) );
  AND2_X2 U14409 ( .A1(n9654), .A2(n11376), .ZN(n12108) );
  AOI22_X1 U14410 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11553) );
  AND2_X1 U14411 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14412 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12160), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14413 ( .A1(n12181), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11551) );
  AND2_X2 U14414 ( .A1(n9641), .A2(n11376), .ZN(n12189) );
  AND2_X1 U14415 ( .A1(n12037), .A2(n11376), .ZN(n12175) );
  AOI22_X1 U14416 ( .A1(n12189), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11550) );
  NAND4_X1 U14417 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11554) );
  AOI22_X1 U14418 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14419 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14420 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11874), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14421 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n11703), .B1(
        n11589), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11557) );
  NAND4_X1 U14422 ( .A1(n11560), .A2(n11559), .A3(n11558), .A4(n11557), .ZN(
        n11566) );
  AOI22_X1 U14423 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14424 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14425 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14426 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12160), .ZN(n11561) );
  NAND4_X1 U14427 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11565) );
  NOR2_X1 U14428 ( .A1(n11566), .A2(n11565), .ZN(n19132) );
  AOI22_X1 U14429 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14430 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14431 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14432 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11567) );
  NAND4_X1 U14433 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11576) );
  AOI22_X1 U14434 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n12175), .ZN(n11574) );
  AOI22_X1 U14435 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14436 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12160), .ZN(n11572) );
  AOI22_X1 U14437 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11571) );
  NAND4_X1 U14438 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11575) );
  AOI22_X1 U14439 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14440 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14441 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14442 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11579) );
  NAND4_X1 U14443 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11588) );
  AOI22_X1 U14444 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14445 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14446 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12160), .ZN(n11584) );
  AOI22_X1 U14447 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11583) );
  NAND4_X1 U14448 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n11587) );
  AOI22_X1 U14449 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11621), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14450 ( .A1(n11578), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14451 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11703), .B1(
        n11589), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14452 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11874), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11590) );
  NAND4_X1 U14453 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n11599) );
  AOI22_X1 U14454 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__4__SCAN_IN), .B2(n12175), .ZN(n11597) );
  AOI22_X1 U14455 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12180), .B1(
        n12189), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14456 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12160), .ZN(n11595) );
  AOI22_X1 U14457 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12181), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11594) );
  NAND4_X1 U14458 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11598) );
  AND2_X2 U14459 ( .A1(n13468), .A2(n12220), .ZN(n13478) );
  AOI22_X1 U14460 ( .A1(n12103), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11578), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14461 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14462 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11589), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14463 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11874), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11600) );
  NAND4_X1 U14464 ( .A1(n11603), .A2(n11602), .A3(n11601), .A4(n11600), .ZN(
        n11609) );
  AOI22_X1 U14465 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14466 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U14467 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12160), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14468 ( .A1(n12189), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11604) );
  NAND4_X1 U14469 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n11608) );
  NOR2_X1 U14470 ( .A1(n11609), .A2(n11608), .ZN(n13476) );
  INV_X1 U14471 ( .A(n13476), .ZN(n11610) );
  AOI22_X1 U14472 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11614) );
  BUF_X1 U14473 ( .A(n11621), .Z(n12119) );
  AOI22_X1 U14474 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14475 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14476 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11611) );
  NAND4_X1 U14477 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(
        n11620) );
  AOI22_X1 U14478 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n12175), .ZN(n11618) );
  AOI22_X1 U14479 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12189), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14480 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12160), .ZN(n11616) );
  AOI22_X1 U14481 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11615) );
  NAND4_X1 U14482 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11619) );
  AOI22_X1 U14483 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14484 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14485 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14486 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14487 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11632) );
  AOI22_X1 U14488 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n12175), .ZN(n11630) );
  AOI22_X1 U14489 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14490 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12160), .ZN(n11628) );
  AOI22_X1 U14491 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11627) );
  NAND4_X1 U14492 ( .A1(n11630), .A2(n11629), .A3(n11628), .A4(n11627), .ZN(
        n11631) );
  OR2_X1 U14493 ( .A1(n11632), .A2(n11631), .ZN(n12229) );
  AOI22_X1 U14494 ( .A1(n12103), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11578), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14495 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14496 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11589), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14497 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11874), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11633) );
  NAND4_X1 U14498 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n11642) );
  AOI22_X1 U14499 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14500 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14501 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12160), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14502 ( .A1(n12189), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11637) );
  NAND4_X1 U14503 ( .A1(n11640), .A2(n11639), .A3(n11638), .A4(n11637), .ZN(
        n11641) );
  OR2_X1 U14504 ( .A1(n11642), .A2(n11641), .ZN(n13961) );
  AOI22_X1 U14505 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14506 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14507 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14508 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11643) );
  NAND4_X1 U14509 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11652) );
  AOI22_X1 U14510 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n12175), .ZN(n11650) );
  AOI22_X1 U14511 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14512 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n12160), .ZN(n11648) );
  AOI22_X1 U14513 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14514 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11651) );
  AOI22_X1 U14515 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14516 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14517 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14518 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11653) );
  NAND4_X1 U14519 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11662) );
  AOI22_X1 U14520 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__2__SCAN_IN), .B2(n12175), .ZN(n11660) );
  AOI22_X1 U14521 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14522 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n12160), .ZN(n11658) );
  AOI22_X1 U14523 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11657) );
  NAND4_X1 U14524 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n11661) );
  NOR2_X1 U14525 ( .A1(n11662), .A2(n11661), .ZN(n16109) );
  AOI22_X1 U14526 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n12103), .B1(
        n11578), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14527 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14528 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n11622), .B1(
        n11589), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14529 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11663) );
  NAND4_X1 U14530 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n11672) );
  AOI22_X1 U14531 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__3__SCAN_IN), .B2(n12175), .ZN(n11670) );
  AOI22_X1 U14532 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14533 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n12160), .ZN(n11668) );
  AOI22_X1 U14534 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11667) );
  NAND4_X1 U14535 ( .A1(n11670), .A2(n11669), .A3(n11668), .A4(n11667), .ZN(
        n11671) );
  NOR2_X1 U14536 ( .A1(n11672), .A2(n11671), .ZN(n15087) );
  AOI22_X1 U14537 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14538 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14539 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14540 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11673) );
  NAND4_X1 U14541 ( .A1(n11676), .A2(n11675), .A3(n11674), .A4(n11673), .ZN(
        n11682) );
  AOI22_X1 U14542 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__4__SCAN_IN), .B2(n12175), .ZN(n11680) );
  AOI22_X1 U14543 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14544 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n12160), .ZN(n11678) );
  AOI22_X1 U14545 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U14546 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11681) );
  OR2_X1 U14547 ( .A1(n11682), .A2(n11681), .ZN(n16105) );
  AOI22_X1 U14548 ( .A1(n12103), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11578), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14549 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14550 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11589), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14551 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11874), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11683) );
  NAND4_X1 U14552 ( .A1(n11686), .A2(n11685), .A3(n11684), .A4(n11683), .ZN(
        n11692) );
  AOI22_X1 U14553 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14554 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14555 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12160), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14556 ( .A1(n12189), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11687) );
  NAND4_X1 U14557 ( .A1(n11690), .A2(n11689), .A3(n11688), .A4(n11687), .ZN(
        n11691) );
  OR2_X1 U14558 ( .A1(n11692), .A2(n11691), .ZN(n15080) );
  AOI22_X1 U14559 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14560 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14561 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14562 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U14563 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11702) );
  AOI22_X1 U14564 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__6__SCAN_IN), .B2(n12175), .ZN(n11700) );
  AOI22_X1 U14565 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14566 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n12160), .ZN(n11698) );
  AOI22_X1 U14567 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11697) );
  NAND4_X1 U14568 ( .A1(n11700), .A2(n11699), .A3(n11698), .A4(n11697), .ZN(
        n11701) );
  NOR2_X1 U14569 ( .A1(n11702), .A2(n11701), .ZN(n16102) );
  AOI22_X1 U14570 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14571 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14572 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14573 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11704) );
  NAND4_X1 U14574 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n11713) );
  AOI22_X1 U14575 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14576 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12160), .ZN(n11710) );
  AOI22_X1 U14577 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12181), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14578 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12189), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11708) );
  NAND4_X1 U14579 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11712) );
  NOR2_X1 U14580 ( .A1(n11713), .A2(n11712), .ZN(n11743) );
  AOI22_X1 U14581 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11714) );
  AND2_X1 U14582 ( .A1(n11715), .A2(n11714), .ZN(n11719) );
  AOI22_X1 U14583 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14584 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11717) );
  XNOR2_X1 U14585 ( .A(n16308), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12030) );
  NAND4_X1 U14586 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n12030), .ZN(
        n11726) );
  AOI22_X1 U14587 ( .A1(n12036), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9639), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11720) );
  AND2_X1 U14588 ( .A1(n11721), .A2(n11720), .ZN(n11724) );
  INV_X1 U14589 ( .A(n12030), .ZN(n12039) );
  AOI22_X1 U14590 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11544), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11723) );
  AOI22_X1 U14591 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11722) );
  NAND4_X1 U14592 ( .A1(n11724), .A2(n12039), .A3(n11723), .A4(n11722), .ZN(
        n11725) );
  NAND2_X1 U14593 ( .A1(n11726), .A2(n11725), .ZN(n11749) );
  NOR2_X1 U14594 ( .A1(n19282), .A2(n11749), .ZN(n11727) );
  XOR2_X1 U14595 ( .A(n11743), .B(n11727), .Z(n11750) );
  XNOR2_X1 U14596 ( .A(n11728), .B(n11729), .ZN(n15125) );
  INV_X1 U14597 ( .A(n11749), .ZN(n11744) );
  NAND2_X1 U14598 ( .A1(n19282), .A2(n11744), .ZN(n15128) );
  INV_X1 U14599 ( .A(n11750), .ZN(n11729) );
  AOI22_X1 U14600 ( .A1(n9654), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14601 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11731) );
  AND2_X1 U14602 ( .A1(n11732), .A2(n11731), .ZN(n11735) );
  AOI22_X1 U14603 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9663), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14604 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11733) );
  NAND4_X1 U14605 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n12030), .ZN(
        n11742) );
  AOI22_X1 U14606 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11736) );
  AND2_X1 U14607 ( .A1(n11737), .A2(n11736), .ZN(n11740) );
  AOI22_X1 U14608 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9662), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14609 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11738) );
  NAND4_X1 U14610 ( .A1(n11740), .A2(n12039), .A3(n11739), .A4(n11738), .ZN(
        n11741) );
  NAND2_X1 U14611 ( .A1(n11742), .A2(n11741), .ZN(n11752) );
  INV_X1 U14612 ( .A(n11743), .ZN(n11745) );
  NAND2_X1 U14613 ( .A1(n11745), .A2(n11744), .ZN(n11753) );
  XOR2_X1 U14614 ( .A(n11752), .B(n11753), .Z(n11746) );
  NAND2_X1 U14615 ( .A1(n11746), .A2(n11804), .ZN(n15073) );
  INV_X1 U14616 ( .A(n15073), .ZN(n11747) );
  INV_X1 U14617 ( .A(n11752), .ZN(n11748) );
  NAND2_X1 U14618 ( .A1(n19282), .A2(n11748), .ZN(n15075) );
  NOR3_X1 U14619 ( .A1(n11750), .A2(n11749), .A3(n15075), .ZN(n11751) );
  NOR2_X1 U14620 ( .A1(n11753), .A2(n11752), .ZN(n11766) );
  AOI22_X1 U14621 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11754) );
  AND2_X1 U14622 ( .A1(n11755), .A2(n11754), .ZN(n11758) );
  AOI22_X1 U14623 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9662), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14624 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11756) );
  NAND4_X1 U14625 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n12030), .ZN(
        n11765) );
  AOI22_X1 U14626 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11759) );
  AND2_X1 U14627 ( .A1(n11760), .A2(n11759), .ZN(n11763) );
  AOI22_X1 U14628 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9663), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14629 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11761) );
  NAND4_X1 U14630 ( .A1(n11763), .A2(n12039), .A3(n11762), .A4(n11761), .ZN(
        n11764) );
  AND2_X1 U14631 ( .A1(n11765), .A2(n11764), .ZN(n11768) );
  NAND2_X1 U14632 ( .A1(n11766), .A2(n11768), .ZN(n11801) );
  OAI211_X1 U14633 ( .C1(n11766), .C2(n11768), .A(n11804), .B(n11801), .ZN(
        n11770) );
  INV_X1 U14634 ( .A(n11770), .ZN(n11767) );
  XNOR2_X1 U14635 ( .A(n11771), .B(n11767), .ZN(n15065) );
  INV_X1 U14636 ( .A(n11768), .ZN(n11769) );
  NOR2_X1 U14637 ( .A1(n13398), .A2(n11769), .ZN(n15067) );
  OR2_X1 U14638 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  AOI22_X1 U14639 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11773) );
  AND2_X1 U14640 ( .A1(n11774), .A2(n11773), .ZN(n11777) );
  AOI22_X1 U14641 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11776) );
  INV_X1 U14642 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n19522) );
  AOI22_X1 U14643 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11775) );
  NAND4_X1 U14644 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n12030), .ZN(
        n11784) );
  AOI22_X1 U14645 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11778) );
  AND2_X1 U14646 ( .A1(n11779), .A2(n11778), .ZN(n11782) );
  AOI22_X1 U14647 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9662), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14648 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11780) );
  NAND4_X1 U14649 ( .A1(n11782), .A2(n12039), .A3(n11781), .A4(n11780), .ZN(
        n11783) );
  AND2_X1 U14650 ( .A1(n11784), .A2(n11783), .ZN(n11799) );
  XNOR2_X1 U14651 ( .A(n11801), .B(n11799), .ZN(n11785) );
  NAND2_X1 U14652 ( .A1(n19282), .A2(n11799), .ZN(n15062) );
  AOI22_X1 U14653 ( .A1(n10149), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14654 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11787) );
  AND2_X1 U14655 ( .A1(n11788), .A2(n11787), .ZN(n11791) );
  AOI22_X1 U14656 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9663), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U14657 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11789) );
  NAND4_X1 U14658 ( .A1(n11791), .A2(n11790), .A3(n11789), .A4(n12030), .ZN(
        n11798) );
  AOI22_X1 U14659 ( .A1(n10149), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11829), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14660 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11792) );
  AND2_X1 U14661 ( .A1(n11793), .A2(n11792), .ZN(n11796) );
  AOI22_X1 U14662 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U14663 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11794) );
  NAND4_X1 U14664 ( .A1(n11796), .A2(n12039), .A3(n11795), .A4(n11794), .ZN(
        n11797) );
  NAND2_X1 U14665 ( .A1(n11798), .A2(n11797), .ZN(n11802) );
  INV_X1 U14666 ( .A(n11802), .ZN(n11810) );
  INV_X1 U14667 ( .A(n11799), .ZN(n11800) );
  OR2_X1 U14668 ( .A1(n11801), .A2(n11800), .ZN(n11803) );
  INV_X1 U14669 ( .A(n11803), .ZN(n11805) );
  OR2_X1 U14670 ( .A1(n11803), .A2(n11802), .ZN(n15046) );
  OAI211_X1 U14671 ( .C1(n11810), .C2(n11805), .A(n15046), .B(n11804), .ZN(
        n11807) );
  INV_X1 U14672 ( .A(n11807), .ZN(n11806) );
  NAND2_X1 U14673 ( .A1(n19282), .A2(n11810), .ZN(n15053) );
  AOI22_X1 U14674 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11811) );
  AND2_X1 U14675 ( .A1(n11812), .A2(n11811), .ZN(n11815) );
  AOI22_X1 U14676 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9631), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14677 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11813) );
  NAND4_X1 U14678 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n12030), .ZN(
        n11822) );
  AOI22_X1 U14679 ( .A1(n10149), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U14680 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11816) );
  AND2_X1 U14681 ( .A1(n11817), .A2(n11816), .ZN(n11820) );
  AOI22_X1 U14682 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14683 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11818) );
  NAND4_X1 U14684 ( .A1(n11820), .A2(n12039), .A3(n11819), .A4(n11818), .ZN(
        n11821) );
  AND2_X1 U14685 ( .A1(n11822), .A2(n11821), .ZN(n15048) );
  NAND2_X1 U14686 ( .A1(n15048), .A2(n13398), .ZN(n11823) );
  NOR2_X1 U14687 ( .A1(n15046), .A2(n11823), .ZN(n11838) );
  AOI22_X1 U14688 ( .A1(n10149), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14689 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11824) );
  AND2_X1 U14690 ( .A1(n11825), .A2(n11824), .ZN(n11828) );
  AOI22_X1 U14691 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11544), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14692 ( .A1(n9662), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11826) );
  NAND4_X1 U14693 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n12030), .ZN(
        n11836) );
  AOI22_X1 U14694 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11830) );
  AND2_X1 U14695 ( .A1(n11831), .A2(n11830), .ZN(n11834) );
  AOI22_X1 U14696 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14697 ( .A1(n9631), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11544), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11832) );
  NAND4_X1 U14698 ( .A1(n11834), .A2(n12039), .A3(n11833), .A4(n11832), .ZN(
        n11835) );
  AND2_X1 U14699 ( .A1(n11836), .A2(n11835), .ZN(n11837) );
  NAND2_X1 U14700 ( .A1(n11838), .A2(n11837), .ZN(n12025) );
  OAI21_X1 U14701 ( .B1(n11838), .B2(n11837), .A(n12025), .ZN(n11840) );
  NAND2_X1 U14702 ( .A1(n11839), .A2(n11840), .ZN(n14268) );
  NAND2_X1 U14703 ( .A1(n19959), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11842) );
  NAND2_X1 U14704 ( .A1(n13812), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11841) );
  NAND2_X1 U14705 ( .A1(n11842), .A2(n11841), .ZN(n11851) );
  NAND2_X1 U14706 ( .A1(n19966), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11850) );
  NAND2_X1 U14707 ( .A1(n16308), .A2(n19950), .ZN(n11843) );
  XNOR2_X1 U14708 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11870) );
  XNOR2_X1 U14709 ( .A(n11871), .B(n11870), .ZN(n12058) );
  OAI21_X1 U14710 ( .B1(n19966), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11850), .ZN(n11849) );
  OAI21_X1 U14711 ( .B1(n11849), .B2(n11851), .A(n12757), .ZN(n11858) );
  INV_X1 U14712 ( .A(n11844), .ZN(n11845) );
  OAI21_X1 U14713 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n11846), .A(
        n11845), .ZN(n11847) );
  XNOR2_X1 U14714 ( .A(n11848), .B(n11847), .ZN(n12059) );
  INV_X1 U14715 ( .A(n11849), .ZN(n12710) );
  NAND2_X1 U14716 ( .A1(n11851), .A2(n11850), .ZN(n12702) );
  AND2_X1 U14717 ( .A1(n11852), .A2(n12702), .ZN(n12061) );
  OAI21_X1 U14718 ( .B1(n13398), .B2(n12710), .A(n12061), .ZN(n11853) );
  OAI21_X1 U14719 ( .B1(n12059), .B2(n13398), .A(n11853), .ZN(n11854) );
  NAND2_X1 U14720 ( .A1(n11854), .A2(n11415), .ZN(n11857) );
  OAI21_X1 U14721 ( .B1(n12774), .B2(n19282), .A(n12059), .ZN(n11856) );
  INV_X1 U14722 ( .A(n12059), .ZN(n11855) );
  AOI22_X1 U14723 ( .A1(n11858), .A2(n11857), .B1(n11856), .B2(n12634), .ZN(
        n11887) );
  AOI22_X1 U14724 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14725 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14726 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14727 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11703), .B1(
        n11874), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11859) );
  NAND4_X1 U14728 ( .A1(n11862), .A2(n11861), .A3(n11860), .A4(n11859), .ZN(
        n11868) );
  AOI22_X1 U14729 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12160), .ZN(n11866) );
  AOI22_X1 U14730 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n12175), .ZN(n11865) );
  AOI22_X1 U14731 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14732 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11863) );
  NAND4_X1 U14733 ( .A1(n11866), .A2(n11865), .A3(n11864), .A4(n11863), .ZN(
        n11867) );
  NOR2_X1 U14734 ( .A1(n11376), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11869) );
  NOR2_X1 U14735 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15862), .ZN(
        n11872) );
  INV_X1 U14736 ( .A(n12060), .ZN(n11873) );
  AOI22_X1 U14737 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14738 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14739 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14740 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n11874), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11875) );
  NAND4_X1 U14741 ( .A1(n11878), .A2(n11877), .A3(n11876), .A4(n11875), .ZN(
        n11884) );
  AOI22_X1 U14742 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12160), .ZN(n11882) );
  AOI22_X1 U14743 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n12175), .ZN(n11881) );
  AOI22_X1 U14744 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14745 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11879) );
  NAND4_X1 U14746 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n11883) );
  INV_X1 U14747 ( .A(n12633), .ZN(n11885) );
  NAND2_X1 U14748 ( .A1(n12639), .A2(n11885), .ZN(n12704) );
  OAI21_X1 U14749 ( .B1(n12058), .B2(n11887), .A(n11886), .ZN(n11893) );
  NAND2_X1 U14750 ( .A1(n12060), .A2(n12757), .ZN(n11892) );
  NAND2_X1 U14751 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15862), .ZN(
        n11888) );
  NAND2_X1 U14752 ( .A1(n11889), .A2(n11888), .ZN(n11891) );
  NAND2_X1 U14753 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12751), .ZN(
        n11890) );
  NAND3_X1 U14754 ( .A1(n11893), .A2(n11892), .A3(n12705), .ZN(n11894) );
  INV_X1 U14755 ( .A(n12705), .ZN(n11895) );
  NAND2_X1 U14756 ( .A1(n11895), .A2(n12774), .ZN(n11896) );
  INV_X1 U14757 ( .A(n16327), .ZN(n11899) );
  INV_X1 U14758 ( .A(n13809), .ZN(n11897) );
  AND2_X1 U14759 ( .A1(n11898), .A2(n11897), .ZN(n16321) );
  NAND2_X1 U14760 ( .A1(n11899), .A2(n16321), .ZN(n12743) );
  INV_X1 U14761 ( .A(n13132), .ZN(n12939) );
  NAND2_X1 U14762 ( .A1(n12743), .A2(n12939), .ZN(n11901) );
  NAND2_X1 U14763 ( .A1(n15593), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19854) );
  INV_X1 U14764 ( .A(n19854), .ZN(n11900) );
  NAND2_X1 U14765 ( .A1(n19148), .A2(n12259), .ZN(n19145) );
  INV_X1 U14766 ( .A(n11908), .ZN(n14261) );
  INV_X1 U14767 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n15199) );
  INV_X1 U14768 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15198) );
  OAI22_X1 U14769 ( .A1(n14261), .A2(n15199), .B1(n15593), .B2(n15198), .ZN(
        n11902) );
  INV_X1 U14770 ( .A(n11902), .ZN(n11906) );
  INV_X1 U14771 ( .A(n11903), .ZN(n11907) );
  INV_X2 U14772 ( .A(n11907), .ZN(n12008) );
  NAND2_X1 U14773 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U14774 ( .A1(n11966), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11904) );
  AND3_X1 U14775 ( .A1(n11906), .A2(n11905), .A3(n11904), .ZN(n14982) );
  NAND2_X1 U14776 ( .A1(n11962), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U14777 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11911) );
  NAND2_X1 U14778 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11910) );
  NAND2_X1 U14779 ( .A1(n14959), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11909) );
  NAND4_X1 U14780 ( .A1(n11912), .A2(n11911), .A3(n11910), .A4(n11909), .ZN(
        n15766) );
  NAND2_X1 U14781 ( .A1(n11962), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11916) );
  NAND2_X1 U14782 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11915) );
  NAND2_X1 U14783 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11914) );
  NAND2_X1 U14784 ( .A1(n14959), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11913) );
  NAND4_X1 U14785 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n16207) );
  NAND2_X1 U14786 ( .A1(n11962), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11926) );
  NAND2_X1 U14787 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11925) );
  NAND2_X1 U14788 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U14789 ( .A1(n14959), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U14790 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n19103) );
  NAND2_X1 U14791 ( .A1(n19104), .A2(n19103), .ZN(n19105) );
  AND2_X1 U14792 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11927) );
  AOI21_X1 U14793 ( .B1(n14959), .B2(P2_REIP_REG_5__SCAN_IN), .A(n11927), .ZN(
        n11930) );
  NAND2_X1 U14794 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11929) );
  NAND2_X1 U14795 ( .A1(n11962), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U14796 ( .A1(n11962), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11934) );
  NAND2_X1 U14797 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U14798 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11932) );
  NAND2_X1 U14799 ( .A1(n14959), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11931) );
  NAND4_X1 U14800 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n13018) );
  AND2_X1 U14801 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11935) );
  AOI21_X1 U14802 ( .B1(n14959), .B2(P2_REIP_REG_7__SCAN_IN), .A(n11935), .ZN(
        n11938) );
  NAND2_X1 U14803 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U14804 ( .A1(n11962), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11936) );
  NAND2_X1 U14805 ( .A1(n11962), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11942) );
  NAND2_X1 U14806 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U14807 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11940) );
  NAND2_X1 U14808 ( .A1(n14959), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11939) );
  NAND4_X1 U14809 ( .A1(n11942), .A2(n11941), .A3(n11940), .A4(n11939), .ZN(
        n13608) );
  AND2_X1 U14810 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11943) );
  AOI21_X1 U14811 ( .B1(n14959), .B2(P2_REIP_REG_9__SCAN_IN), .A(n11943), .ZN(
        n11946) );
  NAND2_X1 U14812 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11945) );
  NAND2_X1 U14813 ( .A1(n11962), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11944) );
  NAND2_X1 U14814 ( .A1(n11962), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11950) );
  NAND2_X1 U14815 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11949) );
  NAND2_X1 U14816 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U14817 ( .A1(n14959), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U14818 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n13465) );
  AND2_X1 U14819 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11951) );
  AOI21_X1 U14820 ( .B1(n14959), .B2(P2_REIP_REG_12__SCAN_IN), .A(n11951), 
        .ZN(n11954) );
  NAND2_X1 U14821 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11953) );
  NAND2_X1 U14822 ( .A1(n11962), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11952) );
  AND2_X1 U14823 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11955) );
  AOI21_X1 U14824 ( .B1(n14959), .B2(P2_REIP_REG_13__SCAN_IN), .A(n11955), 
        .ZN(n11958) );
  NAND2_X1 U14825 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11957) );
  NAND2_X1 U14826 ( .A1(n11962), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11956) );
  INV_X1 U14827 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14171) );
  AOI22_X1 U14828 ( .A1(n14959), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11960) );
  NAND2_X1 U14829 ( .A1(n11962), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11959) );
  OAI211_X1 U14830 ( .C1(n11907), .C2(n14171), .A(n11960), .B(n11959), .ZN(
        n13933) );
  AND2_X1 U14831 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11961) );
  AOI21_X1 U14832 ( .B1(n14959), .B2(P2_REIP_REG_15__SCAN_IN), .A(n11961), 
        .ZN(n11965) );
  NAND2_X1 U14833 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11964) );
  NAND2_X1 U14834 ( .A1(n11962), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11963) );
  NAND2_X1 U14835 ( .A1(n11962), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11970) );
  NAND2_X1 U14836 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11969) );
  NAND2_X1 U14837 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11968) );
  NAND2_X1 U14838 ( .A1(n14959), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11967) );
  NAND4_X1 U14839 ( .A1(n11970), .A2(n11969), .A3(n11968), .A4(n11967), .ZN(
        n13841) );
  INV_X1 U14840 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n11972) );
  INV_X1 U14841 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11971) );
  OAI22_X1 U14842 ( .A1(n14261), .A2(n11972), .B1(n15593), .B2(n11971), .ZN(
        n11973) );
  INV_X1 U14843 ( .A(n11973), .ZN(n11976) );
  NAND2_X1 U14844 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11975) );
  NAND2_X1 U14845 ( .A1(n11962), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11974) );
  INV_X1 U14846 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19899) );
  INV_X1 U14847 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15269) );
  OAI22_X1 U14848 ( .A1(n14261), .A2(n19899), .B1(n15593), .B2(n15269), .ZN(
        n11977) );
  INV_X1 U14849 ( .A(n11977), .ZN(n11980) );
  NAND2_X1 U14850 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11979) );
  NAND2_X1 U14851 ( .A1(n11962), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U14852 ( .A1(n11962), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11984) );
  NAND2_X1 U14853 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11983) );
  NAND2_X1 U14854 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U14855 ( .A1(n14959), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11981) );
  NAND4_X1 U14856 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n15261) );
  INV_X1 U14857 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n11985) );
  INV_X1 U14858 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15246) );
  OAI22_X1 U14859 ( .A1(n14261), .A2(n11985), .B1(n15593), .B2(n15246), .ZN(
        n11986) );
  INV_X1 U14860 ( .A(n11986), .ZN(n11989) );
  NAND2_X1 U14861 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11988) );
  NAND2_X1 U14862 ( .A1(n11962), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11987) );
  INV_X1 U14863 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12243) );
  INV_X1 U14864 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11990) );
  OAI22_X1 U14865 ( .A1(n14261), .A2(n12243), .B1(n15593), .B2(n11990), .ZN(
        n11991) );
  INV_X1 U14866 ( .A(n11991), .ZN(n11994) );
  NAND2_X1 U14867 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11993) );
  NAND2_X1 U14868 ( .A1(n11962), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11992) );
  NAND2_X1 U14869 ( .A1(n11962), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11998) );
  NAND2_X1 U14870 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11997) );
  NAND2_X1 U14871 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U14872 ( .A1(n14959), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11995) );
  NAND2_X1 U14873 ( .A1(n11966), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12002) );
  NAND2_X1 U14874 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12001) );
  NAND2_X1 U14875 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12000) );
  NAND2_X1 U14876 ( .A1(n14959), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11999) );
  NAND4_X1 U14877 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n15000) );
  INV_X1 U14878 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19908) );
  INV_X1 U14879 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16083) );
  OAI22_X1 U14880 ( .A1(n14261), .A2(n19908), .B1(n15593), .B2(n16083), .ZN(
        n12003) );
  INV_X1 U14881 ( .A(n12003), .ZN(n12006) );
  NAND2_X1 U14882 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12005) );
  NAND2_X1 U14883 ( .A1(n11962), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12004) );
  AND3_X1 U14884 ( .A1(n12006), .A2(n12005), .A3(n12004), .ZN(n15068) );
  INV_X1 U14885 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19910) );
  OAI22_X1 U14886 ( .A1(n14261), .A2(n19910), .B1(n15593), .B2(n10124), .ZN(
        n12007) );
  INV_X1 U14887 ( .A(n12007), .ZN(n12011) );
  NAND2_X1 U14888 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12010) );
  NAND2_X1 U14889 ( .A1(n11962), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12009) );
  NAND2_X1 U14890 ( .A1(n11962), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12015) );
  NAND2_X1 U14891 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12014) );
  NAND2_X1 U14892 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12013) );
  NAND2_X1 U14893 ( .A1(n14959), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U14894 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12665) );
  INV_X1 U14895 ( .A(n12020), .ZN(n14985) );
  INV_X1 U14896 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19915) );
  OAI22_X1 U14897 ( .A1(n14261), .A2(n19915), .B1(n15593), .B2(n10125), .ZN(
        n12016) );
  INV_X1 U14898 ( .A(n12016), .ZN(n12019) );
  NAND2_X1 U14899 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12018) );
  NAND2_X1 U14900 ( .A1(n9633), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12017) );
  NAND2_X1 U14901 ( .A1(n12991), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12021) );
  INV_X1 U14902 ( .A(n12025), .ZN(n12026) );
  AOI22_X1 U14903 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9631), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U14904 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12028) );
  NAND2_X1 U14905 ( .A1(n12029), .A2(n12028), .ZN(n12044) );
  AOI22_X1 U14906 ( .A1(n10149), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U14907 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12031) );
  NAND3_X1 U14908 ( .A1(n12032), .A2(n12031), .A3(n12030), .ZN(n12043) );
  AOI22_X1 U14909 ( .A1(n12033), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9663), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U14910 ( .A1(n11544), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11716), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12034) );
  NAND2_X1 U14911 ( .A1(n12035), .A2(n12034), .ZN(n12042) );
  AOI22_X1 U14912 ( .A1(n10149), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U14913 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12038) );
  NAND3_X1 U14914 ( .A1(n12040), .A2(n12039), .A3(n12038), .ZN(n12041) );
  OAI22_X1 U14915 ( .A1(n12044), .A2(n12043), .B1(n12042), .B2(n12041), .ZN(
        n12045) );
  XNOR2_X1 U14916 ( .A(n12046), .B(n12045), .ZN(n14267) );
  NAND2_X1 U14917 ( .A1(n12048), .A2(n19287), .ZN(n12049) );
  NAND2_X1 U14918 ( .A1(n12047), .A2(n12049), .ZN(n12053) );
  NAND2_X1 U14919 ( .A1(n11479), .A2(n12259), .ZN(n12888) );
  NAND2_X1 U14920 ( .A1(n19282), .A2(n19988), .ZN(n12947) );
  INV_X1 U14921 ( .A(n12947), .ZN(n12763) );
  OAI21_X1 U14922 ( .B1(n12888), .B2(n11439), .A(n12763), .ZN(n12935) );
  NOR2_X1 U14923 ( .A1(n11430), .A2(n13398), .ZN(n12054) );
  OAI211_X1 U14924 ( .C1(n12054), .C2(n19988), .A(n19291), .B(n12259), .ZN(
        n12050) );
  NAND2_X1 U14925 ( .A1(n12050), .A2(n19287), .ZN(n12051) );
  NAND4_X1 U14926 ( .A1(n12053), .A2(n12052), .A3(n12935), .A4(n12051), .ZN(
        n12738) );
  INV_X1 U14927 ( .A(n12054), .ZN(n12055) );
  NAND2_X1 U14928 ( .A1(n16327), .A2(n16320), .ZN(n12742) );
  NAND2_X1 U14929 ( .A1(n12927), .A2(n12056), .ZN(n12930) );
  NAND2_X1 U14930 ( .A1(n12742), .A2(n12930), .ZN(n12057) );
  NAND2_X1 U14931 ( .A1(n12057), .A2(n16345), .ZN(n12064) );
  NAND2_X1 U14932 ( .A1(n16348), .A2(n19988), .ZN(n12942) );
  NAND2_X1 U14933 ( .A1(n12942), .A2(n12047), .ZN(n16323) );
  NOR3_X1 U14934 ( .A1(n12060), .A2(n12059), .A3(n12058), .ZN(n12709) );
  NAND2_X1 U14935 ( .A1(n12061), .A2(n12709), .ZN(n12062) );
  NAND2_X1 U14936 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19990) );
  INV_X1 U14937 ( .A(n19990), .ZN(n19985) );
  NOR2_X1 U14938 ( .A1(n12925), .A2(n19985), .ZN(n12739) );
  NAND2_X1 U14939 ( .A1(n18906), .A2(n12739), .ZN(n12063) );
  INV_X1 U14940 ( .A(n12078), .ZN(n12065) );
  NOR4_X1 U14941 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12069) );
  NOR4_X1 U14942 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12068) );
  NOR4_X1 U14943 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12067) );
  NOR4_X1 U14944 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12066) );
  NAND4_X1 U14945 ( .A1(n12069), .A2(n12068), .A3(n12067), .A4(n12066), .ZN(
        n12074) );
  NOR4_X1 U14946 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12072) );
  NOR4_X1 U14947 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12071) );
  NOR4_X1 U14948 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12070) );
  INV_X1 U14949 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19874) );
  NAND4_X1 U14950 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n19874), .ZN(
        n12073) );
  OAI21_X1 U14951 ( .B1(n12074), .B2(n12073), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12075) );
  INV_X1 U14952 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16446) );
  OR2_X1 U14953 ( .A1(n19267), .A2(n16446), .ZN(n12077) );
  NAND2_X1 U14954 ( .A1(n19267), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12076) );
  NAND2_X1 U14955 ( .A1(n12077), .A2(n12076), .ZN(n13744) );
  INV_X1 U14956 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13692) );
  INV_X2 U14957 ( .A(n10263), .ZN(n12211) );
  AND2_X2 U14958 ( .A1(n13398), .A2(n19979), .ZN(n12115) );
  AOI22_X1 U14959 ( .A1(n12211), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12115), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12093) );
  NAND2_X2 U14960 ( .A1(n12079), .A2(n15154), .ZN(n12232) );
  AOI22_X1 U14961 ( .A1(n12103), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11578), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U14962 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U14963 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11589), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U14964 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11874), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12080) );
  NAND4_X1 U14965 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(
        n12091) );
  AOI22_X1 U14966 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U14967 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12088) );
  INV_X1 U14968 ( .A(n12160), .ZN(n12195) );
  INV_X1 U14969 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12084) );
  NOR2_X1 U14970 ( .A1(n12195), .A2(n12084), .ZN(n12085) );
  AOI21_X1 U14971 ( .B1(n12194), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n12085), .ZN(n12087) );
  AOI22_X1 U14972 ( .A1(n12189), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12086) );
  NAND4_X1 U14973 ( .A1(n12089), .A2(n12088), .A3(n12087), .A4(n12086), .ZN(
        n12090) );
  INV_X1 U14974 ( .A(n12641), .ZN(n13672) );
  OR2_X1 U14975 ( .A1(n12232), .A2(n13672), .ZN(n12092) );
  OAI211_X1 U14976 ( .C1(n12257), .C2(n13692), .A(n12093), .B(n12092), .ZN(
        n13689) );
  INV_X1 U14977 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U14978 ( .A1(n12211), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12115), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12096) );
  INV_X1 U14979 ( .A(n13679), .ZN(n12094) );
  OR2_X1 U14980 ( .A1(n12232), .A2(n12094), .ZN(n12095) );
  OAI211_X1 U14981 ( .C1(n12257), .C2(n12097), .A(n12096), .B(n12095), .ZN(
        n13456) );
  INV_X1 U14982 ( .A(n13456), .ZN(n12155) );
  INV_X1 U14983 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13805) );
  INV_X1 U14984 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19210) );
  INV_X1 U14985 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19870) );
  OAI222_X1 U14986 ( .A1(n12146), .A2(n13805), .B1(n10263), .B2(n19210), .C1(
        n12257), .C2(n19870), .ZN(n12131) );
  INV_X1 U14987 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18922) );
  INV_X1 U14988 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12100) );
  INV_X1 U14989 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U14990 ( .A1(n13398), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12099) );
  OAI211_X1 U14991 ( .C1(n12259), .C2(n12100), .A(n19979), .B(n12099), .ZN(
        n12101) );
  INV_X1 U14992 ( .A(n12101), .ZN(n12102) );
  AOI22_X1 U14993 ( .A1(n12103), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11578), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U14994 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U14995 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11589), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U14996 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11874), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12104) );
  NAND4_X1 U14997 ( .A1(n12107), .A2(n12106), .A3(n12105), .A4(n12104), .ZN(
        n12114) );
  AOI22_X1 U14998 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U14999 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U15000 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12160), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15001 ( .A1(n12189), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12109) );
  NAND4_X1 U15002 ( .A1(n12112), .A2(n12111), .A3(n12110), .A4(n12109), .ZN(
        n12113) );
  INV_X1 U15003 ( .A(n12848), .ZN(n12118) );
  MUX2_X1 U15004 ( .A(n12259), .B(n19966), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12117) );
  NAND2_X1 U15005 ( .A1(n12116), .A2(n12115), .ZN(n12144) );
  OAI211_X1 U15006 ( .C1(n12232), .C2(n12118), .A(n12117), .B(n12144), .ZN(
        n12886) );
  XNOR2_X1 U15007 ( .A(n12131), .B(n12132), .ZN(n13151) );
  AOI22_X1 U15008 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11578), .B1(
        n12119), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15009 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15010 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15011 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11703), .B1(
        n11874), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15012 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12129) );
  AOI22_X1 U15013 ( .A1(n12103), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n12188), .ZN(n12127) );
  AOI22_X1 U15014 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12189), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15015 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12160), .ZN(n12125) );
  AOI22_X1 U15016 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12124) );
  NAND4_X1 U15017 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(
        n12128) );
  INV_X1 U15018 ( .A(n12844), .ZN(n12847) );
  MUX2_X1 U15019 ( .A(n12888), .B(n19959), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12130) );
  OAI21_X1 U15020 ( .B1(n12847), .B2(n12232), .A(n12130), .ZN(n13152) );
  NOR2_X1 U15021 ( .A1(n13151), .A2(n13152), .ZN(n13153) );
  NOR2_X1 U15022 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  AOI22_X1 U15023 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15024 ( .A1(n12119), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15025 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n11589), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15026 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11703), .B1(
        n11874), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12134) );
  NAND4_X1 U15027 ( .A1(n12137), .A2(n12136), .A3(n12135), .A4(n12134), .ZN(
        n12143) );
  AOI22_X1 U15028 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n12175), .ZN(n12141) );
  AOI22_X1 U15029 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15030 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12160), .ZN(n12139) );
  AOI22_X1 U15031 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12189), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12138) );
  NAND4_X1 U15032 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n12142) );
  INV_X1 U15033 ( .A(n12846), .ZN(n13422) );
  NAND2_X1 U15034 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12145) );
  OAI211_X1 U15035 ( .C1(n12232), .C2(n13422), .A(n12145), .B(n12144), .ZN(
        n12148) );
  XNOR2_X1 U15036 ( .A(n12149), .B(n12148), .ZN(n13277) );
  INV_X1 U15037 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19872) );
  AOI22_X1 U15038 ( .A1(n12211), .A2(P2_EAX_REG_2__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n12115), .ZN(n12147) );
  OAI21_X1 U15039 ( .B1(n12257), .B2(n19872), .A(n12147), .ZN(n13276) );
  NOR2_X1 U15040 ( .A1(n13277), .A2(n13276), .ZN(n13278) );
  NOR2_X1 U15041 ( .A1(n12149), .A2(n12148), .ZN(n12150) );
  INV_X1 U15042 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13432) );
  NAND2_X1 U15043 ( .A1(n12211), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15044 ( .A1(n12115), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12151) );
  AND2_X1 U15045 ( .A1(n12152), .A2(n12151), .ZN(n12154) );
  OR2_X1 U15046 ( .A1(n12232), .A2(n13354), .ZN(n12153) );
  OAI211_X1 U15047 ( .C1(n12257), .C2(n13432), .A(n12154), .B(n12153), .ZN(
        n13338) );
  AOI22_X1 U15048 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11578), .B1(
        n12103), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15049 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15050 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n11874), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15051 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11703), .B1(
        n11589), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12156) );
  NAND4_X1 U15052 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12167) );
  AOI22_X1 U15053 ( .A1(n12194), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12160), .ZN(n12165) );
  AOI22_X1 U15054 ( .A1(n12108), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12189), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15055 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12180), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15056 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12175), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12162) );
  NAND4_X1 U15057 ( .A1(n12165), .A2(n12164), .A3(n12163), .A4(n12162), .ZN(
        n12166) );
  NOR2_X1 U15058 ( .A1(n12232), .A2(n13888), .ZN(n12168) );
  NAND2_X1 U15059 ( .A1(n14968), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15060 ( .A1(n12211), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12115), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12169) );
  NAND2_X1 U15061 ( .A1(n12103), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12174) );
  NAND2_X1 U15062 ( .A1(n11578), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12173) );
  NAND2_X1 U15063 ( .A1(n11621), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12172) );
  NAND2_X1 U15064 ( .A1(n11556), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12171) );
  INV_X1 U15065 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12178) );
  INV_X1 U15066 ( .A(n12175), .ZN(n12177) );
  INV_X1 U15067 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12176) );
  OAI22_X1 U15068 ( .A1(n12179), .A2(n12178), .B1(n12177), .B2(n12176), .ZN(
        n12187) );
  INV_X1 U15069 ( .A(n12180), .ZN(n12185) );
  INV_X1 U15070 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12184) );
  INV_X1 U15071 ( .A(n12181), .ZN(n12183) );
  INV_X1 U15072 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12182) );
  OAI22_X1 U15073 ( .A1(n12185), .A2(n12184), .B1(n12183), .B2(n12182), .ZN(
        n12186) );
  NOR2_X1 U15074 ( .A1(n12187), .A2(n12186), .ZN(n12206) );
  INV_X1 U15075 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12193) );
  INV_X1 U15076 ( .A(n12188), .ZN(n12192) );
  INV_X1 U15077 ( .A(n12189), .ZN(n12191) );
  INV_X1 U15078 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12190) );
  OAI22_X1 U15079 ( .A1(n12193), .A2(n12192), .B1(n12191), .B2(n12190), .ZN(
        n12200) );
  INV_X1 U15080 ( .A(n12194), .ZN(n12198) );
  INV_X1 U15081 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12197) );
  OAI22_X1 U15082 ( .A1(n12198), .A2(n12197), .B1(n12196), .B2(n12195), .ZN(
        n12199) );
  NOR2_X1 U15083 ( .A1(n12200), .A2(n12199), .ZN(n12205) );
  NAND2_X1 U15084 ( .A1(n11874), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12204) );
  NAND2_X1 U15085 ( .A1(n11589), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12203) );
  NAND2_X1 U15086 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12202) );
  NAND2_X1 U15087 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12201) );
  INV_X1 U15088 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15568) );
  INV_X1 U15089 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19197) );
  INV_X1 U15090 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19879) );
  OAI222_X1 U15091 ( .A1(n12146), .A2(n15568), .B1(n10263), .B2(n19197), .C1(
        n12257), .C2(n19879), .ZN(n13032) );
  INV_X1 U15092 ( .A(n12208), .ZN(n19140) );
  AOI22_X1 U15093 ( .A1(n12211), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12115), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12209) );
  OAI21_X1 U15094 ( .B1(n19140), .B2(n12232), .A(n12209), .ZN(n12210) );
  AOI21_X1 U15095 ( .B1(n14968), .B2(P2_REIP_REG_8__SCAN_IN), .A(n12210), .ZN(
        n13606) );
  AOI22_X1 U15096 ( .A1(n14968), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n12211), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12214) );
  INV_X1 U15097 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15558) );
  OAI22_X1 U15098 ( .A1(n12232), .A2(n19133), .B1(n12146), .B2(n15558), .ZN(
        n12212) );
  INV_X1 U15099 ( .A(n12212), .ZN(n12213) );
  NAND2_X1 U15100 ( .A1(n12214), .A2(n12213), .ZN(n15556) );
  AOI22_X1 U15101 ( .A1(n12211), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12115), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12215) );
  OAI21_X1 U15102 ( .B1(n19132), .B2(n12232), .A(n12215), .ZN(n12216) );
  AOI21_X1 U15103 ( .B1(n14968), .B2(P2_REIP_REG_10__SCAN_IN), .A(n12216), 
        .ZN(n16264) );
  INV_X1 U15104 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15105 ( .A1(n12211), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12115), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12218) );
  OR2_X1 U15106 ( .A1(n12232), .A2(n13470), .ZN(n12217) );
  OAI211_X1 U15107 ( .C1(n12257), .C2(n12219), .A(n12218), .B(n12217), .ZN(
        n13298) );
  INV_X1 U15108 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15109 ( .A1(n12211), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12115), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12222) );
  INV_X1 U15110 ( .A(n12220), .ZN(n19125) );
  OR2_X1 U15111 ( .A1(n12232), .A2(n19125), .ZN(n12221) );
  OAI211_X1 U15112 ( .C1(n12257), .C2(n12223), .A(n12222), .B(n12221), .ZN(
        n15038) );
  INV_X1 U15113 ( .A(n15038), .ZN(n12224) );
  NAND2_X1 U15114 ( .A1(n14968), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15115 ( .A1(n12211), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12115), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12225) );
  OAI211_X1 U15116 ( .C1(n13476), .C2(n12232), .A(n12226), .B(n12225), .ZN(
        n13544) );
  INV_X1 U15117 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U15118 ( .A1(n12211), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12115), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12228) );
  INV_X1 U15119 ( .A(n19121), .ZN(n13632) );
  OR2_X1 U15120 ( .A1(n12232), .A2(n13632), .ZN(n12227) );
  OAI211_X1 U15121 ( .C1(n12257), .C2(n13936), .A(n12228), .B(n12227), .ZN(
        n13747) );
  INV_X1 U15122 ( .A(n12229), .ZN(n13631) );
  NAND2_X1 U15123 ( .A1(n14968), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15124 ( .A1(n12211), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12115), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12230) );
  OAI211_X1 U15125 ( .C1(n13631), .C2(n12232), .A(n12231), .B(n12230), .ZN(
        n13820) );
  NAND2_X1 U15126 ( .A1(n14968), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15127 ( .A1(n12211), .A2(P2_EAX_REG_16__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n12115), .ZN(n12233) );
  INV_X1 U15128 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19896) );
  AOI22_X1 U15129 ( .A1(n12211), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12115), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12235) );
  OAI21_X1 U15130 ( .B1(n12257), .B2(n19896), .A(n12235), .ZN(n13953) );
  NAND2_X1 U15131 ( .A1(n13952), .A2(n13953), .ZN(n15487) );
  NAND2_X1 U15132 ( .A1(n14968), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15133 ( .A1(n12211), .A2(P2_EAX_REG_18__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n12115), .ZN(n12236) );
  AOI22_X1 U15134 ( .A1(n12211), .A2(P2_EAX_REG_19__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n12115), .ZN(n12238) );
  OAI21_X1 U15135 ( .B1(n12257), .B2(n19899), .A(n12238), .ZN(n15143) );
  INV_X1 U15136 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15137 ( .A1(n12211), .A2(P2_EAX_REG_20__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n12115), .ZN(n12239) );
  OAI21_X1 U15138 ( .B1(n12257), .B2(n12240), .A(n12239), .ZN(n15441) );
  AOI22_X1 U15139 ( .A1(n12211), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12115), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12241) );
  OAI21_X1 U15140 ( .B1(n12257), .B2(n11985), .A(n12241), .ZN(n12686) );
  AOI22_X1 U15141 ( .A1(n12211), .A2(P2_EAX_REG_22__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n12115), .ZN(n12242) );
  OAI21_X1 U15142 ( .B1(n12257), .B2(n12243), .A(n12242), .ZN(n15416) );
  INV_X1 U15143 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19904) );
  AOI22_X1 U15144 ( .A1(n12211), .A2(P2_EAX_REG_23__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n12115), .ZN(n12244) );
  OAI21_X1 U15145 ( .B1(n12257), .B2(n19904), .A(n12244), .ZN(n15013) );
  NAND2_X1 U15146 ( .A1(n14968), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15147 ( .A1(n12211), .A2(P2_EAX_REG_24__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n12115), .ZN(n12245) );
  AND2_X1 U15148 ( .A1(n12246), .A2(n12245), .ZN(n15003) );
  NAND2_X1 U15149 ( .A1(n14968), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15150 ( .A1(n12211), .A2(P2_EAX_REG_25__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n12115), .ZN(n12247) );
  AND2_X1 U15151 ( .A1(n12248), .A2(n12247), .ZN(n15110) );
  AOI22_X1 U15152 ( .A1(n12211), .A2(P2_EAX_REG_26__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n12115), .ZN(n12249) );
  OAI21_X1 U15153 ( .B1(n12257), .B2(n19910), .A(n12249), .ZN(n15103) );
  NAND2_X1 U15154 ( .A1(n14968), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15155 ( .A1(n12211), .A2(P2_EAX_REG_27__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n12115), .ZN(n12250) );
  AND2_X1 U15156 ( .A1(n12251), .A2(n12250), .ZN(n12671) );
  NAND2_X1 U15157 ( .A1(n14968), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15158 ( .A1(n12211), .A2(P2_EAX_REG_28__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n12115), .ZN(n12252) );
  AND2_X1 U15159 ( .A1(n12253), .A2(n12252), .ZN(n14986) );
  NAND2_X1 U15160 ( .A1(n14968), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15161 ( .A1(n12211), .A2(P2_EAX_REG_29__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n12115), .ZN(n12254) );
  AND2_X1 U15162 ( .A1(n12255), .A2(n12254), .ZN(n14239) );
  INV_X1 U15163 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19918) );
  AOI22_X1 U15164 ( .A1(n12211), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12115), .ZN(n12256) );
  OAI21_X1 U15165 ( .B1(n12257), .B2(n19918), .A(n12256), .ZN(n14966) );
  XNOR2_X1 U15166 ( .A(n14967), .B(n14966), .ZN(n16057) );
  OR2_X1 U15167 ( .A1(n19169), .A2(n12259), .ZN(n16119) );
  INV_X1 U15168 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12777) );
  OAI22_X1 U15169 ( .A1(n16057), .A2(n16119), .B1(n15130), .B2(n12777), .ZN(
        n12258) );
  AOI21_X1 U15170 ( .B1(n16127), .B2(n13744), .A(n12258), .ZN(n12263) );
  NAND3_X1 U15171 ( .A1(n15130), .A2(n12260), .A3(n12259), .ZN(n12261) );
  NOR2_X2 U15172 ( .A1(n12261), .A2(n19267), .ZN(n19153) );
  NOR2_X2 U15173 ( .A1(n12261), .A2(n19269), .ZN(n19152) );
  AOI22_X1 U15174 ( .A1(n19153), .A2(BUF1_REG_30__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n12262) );
  OAI21_X1 U15175 ( .B1(n14267), .B2(n16120), .A(n12264), .ZN(P2_U2889) );
  INV_X1 U15176 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16944) );
  AOI22_X1 U15177 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12265) );
  OAI21_X1 U15178 ( .B1(n10251), .B2(n16944), .A(n12265), .ZN(n12282) );
  INV_X1 U15180 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12280) );
  INV_X1 U15181 ( .A(n12266), .ZN(n12296) );
  AOI22_X1 U15182 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12279) );
  NAND2_X1 U15183 ( .A1(n18852), .A2(n18841), .ZN(n12267) );
  INV_X1 U15184 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17098) );
  INV_X1 U15185 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16933) );
  OAI22_X1 U15186 ( .A1(n21028), .A2(n17098), .B1(n17133), .B2(n16933), .ZN(
        n12277) );
  AOI22_X1 U15187 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15188 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15190 ( .A1(n9659), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12273) );
  NAND3_X1 U15191 ( .A1(n12275), .A2(n12274), .A3(n12273), .ZN(n12276) );
  AOI211_X1 U15192 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n12277), .B(n12276), .ZN(n12278) );
  OAI211_X1 U15193 ( .C1(n12307), .C2(n12280), .A(n12279), .B(n12278), .ZN(
        n12281) );
  INV_X1 U15194 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U15195 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15196 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12284) );
  OAI211_X1 U15197 ( .C1(n15668), .C2(n16999), .A(n12285), .B(n12284), .ZN(
        n12294) );
  INV_X1 U15198 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17008) );
  INV_X4 U15199 ( .A(n9695), .ZN(n15698) );
  AOI22_X1 U15200 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12292) );
  INV_X1 U15201 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U15202 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12287) );
  OAI21_X1 U15203 ( .B1(n17168), .B2(n17242), .A(n12287), .ZN(n12290) );
  INV_X1 U15204 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15205 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12288) );
  OAI21_X1 U15206 ( .B1(n17133), .B2(n12481), .A(n12288), .ZN(n12289) );
  AOI211_X1 U15207 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n12290), .B(n12289), .ZN(n12291) );
  OAI211_X1 U15208 ( .C1(n10251), .C2(n17008), .A(n12292), .B(n12291), .ZN(
        n12293) );
  INV_X1 U15209 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17032) );
  INV_X2 U15210 ( .A(n10251), .ZN(n17030) );
  AOI22_X1 U15211 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12266), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15212 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12297) );
  OAI211_X1 U15213 ( .C1(n15668), .C2(n17032), .A(n12298), .B(n12297), .ZN(
        n12306) );
  INV_X2 U15214 ( .A(n17080), .ZN(n17044) );
  AOI22_X1 U15215 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15216 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12304) );
  INV_X2 U15217 ( .A(n10258), .ZN(n17192) );
  INV_X1 U15218 ( .A(n12299), .ZN(n12302) );
  INV_X1 U15219 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U15220 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12300) );
  OAI21_X1 U15221 ( .B1(n17181), .B2(n17034), .A(n12300), .ZN(n12301) );
  AOI211_X1 U15222 ( .C1(n17186), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n12302), .B(n12301), .ZN(n12303) );
  INV_X1 U15223 ( .A(n12307), .ZN(n17086) );
  AOI22_X1 U15224 ( .A1(n15626), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12309), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12310) );
  INV_X1 U15225 ( .A(n12310), .ZN(n12315) );
  AOI22_X1 U15226 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12323), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15227 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15228 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12311) );
  NAND3_X1 U15229 ( .A1(n12313), .A2(n12312), .A3(n12311), .ZN(n12314) );
  AOI211_X1 U15230 ( .C1(n17086), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n12315), .B(n12314), .ZN(n12322) );
  INV_X1 U15231 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17261) );
  INV_X2 U15232 ( .A(n10260), .ZN(n17216) );
  AOI22_X1 U15233 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12316) );
  OAI21_X1 U15234 ( .B1(n17168), .B2(n17261), .A(n12316), .ZN(n12320) );
  AOI22_X1 U15235 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12318) );
  NAND3_X1 U15236 ( .A1(n12318), .A2(n10254), .A3(n12317), .ZN(n12319) );
  INV_X1 U15237 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15625) );
  AOI22_X1 U15238 ( .A1(n15626), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12333) );
  INV_X1 U15239 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15240 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12323), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15241 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12324) );
  OAI211_X1 U15242 ( .C1(n15668), .C2(n12326), .A(n12325), .B(n12324), .ZN(
        n12332) );
  AOI22_X1 U15243 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15244 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15245 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U15246 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12327) );
  NAND4_X1 U15247 ( .A1(n12330), .A2(n12329), .A3(n12328), .A4(n12327), .ZN(
        n12331) );
  NAND2_X1 U15248 ( .A1(n17418), .A2(n12536), .ZN(n12374) );
  INV_X1 U15249 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15250 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12344) );
  INV_X1 U15251 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U15252 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15253 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12266), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12335) );
  OAI211_X1 U15254 ( .C1(n17215), .C2(n17132), .A(n12336), .B(n12335), .ZN(
        n12342) );
  INV_X2 U15255 ( .A(n10251), .ZN(n17173) );
  AOI22_X1 U15256 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15257 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15258 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12338) );
  NAND2_X1 U15259 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12337) );
  NAND4_X1 U15260 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(
        n12341) );
  AOI211_X1 U15261 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n12342), .B(n12341), .ZN(n12343) );
  OAI211_X1 U15262 ( .C1(n16984), .C2(n12345), .A(n12344), .B(n12343), .ZN(
        n12537) );
  NAND2_X1 U15263 ( .A1(n12376), .A2(n12537), .ZN(n12357) );
  INV_X1 U15264 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U15265 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15266 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15267 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12346) );
  OAI211_X1 U15268 ( .C1(n17215), .C2(n17123), .A(n12347), .B(n12346), .ZN(
        n12353) );
  AOI22_X1 U15269 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15270 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9657), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15271 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12349) );
  NAND2_X1 U15272 ( .A1(n9659), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12348) );
  NAND4_X1 U15273 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12352) );
  AOI211_X1 U15274 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n12353), .B(n12352), .ZN(n12354) );
  OAI211_X1 U15275 ( .C1(n12307), .C2(n17114), .A(n12355), .B(n12354), .ZN(
        n12538) );
  NAND2_X1 U15276 ( .A1(n12383), .A2(n12538), .ZN(n12386) );
  NAND3_X1 U15277 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17813), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12356) );
  INV_X1 U15278 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18843) );
  NAND2_X1 U15279 ( .A1(n18843), .A2(n10010), .ZN(n12409) );
  NAND2_X1 U15280 ( .A1(n12356), .A2(n12409), .ZN(n12412) );
  INV_X1 U15281 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18029) );
  INV_X1 U15282 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18048) );
  INV_X1 U15283 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18057) );
  INV_X1 U15284 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18120) );
  INV_X1 U15285 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18104) );
  NOR2_X1 U15286 ( .A1(n18120), .A2(n18104), .ZN(n17772) );
  NAND2_X1 U15287 ( .A1(n17772), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18077) );
  INV_X1 U15288 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18081) );
  NOR2_X1 U15289 ( .A1(n18077), .A2(n18081), .ZN(n17734) );
  NAND2_X1 U15290 ( .A1(n17734), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18053) );
  OR2_X1 U15291 ( .A1(n18057), .A2(n18053), .ZN(n18037) );
  NOR2_X1 U15292 ( .A1(n18048), .A2(n18037), .ZN(n16406) );
  INV_X1 U15293 ( .A(n16406), .ZN(n18011) );
  XOR2_X1 U15294 ( .A(n12357), .B(n17401), .Z(n12379) );
  INV_X1 U15295 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18201) );
  OR2_X1 U15296 ( .A1(n18201), .A2(n12358), .ZN(n12372) );
  NAND2_X1 U15297 ( .A1(n12535), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12371) );
  INV_X2 U15298 ( .A(n10260), .ZN(n17194) );
  AOI22_X1 U15299 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12359) );
  OAI21_X1 U15300 ( .B1(n17168), .B2(n17214), .A(n12359), .ZN(n12364) );
  AOI22_X1 U15301 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15302 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15303 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12360) );
  NAND3_X1 U15304 ( .A1(n12362), .A2(n12361), .A3(n12360), .ZN(n12363) );
  AOI211_X1 U15305 ( .C1(n12266), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n12364), .B(n12363), .ZN(n12370) );
  INV_X1 U15306 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15638) );
  INV_X1 U15307 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17078) );
  OAI22_X1 U15308 ( .A1(n17133), .A2(n15638), .B1(n15668), .B2(n17078), .ZN(
        n12368) );
  AOI22_X1 U15309 ( .A1(n17086), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12366) );
  INV_X1 U15310 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17226) );
  NAND3_X1 U15311 ( .A1(n12366), .A2(n10253), .A3(n12365), .ZN(n12367) );
  INV_X1 U15312 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18863) );
  NOR2_X1 U15313 ( .A1(n17899), .A2(n18863), .ZN(n17898) );
  INV_X1 U15314 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18842) );
  NAND2_X1 U15315 ( .A1(n12371), .A2(n17889), .ZN(n17878) );
  NAND2_X1 U15316 ( .A1(n17879), .A2(n17878), .ZN(n17877) );
  NAND2_X1 U15317 ( .A1(n12372), .A2(n17877), .ZN(n12373) );
  NAND2_X1 U15318 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12373), .ZN(
        n12375) );
  INV_X1 U15319 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18177) );
  XNOR2_X1 U15320 ( .A(n18177), .B(n12373), .ZN(n17871) );
  XOR2_X1 U15321 ( .A(n12374), .B(n17408), .Z(n17870) );
  NAND2_X1 U15322 ( .A1(n17871), .A2(n17870), .ZN(n17869) );
  NAND2_X1 U15323 ( .A1(n12375), .A2(n17869), .ZN(n17856) );
  INV_X1 U15324 ( .A(n12537), .ZN(n17405) );
  XOR2_X1 U15325 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12377), .Z(
        n17857) );
  NAND2_X1 U15326 ( .A1(n17856), .A2(n17857), .ZN(n17855) );
  NAND2_X1 U15327 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12377), .ZN(
        n12378) );
  NAND2_X1 U15328 ( .A1(n12379), .A2(n12381), .ZN(n12382) );
  NAND2_X1 U15329 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17849), .ZN(
        n17848) );
  NAND2_X1 U15330 ( .A1(n12382), .A2(n17848), .ZN(n17834) );
  INV_X1 U15331 ( .A(n12538), .ZN(n17398) );
  XNOR2_X1 U15332 ( .A(n12383), .B(n17398), .ZN(n12384) );
  XOR2_X1 U15333 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12384), .Z(
        n17835) );
  NAND2_X1 U15334 ( .A1(n17834), .A2(n17835), .ZN(n17833) );
  NAND2_X1 U15335 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12384), .ZN(
        n12385) );
  AOI21_X1 U15336 ( .B1(n17394), .B2(n12386), .A(n17813), .ZN(n12389) );
  NAND2_X1 U15337 ( .A1(n12389), .A2(n12388), .ZN(n12390) );
  NOR4_X1 U15338 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12393) );
  INV_X1 U15339 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17747) );
  NAND4_X1 U15340 ( .A1(n12393), .A2(n18081), .A3(n17747), .A4(n18048), .ZN(
        n12394) );
  OAI221_X2 U15341 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n10010), 
        .C1(n18029), .C2(n12396), .A(n12398), .ZN(n17685) );
  INV_X1 U15342 ( .A(n12396), .ZN(n12397) );
  NAND2_X1 U15343 ( .A1(n12398), .A2(n12397), .ZN(n17694) );
  INV_X1 U15344 ( .A(n17694), .ZN(n17631) );
  INV_X1 U15345 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18008) );
  NOR2_X1 U15346 ( .A1(n18029), .A2(n18008), .ZN(n16369) );
  INV_X1 U15347 ( .A(n16369), .ZN(n18005) );
  INV_X1 U15348 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17618) );
  INV_X1 U15349 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18017) );
  NAND2_X1 U15350 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17981) );
  INV_X1 U15351 ( .A(n17981), .ZN(n17641) );
  NAND2_X1 U15352 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17641), .ZN(
        n17969) );
  NOR2_X1 U15353 ( .A1(n18017), .A2(n17969), .ZN(n16368) );
  NAND2_X1 U15354 ( .A1(n16368), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17606) );
  OR2_X1 U15355 ( .A1(n17618), .A2(n17606), .ZN(n12402) );
  NOR2_X1 U15356 ( .A1(n18005), .A2(n12402), .ZN(n17951) );
  INV_X1 U15357 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18001) );
  NAND2_X1 U15358 ( .A1(n17675), .A2(n18001), .ZN(n12399) );
  NOR2_X1 U15359 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12399), .ZN(
        n17640) );
  INV_X1 U15360 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17982) );
  NAND2_X1 U15361 ( .A1(n17640), .A2(n17982), .ZN(n17630) );
  NOR2_X1 U15362 ( .A1(n12404), .A2(n10010), .ZN(n17590) );
  INV_X1 U15363 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17927) );
  NAND2_X1 U15364 ( .A1(n10010), .A2(n17591), .ZN(n12403) );
  OAI221_X1 U15365 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n10010), 
        .C1(n17927), .C2(n12404), .A(n12403), .ZN(n17564) );
  INV_X1 U15366 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16416) );
  NAND2_X1 U15367 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15750) );
  INV_X1 U15368 ( .A(n15750), .ZN(n16372) );
  NAND2_X1 U15369 ( .A1(n16372), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15846) );
  INV_X1 U15370 ( .A(n12407), .ZN(n15843) );
  NAND2_X1 U15371 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18843), .ZN(
        n16393) );
  OAI211_X1 U15372 ( .C1(n17813), .C2(n12405), .A(n15843), .B(n16393), .ZN(
        n12411) );
  OAI22_X1 U15373 ( .A1(n18859), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18693), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12522) );
  NAND2_X1 U15374 ( .A1(n18469), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12521) );
  NOR2_X1 U15375 ( .A1(n12522), .A2(n12521), .ZN(n12413) );
  AOI21_X1 U15376 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18693), .A(
        n12413), .ZN(n12419) );
  AOI22_X1 U15377 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18698), .B2(n18852), .ZN(
        n12418) );
  NOR2_X1 U15378 ( .A1(n12419), .A2(n12418), .ZN(n12414) );
  AOI21_X1 U15379 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18698), .A(
        n12414), .ZN(n12415) );
  AOI22_X1 U15380 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18719), .B1(
        n12415), .B2(n18841), .ZN(n12422) );
  NOR2_X1 U15381 ( .A1(n12415), .A2(n18841), .ZN(n12421) );
  NAND2_X1 U15382 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18719), .ZN(
        n12416) );
  OAI22_X1 U15383 ( .A1(n12422), .A2(n18701), .B1(n12421), .B2(n12416), .ZN(
        n12417) );
  INV_X1 U15384 ( .A(n12417), .ZN(n12420) );
  OAI211_X1 U15385 ( .C1(n18469), .C2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12521), .B(n12420), .ZN(n12520) );
  XOR2_X1 U15386 ( .A(n12419), .B(n12418), .Z(n12527) );
  NAND2_X1 U15387 ( .A1(n12420), .A2(n12527), .ZN(n12525) );
  INV_X1 U15388 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18702) );
  OR2_X1 U15389 ( .A1(n12421), .A2(n18701), .ZN(n12423) );
  AOI22_X1 U15390 ( .A1(n18702), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n12423), .B2(n12422), .ZN(n12523) );
  OAI211_X1 U15391 ( .C1(n12522), .C2(n12520), .A(n12525), .B(n12523), .ZN(
        n12424) );
  INV_X1 U15392 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U15393 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9657), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12425) );
  OAI21_X1 U15394 ( .B1(n10251), .B2(n17203), .A(n12425), .ZN(n12430) );
  AOI22_X1 U15395 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12428) );
  INV_X1 U15396 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12426) );
  OAI22_X1 U15397 ( .A1(n17172), .A2(n17063), .B1(n10260), .B2(n12426), .ZN(
        n12427) );
  INV_X4 U15398 ( .A(n17181), .ZN(n17191) );
  INV_X2 U15399 ( .A(n17190), .ZN(n17165) );
  AOI211_X4 U15400 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n12430), .B(n12429), .ZN(n18884) );
  INV_X1 U15401 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U15402 ( .A1(n15626), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n9646), .ZN(n12431) );
  OAI21_X1 U15403 ( .B1(n17104), .B2(n17181), .A(n12431), .ZN(n12438) );
  AOI22_X1 U15404 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12437) );
  INV_X1 U15405 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U15406 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17086), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17151), .ZN(n12432) );
  OAI21_X1 U15407 ( .B1(n17097), .B2(n17168), .A(n12432), .ZN(n12436) );
  INV_X1 U15408 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U15409 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n15698), .ZN(n12434) );
  AOI22_X1 U15410 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17194), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12433) );
  OAI211_X1 U15411 ( .C1(n16934), .C2(n15668), .A(n12434), .B(n12433), .ZN(
        n12435) );
  AOI22_X1 U15412 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12448) );
  INV_X1 U15413 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U15414 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15415 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12439) );
  OAI211_X1 U15416 ( .C1(n15668), .C2(n17079), .A(n12440), .B(n12439), .ZN(
        n12446) );
  AOI22_X1 U15417 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15418 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U15419 ( .A1(n15626), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U15420 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12441) );
  NAND4_X1 U15421 ( .A1(n12444), .A2(n12443), .A3(n12442), .A4(n12441), .ZN(
        n12445) );
  INV_X1 U15422 ( .A(n12506), .ZN(n12503) );
  INV_X1 U15423 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U15424 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17169), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12458) );
  INV_X1 U15425 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U15426 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15427 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12449) );
  OAI211_X1 U15428 ( .C1(n15668), .C2(n17160), .A(n12450), .B(n12449), .ZN(
        n12456) );
  AOI22_X1 U15429 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9657), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15430 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15431 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12452) );
  NAND2_X1 U15432 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12451) );
  NAND4_X1 U15433 ( .A1(n12454), .A2(n12453), .A3(n12452), .A4(n12451), .ZN(
        n12455) );
  AOI211_X1 U15434 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n12456), .B(n12455), .ZN(n12457) );
  INV_X1 U15435 ( .A(n12514), .ZN(n18249) );
  INV_X1 U15436 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U15437 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17169), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12468) );
  INV_X1 U15438 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U15439 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15440 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12459) );
  OAI211_X1 U15441 ( .C1(n17215), .C2(n17180), .A(n12460), .B(n12459), .ZN(
        n12466) );
  AOI22_X1 U15442 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15443 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15444 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U15445 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12461) );
  NAND4_X1 U15446 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(
        n12465) );
  AOI211_X1 U15447 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n12466), .B(n12465), .ZN(n12467) );
  NAND2_X1 U15448 ( .A1(n18249), .A2(n18244), .ZN(n18667) );
  INV_X1 U15449 ( .A(n18667), .ZN(n12490) );
  INV_X1 U15450 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U15451 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12469) );
  OAI21_X1 U15452 ( .B1(n10260), .B2(n17116), .A(n12469), .ZN(n12478) );
  INV_X1 U15453 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16925) );
  AOI22_X1 U15454 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15455 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12470) );
  OAI21_X1 U15456 ( .B1(n17168), .B2(n17123), .A(n12470), .ZN(n12474) );
  INV_X1 U15457 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U15458 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12266), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15459 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12471) );
  OAI211_X1 U15460 ( .C1(n15668), .C2(n16922), .A(n12472), .B(n12471), .ZN(
        n12473) );
  AOI211_X1 U15461 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n12474), .B(n12473), .ZN(n12475) );
  OAI211_X1 U15462 ( .C1(n12307), .C2(n16925), .A(n12476), .B(n12475), .ZN(
        n12477) );
  INV_X1 U15463 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U15464 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15465 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15466 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12479) );
  OAI211_X1 U15467 ( .C1(n17215), .C2(n12481), .A(n12480), .B(n12479), .ZN(
        n12487) );
  AOI22_X1 U15468 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15469 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15470 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12483) );
  NAND2_X1 U15471 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12482) );
  NAND4_X1 U15472 ( .A1(n12485), .A2(n12484), .A3(n12483), .A4(n12482), .ZN(
        n12486) );
  AOI211_X1 U15473 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n12487), .B(n12486), .ZN(n12488) );
  NOR2_X1 U15474 ( .A1(n18262), .A2(n17278), .ZN(n12532) );
  NAND2_X1 U15475 ( .A1(n12490), .A2(n12532), .ZN(n15690) );
  INV_X1 U15476 ( .A(n17278), .ZN(n18257) );
  INV_X1 U15477 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U15478 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12500) );
  INV_X1 U15479 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U15480 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15481 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12491) );
  OAI211_X1 U15482 ( .C1(n17215), .C2(n17131), .A(n12492), .B(n12491), .ZN(
        n12498) );
  AOI22_X1 U15483 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15484 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U15485 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12494) );
  NAND2_X1 U15486 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12493) );
  NAND4_X1 U15487 ( .A1(n12496), .A2(n12495), .A3(n12494), .A4(n12493), .ZN(
        n12497) );
  AOI211_X1 U15488 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n12498), .B(n12497), .ZN(n12499) );
  NAND4_X1 U15489 ( .A1(n12517), .A2(n18257), .A3(n12505), .A4(n17428), .ZN(
        n12501) );
  NAND2_X1 U15490 ( .A1(n12515), .A2(n12528), .ZN(n15717) );
  NAND2_X1 U15491 ( .A1(n12501), .A2(n15717), .ZN(n16522) );
  NAND2_X1 U15492 ( .A1(n17278), .A2(n18244), .ZN(n12519) );
  INV_X1 U15493 ( .A(n12519), .ZN(n15731) );
  NAND2_X1 U15494 ( .A1(n17278), .A2(n18262), .ZN(n15867) );
  NOR2_X1 U15495 ( .A1(n18237), .A2(n16544), .ZN(n12504) );
  OAI21_X1 U15496 ( .B1(n18268), .B2(n18688), .A(n12504), .ZN(n15720) );
  OAI21_X1 U15497 ( .B1(n15731), .B2(n12505), .A(n15720), .ZN(n12513) );
  NOR2_X1 U15498 ( .A1(n12528), .A2(n12508), .ZN(n15736) );
  NOR2_X1 U15499 ( .A1(n12505), .A2(n15736), .ZN(n12512) );
  INV_X1 U15500 ( .A(n15735), .ZN(n18253) );
  AOI22_X1 U15501 ( .A1(n18249), .A2(n12506), .B1(n18253), .B2(n18688), .ZN(
        n12511) );
  NAND2_X1 U15502 ( .A1(n17365), .A2(n12508), .ZN(n12509) );
  NAND2_X1 U15503 ( .A1(n18237), .A2(n16544), .ZN(n12507) );
  NAND2_X1 U15504 ( .A1(n18244), .A2(n12507), .ZN(n12530) );
  AOI22_X1 U15505 ( .A1(n12509), .A2(n15735), .B1(n12530), .B2(n12508), .ZN(
        n12510) );
  OAI211_X1 U15506 ( .C1(n12512), .C2(n17428), .A(n12511), .B(n12510), .ZN(
        n15718) );
  NAND2_X1 U15507 ( .A1(n12515), .A2(n12518), .ZN(n15715) );
  NAND2_X1 U15508 ( .A1(n18262), .A2(n15735), .ZN(n18668) );
  INV_X1 U15509 ( .A(n12520), .ZN(n12526) );
  XNOR2_X1 U15510 ( .A(n12522), .B(n12521), .ZN(n12524) );
  AOI21_X1 U15511 ( .B1(n12527), .B2(n12526), .A(n16517), .ZN(n18712) );
  NOR2_X1 U15512 ( .A1(n18884), .A2(n12528), .ZN(n15730) );
  NAND2_X1 U15513 ( .A1(n15730), .A2(n12529), .ZN(n15728) );
  INV_X1 U15514 ( .A(n12530), .ZN(n12534) );
  AOI211_X1 U15515 ( .C1(n15735), .C2(n15867), .A(n12532), .B(n12531), .ZN(
        n12533) );
  NAND2_X1 U15516 ( .A1(n12534), .A2(n12533), .ZN(n15719) );
  NOR3_X1 U15517 ( .A1(n18735), .A2(n18727), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18723) );
  INV_X1 U15518 ( .A(n18723), .ZN(n18732) );
  NOR2_X1 U15519 ( .A1(n12535), .A2(n17899), .ZN(n12546) );
  NOR2_X1 U15520 ( .A1(n12546), .A2(n12536), .ZN(n12544) );
  NOR2_X1 U15521 ( .A1(n17408), .A2(n12544), .ZN(n12543) );
  NAND2_X1 U15522 ( .A1(n12543), .A2(n12537), .ZN(n12541) );
  NOR2_X1 U15523 ( .A1(n17401), .A2(n12541), .ZN(n12540) );
  NAND2_X1 U15524 ( .A1(n12540), .A2(n12538), .ZN(n12539) );
  NOR2_X1 U15525 ( .A1(n17394), .A2(n12539), .ZN(n12563) );
  XOR2_X1 U15526 ( .A(n17394), .B(n12539), .Z(n17826) );
  XNOR2_X1 U15527 ( .A(n17398), .B(n12540), .ZN(n12556) );
  XOR2_X1 U15528 ( .A(n17401), .B(n12541), .Z(n12542) );
  NAND2_X1 U15529 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12542), .ZN(
        n12555) );
  XOR2_X1 U15530 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12542), .Z(
        n17845) );
  XNOR2_X1 U15531 ( .A(n17405), .B(n12543), .ZN(n12553) );
  XOR2_X1 U15532 ( .A(n12544), .B(n17408), .Z(n12545) );
  NAND2_X1 U15533 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12545), .ZN(
        n12551) );
  XOR2_X1 U15534 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12545), .Z(
        n17868) );
  XNOR2_X1 U15535 ( .A(n17413), .B(n12546), .ZN(n12547) );
  OR2_X1 U15536 ( .A1(n18201), .A2(n12547), .ZN(n12550) );
  XOR2_X1 U15537 ( .A(n18201), .B(n12547), .Z(n17882) );
  INV_X1 U15538 ( .A(n17899), .ZN(n15868) );
  AOI21_X1 U15539 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17418), .A(
        n15868), .ZN(n12549) );
  NOR2_X1 U15540 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17418), .ZN(
        n12548) );
  AOI221_X1 U15541 ( .B1(n15868), .B2(n17418), .C1(n12549), .C2(n18863), .A(
        n12548), .ZN(n17881) );
  NAND2_X1 U15542 ( .A1(n17882), .A2(n17881), .ZN(n17880) );
  NAND2_X1 U15543 ( .A1(n12550), .A2(n17880), .ZN(n17867) );
  NAND2_X1 U15544 ( .A1(n17868), .A2(n17867), .ZN(n17866) );
  NAND2_X1 U15545 ( .A1(n12551), .A2(n17866), .ZN(n12552) );
  NAND2_X1 U15546 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  NAND2_X1 U15547 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17859), .ZN(
        n17858) );
  NAND2_X1 U15548 ( .A1(n12554), .A2(n17858), .ZN(n17844) );
  NAND2_X1 U15549 ( .A1(n17845), .A2(n17844), .ZN(n17843) );
  NAND2_X1 U15550 ( .A1(n12555), .A2(n17843), .ZN(n12557) );
  NAND2_X1 U15551 ( .A1(n12556), .A2(n12557), .ZN(n12558) );
  XOR2_X1 U15552 ( .A(n12557), .B(n12556), .Z(n17832) );
  NAND2_X1 U15553 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17832), .ZN(
        n17831) );
  NAND2_X1 U15554 ( .A1(n12563), .A2(n12559), .ZN(n12564) );
  INV_X1 U15555 ( .A(n12559), .ZN(n12562) );
  NAND2_X1 U15556 ( .A1(n17826), .A2(n17825), .ZN(n12561) );
  NAND2_X1 U15557 ( .A1(n12563), .A2(n12562), .ZN(n12560) );
  OAI211_X1 U15558 ( .C1(n12563), .C2(n12562), .A(n12561), .B(n12560), .ZN(
        n17804) );
  NAND2_X1 U15559 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17804), .ZN(
        n17803) );
  INV_X1 U15560 ( .A(n18034), .ZN(n12565) );
  NOR2_X1 U15561 ( .A1(n18005), .A2(n17606), .ZN(n15742) );
  INV_X1 U15562 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17949) );
  NOR2_X1 U15563 ( .A1(n17618), .A2(n17949), .ZN(n17929) );
  NAND2_X1 U15564 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17929), .ZN(
        n17570) );
  INV_X1 U15565 ( .A(n17570), .ZN(n17905) );
  NAND2_X1 U15566 ( .A1(n15742), .A2(n17905), .ZN(n17578) );
  NOR2_X1 U15567 ( .A1(n12565), .A2(n17578), .ZN(n17589) );
  NAND2_X1 U15568 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17589), .ZN(
        n17545) );
  NOR2_X1 U15569 ( .A1(n15846), .A2(n17545), .ZN(n16377) );
  NAND2_X1 U15570 ( .A1(n16377), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12566) );
  XNOR2_X1 U15571 ( .A(n18843), .B(n12566), .ZN(n16402) );
  INV_X1 U15572 ( .A(n12568), .ZN(n16523) );
  NAND2_X1 U15573 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17730), .ZN(
        n17729) );
  NAND2_X1 U15574 ( .A1(n18035), .A2(n17951), .ZN(n17941) );
  NOR2_X1 U15575 ( .A1(n17941), .A2(n17949), .ZN(n17580) );
  NAND2_X1 U15576 ( .A1(n17580), .A2(n9777), .ZN(n17912) );
  NOR2_X1 U15577 ( .A1(n17912), .A2(n15846), .ZN(n16386) );
  NAND2_X1 U15578 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16386), .ZN(
        n12567) );
  XOR2_X1 U15579 ( .A(n12567), .B(n18843), .Z(n16399) );
  INV_X1 U15580 ( .A(n17394), .ZN(n16414) );
  AOI21_X1 U15581 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n15708)
         );
  INV_X1 U15582 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18844) );
  INV_X1 U15583 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18883) );
  NOR2_X1 U15584 ( .A1(n18844), .A2(n18883), .ZN(n17805) );
  INV_X1 U15585 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12574) );
  INV_X1 U15586 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17567) );
  NAND3_X1 U15587 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12569) );
  NAND2_X1 U15588 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17742) );
  INV_X1 U15589 ( .A(n17742), .ZN(n17724) );
  NAND2_X1 U15590 ( .A1(n17724), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16556) );
  INV_X1 U15591 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17680) );
  INV_X1 U15592 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17623) );
  INV_X1 U15593 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17584) );
  NAND3_X1 U15594 ( .A1(n17582), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17566) );
  AND2_X2 U15595 ( .A1(n17534), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16562) );
  INV_X1 U15596 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16378) );
  INV_X1 U15597 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18819) );
  NOR2_X1 U15598 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18862) );
  NAND2_X1 U15599 ( .A1(n18727), .A2(n18862), .ZN(n18896) );
  OR2_X2 U15600 ( .A1(n18896), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18108) );
  NOR2_X1 U15601 ( .A1(n18819), .A2(n18108), .ZN(n16396) );
  NAND2_X1 U15602 ( .A1(n17534), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16376) );
  NOR2_X1 U15603 ( .A1(n16378), .A2(n16376), .ZN(n12571) );
  NAND2_X1 U15604 ( .A1(n18735), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18742) );
  NAND3_X1 U15605 ( .A1(n18727), .A2(n18833), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18574) );
  NAND2_X1 U15606 ( .A1(n18719), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18846) );
  NOR2_X1 U15607 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18888) );
  AOI21_X1 U15608 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18888), .ZN(n18739) );
  OR2_X1 U15609 ( .A1(n18860), .A2(n18739), .ZN(n18235) );
  AOI21_X1 U15610 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17624), .A(
        n18548), .ZN(n17754) );
  NAND2_X1 U15611 ( .A1(n12571), .A2(n17710), .ZN(n16364) );
  XNOR2_X1 U15612 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12575) );
  NOR2_X1 U15613 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17682), .ZN(
        n16379) );
  INV_X1 U15614 ( .A(n12571), .ZN(n12572) );
  INV_X1 U15615 ( .A(n18742), .ZN(n17697) );
  AOI22_X1 U15616 ( .A1(n18548), .A2(n12572), .B1(n17697), .B2(n16561), .ZN(
        n12573) );
  NAND2_X1 U15617 ( .A1(n12573), .A2(n17900), .ZN(n16385) );
  NOR2_X1 U15618 ( .A1(n16379), .A2(n16385), .ZN(n16363) );
  OAI22_X1 U15619 ( .A1(n16364), .A2(n12575), .B1(n16363), .B2(n12574), .ZN(
        n12576) );
  AOI211_X1 U15620 ( .C1(n17756), .C2(n10056), .A(n16396), .B(n12576), .ZN(
        n12577) );
  INV_X1 U15621 ( .A(n12577), .ZN(n12578) );
  NOR2_X1 U15622 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12583) );
  NOR4_X1 U15623 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12582) );
  NAND4_X1 U15624 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12583), .A4(n12582), .ZN(n12586) );
  NOR2_X1 U15625 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12586), .ZN(n16503)
         );
  INV_X1 U15626 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20923) );
  NOR3_X1 U15627 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        n20923), .ZN(n12585) );
  NOR4_X1 U15628 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12584)
         );
  NAND4_X1 U15629 ( .A1(n14535), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12585), .A4(
        n12584), .ZN(U214) );
  NOR2_X1 U15630 ( .A1(n19267), .A2(n12586), .ZN(n16423) );
  NAND2_X1 U15631 ( .A1(n16423), .A2(U214), .ZN(U212) );
  INV_X1 U15632 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12592) );
  NAND2_X1 U15633 ( .A1(n12617), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12615) );
  INV_X1 U15634 ( .A(n12615), .ZN(n12588) );
  NAND2_X1 U15635 ( .A1(n12588), .A2(n10252), .ZN(n12612) );
  NAND2_X1 U15636 ( .A1(n12608), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12609) );
  INV_X1 U15637 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16176) );
  NAND2_X1 U15638 ( .A1(n12607), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12606) );
  INV_X1 U15639 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18968) );
  OR2_X1 U15640 ( .A1(n11971), .A2(n18968), .ZN(n12589) );
  NAND2_X1 U15641 ( .A1(n12604), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12602) );
  INV_X1 U15642 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16140) );
  NAND2_X1 U15643 ( .A1(n12600), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12599) );
  INV_X1 U15644 ( .A(n14955), .ZN(n12591) );
  AOI21_X1 U15645 ( .B1(n12592), .B2(n12590), .A(n12591), .ZN(n15211) );
  INV_X1 U15646 ( .A(n14952), .ZN(n12593) );
  NAND2_X1 U15647 ( .A1(n12593), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12595) );
  INV_X1 U15648 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12594) );
  INV_X1 U15649 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12596) );
  INV_X1 U15650 ( .A(n13601), .ZN(n12631) );
  OR2_X1 U15651 ( .A1(n12597), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12598) );
  NAND2_X1 U15652 ( .A1(n12590), .A2(n12598), .ZN(n15220) );
  INV_X1 U15653 ( .A(n15220), .ZN(n16073) );
  AOI21_X1 U15654 ( .B1(n16083), .B2(n12601), .A(n12597), .ZN(n16092) );
  OAI21_X1 U15655 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12600), .A(
        n12601), .ZN(n16139) );
  INV_X1 U15656 ( .A(n16139), .ZN(n14998) );
  AOI21_X1 U15657 ( .B1(n16140), .B2(n12603), .A(n12600), .ZN(n16142) );
  OAI21_X1 U15658 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12604), .A(
        n12603), .ZN(n16154) );
  INV_X1 U15659 ( .A(n16154), .ZN(n15778) );
  AOI21_X1 U15660 ( .B1(n15246), .B2(n9680), .A(n12604), .ZN(n15244) );
  OAI21_X1 U15661 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12605), .A(
        n9680), .ZN(n15260) );
  INV_X1 U15662 ( .A(n15260), .ZN(n18935) );
  AOI21_X1 U15663 ( .B1(n9673), .B2(n15269), .A(n12605), .ZN(n18946) );
  NOR2_X1 U15664 ( .A1(n18968), .A2(n12606), .ZN(n12629) );
  OAI21_X1 U15665 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12629), .A(
        n9673), .ZN(n16160) );
  INV_X1 U15666 ( .A(n16160), .ZN(n18958) );
  OAI21_X1 U15667 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12607), .A(
        n12606), .ZN(n18982) );
  INV_X1 U15668 ( .A(n18982), .ZN(n12628) );
  OAI21_X1 U15669 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12608), .A(
        n12609), .ZN(n16186) );
  INV_X1 U15670 ( .A(n16186), .ZN(n12627) );
  OAI21_X1 U15671 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12610), .A(
        n12626), .ZN(n16192) );
  INV_X1 U15672 ( .A(n16192), .ZN(n12625) );
  INV_X1 U15673 ( .A(n12613), .ZN(n12614) );
  AOI21_X1 U15674 ( .B1(n16213), .B2(n12622), .A(n12614), .ZN(n19033) );
  NOR2_X1 U15675 ( .A1(n16235), .A2(n12615), .ZN(n12623) );
  AOI21_X1 U15676 ( .B1(n16235), .B2(n12615), .A(n12623), .ZN(n16220) );
  AOI21_X1 U15677 ( .B1(n19068), .B2(n12616), .A(n12617), .ZN(n19074) );
  AOI21_X1 U15678 ( .B1(n19230), .B2(n12618), .A(n12619), .ZN(n19215) );
  AOI21_X1 U15679 ( .B1(n13827), .B2(n12621), .A(n12620), .ZN(n13616) );
  AOI22_X1 U15680 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19986), .ZN(n13807) );
  AOI22_X1 U15681 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13827), .B2(n19986), .ZN(
        n13804) );
  NAND2_X1 U15682 ( .A1(n13807), .A2(n13804), .ZN(n13803) );
  NOR2_X1 U15683 ( .A1(n13616), .A2(n13803), .ZN(n13724) );
  OAI21_X1 U15684 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12620), .A(
        n12618), .ZN(n13725) );
  NAND2_X1 U15685 ( .A1(n13724), .A2(n13725), .ZN(n19110) );
  NOR2_X1 U15686 ( .A1(n19215), .A2(n19110), .ZN(n19084) );
  OAI21_X1 U15687 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12619), .A(
        n12616), .ZN(n19086) );
  NAND2_X1 U15688 ( .A1(n19084), .A2(n19086), .ZN(n19072) );
  NOR2_X1 U15689 ( .A1(n19074), .A2(n19072), .ZN(n19053) );
  OAI21_X1 U15690 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12617), .A(
        n12615), .ZN(n19055) );
  NAND2_X1 U15691 ( .A1(n19053), .A2(n19055), .ZN(n13602) );
  NOR2_X1 U15692 ( .A1(n16220), .A2(n13602), .ZN(n19045) );
  OAI21_X1 U15693 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n12623), .A(
        n12622), .ZN(n19047) );
  NAND2_X1 U15694 ( .A1(n19045), .A2(n19047), .ZN(n19032) );
  NOR2_X1 U15695 ( .A1(n19033), .A2(n19032), .ZN(n19020) );
  AOI21_X1 U15696 ( .B1(n19017), .B2(n12613), .A(n12610), .ZN(n19023) );
  INV_X1 U15697 ( .A(n19023), .ZN(n12624) );
  NAND2_X1 U15698 ( .A1(n19020), .A2(n12624), .ZN(n15025) );
  NOR2_X1 U15699 ( .A1(n12625), .A2(n15025), .ZN(n19013) );
  AOI21_X1 U15700 ( .B1(n15296), .B2(n12626), .A(n12608), .ZN(n19008) );
  INV_X1 U15701 ( .A(n19008), .ZN(n19012) );
  NAND2_X1 U15702 ( .A1(n19013), .A2(n19012), .ZN(n13930) );
  NOR2_X1 U15703 ( .A1(n12627), .A2(n13930), .ZN(n18997) );
  AOI21_X1 U15704 ( .B1(n16176), .B2(n12609), .A(n12607), .ZN(n16169) );
  INV_X1 U15705 ( .A(n16169), .ZN(n18996) );
  NAND2_X1 U15706 ( .A1(n18997), .A2(n18996), .ZN(n18994) );
  NOR2_X1 U15707 ( .A1(n12628), .A2(n18994), .ZN(n18965) );
  AOI21_X1 U15708 ( .B1(n18968), .B2(n12606), .A(n12629), .ZN(n12630) );
  INV_X1 U15709 ( .A(n12630), .ZN(n18966) );
  NOR2_X1 U15710 ( .A1(n18935), .A2(n18934), .ZN(n18933) );
  NOR2_X1 U15711 ( .A1(n19021), .A2(n15777), .ZN(n15020) );
  NOR2_X1 U15712 ( .A1(n16142), .A2(n15020), .ZN(n15019) );
  NOR2_X1 U15713 ( .A1(n14998), .A2(n14996), .ZN(n14997) );
  NOR2_X1 U15714 ( .A1(n19021), .A2(n14997), .ZN(n16091) );
  NOR2_X1 U15715 ( .A1(n16092), .A2(n16091), .ZN(n16090) );
  NOR2_X1 U15716 ( .A1(n16073), .A2(n16072), .ZN(n16071) );
  NOR2_X1 U15717 ( .A1(n19021), .A2(n16071), .ZN(n12632) );
  NOR2_X1 U15718 ( .A1(n15211), .A2(n12632), .ZN(n14956) );
  INV_X1 U15719 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19980) );
  INV_X1 U15720 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19989) );
  NAND4_X1 U15721 ( .A1(n19980), .A2(n19986), .A3(n19989), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19851) );
  AOI211_X1 U15722 ( .C1(n15211), .C2(n12632), .A(n14956), .B(n19851), .ZN(
        n12677) );
  MUX2_X1 U15723 ( .A(n12633), .B(P2_EBX_REG_3__SCAN_IN), .S(n14206), .Z(
        n13429) );
  NAND2_X1 U15724 ( .A1(n12757), .A2(n12846), .ZN(n12635) );
  NAND2_X1 U15725 ( .A1(n12635), .A2(n12634), .ZN(n12701) );
  INV_X1 U15726 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12636) );
  MUX2_X1 U15727 ( .A(n12701), .B(n12636), .S(n14206), .Z(n12862) );
  NOR2_X1 U15728 ( .A1(n15154), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12759) );
  INV_X1 U15729 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13832) );
  NAND2_X1 U15730 ( .A1(n12759), .A2(n13832), .ZN(n12638) );
  NAND2_X1 U15731 ( .A1(n12844), .A2(n15154), .ZN(n12637) );
  NAND2_X1 U15732 ( .A1(n12638), .A2(n12637), .ZN(n12861) );
  NAND2_X1 U15733 ( .A1(n12862), .A2(n12861), .ZN(n13428) );
  INV_X1 U15734 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12640) );
  MUX2_X1 U15735 ( .A(n12640), .B(n12639), .S(n15154), .Z(n13638) );
  INV_X1 U15736 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12642) );
  MUX2_X1 U15737 ( .A(n12642), .B(n12641), .S(n15154), .Z(n13675) );
  MUX2_X1 U15738 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n13888), .S(n15154), .Z(
        n13902) );
  INV_X1 U15739 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12643) );
  MUX2_X1 U15740 ( .A(n12643), .B(n13426), .S(n15154), .Z(n14105) );
  INV_X1 U15741 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19031) );
  NAND2_X1 U15742 ( .A1(n14206), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13598) );
  INV_X1 U15743 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12644) );
  INV_X1 U15744 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19138) );
  NAND2_X1 U15745 ( .A1(n19031), .A2(n14123), .ZN(n14133) );
  NAND2_X1 U15746 ( .A1(n14206), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12645) );
  INV_X1 U15747 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12646) );
  NOR2_X1 U15748 ( .A1(n15154), .A2(n12646), .ZN(n14139) );
  NOR2_X1 U15749 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n12647) );
  INV_X1 U15750 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U15751 ( .A1(n14206), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14157) );
  INV_X1 U15752 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12649) );
  NOR2_X1 U15753 ( .A1(n15154), .A2(n12649), .ZN(n14152) );
  NAND2_X1 U15754 ( .A1(n14206), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14151) );
  NAND2_X1 U15755 ( .A1(n14206), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14196) );
  NAND2_X1 U15756 ( .A1(n14206), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14201) );
  INV_X1 U15757 ( .A(n14201), .ZN(n12651) );
  INV_X1 U15758 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15070) );
  NAND2_X1 U15759 ( .A1(n14220), .A2(n9699), .ZN(n14951) );
  NAND2_X1 U15760 ( .A1(n14206), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12652) );
  NAND2_X1 U15761 ( .A1(n14951), .A2(n12652), .ZN(n14227) );
  INV_X1 U15762 ( .A(n12652), .ZN(n12653) );
  NAND2_X1 U15763 ( .A1(n12653), .A2(n9699), .ZN(n12654) );
  NAND2_X1 U15764 ( .A1(n14227), .A2(n12654), .ZN(n14217) );
  OR2_X1 U15765 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19985), .ZN(n12667) );
  NAND2_X1 U15766 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12667), .ZN(n12655) );
  INV_X1 U15767 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19913) );
  AND2_X1 U15768 ( .A1(n19981), .A2(n19938), .ZN(n12657) );
  INV_X2 U15769 ( .A(n12657), .ZN(n19066) );
  NOR3_X1 U15770 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19854), .A3(n19979), 
        .ZN(n16344) );
  NOR2_X1 U15771 ( .A1(n15785), .A2(n16344), .ZN(n12658) );
  NAND2_X1 U15772 ( .A1(n19851), .A2(n12658), .ZN(n12659) );
  OAI22_X1 U15773 ( .A1(n14217), .A2(n19099), .B1(n19913), .B2(n19067), .ZN(
        n12676) );
  INV_X1 U15774 ( .A(n12693), .ZN(n12660) );
  INV_X1 U15775 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19858) );
  NAND2_X2 U15776 ( .A1(n19880), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19917) );
  INV_X1 U15777 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19869) );
  NAND2_X1 U15778 ( .A1(n18904), .A2(n19869), .ZN(n19863) );
  NAND3_X1 U15779 ( .A1(n19858), .A2(n19917), .A3(n19863), .ZN(n19987) );
  NOR2_X1 U15780 ( .A1(n19987), .A2(n19985), .ZN(n12907) );
  NAND2_X1 U15781 ( .A1(n19989), .A2(n12907), .ZN(n12669) );
  NAND2_X1 U15782 ( .A1(n12824), .A2(n12669), .ZN(n14973) );
  INV_X1 U15783 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12661) );
  NAND2_X1 U15784 ( .A1(n12661), .A2(n12667), .ZN(n12662) );
  OR2_X1 U15785 ( .A1(n12715), .A2(n12662), .ZN(n12663) );
  NAND2_X1 U15786 ( .A1(n19067), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19093) );
  AOI22_X1 U15787 ( .A1(n19096), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19095), .ZN(n12664) );
  INV_X1 U15788 ( .A(n12664), .ZN(n12675) );
  OR2_X1 U15789 ( .A1(n15058), .A2(n12665), .ZN(n12666) );
  NAND2_X1 U15790 ( .A1(n14983), .A2(n12666), .ZN(n15345) );
  NOR2_X1 U15791 ( .A1(n12947), .A2(n12669), .ZN(n16347) );
  AND2_X1 U15792 ( .A1(n18906), .A2(n16347), .ZN(n18973) );
  INV_X2 U15793 ( .A(n18973), .ZN(n19098) );
  NAND2_X1 U15794 ( .A1(n12670), .A2(n12671), .ZN(n12672) );
  INV_X1 U15795 ( .A(n15343), .ZN(n12673) );
  OAI22_X1 U15796 ( .A1(n15345), .A2(n19107), .B1(n19098), .B2(n12673), .ZN(
        n12674) );
  OR4_X1 U15797 ( .A1(n12677), .A2(n12676), .A3(n12675), .A4(n12674), .ZN(
        P2_U2828) );
  AOI211_X1 U15798 ( .C1(n15244), .C2(n12679), .A(n12678), .B(n19851), .ZN(
        n12692) );
  OAI22_X1 U15799 ( .A1(n15246), .A2(n19093), .B1(n11985), .B2(n19067), .ZN(
        n12691) );
  NAND3_X1 U15800 ( .A1(n14148), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n14206), 
        .ZN(n12680) );
  NAND2_X1 U15801 ( .A1(n12681), .A2(n12680), .ZN(n14180) );
  INV_X1 U15802 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12682) );
  OAI22_X1 U15803 ( .A1(n14180), .A2(n19099), .B1(n19082), .B2(n12682), .ZN(
        n12690) );
  INV_X1 U15804 ( .A(n15412), .ZN(n12684) );
  AOI21_X1 U15805 ( .B1(n12685), .B2(n12683), .A(n12684), .ZN(n15251) );
  INV_X1 U15806 ( .A(n15251), .ZN(n15432) );
  OR2_X1 U15807 ( .A1(n15444), .A2(n12686), .ZN(n12688) );
  INV_X1 U15808 ( .A(n15415), .ZN(n12687) );
  AND2_X1 U15809 ( .A1(n12688), .A2(n12687), .ZN(n15429) );
  INV_X1 U15810 ( .A(n15429), .ZN(n15139) );
  OAI22_X1 U15811 ( .A1(n15432), .A2(n19107), .B1(n19098), .B2(n15139), .ZN(
        n12689) );
  OR4_X1 U15812 ( .A1(n12692), .A2(n12691), .A3(n12690), .A4(n12689), .ZN(
        P2_U2834) );
  INV_X1 U15813 ( .A(n12047), .ZN(n12694) );
  NAND2_X1 U15814 ( .A1(n12694), .A2(n12693), .ZN(n19108) );
  INV_X1 U15815 ( .A(n19108), .ZN(n12696) );
  INV_X1 U15816 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12695) );
  NAND2_X1 U15817 ( .A1(n19938), .A2(n15593), .ZN(n12697) );
  OAI211_X1 U15818 ( .C1(n12696), .C2(n12695), .A(n12715), .B(n12697), .ZN(
        P2_U2814) );
  NOR2_X1 U15819 ( .A1(n18906), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12698)
         );
  AOI22_X1 U15820 ( .A1(n12698), .A2(n12697), .B1(n12925), .B2(n18906), .ZN(
        P2_U3612) );
  INV_X1 U15821 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12746) );
  OR2_X1 U15822 ( .A1(n16322), .A2(n12907), .ZN(n12699) );
  NOR2_X1 U15823 ( .A1(n12739), .A2(n12699), .ZN(n12700) );
  NAND2_X1 U15824 ( .A1(n16323), .A2(n12700), .ZN(n16334) );
  AND2_X1 U15825 ( .A1(n16334), .A2(n16345), .ZN(n19969) );
  AOI21_X1 U15826 ( .B1(n12758), .B2(n12702), .A(n12701), .ZN(n12703) );
  OR2_X1 U15827 ( .A1(n12704), .A2(n12703), .ZN(n12706) );
  NAND2_X1 U15828 ( .A1(n12706), .A2(n12705), .ZN(n19974) );
  NAND2_X1 U15829 ( .A1(n13136), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12707) );
  NAND2_X1 U15830 ( .A1(n12707), .A2(n12751), .ZN(n16330) );
  OAI21_X1 U15831 ( .B1(n12188), .B2(n16330), .A(n12746), .ZN(n12708) );
  AND2_X1 U15832 ( .A1(n12708), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19963) );
  AOI211_X1 U15833 ( .C1(n12710), .C2(n12709), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n16322), .ZN(n12711) );
  NOR2_X1 U15834 ( .A1(n19963), .A2(n12711), .ZN(n19970) );
  OAI22_X1 U15835 ( .A1(n19974), .A2(n12947), .B1(n19282), .B2(n19970), .ZN(
        n12714) );
  NOR2_X1 U15836 ( .A1(n16328), .A2(n12770), .ZN(n12713) );
  NAND2_X1 U15837 ( .A1(n12919), .A2(n19988), .ZN(n12756) );
  OAI21_X1 U15838 ( .B1(n12746), .B2(n19969), .A(n12756), .ZN(P2_U2819) );
  INV_X1 U15839 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19191) );
  NOR2_X1 U15840 ( .A1(n12715), .A2(n19985), .ZN(n12716) );
  NAND2_X1 U15841 ( .A1(n12731), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12721) );
  INV_X1 U15842 ( .A(n12716), .ZN(n12717) );
  INV_X1 U15843 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16453) );
  OR2_X1 U15844 ( .A1(n19267), .A2(n16453), .ZN(n12720) );
  NAND2_X1 U15845 ( .A1(n19267), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12719) );
  NAND2_X1 U15846 ( .A1(n12720), .A2(n12719), .ZN(n19160) );
  NAND2_X1 U15847 ( .A1(n12718), .A2(n19160), .ZN(n12879) );
  OAI211_X1 U15848 ( .C1(n19191), .C2(n12881), .A(n12721), .B(n12879), .ZN(
        P2_U2977) );
  INV_X1 U15849 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13000) );
  NAND2_X1 U15850 ( .A1(n12731), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12722) );
  INV_X1 U15851 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16457) );
  INV_X1 U15852 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17393) );
  MUX2_X1 U15853 ( .A(n16457), .B(n17393), .S(n19267), .Z(n15119) );
  INV_X1 U15854 ( .A(n15119), .ZN(n19166) );
  NAND2_X1 U15855 ( .A1(n12718), .A2(n19166), .ZN(n12723) );
  OAI211_X1 U15856 ( .C1(n13000), .C2(n12881), .A(n12722), .B(n12723), .ZN(
        P2_U2960) );
  INV_X1 U15857 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19195) );
  NAND2_X1 U15858 ( .A1(n12731), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12724) );
  OAI211_X1 U15859 ( .C1(n19195), .C2(n12881), .A(n12724), .B(n12723), .ZN(
        P2_U2975) );
  INV_X1 U15860 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19187) );
  NAND2_X1 U15861 ( .A1(n12731), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12725) );
  INV_X1 U15862 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16450) );
  INV_X1 U15863 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17375) );
  MUX2_X1 U15864 ( .A(n16450), .B(n17375), .S(n19267), .Z(n15091) );
  INV_X1 U15865 ( .A(n15091), .ZN(n19157) );
  NAND2_X1 U15866 ( .A1(n12718), .A2(n19157), .ZN(n12726) );
  OAI211_X1 U15867 ( .C1(n19187), .C2(n12881), .A(n12725), .B(n12726), .ZN(
        P2_U2979) );
  INV_X1 U15868 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12781) );
  NAND2_X1 U15869 ( .A1(n12731), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12727) );
  OAI211_X1 U15870 ( .C1(n12781), .C2(n12881), .A(n12727), .B(n12726), .ZN(
        P2_U2964) );
  INV_X1 U15871 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19193) );
  NAND2_X1 U15872 ( .A1(n12731), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12730) );
  INV_X1 U15873 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16455) );
  OR2_X1 U15874 ( .A1(n19267), .A2(n16455), .ZN(n12729) );
  NAND2_X1 U15875 ( .A1(n19267), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12728) );
  AND2_X1 U15876 ( .A1(n12729), .A2(n12728), .ZN(n15115) );
  INV_X1 U15877 ( .A(n15115), .ZN(n19163) );
  NAND2_X1 U15878 ( .A1(n12718), .A2(n19163), .ZN(n12816) );
  OAI211_X1 U15879 ( .C1(n19193), .C2(n12881), .A(n12730), .B(n12816), .ZN(
        P2_U2976) );
  INV_X1 U15880 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12734) );
  INV_X1 U15881 ( .A(n12731), .ZN(n12784) );
  INV_X1 U15882 ( .A(n12718), .ZN(n12733) );
  AOI22_X1 U15883 ( .A1(n19269), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19267), .ZN(n13821) );
  INV_X1 U15884 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12732) );
  OAI222_X1 U15885 ( .A1(n12734), .A2(n12784), .B1(n12733), .B2(n13821), .C1(
        n12881), .C2(n12732), .ZN(P2_U2982) );
  NOR2_X1 U15886 ( .A1(n12047), .A2(n19282), .ZN(n12735) );
  NAND2_X1 U15887 ( .A1(n16327), .A2(n12735), .ZN(n12771) );
  INV_X1 U15888 ( .A(n12907), .ZN(n12745) );
  NOR2_X1 U15889 ( .A1(n16322), .A2(n12745), .ZN(n12736) );
  AND2_X1 U15890 ( .A1(n16348), .A2(n12736), .ZN(n12737) );
  NOR2_X1 U15891 ( .A1(n12738), .A2(n12737), .ZN(n12916) );
  INV_X1 U15892 ( .A(n16322), .ZN(n12912) );
  NAND3_X1 U15893 ( .A1(n16323), .A2(n12912), .A3(n12739), .ZN(n12740) );
  AND2_X1 U15894 ( .A1(n12916), .A2(n12740), .ZN(n12741) );
  AND2_X1 U15895 ( .A1(n12742), .A2(n12741), .ZN(n12744) );
  OAI211_X1 U15896 ( .C1(n12771), .C2(n12745), .A(n12744), .B(n12743), .ZN(
        n16337) );
  NAND2_X1 U15897 ( .A1(n16337), .A2(n16345), .ZN(n12749) );
  NAND2_X1 U15898 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n15857) );
  NOR2_X1 U15899 ( .A1(n19986), .A2(n15857), .ZN(n16358) );
  INV_X1 U15900 ( .A(n16358), .ZN(n16357) );
  OAI22_X1 U15901 ( .A1(n16357), .A2(n12746), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n19979), .ZN(n12747) );
  INV_X1 U15902 ( .A(n12747), .ZN(n12748) );
  NAND2_X1 U15903 ( .A1(n12749), .A2(n12748), .ZN(n15611) );
  NOR2_X1 U15904 ( .A1(n12047), .A2(n13398), .ZN(n16331) );
  NAND2_X1 U15905 ( .A1(n15593), .A2(n19979), .ZN(n15608) );
  INV_X1 U15906 ( .A(n15608), .ZN(n19933) );
  NAND4_X1 U15907 ( .A1(n15611), .A2(n16331), .A3(n16330), .A4(n19933), .ZN(
        n12750) );
  OAI21_X1 U15908 ( .B1(n12751), .B2(n15611), .A(n12750), .ZN(P2_U3595) );
  NAND2_X1 U15909 ( .A1(n12753), .A2(n12837), .ZN(n12827) );
  NOR2_X1 U15910 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20664), .ZN(n12883) );
  AOI21_X1 U15911 ( .B1(n12882), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n12883), 
        .ZN(n12754) );
  NAND2_X1 U15912 ( .A1(n13036), .A2(n12754), .ZN(P1_U2801) );
  OR2_X1 U15913 ( .A1(n19938), .A2(n19933), .ZN(n19951) );
  NAND2_X1 U15914 ( .A1(n19951), .A2(n19986), .ZN(n12755) );
  AND2_X1 U15915 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19952) );
  AND2_X1 U15916 ( .A1(n12919), .A2(n12757), .ZN(n16240) );
  INV_X1 U15917 ( .A(n12758), .ZN(n12760) );
  AOI21_X1 U15918 ( .B1(n12760), .B2(n15154), .A(n12759), .ZN(n13943) );
  INV_X1 U15919 ( .A(n13943), .ZN(n12762) );
  NAND2_X1 U15920 ( .A1(n13943), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12869) );
  INV_X1 U15921 ( .A(n12869), .ZN(n12761) );
  AOI21_X1 U15922 ( .B1(n12098), .B2(n12762), .A(n12761), .ZN(n12955) );
  AND2_X1 U15923 ( .A1(n12657), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12953) );
  AND2_X1 U15924 ( .A1(n19282), .A2(n12848), .ZN(n12845) );
  INV_X1 U15925 ( .A(n12845), .ZN(n12764) );
  NAND2_X1 U15926 ( .A1(n12764), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12850) );
  OAI21_X1 U15927 ( .B1(n12764), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12850), .ZN(n12951) );
  NOR2_X1 U15928 ( .A1(n16251), .A2(n12951), .ZN(n12765) );
  AOI211_X1 U15929 ( .C1(n16240), .C2(n12955), .A(n12953), .B(n12765), .ZN(
        n12769) );
  INV_X1 U15930 ( .A(n19231), .ZN(n16187) );
  NAND2_X1 U15931 ( .A1(n19989), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12766) );
  NAND2_X1 U15932 ( .A1(n12767), .A2(n12766), .ZN(n12854) );
  OAI21_X1 U15933 ( .B1(n16187), .B2(n12854), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12768) );
  OAI211_X1 U15934 ( .C1(n19223), .C2(n13374), .A(n12769), .B(n12768), .ZN(
        P2_U3014) );
  OAI21_X1 U15935 ( .B1(n12771), .B2(n12770), .A(n12881), .ZN(n12773) );
  INV_X1 U15936 ( .A(n19987), .ZN(n12772) );
  AND2_X1 U15937 ( .A1(n12773), .A2(n12772), .ZN(n19180) );
  NAND2_X1 U15938 ( .A1(n19180), .A2(n12774), .ZN(n13014) );
  INV_X1 U15939 ( .A(n15857), .ZN(n12775) );
  NAND2_X1 U15940 ( .A1(n19986), .A2(n12775), .ZN(n19984) );
  INV_X2 U15941 ( .A(n19984), .ZN(n19212) );
  AOI22_X1 U15942 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19198), .B1(n19212), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12776) );
  OAI21_X1 U15943 ( .B1(n12777), .B2(n13014), .A(n12776), .ZN(P2_U2921) );
  INV_X1 U15944 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U15945 ( .A1(n19212), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19198), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12778) );
  OAI21_X1 U15946 ( .B1(n12779), .B2(n13014), .A(n12778), .ZN(P2_U2926) );
  AOI22_X1 U15947 ( .A1(n19212), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19198), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12780) );
  OAI21_X1 U15948 ( .B1(n12781), .B2(n13014), .A(n12780), .ZN(P2_U2923) );
  INV_X1 U15949 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U15950 ( .A1(n19212), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19198), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12782) );
  OAI21_X1 U15951 ( .B1(n12783), .B2(n13014), .A(n12782), .ZN(P2_U2924) );
  AOI22_X1 U15952 ( .A1(n12878), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12787) );
  INV_X1 U15953 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16448) );
  OR2_X1 U15954 ( .A1(n19267), .A2(n16448), .ZN(n12786) );
  NAND2_X1 U15955 ( .A1(n19267), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12785) );
  NAND2_X1 U15956 ( .A1(n12786), .A2(n12785), .ZN(n14271) );
  NAND2_X1 U15957 ( .A1(n12718), .A2(n14271), .ZN(n12809) );
  NAND2_X1 U15958 ( .A1(n12787), .A2(n12809), .ZN(P2_U2980) );
  AOI22_X1 U15959 ( .A1(n12878), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12788) );
  INV_X1 U15960 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16465) );
  INV_X1 U15961 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18252) );
  AOI22_X1 U15962 ( .A1(n19269), .A2(n16465), .B1(n18252), .B2(n19267), .ZN(
        n16117) );
  NAND2_X1 U15963 ( .A1(n12718), .A2(n16117), .ZN(n12825) );
  NAND2_X1 U15964 ( .A1(n12788), .A2(n12825), .ZN(P2_U2971) );
  AOI22_X1 U15965 ( .A1(n12878), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U15966 ( .A1(n19269), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19267), .ZN(n19290) );
  INV_X1 U15967 ( .A(n19290), .ZN(n15145) );
  NAND2_X1 U15968 ( .A1(n12718), .A2(n15145), .ZN(n12811) );
  NAND2_X1 U15969 ( .A1(n12789), .A2(n12811), .ZN(P2_U2970) );
  AOI22_X1 U15970 ( .A1(n12878), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12790) );
  NAND2_X1 U15971 ( .A1(n12718), .A2(n13744), .ZN(n12793) );
  NAND2_X1 U15972 ( .A1(n12790), .A2(n12793), .ZN(P2_U2981) );
  AOI22_X1 U15973 ( .A1(n12878), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U15974 ( .A1(n19269), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19267), .ZN(n19274) );
  INV_X1 U15975 ( .A(n19274), .ZN(n12791) );
  NAND2_X1 U15976 ( .A1(n12718), .A2(n12791), .ZN(n12818) );
  NAND2_X1 U15977 ( .A1(n12792), .A2(n12818), .ZN(P2_U2967) );
  AOI22_X1 U15978 ( .A1(n12731), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n12824), .ZN(n12794) );
  NAND2_X1 U15979 ( .A1(n12794), .A2(n12793), .ZN(P2_U2966) );
  AOI22_X1 U15980 ( .A1(n12878), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U15981 ( .A1(n19269), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19267), .ZN(n19281) );
  INV_X1 U15982 ( .A(n19281), .ZN(n13955) );
  NAND2_X1 U15983 ( .A1(n12718), .A2(n13955), .ZN(n12800) );
  NAND2_X1 U15984 ( .A1(n12795), .A2(n12800), .ZN(P2_U2968) );
  AOI22_X1 U15985 ( .A1(n12878), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12796) );
  INV_X1 U15986 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16462) );
  INV_X1 U15987 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18261) );
  AOI22_X1 U15988 ( .A1(n19269), .A2(n16462), .B1(n18261), .B2(n19267), .ZN(
        n16111) );
  NAND2_X1 U15989 ( .A1(n12718), .A2(n16111), .ZN(n12804) );
  NAND2_X1 U15990 ( .A1(n12796), .A2(n12804), .ZN(P2_U2973) );
  AOI22_X1 U15991 ( .A1(n12878), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12798) );
  AOI22_X1 U15992 ( .A1(n19269), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19267), .ZN(n19308) );
  INV_X1 U15993 ( .A(n19308), .ZN(n12797) );
  NAND2_X1 U15994 ( .A1(n12718), .A2(n12797), .ZN(n12802) );
  NAND2_X1 U15995 ( .A1(n12798), .A2(n12802), .ZN(P2_U2974) );
  AOI22_X1 U15996 ( .A1(n12878), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U15997 ( .A1(n19269), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19267), .ZN(n19300) );
  INV_X1 U15998 ( .A(n19300), .ZN(n19170) );
  NAND2_X1 U15999 ( .A1(n12718), .A2(n19170), .ZN(n12822) );
  NAND2_X1 U16000 ( .A1(n12799), .A2(n12822), .ZN(P2_U2972) );
  AOI22_X1 U16001 ( .A1(n12878), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U16002 ( .A1(n12801), .A2(n12800), .ZN(P2_U2953) );
  AOI22_X1 U16003 ( .A1(n12878), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12803) );
  NAND2_X1 U16004 ( .A1(n12803), .A2(n12802), .ZN(P2_U2959) );
  AOI22_X1 U16005 ( .A1(n12878), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n12824), .ZN(n12805) );
  NAND2_X1 U16006 ( .A1(n12805), .A2(n12804), .ZN(P2_U2958) );
  AOI22_X1 U16007 ( .A1(n12878), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12808) );
  INV_X1 U16008 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13220) );
  OR2_X1 U16009 ( .A1(n19267), .A2(n13220), .ZN(n12807) );
  NAND2_X1 U16010 ( .A1(n19267), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12806) );
  NAND2_X1 U16011 ( .A1(n12807), .A2(n12806), .ZN(n15097) );
  NAND2_X1 U16012 ( .A1(n12718), .A2(n15097), .ZN(n12814) );
  NAND2_X1 U16013 ( .A1(n12808), .A2(n12814), .ZN(P2_U2978) );
  AOI22_X1 U16014 ( .A1(n12878), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n12824), .ZN(n12810) );
  NAND2_X1 U16015 ( .A1(n12810), .A2(n12809), .ZN(P2_U2965) );
  AOI22_X1 U16016 ( .A1(n12878), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12812) );
  NAND2_X1 U16017 ( .A1(n12812), .A2(n12811), .ZN(P2_U2955) );
  AOI22_X1 U16018 ( .A1(n12878), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12813) );
  OAI22_X1 U16019 ( .A1(n19267), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19269), .ZN(n19286) );
  INV_X1 U16020 ( .A(n19286), .ZN(n16126) );
  NAND2_X1 U16021 ( .A1(n12718), .A2(n16126), .ZN(n12820) );
  NAND2_X1 U16022 ( .A1(n12813), .A2(n12820), .ZN(P2_U2954) );
  AOI22_X1 U16023 ( .A1(n12878), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n12824), .ZN(n12815) );
  NAND2_X1 U16024 ( .A1(n12815), .A2(n12814), .ZN(P2_U2963) );
  AOI22_X1 U16025 ( .A1(n12878), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n12824), .ZN(n12817) );
  NAND2_X1 U16026 ( .A1(n12817), .A2(n12816), .ZN(P2_U2961) );
  AOI22_X1 U16027 ( .A1(n12878), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n12819) );
  NAND2_X1 U16028 ( .A1(n12819), .A2(n12818), .ZN(P2_U2952) );
  AOI22_X1 U16029 ( .A1(n12878), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12821) );
  NAND2_X1 U16030 ( .A1(n12821), .A2(n12820), .ZN(P2_U2969) );
  AOI22_X1 U16031 ( .A1(n12878), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12823) );
  NAND2_X1 U16032 ( .A1(n12823), .A2(n12822), .ZN(P2_U2957) );
  AOI22_X1 U16033 ( .A1(n12878), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n12824), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U16034 ( .A1(n12826), .A2(n12825), .ZN(P2_U2956) );
  AND2_X1 U16035 ( .A1(n12752), .A2(n12827), .ZN(n12828) );
  AOI21_X1 U16036 ( .B1(n13126), .B2(n13565), .A(n12828), .ZN(n20000) );
  OR2_X1 U16037 ( .A1(n20184), .A2(n20192), .ZN(n13171) );
  INV_X1 U16038 ( .A(n12829), .ZN(n12830) );
  NAND2_X1 U16039 ( .A1(n12830), .A2(n20739), .ZN(n15853) );
  NAND3_X1 U16040 ( .A1(n13171), .A2(n13565), .A3(n15853), .ZN(n12831) );
  NAND2_X1 U16041 ( .A1(n12831), .A2(n20738), .ZN(n12832) );
  AND2_X1 U16042 ( .A1(n20000), .A2(n12832), .ZN(n15813) );
  NOR2_X1 U16043 ( .A1(n15813), .A2(n20001), .ZN(n20008) );
  INV_X1 U16044 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n20944) );
  INV_X1 U16045 ( .A(n12753), .ZN(n13061) );
  NAND2_X1 U16046 ( .A1(n15808), .A2(n13102), .ZN(n12833) );
  OAI21_X1 U16047 ( .B1(n11283), .B2(n12833), .A(n13126), .ZN(n12836) );
  NAND2_X1 U16048 ( .A1(n13291), .A2(n13080), .ZN(n12834) );
  NOR2_X1 U16049 ( .A1(n12834), .A2(n13179), .ZN(n13103) );
  INV_X1 U16050 ( .A(n13103), .ZN(n13088) );
  OR2_X1 U16051 ( .A1(n13126), .A2(n13088), .ZN(n12835) );
  OAI211_X1 U16052 ( .C1(n12837), .C2(n13061), .A(n12836), .B(n12835), .ZN(
        n15810) );
  NAND2_X1 U16053 ( .A1(n20008), .A2(n15810), .ZN(n12838) );
  OAI21_X1 U16054 ( .B1(n20008), .B2(n20944), .A(n12838), .ZN(P1_U3484) );
  NAND2_X1 U16055 ( .A1(n13398), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12839) );
  AND4_X1 U16056 ( .A1(n19305), .A2(n12839), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19979), .ZN(n12840) );
  NOR2_X1 U16057 ( .A1(n13374), .A2(n12991), .ZN(n12841) );
  AOI21_X1 U16058 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n12991), .A(n12841), .ZN(
        n12842) );
  OAI21_X1 U16059 ( .B1(n19145), .B2(n19961), .A(n12842), .ZN(P2_U2887) );
  AND2_X1 U16060 ( .A1(n12845), .A2(n12844), .ZN(n13421) );
  XOR2_X1 U16061 ( .A(n12846), .B(n13421), .Z(n12853) );
  XOR2_X1 U16062 ( .A(n12848), .B(n12847), .Z(n12849) );
  NOR2_X1 U16063 ( .A1(n12850), .A2(n12849), .ZN(n12851) );
  XNOR2_X1 U16064 ( .A(n12850), .B(n12849), .ZN(n12872) );
  NOR2_X1 U16065 ( .A1(n13805), .A2(n12872), .ZN(n12871) );
  NOR2_X1 U16066 ( .A1(n12851), .A2(n12871), .ZN(n13434) );
  XOR2_X1 U16067 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13434), .Z(
        n12852) );
  NOR2_X1 U16068 ( .A1(n12853), .A2(n12852), .ZN(n13435) );
  AOI21_X1 U16069 ( .B1(n12853), .B2(n12852), .A(n13435), .ZN(n19251) );
  INV_X1 U16070 ( .A(n13616), .ZN(n12856) );
  AND2_X1 U16071 ( .A1(n12657), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19249) );
  AOI21_X1 U16072 ( .B1(n16187), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n19249), .ZN(n12855) );
  OAI21_X1 U16073 ( .B1(n16236), .B2(n12856), .A(n12855), .ZN(n12857) );
  AOI21_X1 U16074 ( .B1(n19251), .B2(n19227), .A(n12857), .ZN(n12866) );
  NAND2_X1 U16075 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12858) );
  NOR2_X1 U16076 ( .A1(n15154), .A2(n12858), .ZN(n12859) );
  OR2_X1 U16077 ( .A1(n12861), .A2(n12859), .ZN(n13826) );
  NOR2_X1 U16078 ( .A1(n12869), .A2(n13826), .ZN(n12860) );
  NAND2_X1 U16079 ( .A1(n12869), .A2(n13826), .ZN(n12868) );
  OAI21_X1 U16080 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12860), .A(
        n12868), .ZN(n12864) );
  OAI21_X1 U16081 ( .B1(n12862), .B2(n12861), .A(n13428), .ZN(n13620) );
  INV_X1 U16082 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19265) );
  XNOR2_X1 U16083 ( .A(n13620), .B(n19265), .ZN(n12863) );
  OR2_X1 U16084 ( .A1(n12864), .A2(n12863), .ZN(n19256) );
  NAND2_X1 U16085 ( .A1(n12864), .A2(n12863), .ZN(n19254) );
  NAND3_X1 U16086 ( .A1(n19256), .A2(n16240), .A3(n19254), .ZN(n12865) );
  OAI211_X1 U16087 ( .C1(n13355), .C2(n19223), .A(n12866), .B(n12865), .ZN(
        P2_U3012) );
  INV_X1 U16088 ( .A(n12867), .ZN(n12877) );
  OAI21_X1 U16089 ( .B1(n13826), .B2(n12869), .A(n12868), .ZN(n12870) );
  XOR2_X1 U16090 ( .A(n12870), .B(n13805), .Z(n15580) );
  AOI21_X1 U16091 ( .B1(n13805), .B2(n12872), .A(n12871), .ZN(n15582) );
  AND2_X1 U16092 ( .A1(n12657), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15581) );
  AOI21_X1 U16093 ( .B1(n19227), .B2(n15582), .A(n15581), .ZN(n12874) );
  NAND2_X1 U16094 ( .A1(n16187), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12873) );
  OAI211_X1 U16095 ( .C1(n16236), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n12874), .B(n12873), .ZN(n12875) );
  AOI21_X1 U16096 ( .B1(n16240), .B2(n15580), .A(n12875), .ZN(n12876) );
  OAI21_X1 U16097 ( .B1(n12877), .B2(n19223), .A(n12876), .ZN(P2_U3013) );
  INV_X1 U16098 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U16099 ( .A1(n12878), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12880) );
  OAI211_X1 U16100 ( .C1(n12996), .C2(n12881), .A(n12880), .B(n12879), .ZN(
        P2_U2962) );
  INV_X1 U16101 ( .A(n13583), .ZN(n13564) );
  OAI21_X1 U16102 ( .B1(n12883), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13564), 
        .ZN(n12884) );
  OAI21_X1 U16103 ( .B1(n12885), .B2(n13564), .A(n12884), .ZN(P1_U3487) );
  AOI21_X1 U16104 ( .B1(n19961), .B2(n19173), .A(n19150), .ZN(n12892) );
  XNOR2_X1 U16105 ( .A(n12887), .B(n12886), .ZN(n13948) );
  NOR2_X1 U16106 ( .A1(n13822), .A2(n19274), .ZN(n12890) );
  INV_X1 U16107 ( .A(n13948), .ZN(n13156) );
  NOR3_X1 U16108 ( .A1(n19961), .A2(n13156), .A3(n16120), .ZN(n12889) );
  AOI211_X1 U16109 ( .C1(P2_EAX_REG_0__SCAN_IN), .C2(n19169), .A(n12890), .B(
        n12889), .ZN(n12891) );
  OAI21_X1 U16110 ( .B1(n12892), .B2(n13948), .A(n12891), .ZN(P2_U2919) );
  INV_X1 U16111 ( .A(n20738), .ZN(n20731) );
  NOR2_X1 U16112 ( .A1(n20731), .A2(n20728), .ZN(n12895) );
  NAND3_X1 U16113 ( .A1(n16039), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n12895), 
        .ZN(n12893) );
  AND4_X1 U16114 ( .A1(n13564), .A2(n20664), .A3(n12894), .A4(n12893), .ZN(
        n12900) );
  NOR2_X1 U16115 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15828) );
  NOR2_X1 U16116 ( .A1(n12900), .A2(n15828), .ZN(n12902) );
  INV_X1 U16117 ( .A(n15853), .ZN(n13118) );
  OR2_X1 U16118 ( .A1(n20192), .A2(n13118), .ZN(n13052) );
  INV_X1 U16119 ( .A(n13052), .ZN(n12899) );
  OAI21_X1 U16120 ( .B1(n20974), .B2(n15853), .A(n13034), .ZN(n12896) );
  AOI21_X1 U16121 ( .B1(n12896), .B2(n12895), .A(n16039), .ZN(n12897) );
  AOI21_X1 U16122 ( .B1(n12899), .B2(n12898), .A(n12897), .ZN(n12901) );
  INV_X1 U16123 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20953) );
  AOI22_X1 U16124 ( .A1(n12902), .A2(n12901), .B1(n12900), .B2(n20953), .ZN(
        P1_U3485) );
  NOR2_X1 U16125 ( .A1(n19148), .A2(n13832), .ZN(n12905) );
  AOI21_X1 U16126 ( .B1(n12867), .B2(n19148), .A(n12905), .ZN(n12906) );
  OAI21_X1 U16127 ( .B1(n19275), .B2(n19145), .A(n12906), .ZN(P2_U2886) );
  AND2_X1 U16128 ( .A1(n16327), .A2(n13398), .ZN(n12908) );
  NAND3_X1 U16129 ( .A1(n12908), .A2(n12907), .A3(n12922), .ZN(n12917) );
  INV_X1 U16130 ( .A(n12908), .ZN(n12911) );
  AOI21_X1 U16131 ( .B1(n12909), .B2(n11415), .A(n11430), .ZN(n12910) );
  NAND2_X1 U16132 ( .A1(n12911), .A2(n12910), .ZN(n12915) );
  MUX2_X1 U16133 ( .A(n12922), .B(n16348), .S(n13398), .Z(n12913) );
  NAND3_X1 U16134 ( .A1(n12913), .A2(n12912), .A3(n19990), .ZN(n12914) );
  NAND4_X1 U16135 ( .A1(n12917), .A2(n12916), .A3(n12915), .A4(n12914), .ZN(
        n12918) );
  NAND2_X1 U16136 ( .A1(n12918), .A2(n16345), .ZN(n12921) );
  INV_X1 U16137 ( .A(n12919), .ZN(n12920) );
  AOI22_X1 U16138 ( .A1(n12925), .A2(n12923), .B1(n19988), .B2(n12922), .ZN(
        n12932) );
  INV_X1 U16139 ( .A(n12924), .ZN(n12926) );
  INV_X1 U16140 ( .A(n12925), .ZN(n19992) );
  OAI21_X1 U16141 ( .B1(n12927), .B2(n12926), .A(n19992), .ZN(n12929) );
  NAND2_X1 U16142 ( .A1(n12929), .A2(n12928), .ZN(n12931) );
  AND4_X1 U16143 ( .A1(n12933), .A2(n12932), .A3(n12931), .A4(n12930), .ZN(
        n12938) );
  NAND2_X1 U16144 ( .A1(n12934), .A2(n13398), .ZN(n13810) );
  NAND2_X1 U16145 ( .A1(n13810), .A2(n12935), .ZN(n12936) );
  NAND2_X1 U16146 ( .A1(n12936), .A2(n19291), .ZN(n12937) );
  AND2_X1 U16147 ( .A1(n12938), .A2(n12937), .ZN(n13808) );
  NAND2_X1 U16148 ( .A1(n13808), .A2(n12939), .ZN(n12940) );
  INV_X1 U16149 ( .A(n13133), .ZN(n12945) );
  INV_X1 U16150 ( .A(n12941), .ZN(n12943) );
  NAND2_X1 U16151 ( .A1(n12943), .A2(n12942), .ZN(n15587) );
  NAND2_X1 U16152 ( .A1(n15587), .A2(n19282), .ZN(n12944) );
  NAND2_X1 U16153 ( .A1(n12945), .A2(n12944), .ZN(n12946) );
  NOR2_X1 U16154 ( .A1(n16328), .A2(n12947), .ZN(n19975) );
  INV_X1 U16155 ( .A(n16321), .ZN(n12949) );
  NAND2_X1 U16156 ( .A1(n16323), .A2(n13398), .ZN(n12948) );
  NAND2_X1 U16157 ( .A1(n12949), .A2(n12948), .ZN(n12950) );
  NAND2_X1 U16158 ( .A1(n12954), .A2(n12950), .ZN(n16290) );
  OAI22_X1 U16159 ( .A1(n16292), .A2(n12951), .B1(n16290), .B2(n13948), .ZN(
        n12952) );
  AOI211_X1 U16160 ( .C1(n19248), .C2(n15590), .A(n12953), .B(n12952), .ZN(
        n12957) );
  NOR2_X1 U16161 ( .A1(n12954), .A2(n15785), .ZN(n19244) );
  AOI22_X1 U16162 ( .A1(n19244), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19255), .B2(n12955), .ZN(n12956) );
  OAI211_X1 U16163 ( .C1(n15787), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12957), .B(n12956), .ZN(P2_U3046) );
  MUX2_X1 U16164 ( .A(n12636), .B(n13355), .S(n19148), .Z(n12960) );
  OAI21_X1 U16165 ( .B1(n19412), .B2(n19145), .A(n12960), .ZN(P2_U2885) );
  XOR2_X1 U16166 ( .A(n12961), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n12964)
         );
  AOI21_X1 U16167 ( .B1(n12962), .B2(n19105), .A(n13017), .ZN(n13702) );
  INV_X1 U16168 ( .A(n13702), .ZN(n19087) );
  MUX2_X1 U16169 ( .A(n12642), .B(n19087), .S(n19148), .Z(n12963) );
  OAI21_X1 U16170 ( .B1(n12964), .B2(n19145), .A(n12963), .ZN(P2_U2882) );
  INV_X1 U16171 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12969) );
  NAND2_X1 U16172 ( .A1(n12753), .A2(n10412), .ZN(n15795) );
  OR2_X1 U16173 ( .A1(n15795), .A2(n15853), .ZN(n13120) );
  NAND2_X1 U16174 ( .A1(n12965), .A2(n13034), .ZN(n13073) );
  NAND2_X1 U16175 ( .A1(n20104), .A2(n13581), .ZN(n13274) );
  NOR2_X1 U16176 ( .A1(n20728), .A2(n15823), .ZN(n20726) );
  INV_X1 U16177 ( .A(n20726), .ZN(n12967) );
  NOR2_X1 U16178 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12967), .ZN(n20120) );
  AOI22_X1 U16179 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20120), .B1(n15855), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12968) );
  OAI21_X1 U16180 ( .B1(n12969), .B2(n13274), .A(n12968), .ZN(P1_U2918) );
  INV_X1 U16181 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14576) );
  AOI22_X1 U16182 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20120), .B1(n15855), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12970) );
  OAI21_X1 U16183 ( .B1(n14576), .B2(n13274), .A(n12970), .ZN(P1_U2917) );
  INV_X1 U16184 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16185 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20120), .B1(n15855), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12971) );
  OAI21_X1 U16186 ( .B1(n12972), .B2(n13274), .A(n12971), .ZN(P1_U2919) );
  INV_X1 U16187 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U16188 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20120), .B1(n15855), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12973) );
  OAI21_X1 U16189 ( .B1(n12974), .B2(n13274), .A(n12973), .ZN(P1_U2920) );
  INV_X1 U16190 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12976) );
  AOI22_X1 U16191 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20130), .B1(n15855), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12975) );
  OAI21_X1 U16192 ( .B1(n12976), .B2(n13274), .A(n12975), .ZN(P1_U2912) );
  AOI22_X1 U16193 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20130), .B1(n15855), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12977) );
  OAI21_X1 U16194 ( .B1(n14548), .B2(n13274), .A(n12977), .ZN(P1_U2911) );
  INV_X1 U16195 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12979) );
  AOI22_X1 U16196 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20130), .B1(n15855), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12978) );
  OAI21_X1 U16197 ( .B1(n12979), .B2(n13274), .A(n12978), .ZN(P1_U2909) );
  INV_X1 U16198 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12981) );
  AOI22_X1 U16199 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20130), .B1(n15855), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12980) );
  OAI21_X1 U16200 ( .B1(n12981), .B2(n13274), .A(n12980), .ZN(P1_U2915) );
  INV_X1 U16201 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12983) );
  AOI22_X1 U16202 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20130), .B1(n15855), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12982) );
  OAI21_X1 U16203 ( .B1(n12983), .B2(n13274), .A(n12982), .ZN(P1_U2916) );
  INV_X1 U16204 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16205 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20130), .B1(n15855), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12984) );
  OAI21_X1 U16206 ( .B1(n12985), .B2(n13274), .A(n12984), .ZN(P1_U2914) );
  BUF_X2 U16207 ( .A(n12990), .Z(n13361) );
  INV_X1 U16208 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13729) );
  MUX2_X1 U16209 ( .A(n12990), .B(n13729), .S(n12991), .Z(n12992) );
  OAI21_X1 U16210 ( .B1(n19566), .B2(n19145), .A(n12992), .ZN(P2_U2884) );
  INV_X1 U16211 ( .A(n16111), .ZN(n19304) );
  XNOR2_X1 U16212 ( .A(n12994), .B(n12993), .ZN(n19080) );
  INV_X1 U16213 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19200) );
  OAI222_X1 U16214 ( .A1(n13822), .A2(n19304), .B1(n19080), .B2(n19179), .C1(
        n15130), .C2(n19200), .ZN(P2_U2913) );
  AOI22_X1 U16215 ( .A1(n19212), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12995) );
  OAI21_X1 U16216 ( .B1(n12996), .B2(n13014), .A(n12995), .ZN(P2_U2925) );
  INV_X1 U16217 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16218 ( .A1(n19212), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12997) );
  OAI21_X1 U16219 ( .B1(n12998), .B2(n13014), .A(n12997), .ZN(P2_U2931) );
  AOI22_X1 U16220 ( .A1(n19212), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12999) );
  OAI21_X1 U16221 ( .B1(n13000), .B2(n13014), .A(n12999), .ZN(P2_U2927) );
  INV_X1 U16222 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U16223 ( .A1(n19212), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13001) );
  OAI21_X1 U16224 ( .B1(n13002), .B2(n13014), .A(n13001), .ZN(P2_U2933) );
  INV_X1 U16225 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13965) );
  AOI22_X1 U16226 ( .A1(n19212), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13003) );
  OAI21_X1 U16227 ( .B1(n13965), .B2(n13014), .A(n13003), .ZN(P2_U2935) );
  INV_X1 U16228 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U16229 ( .A1(n19212), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13004) );
  OAI21_X1 U16230 ( .B1(n13005), .B2(n13014), .A(n13004), .ZN(P2_U2929) );
  INV_X1 U16231 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U16232 ( .A1(n19212), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13006) );
  OAI21_X1 U16233 ( .B1(n13007), .B2(n13014), .A(n13006), .ZN(P2_U2934) );
  INV_X1 U16234 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14269) );
  AOI22_X1 U16235 ( .A1(n19212), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13008) );
  OAI21_X1 U16236 ( .B1(n14269), .B2(n13014), .A(n13008), .ZN(P2_U2922) );
  INV_X1 U16237 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13010) );
  AOI22_X1 U16238 ( .A1(n19212), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13009) );
  OAI21_X1 U16239 ( .B1(n13010), .B2(n13014), .A(n13009), .ZN(P2_U2932) );
  INV_X1 U16240 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U16241 ( .A1(n19212), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13011) );
  OAI21_X1 U16242 ( .B1(n13012), .B2(n13014), .A(n13011), .ZN(P2_U2930) );
  INV_X1 U16243 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U16244 ( .A1(n19212), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13013) );
  OAI21_X1 U16245 ( .B1(n15129), .B2(n13014), .A(n13013), .ZN(P2_U2928) );
  INV_X1 U16246 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13022) );
  NOR2_X1 U16247 ( .A1(n12961), .A2(n12084), .ZN(n13016) );
  OAI211_X1 U16248 ( .C1(n13016), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19127), .B(n13015), .ZN(n13021) );
  OR2_X1 U16249 ( .A1(n13018), .A2(n13017), .ZN(n13019) );
  NAND2_X1 U16250 ( .A1(n13019), .A2(n13042), .ZN(n16245) );
  INV_X1 U16251 ( .A(n16245), .ZN(n19075) );
  NAND2_X1 U16252 ( .A1(n19148), .A2(n19075), .ZN(n13020) );
  OAI211_X1 U16253 ( .C1(n19148), .C2(n13022), .A(n13021), .B(n13020), .ZN(
        P2_U2881) );
  INV_X1 U16254 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20166) );
  NAND2_X1 U16255 ( .A1(n14058), .A2(n20166), .ZN(n13025) );
  NAND2_X1 U16256 ( .A1(n14066), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13024) );
  OAI21_X1 U16257 ( .B1(n10265), .B2(P1_EBX_REG_0__SCAN_IN), .A(n13024), .ZN(
        n13174) );
  NAND2_X1 U16258 ( .A1(n13025), .A2(n13174), .ZN(n13719) );
  NAND2_X1 U16259 ( .A1(n13126), .A2(n13103), .ZN(n13117) );
  OR2_X1 U16260 ( .A1(n13026), .A2(n14068), .ZN(n13027) );
  NAND2_X1 U16261 ( .A1(n13117), .A2(n13027), .ZN(n13028) );
  INV_X1 U16262 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13031) );
  NAND2_X2 U16263 ( .A1(n20103), .A2(n14525), .ZN(n14524) );
  XNOR2_X1 U16264 ( .A(n13030), .B(n13029), .ZN(n13723) );
  OAI222_X1 U16265 ( .A1(n13719), .A2(n14523), .B1(n13031), .B2(n20103), .C1(
        n14524), .C2(n13723), .ZN(P1_U2872) );
  OAI21_X1 U16266 ( .B1(n13033), .B2(n13032), .A(n13605), .ZN(n19060) );
  OAI222_X1 U16267 ( .A1(n13822), .A2(n19308), .B1(n19060), .B2(n19179), .C1(
        n15130), .C2(n19197), .ZN(P2_U2912) );
  NOR2_X1 U16268 ( .A1(n13034), .A2(n20738), .ZN(n13035) );
  OR2_X1 U16269 ( .A1(n9650), .A2(n10412), .ZN(n13194) );
  INV_X1 U16270 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13040) );
  NOR2_X2 U16271 ( .A1(n9650), .A2(n20192), .ZN(n20149) );
  INV_X1 U16272 ( .A(n20149), .ZN(n13039) );
  NOR2_X1 U16273 ( .A1(n14535), .A2(n20906), .ZN(n13037) );
  AOI21_X1 U16274 ( .B1(n14535), .B2(BUF1_REG_15__SCAN_IN), .A(n13037), .ZN(
        n14597) );
  INV_X1 U16275 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13038) );
  OAI222_X1 U16276 ( .A1(n13194), .A2(n13040), .B1(n13039), .B2(n14597), .C1(
        n13038), .C2(n13224), .ZN(P1_U2967) );
  XOR2_X1 U16277 ( .A(n13015), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13046)
         );
  AOI21_X1 U16278 ( .B1(n13043), .B2(n13042), .A(n13041), .ZN(n19059) );
  NOR2_X1 U16279 ( .A1(n19148), .A2(n12643), .ZN(n13044) );
  AOI21_X1 U16280 ( .B1(n19059), .B2(n19148), .A(n13044), .ZN(n13045) );
  OAI21_X1 U16281 ( .B1(n13046), .B2(n19145), .A(n13045), .ZN(P2_U2880) );
  INV_X1 U16282 ( .A(n13047), .ZN(n13049) );
  AOI21_X1 U16283 ( .B1(n13049), .B2(n20166), .A(n13048), .ZN(n13264) );
  INV_X1 U16284 ( .A(n13264), .ZN(n13094) );
  INV_X1 U16285 ( .A(n13050), .ZN(n13051) );
  NAND2_X1 U16286 ( .A1(n13052), .A2(n13051), .ZN(n13057) );
  NAND2_X1 U16287 ( .A1(n20192), .A2(n15853), .ZN(n13580) );
  AND2_X1 U16288 ( .A1(n13580), .A2(n20738), .ZN(n13054) );
  NAND2_X1 U16289 ( .A1(n13581), .A2(n10409), .ZN(n13053) );
  AOI21_X1 U16290 ( .B1(n12965), .B2(n13054), .A(n13053), .ZN(n13055) );
  OR2_X1 U16291 ( .A1(n13126), .A2(n13055), .ZN(n13056) );
  MUX2_X1 U16292 ( .A(n13057), .B(n13056), .S(n10359), .Z(n13063) );
  OAI211_X1 U16293 ( .C1(n20192), .C2(n10415), .A(n13058), .B(n13581), .ZN(
        n13079) );
  NAND2_X1 U16294 ( .A1(n13059), .A2(n13079), .ZN(n13060) );
  NAND2_X1 U16295 ( .A1(n13061), .A2(n13060), .ZN(n13124) );
  NAND3_X1 U16296 ( .A1(n13126), .A2(n15793), .A3(n10412), .ZN(n13062) );
  NAND3_X1 U16297 ( .A1(n13063), .A2(n13124), .A3(n13062), .ZN(n13065) );
  OAI211_X1 U16298 ( .C1(n13070), .C2(n13066), .A(n15808), .B(n13102), .ZN(
        n13067) );
  NOR2_X1 U16299 ( .A1(n13068), .A2(n13067), .ZN(n13069) );
  INV_X1 U16300 ( .A(n13066), .ZN(n13071) );
  NAND2_X1 U16301 ( .A1(n13071), .A2(n13070), .ZN(n13072) );
  AND2_X1 U16302 ( .A1(n13073), .A2(n13072), .ZN(n13074) );
  INV_X1 U16303 ( .A(n13719), .ZN(n13090) );
  INV_X1 U16304 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13075) );
  NOR2_X1 U16305 ( .A1(n20073), .A2(n13075), .ZN(n13263) );
  OAI21_X1 U16306 ( .B1(n13076), .B2(n13581), .A(n13304), .ZN(n13077) );
  OAI211_X1 U16307 ( .C1(n13080), .C2(n14058), .A(n13079), .B(n13078), .ZN(
        n13081) );
  INV_X1 U16308 ( .A(n13081), .ZN(n13083) );
  OAI211_X1 U16309 ( .C1(n13084), .C2(n20192), .A(n13083), .B(n13082), .ZN(
        n13096) );
  OAI21_X1 U16310 ( .B1(n13097), .B2(n13581), .A(n13085), .ZN(n13086) );
  NOR2_X1 U16311 ( .A1(n13096), .A2(n13086), .ZN(n13087) );
  NAND2_X1 U16312 ( .A1(n14892), .A2(n20168), .ZN(n13189) );
  AND2_X1 U16313 ( .A1(n20166), .A2(n13189), .ZN(n13089) );
  AOI211_X1 U16314 ( .C1(n16032), .C2(n13090), .A(n13263), .B(n13089), .ZN(
        n13093) );
  NAND2_X1 U16315 ( .A1(n20073), .A2(n13091), .ZN(n13351) );
  INV_X1 U16316 ( .A(n13351), .ZN(n13187) );
  OAI21_X1 U16317 ( .B1(n13349), .B2(n13187), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13092) );
  OAI211_X1 U16318 ( .C1(n13094), .C2(n20164), .A(n13093), .B(n13092), .ZN(
        P1_U3031) );
  INV_X1 U16319 ( .A(n13096), .ZN(n13101) );
  NAND2_X1 U16320 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  NOR2_X1 U16321 ( .A1(n12965), .A2(n13099), .ZN(n13100) );
  NAND3_X1 U16322 ( .A1(n13101), .A2(n13100), .A3(n13326), .ZN(n15794) );
  INV_X1 U16323 ( .A(n15794), .ZN(n13315) );
  INV_X1 U16324 ( .A(n13102), .ZN(n13104) );
  NOR2_X1 U16325 ( .A1(n13104), .A2(n13103), .ZN(n13311) );
  INV_X1 U16326 ( .A(n13311), .ZN(n13109) );
  NOR2_X1 U16327 ( .A1(n13307), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13309) );
  INV_X1 U16328 ( .A(n13309), .ZN(n13106) );
  INV_X1 U16329 ( .A(n13302), .ZN(n13105) );
  NAND2_X1 U16330 ( .A1(n13106), .A2(n13105), .ZN(n13110) );
  NOR3_X1 U16331 ( .A1(n15795), .A2(n13305), .A3(n13107), .ZN(n13108) );
  AOI21_X1 U16332 ( .B1(n13109), .B2(n13110), .A(n13108), .ZN(n13113) );
  INV_X1 U16333 ( .A(n13110), .ZN(n13116) );
  NAND3_X1 U16334 ( .A1(n13315), .A2(n13111), .A3(n13116), .ZN(n13112) );
  OAI211_X1 U16335 ( .C1(n13095), .C2(n13315), .A(n13113), .B(n13112), .ZN(
        n13301) );
  INV_X1 U16336 ( .A(n20809), .ZN(n13148) );
  NAND2_X1 U16337 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13181) );
  INV_X1 U16338 ( .A(n13181), .ZN(n20803) );
  INV_X1 U16339 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16340 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n14093), .B2(n13114), .ZN(
        n13182) );
  INV_X1 U16341 ( .A(n20801), .ZN(n15829) );
  AOI222_X1 U16342 ( .A1(n13301), .A2(n13148), .B1(n20803), .B2(n13182), .C1(
        n15829), .C2(n13116), .ZN(n13131) );
  INV_X1 U16343 ( .A(n13117), .ZN(n13128) );
  OAI21_X1 U16344 ( .B1(n13291), .B2(n13118), .A(n12965), .ZN(n13119) );
  NAND2_X1 U16345 ( .A1(n13120), .A2(n13119), .ZN(n13121) );
  NAND2_X1 U16346 ( .A1(n13121), .A2(n20738), .ZN(n13125) );
  OR2_X1 U16347 ( .A1(n13572), .A2(n13122), .ZN(n13123) );
  OAI211_X1 U16348 ( .C1(n13126), .C2(n13125), .A(n13124), .B(n13123), .ZN(
        n13127) );
  INV_X1 U16349 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20968) );
  NAND2_X1 U16350 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20726), .ZN(n16045) );
  OAI22_X1 U16351 ( .A1(n15798), .A2(n20001), .B1(n20968), .B2(n16045), .ZN(
        n13147) );
  AOI21_X1 U16352 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n16039), .A(n13147), 
        .ZN(n20806) );
  NAND2_X1 U16353 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20806), .ZN(
        n13130) );
  OAI21_X1 U16354 ( .B1(n13131), .B2(n20806), .A(n13130), .ZN(P1_U3472) );
  INV_X1 U16355 ( .A(n19566), .ZN(n19935) );
  INV_X1 U16356 ( .A(n15860), .ZN(n16350) );
  OR2_X1 U16357 ( .A1(n13361), .A2(n13808), .ZN(n13142) );
  OAI21_X1 U16358 ( .B1(n13133), .B2(n13132), .A(n11319), .ZN(n15600) );
  NOR2_X1 U16359 ( .A1(n13134), .A2(n16308), .ZN(n15598) );
  INV_X1 U16360 ( .A(n15598), .ZN(n15599) );
  INV_X1 U16361 ( .A(n13136), .ZN(n13135) );
  NAND2_X1 U16362 ( .A1(n15587), .A2(n13135), .ZN(n15604) );
  NAND3_X1 U16363 ( .A1(n15600), .A2(n15599), .A3(n15604), .ZN(n13139) );
  NOR2_X1 U16364 ( .A1(n16320), .A2(n16321), .ZN(n15597) );
  AOI21_X1 U16365 ( .B1(n15587), .B2(n13136), .A(n9662), .ZN(n13137) );
  OAI21_X1 U16366 ( .B1(n15597), .B2(n15598), .A(n13137), .ZN(n13138) );
  MUX2_X1 U16367 ( .A(n13139), .B(n13138), .S(n11376), .Z(n13140) );
  INV_X1 U16368 ( .A(n13140), .ZN(n13141) );
  NAND2_X1 U16369 ( .A1(n13142), .A2(n13141), .ZN(n16314) );
  AOI22_X1 U16370 ( .A1(n19935), .A2(n16350), .B1(n19933), .B2(n16314), .ZN(
        n13144) );
  INV_X1 U16371 ( .A(n15611), .ZN(n13817) );
  NAND2_X1 U16372 ( .A1(n13817), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13143) );
  OAI21_X1 U16373 ( .B1(n13144), .B2(n13817), .A(n13143), .ZN(P2_U3596) );
  INV_X1 U16374 ( .A(n20806), .ZN(n20804) );
  INV_X1 U16375 ( .A(n20325), .ZN(n20550) );
  OR2_X1 U16376 ( .A1(n13145), .A2(n20550), .ZN(n13146) );
  XNOR2_X1 U16377 ( .A(n13146), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20090) );
  INV_X1 U16378 ( .A(n13326), .ZN(n13149) );
  NAND4_X1 U16379 ( .A1(n20090), .A2(n13149), .A3(n13148), .A4(n13147), .ZN(
        n13150) );
  OAI21_X1 U16380 ( .B1(n11134), .B2(n20804), .A(n13150), .ZN(P1_U3468) );
  NAND2_X1 U16381 ( .A1(n13152), .A2(n13151), .ZN(n13155) );
  INV_X1 U16382 ( .A(n13153), .ZN(n13154) );
  NAND2_X1 U16383 ( .A1(n13155), .A2(n13154), .ZN(n19957) );
  INV_X1 U16384 ( .A(n19957), .ZN(n13162) );
  NOR2_X1 U16385 ( .A1(n19953), .A2(n19957), .ZN(n13280) );
  AOI21_X1 U16386 ( .B1(n19953), .B2(n19957), .A(n13280), .ZN(n13158) );
  NAND2_X1 U16387 ( .A1(n19536), .A2(n13156), .ZN(n13157) );
  NAND2_X1 U16388 ( .A1(n13158), .A2(n13157), .ZN(n13282) );
  OAI21_X1 U16389 ( .B1(n13158), .B2(n13157), .A(n13282), .ZN(n13159) );
  NAND2_X1 U16390 ( .A1(n13159), .A2(n19173), .ZN(n13161) );
  INV_X1 U16391 ( .A(n13822), .ZN(n19171) );
  AOI22_X1 U16392 ( .A1(n19171), .A2(n13955), .B1(n19169), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13160) );
  OAI211_X1 U16393 ( .C1(n13162), .C2(n16119), .A(n13161), .B(n13160), .ZN(
        P2_U2918) );
  NAND2_X1 U16394 ( .A1(n10415), .A2(n14525), .ZN(n13165) );
  NAND2_X1 U16395 ( .A1(n13519), .A2(DATAI_1_), .ZN(n13164) );
  NAND2_X1 U16396 ( .A1(n14535), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13163) );
  AND2_X1 U16397 ( .A1(n13164), .A2(n13163), .ZN(n20193) );
  XNOR2_X1 U16398 ( .A(n13167), .B(n13166), .ZN(n13590) );
  INV_X1 U16399 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20128) );
  OAI222_X1 U16400 ( .A1(n14602), .A2(n20193), .B1(n14605), .B2(n13590), .C1(
        n20128), .C2(n14603), .ZN(P1_U2903) );
  NAND2_X1 U16401 ( .A1(n13519), .A2(DATAI_0_), .ZN(n13169) );
  NAND2_X1 U16402 ( .A1(n14535), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13168) );
  AND2_X1 U16403 ( .A1(n13169), .A2(n13168), .ZN(n20185) );
  INV_X1 U16404 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20133) );
  OAI222_X1 U16405 ( .A1(n14602), .A2(n20185), .B1(n14605), .B2(n13723), .C1(
        n20133), .C2(n14603), .ZN(P1_U2904) );
  NAND2_X1 U16406 ( .A1(n14066), .A2(n13114), .ZN(n13170) );
  INV_X1 U16407 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13575) );
  NAND2_X1 U16408 ( .A1(n10265), .A2(n13575), .ZN(n13172) );
  NAND2_X1 U16409 ( .A1(n13173), .A2(n13172), .ZN(n13247) );
  XNOR2_X1 U16410 ( .A(n13247), .B(n13174), .ZN(n13578) );
  XNOR2_X1 U16411 ( .A(n13578), .B(n13291), .ZN(n13192) );
  AOI22_X1 U16412 ( .A1(n20098), .A2(n13192), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14485), .ZN(n13175) );
  OAI21_X1 U16413 ( .B1(n13590), .B2(n14524), .A(n13175), .ZN(P1_U2871) );
  INV_X1 U16414 ( .A(n9637), .ZN(n20625) );
  INV_X1 U16415 ( .A(n13177), .ZN(n13323) );
  INV_X1 U16416 ( .A(n13307), .ZN(n13178) );
  NAND2_X1 U16417 ( .A1(n13323), .A2(n13178), .ZN(n13183) );
  OAI22_X1 U16418 ( .A1(n15795), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n13183), .B2(n13179), .ZN(n13180) );
  AOI21_X1 U16419 ( .B1(n20625), .B2(n15794), .A(n13180), .ZN(n15797) );
  NOR2_X1 U16420 ( .A1(n15797), .A2(n20809), .ZN(n13185) );
  OAI22_X1 U16421 ( .A1(n20801), .A2(n13183), .B1(n13182), .B2(n13181), .ZN(
        n13184) );
  OAI21_X1 U16422 ( .B1(n13185), .B2(n13184), .A(n20804), .ZN(n13186) );
  OAI21_X1 U16423 ( .B1(n20804), .B2(n10469), .A(n13186), .ZN(P1_U3473) );
  INV_X1 U16424 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20824) );
  OAI221_X1 U16425 ( .B1(n13187), .B2(n20166), .C1(n13187), .C2(n13189), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13188) );
  OAI21_X1 U16426 ( .B1(n20073), .B2(n20824), .A(n13188), .ZN(n13191) );
  NOR2_X2 U16427 ( .A1(n13189), .A2(n13349), .ZN(n14939) );
  AOI211_X1 U16428 ( .C1(n20166), .C2(n14890), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n14939), .ZN(n13190) );
  AOI211_X1 U16429 ( .C1(n16032), .C2(n13192), .A(n13191), .B(n13190), .ZN(
        n13193) );
  OAI21_X1 U16430 ( .B1(n13557), .B2(n20164), .A(n13193), .ZN(P1_U3030) );
  AOI22_X1 U16431 ( .A1(n20161), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n9650), .ZN(n13196) );
  INV_X1 U16432 ( .A(n20185), .ZN(n13195) );
  NAND2_X1 U16433 ( .A1(n20149), .A2(n13195), .ZN(n13227) );
  NAND2_X1 U16434 ( .A1(n13196), .A2(n13227), .ZN(P1_U2952) );
  AOI22_X1 U16435 ( .A1(n20161), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n9650), .ZN(n13198) );
  INV_X1 U16436 ( .A(n20193), .ZN(n13197) );
  NAND2_X1 U16437 ( .A1(n20149), .A2(n13197), .ZN(n13229) );
  NAND2_X1 U16438 ( .A1(n13198), .A2(n13229), .ZN(P1_U2953) );
  AOI22_X1 U16439 ( .A1(n20161), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n9650), .ZN(n13202) );
  NAND2_X1 U16440 ( .A1(n13519), .A2(DATAI_2_), .ZN(n13200) );
  NAND2_X1 U16441 ( .A1(n14535), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13199) );
  AND2_X1 U16442 ( .A1(n13200), .A2(n13199), .ZN(n20199) );
  INV_X1 U16443 ( .A(n20199), .ZN(n13201) );
  NAND2_X1 U16444 ( .A1(n20149), .A2(n13201), .ZN(n13241) );
  NAND2_X1 U16445 ( .A1(n13202), .A2(n13241), .ZN(P1_U2954) );
  AOI22_X1 U16446 ( .A1(n20161), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n9650), .ZN(n13206) );
  NAND2_X1 U16447 ( .A1(n13519), .A2(DATAI_3_), .ZN(n13204) );
  NAND2_X1 U16448 ( .A1(n14535), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13203) );
  AND2_X1 U16449 ( .A1(n13204), .A2(n13203), .ZN(n20206) );
  INV_X1 U16450 ( .A(n20206), .ZN(n13205) );
  NAND2_X1 U16451 ( .A1(n20149), .A2(n13205), .ZN(n13231) );
  NAND2_X1 U16452 ( .A1(n13206), .A2(n13231), .ZN(P1_U2955) );
  AOI22_X1 U16453 ( .A1(n20161), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n9650), .ZN(n13210) );
  INV_X1 U16454 ( .A(DATAI_5_), .ZN(n13208) );
  INV_X1 U16455 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13207) );
  MUX2_X1 U16456 ( .A(n13208), .B(n13207), .S(n14535), .Z(n20214) );
  INV_X1 U16457 ( .A(n20214), .ZN(n13209) );
  NAND2_X1 U16458 ( .A1(n20149), .A2(n13209), .ZN(n13225) );
  NAND2_X1 U16459 ( .A1(n13210), .A2(n13225), .ZN(P1_U2957) );
  AOI22_X1 U16460 ( .A1(n20161), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n9650), .ZN(n13213) );
  INV_X1 U16461 ( .A(DATAI_4_), .ZN(n13212) );
  NAND2_X1 U16462 ( .A1(n14535), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13211) );
  OAI21_X1 U16463 ( .B1(n14535), .B2(n13212), .A(n13211), .ZN(n14570) );
  NAND2_X1 U16464 ( .A1(n20149), .A2(n14570), .ZN(n13235) );
  NAND2_X1 U16465 ( .A1(n13213), .A2(n13235), .ZN(P1_U2956) );
  AOI22_X1 U16466 ( .A1(n20161), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n9650), .ZN(n13216) );
  INV_X1 U16467 ( .A(DATAI_7_), .ZN(n13215) );
  NAND2_X1 U16468 ( .A1(n14535), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13214) );
  OAI21_X1 U16469 ( .B1(n14535), .B2(n13215), .A(n13214), .ZN(n14555) );
  NAND2_X1 U16470 ( .A1(n20149), .A2(n14555), .ZN(n13239) );
  NAND2_X1 U16471 ( .A1(n13216), .A2(n13239), .ZN(P1_U2959) );
  AOI22_X1 U16472 ( .A1(n20161), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n9650), .ZN(n13219) );
  INV_X1 U16473 ( .A(DATAI_6_), .ZN(n13218) );
  NAND2_X1 U16474 ( .A1(n14535), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13217) );
  OAI21_X1 U16475 ( .B1(n14535), .B2(n13218), .A(n13217), .ZN(n14559) );
  NAND2_X1 U16476 ( .A1(n20149), .A2(n14559), .ZN(n13237) );
  NAND2_X1 U16477 ( .A1(n13219), .A2(n13237), .ZN(P1_U2958) );
  AOI22_X1 U16478 ( .A1(n20161), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n9650), .ZN(n13223) );
  INV_X1 U16479 ( .A(DATAI_11_), .ZN(n13221) );
  MUX2_X1 U16480 ( .A(n13221), .B(n13220), .S(n14535), .Z(n14541) );
  INV_X1 U16481 ( .A(n14541), .ZN(n13222) );
  NAND2_X1 U16482 ( .A1(n20149), .A2(n13222), .ZN(n13233) );
  NAND2_X1 U16483 ( .A1(n13223), .A2(n13233), .ZN(P1_U2948) );
  AOI22_X1 U16484 ( .A1(n20161), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n9650), .ZN(n13226) );
  NAND2_X1 U16485 ( .A1(n13226), .A2(n13225), .ZN(P1_U2942) );
  AOI22_X1 U16486 ( .A1(n20161), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n9650), .ZN(n13228) );
  NAND2_X1 U16487 ( .A1(n13228), .A2(n13227), .ZN(P1_U2937) );
  AOI22_X1 U16488 ( .A1(n20161), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n9650), .ZN(n13230) );
  NAND2_X1 U16489 ( .A1(n13230), .A2(n13229), .ZN(P1_U2938) );
  AOI22_X1 U16490 ( .A1(n20161), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n9650), .ZN(n13232) );
  NAND2_X1 U16491 ( .A1(n13232), .A2(n13231), .ZN(P1_U2940) );
  AOI22_X1 U16492 ( .A1(n20161), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n9650), .ZN(n13234) );
  NAND2_X1 U16493 ( .A1(n13234), .A2(n13233), .ZN(P1_U2963) );
  AOI22_X1 U16494 ( .A1(n20161), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n9650), .ZN(n13236) );
  NAND2_X1 U16495 ( .A1(n13236), .A2(n13235), .ZN(P1_U2941) );
  AOI22_X1 U16496 ( .A1(n20161), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n9650), .ZN(n13238) );
  NAND2_X1 U16497 ( .A1(n13238), .A2(n13237), .ZN(P1_U2943) );
  AOI22_X1 U16498 ( .A1(n20161), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n9650), .ZN(n13240) );
  NAND2_X1 U16499 ( .A1(n13240), .A2(n13239), .ZN(P1_U2944) );
  AOI22_X1 U16500 ( .A1(n20161), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n9650), .ZN(n13242) );
  NAND2_X1 U16501 ( .A1(n13242), .A2(n13241), .ZN(P1_U2939) );
  NAND2_X1 U16502 ( .A1(n13244), .A2(n13243), .ZN(n13245) );
  NAND2_X1 U16503 ( .A1(n13246), .A2(n13245), .ZN(n13774) );
  INV_X1 U16504 ( .A(n13247), .ZN(n13248) );
  AOI21_X1 U16505 ( .B1(n13578), .B2(n13291), .A(n13248), .ZN(n13253) );
  NAND2_X1 U16506 ( .A1(n14066), .A2(n20180), .ZN(n13249) );
  OAI211_X1 U16507 ( .C1(n14068), .C2(P1_EBX_REG_2__SCAN_IN), .A(n13249), .B(
        n14293), .ZN(n13251) );
  INV_X1 U16508 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13765) );
  NAND2_X1 U16509 ( .A1(n10265), .A2(n13765), .ZN(n13250) );
  NAND2_X1 U16510 ( .A1(n13251), .A2(n13250), .ZN(n13252) );
  NAND2_X1 U16511 ( .A1(n13253), .A2(n13252), .ZN(n13295) );
  OAI21_X1 U16512 ( .B1(n13253), .B2(n13252), .A(n13295), .ZN(n20172) );
  INV_X1 U16513 ( .A(n20172), .ZN(n13254) );
  AOI22_X1 U16514 ( .A1(n20098), .A2(n13254), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14485), .ZN(n13255) );
  OAI21_X1 U16515 ( .B1(n13774), .B2(n14524), .A(n13255), .ZN(P1_U2870) );
  XNOR2_X1 U16516 ( .A(n13256), .B(n19133), .ZN(n13259) );
  AOI21_X1 U16517 ( .B1(n13257), .B2(n13609), .A(n9759), .ZN(n16215) );
  INV_X1 U16518 ( .A(n16215), .ZN(n19048) );
  MUX2_X1 U16519 ( .A(n12644), .B(n19048), .S(n19148), .Z(n13258) );
  OAI21_X1 U16520 ( .B1(n13259), .B2(n19145), .A(n13258), .ZN(P2_U2878) );
  INV_X1 U16521 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13260) );
  AOI21_X1 U16522 ( .B1(n14772), .B2(n13261), .A(n13260), .ZN(n13262) );
  AOI211_X1 U16523 ( .C1(n13264), .C2(n15959), .A(n13263), .B(n13262), .ZN(
        n13265) );
  OAI21_X1 U16524 ( .B1(n13723), .B2(n15934), .A(n13265), .ZN(P1_U2999) );
  INV_X1 U16525 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20126) );
  OAI222_X1 U16526 ( .A1(n14605), .A2(n13774), .B1(n14603), .B2(n20126), .C1(
        n14602), .C2(n20199), .ZN(P1_U2902) );
  INV_X1 U16527 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13267) );
  AOI22_X1 U16528 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13266) );
  OAI21_X1 U16529 ( .B1(n13267), .B2(n13274), .A(n13266), .ZN(P1_U2910) );
  AOI22_X1 U16530 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13268) );
  OAI21_X1 U16531 ( .B1(n14537), .B2(n13274), .A(n13268), .ZN(P1_U2908) );
  INV_X1 U16532 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13270) );
  AOI22_X1 U16533 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13269) );
  OAI21_X1 U16534 ( .B1(n13270), .B2(n13274), .A(n13269), .ZN(P1_U2907) );
  INV_X1 U16535 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13272) );
  AOI22_X1 U16536 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13271) );
  OAI21_X1 U16537 ( .B1(n13272), .B2(n13274), .A(n13271), .ZN(P1_U2913) );
  INV_X1 U16538 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13275) );
  AOI22_X1 U16539 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20130), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20129), .ZN(n13273) );
  OAI21_X1 U16540 ( .B1(n13275), .B2(n13274), .A(n13273), .ZN(P1_U2906) );
  NAND2_X1 U16541 ( .A1(n13277), .A2(n13276), .ZN(n13279) );
  AND2_X1 U16542 ( .A1(n13279), .A2(n10134), .ZN(n19943) );
  INV_X1 U16543 ( .A(n19412), .ZN(n19948) );
  INV_X1 U16544 ( .A(n19943), .ZN(n19263) );
  NOR2_X1 U16545 ( .A1(n19948), .A2(n19263), .ZN(n13339) );
  AOI21_X1 U16546 ( .B1(n19948), .B2(n19263), .A(n13339), .ZN(n13284) );
  INV_X1 U16547 ( .A(n13280), .ZN(n13281) );
  NAND2_X1 U16548 ( .A1(n13282), .A2(n13281), .ZN(n13283) );
  NAND2_X1 U16549 ( .A1(n13284), .A2(n13283), .ZN(n13341) );
  OAI21_X1 U16550 ( .B1(n13284), .B2(n13283), .A(n13341), .ZN(n13285) );
  NAND2_X1 U16551 ( .A1(n13285), .A2(n19173), .ZN(n13287) );
  AOI22_X1 U16552 ( .A1(n19171), .A2(n16126), .B1(n19169), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13286) );
  OAI211_X1 U16553 ( .C1(n19943), .C2(n16119), .A(n13287), .B(n13286), .ZN(
        P2_U2917) );
  NOR2_X1 U16554 ( .A1(n13289), .A2(n13288), .ZN(n13290) );
  OR2_X1 U16555 ( .A1(n13441), .A2(n13290), .ZN(n13794) );
  MUX2_X1 U16556 ( .A(n14057), .B(n14293), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13293) );
  NAND2_X1 U16557 ( .A1(n14058), .A2(n11188), .ZN(n13292) );
  NAND2_X1 U16558 ( .A1(n13293), .A2(n13292), .ZN(n13294) );
  NAND2_X1 U16559 ( .A1(n13295), .A2(n13294), .ZN(n13296) );
  AND2_X1 U16560 ( .A1(n13447), .A2(n13296), .ZN(n13785) );
  AOI22_X1 U16561 ( .A1(n20098), .A2(n13785), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14485), .ZN(n13297) );
  OAI21_X1 U16562 ( .B1(n13794), .B2(n14524), .A(n13297), .ZN(P1_U2869) );
  INV_X1 U16563 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20124) );
  OAI222_X1 U16564 ( .A1(n14605), .A2(n13794), .B1(n14603), .B2(n20124), .C1(
        n14602), .C2(n20206), .ZN(P1_U2901) );
  INV_X1 U16565 ( .A(n15097), .ZN(n13300) );
  OR2_X1 U16566 ( .A1(n13298), .A2(n9750), .ZN(n13299) );
  NAND2_X1 U16567 ( .A1(n13299), .A2(n15036), .ZN(n19025) );
  INV_X1 U16568 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19189) );
  OAI222_X1 U16569 ( .A1(n13822), .A2(n13300), .B1(n19025), .B2(n19179), .C1(
        n15130), .C2(n19189), .ZN(P2_U2908) );
  NOR2_X1 U16570 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15823), .ZN(n13319) );
  MUX2_X1 U16571 ( .A(n13301), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15798), .Z(n15803) );
  AOI22_X1 U16572 ( .A1(n13319), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15823), .B2(n15803), .ZN(n13322) );
  NAND2_X1 U16573 ( .A1(n20813), .A2(n15794), .ZN(n13317) );
  NOR2_X1 U16574 ( .A1(n13302), .A2(n10613), .ZN(n13303) );
  NOR2_X1 U16575 ( .A1(n10396), .A2(n13303), .ZN(n20796) );
  NOR2_X1 U16576 ( .A1(n13304), .A2(n20796), .ZN(n13314) );
  XNOR2_X1 U16577 ( .A(n13305), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13312) );
  INV_X1 U16578 ( .A(n13306), .ZN(n13308) );
  OAI22_X1 U16579 ( .A1(n13309), .A2(n10613), .B1(n13308), .B2(n13307), .ZN(
        n13310) );
  OAI22_X1 U16580 ( .A1(n15795), .A2(n13312), .B1(n13311), .B2(n13310), .ZN(
        n13313) );
  AOI21_X1 U16581 ( .B1(n13315), .B2(n13314), .A(n13313), .ZN(n13316) );
  NAND2_X1 U16582 ( .A1(n13317), .A2(n13316), .ZN(n20795) );
  NOR2_X1 U16583 ( .A1(n13325), .A2(n10613), .ZN(n13318) );
  AOI21_X1 U16584 ( .B1(n20795), .B2(n13325), .A(n13318), .ZN(n15804) );
  INV_X1 U16585 ( .A(n15804), .ZN(n13320) );
  AOI22_X1 U16586 ( .A1(n13320), .A2(n15823), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13319), .ZN(n13321) );
  INV_X1 U16587 ( .A(n15814), .ZN(n13324) );
  NAND2_X1 U16588 ( .A1(n13324), .A2(n13323), .ZN(n13333) );
  NAND2_X1 U16589 ( .A1(n13325), .A2(n15823), .ZN(n13327) );
  NOR2_X1 U16590 ( .A1(n13327), .A2(n13326), .ZN(n13330) );
  NAND2_X1 U16591 ( .A1(n13327), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13328) );
  NOR2_X1 U16592 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13328), .ZN(n13329) );
  AOI21_X1 U16593 ( .B1(n20090), .B2(n13330), .A(n13329), .ZN(n15816) );
  AND3_X1 U16594 ( .A1(n13333), .A2(n15816), .A3(n20968), .ZN(n13331) );
  AND2_X1 U16595 ( .A1(n15816), .A2(n20726), .ZN(n13332) );
  AND2_X1 U16596 ( .A1(n13333), .A2(n13332), .ZN(n15824) );
  INV_X1 U16597 ( .A(n9664), .ZN(n13334) );
  NAND2_X1 U16598 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n13115), .ZN(n20814) );
  INV_X1 U16599 ( .A(n20814), .ZN(n14947) );
  OAI22_X1 U16600 ( .A1(n20261), .A2(n20664), .B1(n13334), .B2(n14947), .ZN(
        n13335) );
  OAI21_X1 U16601 ( .B1(n15824), .B2(n13335), .A(n20823), .ZN(n13336) );
  OAI21_X1 U16602 ( .B1(n20823), .B2(n20588), .A(n13336), .ZN(P1_U3478) );
  XNOR2_X1 U16603 ( .A(n13337), .B(n13338), .ZN(n16291) );
  XOR2_X1 U16604 ( .A(n16291), .B(n19566), .Z(n13343) );
  INV_X1 U16605 ( .A(n13339), .ZN(n13340) );
  NAND2_X1 U16606 ( .A1(n13341), .A2(n13340), .ZN(n13342) );
  NAND2_X1 U16607 ( .A1(n13342), .A2(n13343), .ZN(n13455) );
  OAI21_X1 U16608 ( .B1(n13343), .B2(n13342), .A(n13455), .ZN(n13344) );
  NAND2_X1 U16609 ( .A1(n13344), .A2(n19173), .ZN(n13346) );
  AOI22_X1 U16610 ( .A1(n19171), .A2(n15145), .B1(n19169), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n13345) );
  OAI211_X1 U16611 ( .C1(n16291), .C2(n16119), .A(n13346), .B(n13345), .ZN(
        P2_U2916) );
  XNOR2_X1 U16612 ( .A(n13348), .B(n13347), .ZN(n13506) );
  NAND2_X1 U16613 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20167) );
  INV_X1 U16614 ( .A(n14892), .ZN(n13350) );
  OAI21_X1 U16615 ( .B1(n14892), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13351), .ZN(n14894) );
  AOI21_X1 U16616 ( .B1(n20167), .B2(n14913), .A(n14894), .ZN(n20179) );
  AOI21_X1 U16617 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14012) );
  NAND2_X1 U16618 ( .A1(n14916), .A2(n14012), .ZN(n20169) );
  NAND2_X1 U16619 ( .A1(n20179), .A2(n20169), .ZN(n13547) );
  OAI21_X1 U16620 ( .B1(n14892), .B2(n20166), .A(n14890), .ZN(n14838) );
  NAND2_X1 U16621 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14838), .ZN(
        n20181) );
  NOR2_X1 U16622 ( .A1(n20180), .A2(n20181), .ZN(n14920) );
  NOR2_X1 U16623 ( .A1(n14916), .A2(n14920), .ZN(n14912) );
  AOI22_X1 U16624 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13547), .B1(
        n15998), .B2(n11188), .ZN(n13353) );
  AND2_X1 U16625 ( .A1(n9645), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13501) );
  AOI21_X1 U16626 ( .B1(n16032), .B2(n13785), .A(n13501), .ZN(n13352) );
  OAI211_X1 U16627 ( .C1(n20164), .C2(n13506), .A(n13353), .B(n13352), .ZN(
        P1_U3028) );
  INV_X1 U16628 ( .A(n13354), .ZN(n13400) );
  INV_X1 U16629 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13357) );
  NAND2_X2 U16630 ( .A1(n13355), .A2(n13361), .ZN(n13388) );
  INV_X1 U16631 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13356) );
  OAI22_X1 U16632 ( .A1(n13357), .A2(n19677), .B1(n13658), .B2(n13356), .ZN(
        n13365) );
  OR2_X2 U16633 ( .A1(n13361), .A2(n12843), .ZN(n13384) );
  INV_X1 U16634 ( .A(n13359), .ZN(n13360) );
  NOR2_X1 U16635 ( .A1(n13358), .A2(n13360), .ZN(n13367) );
  INV_X1 U16636 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13363) );
  NAND2_X1 U16637 ( .A1(n13361), .A2(n12843), .ZN(n13390) );
  INV_X1 U16638 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13362) );
  OAI22_X1 U16639 ( .A1(n19640), .A2(n13363), .B1(n19411), .B2(n13362), .ZN(
        n13364) );
  NOR2_X1 U16640 ( .A1(n13365), .A2(n13364), .ZN(n13397) );
  INV_X1 U16641 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13369) );
  NAND2_X1 U16642 ( .A1(n15590), .A2(n13366), .ZN(n13387) );
  INV_X1 U16643 ( .A(n13367), .ZN(n13389) );
  INV_X1 U16645 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13368) );
  OAI22_X1 U16646 ( .A1(n13369), .A2(n13866), .B1(n19380), .B2(n13368), .ZN(
        n13373) );
  INV_X1 U16647 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13371) );
  OR2_X2 U16648 ( .A1(n13390), .A2(n13387), .ZN(n19440) );
  INV_X1 U16649 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13370) );
  OAI22_X1 U16650 ( .A1(n19785), .A2(n13371), .B1(n19440), .B2(n13370), .ZN(
        n13372) );
  NOR2_X1 U16651 ( .A1(n13373), .A2(n13372), .ZN(n13396) );
  INV_X1 U16652 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13376) );
  INV_X1 U16653 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13375) );
  OAI22_X1 U16654 ( .A1(n13376), .A2(n13654), .B1(n19351), .B2(n13375), .ZN(
        n13381) );
  INV_X1 U16655 ( .A(n13377), .ZN(n13378) );
  OR2_X2 U16656 ( .A1(n13390), .A2(n13383), .ZN(n19469) );
  INV_X1 U16657 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13379) );
  NOR2_X1 U16658 ( .A1(n13381), .A2(n13380), .ZN(n13395) );
  INV_X1 U16659 ( .A(n13387), .ZN(n13382) );
  INV_X1 U16660 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13386) );
  NOR2_X2 U16661 ( .A1(n13384), .A2(n13383), .ZN(n19606) );
  NAND2_X1 U16662 ( .A1(n19606), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13385) );
  OAI21_X1 U16663 ( .B1(n19572), .B2(n13386), .A(n13385), .ZN(n13393) );
  INV_X1 U16664 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13391) );
  OR2_X2 U16665 ( .A1(n13390), .A2(n13389), .ZN(n19504) );
  OAI22_X1 U16666 ( .A1(n13881), .A2(n13391), .B1(n19504), .B2(n19522), .ZN(
        n13392) );
  NOR2_X1 U16667 ( .A1(n13393), .A2(n13392), .ZN(n13394) );
  NAND4_X1 U16668 ( .A1(n13397), .A2(n13396), .A3(n13395), .A4(n13394), .ZN(
        n13399) );
  INV_X1 U16669 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13402) );
  INV_X1 U16670 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13401) );
  INV_X1 U16671 ( .A(n13403), .ZN(n13407) );
  INV_X1 U16672 ( .A(n19351), .ZN(n19346) );
  AOI22_X1 U16673 ( .A1(n19346), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n19606), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13405) );
  INV_X1 U16674 ( .A(n19640), .ZN(n13648) );
  AOI22_X1 U16675 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n13648), .B1(
        n13649), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13404) );
  INV_X1 U16676 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13409) );
  INV_X1 U16677 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13408) );
  OAI22_X1 U16678 ( .A1(n19785), .A2(n13409), .B1(n19411), .B2(n13408), .ZN(
        n13413) );
  INV_X1 U16679 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13411) );
  INV_X1 U16680 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13410) );
  OAI22_X1 U16681 ( .A1(n13411), .A2(n19504), .B1(n19440), .B2(n13410), .ZN(
        n13412) );
  NOR2_X1 U16682 ( .A1(n13413), .A2(n13412), .ZN(n13420) );
  INV_X1 U16683 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13415) );
  INV_X1 U16684 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13414) );
  OAI22_X1 U16685 ( .A1(n13881), .A2(n13415), .B1(n19469), .B2(n13414), .ZN(
        n13416) );
  INV_X1 U16686 ( .A(n13416), .ZN(n13419) );
  INV_X1 U16687 ( .A(n19677), .ZN(n19671) );
  AOI21_X1 U16688 ( .B1(n19671), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n19282), .ZN(n13418) );
  INV_X1 U16689 ( .A(n13654), .ZN(n19743) );
  NAND2_X1 U16690 ( .A1(n19743), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13417) );
  INV_X1 U16691 ( .A(n13421), .ZN(n13423) );
  NAND2_X1 U16692 ( .A1(n13423), .A2(n13422), .ZN(n13424) );
  INV_X1 U16693 ( .A(n13427), .ZN(n13640) );
  NAND2_X1 U16694 ( .A1(n13429), .A2(n13428), .ZN(n13430) );
  NAND2_X1 U16695 ( .A1(n13640), .A2(n13430), .ZN(n13728) );
  OAI21_X1 U16696 ( .B1(n13620), .B2(n19265), .A(n19256), .ZN(n13636) );
  XNOR2_X1 U16697 ( .A(n13636), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13431) );
  XNOR2_X1 U16698 ( .A(n13637), .B(n13431), .ZN(n16297) );
  INV_X1 U16699 ( .A(n16297), .ZN(n13439) );
  INV_X1 U16700 ( .A(n13361), .ZN(n16288) );
  NOR2_X1 U16701 ( .A1(n19066), .A2(n13432), .ZN(n16287) );
  INV_X1 U16702 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13727) );
  OAI22_X1 U16703 ( .A1(n13727), .A2(n19231), .B1(n16236), .B2(n13725), .ZN(
        n13433) );
  AOI211_X1 U16704 ( .C1(n16239), .C2(n16288), .A(n16287), .B(n13433), .ZN(
        n13438) );
  NOR2_X1 U16705 ( .A1(n13434), .A2(n19265), .ZN(n13436) );
  NOR2_X1 U16706 ( .A1(n13436), .A2(n13435), .ZN(n13677) );
  OR3_X1 U16707 ( .A1(n16293), .A2(n16294), .A3(n16251), .ZN(n13437) );
  OAI211_X1 U16708 ( .C1(n13439), .C2(n19224), .A(n13438), .B(n13437), .ZN(
        P2_U3011) );
  OAI21_X1 U16709 ( .B1(n13441), .B2(n13440), .A(n13496), .ZN(n13481) );
  INV_X1 U16710 ( .A(n14570), .ZN(n13540) );
  OAI222_X1 U16711 ( .A1(n13481), .A2(n14605), .B1(n20122), .B2(n14603), .C1(
        n14602), .C2(n13540), .ZN(P1_U2900) );
  INV_X1 U16712 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13449) );
  OAI21_X1 U16713 ( .B1(n10265), .B2(n13442), .A(n14066), .ZN(n13443) );
  OAI21_X1 U16714 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n14068), .A(n13443), .ZN(
        n13445) );
  NAND2_X1 U16715 ( .A1(n10265), .A2(n13449), .ZN(n13444) );
  AND2_X1 U16716 ( .A1(n13445), .A2(n13444), .ZN(n13446) );
  AND2_X1 U16717 ( .A1(n13447), .A2(n13446), .ZN(n13448) );
  OR2_X1 U16718 ( .A1(n13448), .A2(n13531), .ZN(n20085) );
  OAI222_X1 U16719 ( .A1(n13481), .A2(n14524), .B1(n13449), .B2(n20103), .C1(
        n20085), .C2(n14523), .ZN(P1_U2868) );
  XNOR2_X1 U16720 ( .A(n13451), .B(n13450), .ZN(n13485) );
  NAND2_X1 U16721 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13546) );
  OAI211_X1 U16722 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n15998), .B(n13546), .ZN(n13454) );
  INV_X1 U16723 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20748) );
  OAI22_X1 U16724 ( .A1(n20173), .A2(n20085), .B1(n20748), .B2(n20073), .ZN(
        n13452) );
  AOI21_X1 U16725 ( .B1(n13547), .B2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13452), .ZN(n13453) );
  OAI211_X1 U16726 ( .C1(n20164), .C2(n13485), .A(n13454), .B(n13453), .ZN(
        P1_U3027) );
  INV_X1 U16727 ( .A(n16117), .ZN(n19294) );
  INV_X1 U16728 ( .A(n16291), .ZN(n19939) );
  OAI21_X1 U16729 ( .B1(n19935), .B2(n19939), .A(n13455), .ZN(n13458) );
  OR2_X1 U16730 ( .A1(n13456), .A2(n9767), .ZN(n13457) );
  NAND2_X1 U16731 ( .A1(n13457), .A2(n10136), .ZN(n19097) );
  NAND2_X1 U16732 ( .A1(n13458), .A2(n19097), .ZN(n19175) );
  OR2_X1 U16733 ( .A1(n13460), .A2(n13459), .ZN(n13461) );
  NAND2_X1 U16734 ( .A1(n12961), .A2(n13461), .ZN(n19172) );
  XNOR2_X1 U16735 ( .A(n19175), .B(n19172), .ZN(n13462) );
  NAND2_X1 U16736 ( .A1(n13462), .A2(n19173), .ZN(n13464) );
  INV_X1 U16737 ( .A(n19097), .ZN(n19236) );
  AOI22_X1 U16738 ( .A1(n19150), .A2(n19236), .B1(n19169), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13463) );
  OAI211_X1 U16739 ( .C1(n19294), .C2(n13822), .A(n13464), .B(n13463), .ZN(
        P2_U2915) );
  OR2_X1 U16740 ( .A1(n16209), .A2(n13465), .ZN(n13466) );
  AND2_X1 U16741 ( .A1(n13466), .A2(n15033), .ZN(n19024) );
  NOR2_X1 U16742 ( .A1(n19148), .A2(n19031), .ZN(n13472) );
  AOI211_X1 U16743 ( .C1(n13470), .C2(n13467), .A(n19145), .B(n13469), .ZN(
        n13471) );
  AOI211_X1 U16744 ( .C1(n19024), .C2(n19148), .A(n13472), .B(n13471), .ZN(
        n13473) );
  INV_X1 U16745 ( .A(n13473), .ZN(P2_U2876) );
  AND2_X1 U16746 ( .A1(n15035), .A2(n13474), .ZN(n13475) );
  OR2_X1 U16747 ( .A1(n13475), .A2(n13934), .ZN(n19001) );
  OAI211_X1 U16748 ( .C1(n13478), .C2(n11610), .A(n19127), .B(n13477), .ZN(
        n13480) );
  NAND2_X1 U16749 ( .A1(n12991), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13479) );
  OAI211_X1 U16750 ( .C1(n19001), .C2(n12991), .A(n13480), .B(n13479), .ZN(
        P2_U2874) );
  INV_X1 U16751 ( .A(n13481), .ZN(n20093) );
  AOI22_X1 U16752 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n9645), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n13482) );
  OAI21_X1 U16753 ( .B1(n15963), .B2(n20086), .A(n13482), .ZN(n13483) );
  AOI21_X1 U16754 ( .B1(n20093), .B2(n15960), .A(n13483), .ZN(n13484) );
  OAI21_X1 U16755 ( .B1(n20007), .B2(n13485), .A(n13484), .ZN(P1_U2995) );
  XNOR2_X1 U16756 ( .A(n13487), .B(n13486), .ZN(n20165) );
  INV_X1 U16757 ( .A(n13774), .ZN(n13490) );
  AND2_X1 U16758 ( .A1(n9645), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20170) );
  AOI21_X1 U16759 ( .B1(n15948), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n20170), .ZN(n13488) );
  OAI21_X1 U16760 ( .B1(n15963), .B2(n13769), .A(n13488), .ZN(n13489) );
  AOI21_X1 U16761 ( .B1(n13490), .B2(n15960), .A(n13489), .ZN(n13491) );
  OAI21_X1 U16762 ( .B1(n20007), .B2(n20165), .A(n13491), .ZN(P1_U2997) );
  XNOR2_X1 U16763 ( .A(n13492), .B(n13493), .ZN(n13553) );
  INV_X1 U16764 ( .A(n13494), .ZN(n13495) );
  AOI21_X1 U16765 ( .B1(n13497), .B2(n13496), .A(n13495), .ZN(n20070) );
  AND2_X1 U16766 ( .A1(n9645), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n13550) );
  AOI21_X1 U16767 ( .B1(n15948), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13550), .ZN(n13498) );
  OAI21_X1 U16768 ( .B1(n15963), .B2(n20068), .A(n13498), .ZN(n13499) );
  AOI21_X1 U16769 ( .B1(n20070), .B2(n15960), .A(n13499), .ZN(n13500) );
  OAI21_X1 U16770 ( .B1(n20007), .B2(n13553), .A(n13500), .ZN(P1_U2994) );
  INV_X1 U16771 ( .A(n13794), .ZN(n13504) );
  AOI21_X1 U16772 ( .B1(n15948), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13501), .ZN(n13502) );
  OAI21_X1 U16773 ( .B1(n15963), .B2(n13789), .A(n13502), .ZN(n13503) );
  AOI21_X1 U16774 ( .B1(n13504), .B2(n15960), .A(n13503), .ZN(n13505) );
  OAI21_X1 U16775 ( .B1(n20007), .B2(n13506), .A(n13505), .ZN(P1_U2996) );
  NAND2_X1 U16776 ( .A1(n13507), .A2(n10610), .ZN(n20624) );
  AOI21_X1 U16777 ( .B1(n20233), .B2(n20724), .A(n20974), .ZN(n13511) );
  NOR2_X1 U16778 ( .A1(n13511), .A2(n20664), .ZN(n13514) );
  INV_X1 U16779 ( .A(n13095), .ZN(n13772) );
  OR2_X1 U16780 ( .A1(n20813), .A2(n13772), .ZN(n20293) );
  OR2_X1 U16781 ( .A1(n20293), .A2(n20625), .ZN(n13517) );
  INV_X1 U16782 ( .A(n13516), .ZN(n13512) );
  NOR2_X1 U16783 ( .A1(n13512), .A2(n20728), .ZN(n20552) );
  NOR2_X1 U16784 ( .A1(n20330), .A2(n20552), .ZN(n20491) );
  INV_X1 U16785 ( .A(n20491), .ZN(n20265) );
  AND2_X1 U16786 ( .A1(n20431), .A2(n20486), .ZN(n13515) );
  NOR3_X1 U16787 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20239) );
  INV_X1 U16788 ( .A(n20239), .ZN(n20236) );
  NOR2_X1 U16789 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20236), .ZN(
        n20226) );
  OAI22_X1 U16790 ( .A1(n13515), .A2(n20728), .B1(n20226), .B2(n13115), .ZN(
        n13513) );
  AOI211_X2 U16791 ( .C1(n13514), .C2(n13517), .A(n20265), .B(n13513), .ZN(
        n20227) );
  INV_X1 U16792 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13526) );
  INV_X1 U16793 ( .A(n13514), .ZN(n13518) );
  INV_X1 U16794 ( .A(n13515), .ZN(n20326) );
  NOR2_X1 U16795 ( .A1(n13516), .A2(n20728), .ZN(n20488) );
  INV_X1 U16796 ( .A(n20488), .ZN(n20433) );
  OAI22_X1 U16797 ( .A1(n13518), .A2(n13517), .B1(n20326), .B2(n20433), .ZN(
        n20229) );
  INV_X1 U16798 ( .A(n14559), .ZN(n13625) );
  INV_X1 U16799 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16425) );
  INV_X1 U16800 ( .A(DATAI_30_), .ZN(n20933) );
  INV_X1 U16801 ( .A(n20651), .ZN(n20714) );
  INV_X1 U16802 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16435) );
  INV_X1 U16803 ( .A(DATAI_22_), .ZN(n13520) );
  OAI22_X1 U16804 ( .A1(n16435), .A2(n20222), .B1(n13520), .B2(n20221), .ZN(
        n20709) );
  AOI22_X1 U16805 ( .A1(n20257), .A2(n9780), .B1(n20226), .B2(n20707), .ZN(
        n13523) );
  OAI21_X1 U16806 ( .B1(n20724), .B2(n20714), .A(n13523), .ZN(n13524) );
  AOI21_X1 U16807 ( .B1(n20229), .B2(n20708), .A(n13524), .ZN(n13525) );
  OAI21_X1 U16808 ( .B1(n20227), .B2(n13526), .A(n13525), .ZN(P1_U3039) );
  INV_X1 U16809 ( .A(n20070), .ZN(n13534) );
  INV_X1 U16810 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13533) );
  NAND2_X1 U16811 ( .A1(n14048), .A2(n13533), .ZN(n13529) );
  NAND2_X1 U16812 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13527) );
  OAI211_X1 U16813 ( .C1(n14068), .C2(P1_EBX_REG_5__SCAN_IN), .A(n13527), .B(
        n14066), .ZN(n13528) );
  NOR2_X1 U16814 ( .A1(n13531), .A2(n13530), .ZN(n13532) );
  OR2_X1 U16815 ( .A1(n16026), .A2(n13532), .ZN(n20063) );
  OAI222_X1 U16816 ( .A1(n13534), .A2(n14524), .B1(n13533), .B2(n20103), .C1(
        n20063), .C2(n14523), .ZN(P1_U2867) );
  OAI222_X1 U16817 ( .A1(n14605), .A2(n13534), .B1(n14603), .B2(n10634), .C1(
        n14602), .C2(n20214), .ZN(P1_U2899) );
  INV_X1 U16818 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13543) );
  INV_X1 U16819 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16428) );
  INV_X1 U16820 ( .A(DATAI_28_), .ZN(n13535) );
  OAI22_X2 U16821 ( .A1(n16428), .A2(n20222), .B1(n13535), .B2(n20221), .ZN(
        n20643) );
  INV_X1 U16822 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16438) );
  INV_X1 U16823 ( .A(DATAI_20_), .ZN(n20886) );
  OAI22_X1 U16824 ( .A1(n16438), .A2(n20222), .B1(n20886), .B2(n20221), .ZN(
        n20697) );
  INV_X1 U16825 ( .A(n20697), .ZN(n20646) );
  INV_X1 U16826 ( .A(n20226), .ZN(n13538) );
  INV_X1 U16827 ( .A(n20225), .ZN(n13537) );
  NAND2_X1 U16828 ( .A1(n13537), .A2(n13536), .ZN(n20248) );
  OAI22_X1 U16829 ( .A1(n20233), .A2(n20646), .B1(n13538), .B2(n20248), .ZN(
        n13539) );
  AOI21_X1 U16830 ( .B1(n20710), .B2(n20643), .A(n13539), .ZN(n13542) );
  NAND2_X1 U16831 ( .A1(n20229), .A2(n20695), .ZN(n13541) );
  OAI211_X1 U16832 ( .C1(n20227), .C2(n13543), .A(n13542), .B(n13541), .ZN(
        P1_U3037) );
  INV_X1 U16833 ( .A(n14271), .ZN(n13545) );
  OAI21_X1 U16834 ( .B1(n13544), .B2(n15039), .A(n13745), .ZN(n19016) );
  INV_X1 U16835 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19185) );
  OAI222_X1 U16836 ( .A1(n13822), .A2(n13545), .B1(n19016), .B2(n19179), .C1(
        n15130), .C2(n19185), .ZN(P2_U2906) );
  INV_X1 U16837 ( .A(n20063), .ZN(n13551) );
  INV_X1 U16838 ( .A(n15998), .ZN(n14935) );
  NOR2_X1 U16839 ( .A1(n13546), .A2(n14935), .ZN(n13548) );
  INV_X1 U16840 ( .A(n14939), .ZN(n14895) );
  NAND3_X1 U16841 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13853) );
  AOI21_X1 U16842 ( .B1(n14895), .B2(n13853), .A(n13547), .ZN(n13852) );
  INV_X1 U16843 ( .A(n13852), .ZN(n13711) );
  MUX2_X1 U16844 ( .A(n13548), .B(n13711), .S(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n13549) );
  AOI211_X1 U16845 ( .C1(n16032), .C2(n13551), .A(n13550), .B(n13549), .ZN(
        n13552) );
  OAI21_X1 U16846 ( .B1(n20164), .B2(n13553), .A(n13552), .ZN(P1_U3026) );
  OAI22_X1 U16847 ( .A1(n14772), .A2(n13588), .B1(n20073), .B2(n20824), .ZN(
        n13555) );
  NOR2_X1 U16848 ( .A1(n13590), .A2(n15934), .ZN(n13554) );
  AOI211_X1 U16849 ( .C1(n15950), .C2(n13588), .A(n13555), .B(n13554), .ZN(
        n13556) );
  OAI21_X1 U16850 ( .B1(n13557), .B2(n20007), .A(n13556), .ZN(P1_U2998) );
  INV_X1 U16851 ( .A(n15828), .ZN(n13558) );
  NOR2_X1 U16852 ( .A1(n13115), .A2(n13558), .ZN(n15827) );
  AND2_X1 U16853 ( .A1(n13559), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13560) );
  MUX2_X1 U16854 ( .A(n15827), .B(n13560), .S(n16039), .Z(n13561) );
  INV_X1 U16855 ( .A(n13561), .ZN(n13562) );
  NAND2_X1 U16856 ( .A1(n13562), .A2(n20073), .ZN(n13563) );
  OAI21_X1 U16857 ( .B1(n13565), .B2(n13564), .A(n15914), .ZN(n20092) );
  INV_X1 U16858 ( .A(n20092), .ZN(n13795) );
  INV_X1 U16859 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14474) );
  NAND2_X1 U16860 ( .A1(n20738), .A2(n20974), .ZN(n15819) );
  INV_X1 U16861 ( .A(n15819), .ZN(n13579) );
  NAND2_X1 U16862 ( .A1(n13580), .A2(n13579), .ZN(n13569) );
  OAI211_X1 U16863 ( .C1(n20192), .C2(n14474), .A(n13569), .B(n13581), .ZN(
        n13570) );
  INV_X1 U16864 ( .A(n13570), .ZN(n13571) );
  INV_X1 U16865 ( .A(n13572), .ZN(n13573) );
  AND2_X1 U16866 ( .A1(n13583), .A2(n13573), .ZN(n20091) );
  INV_X1 U16867 ( .A(n20091), .ZN(n13574) );
  OAI22_X1 U16868 ( .A1(n13575), .A2(n20038), .B1(n13574), .B2(n9637), .ZN(
        n13587) );
  NAND2_X1 U16869 ( .A1(n15819), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13576) );
  NOR2_X1 U16870 ( .A1(n14068), .A2(n13576), .ZN(n13577) );
  AND2_X2 U16871 ( .A1(n13796), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20051) );
  AOI22_X1 U16872 ( .A1(n20053), .A2(n13578), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20051), .ZN(n13585) );
  AND3_X1 U16873 ( .A1(n13581), .A2(n13580), .A3(n13579), .ZN(n13582) );
  NAND2_X1 U16874 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n13796), .ZN(n13763) );
  OAI21_X1 U16875 ( .B1(n20042), .B2(P1_REIP_REG_1__SCAN_IN), .A(n13763), .ZN(
        n13584) );
  NAND2_X1 U16876 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  AOI211_X1 U16877 ( .C1(n20049), .C2(n13588), .A(n13587), .B(n13586), .ZN(
        n13589) );
  OAI21_X1 U16878 ( .B1(n13795), .B2(n13590), .A(n13589), .ZN(P1_U2839) );
  AOI21_X1 U16879 ( .B1(n13591), .B2(n13494), .A(n13915), .ZN(n20056) );
  INV_X1 U16880 ( .A(n20056), .ZN(n13626) );
  OAI21_X1 U16881 ( .B1(n10265), .B2(n13592), .A(n14066), .ZN(n13593) );
  OAI21_X1 U16882 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n14068), .A(n13593), .ZN(
        n13596) );
  INV_X1 U16883 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13594) );
  NAND2_X1 U16884 ( .A1(n10265), .A2(n13594), .ZN(n13595) );
  XNOR2_X1 U16885 ( .A(n16026), .B(n16024), .ZN(n20052) );
  AOI22_X1 U16886 ( .A1(n20098), .A2(n20052), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14485), .ZN(n13597) );
  OAI21_X1 U16887 ( .B1(n13626), .B2(n14524), .A(n13597), .ZN(P1_U2866) );
  INV_X1 U16888 ( .A(n14108), .ZN(n13600) );
  OR2_X1 U16889 ( .A1(n9696), .A2(n13598), .ZN(n13599) );
  NAND2_X1 U16890 ( .A1(n13600), .A2(n13599), .ZN(n14107) );
  NAND2_X1 U16891 ( .A1(n9634), .A2(n13602), .ZN(n13603) );
  XNOR2_X1 U16892 ( .A(n16220), .B(n13603), .ZN(n13604) );
  INV_X1 U16893 ( .A(n19851), .ZN(n19089) );
  NAND2_X1 U16894 ( .A1(n13604), .A2(n19089), .ZN(n13614) );
  AOI21_X1 U16895 ( .B1(n13606), .B2(n13605), .A(n15557), .ZN(n16275) );
  INV_X1 U16896 ( .A(n16275), .ZN(n19168) );
  AOI22_X1 U16897 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19095), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19096), .ZN(n13607) );
  OAI211_X1 U16898 ( .C1(n19168), .C2(n19098), .A(n13607), .B(n19066), .ZN(
        n13612) );
  OR2_X1 U16899 ( .A1(n13608), .A2(n13041), .ZN(n13610) );
  NAND2_X1 U16900 ( .A1(n13610), .A2(n13609), .ZN(n19144) );
  NOR2_X1 U16901 ( .A1(n19144), .A2(n19107), .ZN(n13611) );
  AOI211_X1 U16902 ( .C1(n19102), .C2(P2_REIP_REG_8__SCAN_IN), .A(n13612), .B(
        n13611), .ZN(n13613) );
  OAI211_X1 U16903 ( .C1(n14107), .C2(n19099), .A(n13614), .B(n13613), .ZN(
        P2_U2847) );
  NAND2_X1 U16904 ( .A1(n9634), .A2(n13803), .ZN(n13615) );
  XNOR2_X1 U16905 ( .A(n13616), .B(n13615), .ZN(n13617) );
  NAND2_X1 U16906 ( .A1(n13617), .A2(n19089), .ZN(n13624) );
  OAI22_X1 U16907 ( .A1(n19082), .A2(n12636), .B1(n19872), .B2(n19067), .ZN(
        n13618) );
  AOI21_X1 U16908 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19095), .A(
        n13618), .ZN(n13619) );
  OAI21_X1 U16909 ( .B1(n19099), .B2(n13620), .A(n13619), .ZN(n13622) );
  NOR2_X1 U16910 ( .A1(n19943), .A2(n19098), .ZN(n13621) );
  AOI211_X1 U16911 ( .C1(n19076), .C2(n12843), .A(n13622), .B(n13621), .ZN(
        n13623) );
  OAI211_X1 U16912 ( .C1(n19108), .C2(n19412), .A(n13624), .B(n13623), .ZN(
        P2_U2853) );
  OAI222_X1 U16913 ( .A1(n14605), .A2(n13626), .B1(n14603), .B2(n10645), .C1(
        n14602), .C2(n13625), .ZN(P1_U2898) );
  NAND2_X1 U16914 ( .A1(n13627), .A2(n13932), .ZN(n13630) );
  INV_X1 U16915 ( .A(n13628), .ZN(n13629) );
  INV_X1 U16916 ( .A(n18990), .ZN(n15502) );
  OAI21_X1 U16917 ( .B1(n13477), .B2(n13632), .A(n13631), .ZN(n13633) );
  NAND3_X1 U16918 ( .A1(n9734), .A2(n19127), .A3(n13633), .ZN(n13635) );
  NAND2_X1 U16919 ( .A1(n12991), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n13634) );
  OAI211_X1 U16920 ( .C1(n15502), .C2(n12991), .A(n13635), .B(n13634), .ZN(
        P2_U2872) );
  INV_X1 U16921 ( .A(n13676), .ZN(n13642) );
  INV_X1 U16922 ( .A(n13638), .ZN(n13639) );
  NAND2_X1 U16923 ( .A1(n13640), .A2(n13639), .ZN(n13641) );
  NAND2_X1 U16924 ( .A1(n13642), .A2(n13641), .ZN(n19100) );
  XNOR2_X1 U16925 ( .A(n19100), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19222) );
  INV_X1 U16926 ( .A(n19100), .ZN(n13643) );
  NAND2_X1 U16927 ( .A1(n13643), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13644) );
  INV_X1 U16928 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13646) );
  INV_X1 U16929 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13645) );
  OAI22_X1 U16930 ( .A1(n13646), .A2(n19785), .B1(n19380), .B2(n13645), .ZN(
        n13647) );
  INV_X1 U16931 ( .A(n13647), .ZN(n13653) );
  AOI22_X1 U16932 ( .A1(n19704), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13648), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13652) );
  INV_X1 U16933 ( .A(n13881), .ZN(n19318) );
  AOI22_X1 U16934 ( .A1(n19318), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n19606), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13651) );
  AOI22_X1 U16935 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n13649), .B1(
        n19576), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13650) );
  NAND4_X1 U16936 ( .A1(n13653), .A2(n13652), .A3(n13651), .A4(n13650), .ZN(
        n13671) );
  INV_X1 U16937 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13656) );
  INV_X1 U16938 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13655) );
  INV_X1 U16939 ( .A(n13657), .ZN(n13669) );
  INV_X1 U16940 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13659) );
  OAI22_X1 U16941 ( .A1(n13658), .A2(n12084), .B1(n19411), .B2(n13659), .ZN(
        n13660) );
  INV_X1 U16942 ( .A(n13660), .ZN(n13668) );
  INV_X1 U16943 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13662) );
  INV_X1 U16944 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13661) );
  OAI22_X1 U16945 ( .A1(n19677), .A2(n13662), .B1(n19440), .B2(n13661), .ZN(
        n13663) );
  INV_X1 U16946 ( .A(n13663), .ZN(n13667) );
  INV_X1 U16947 ( .A(n19504), .ZN(n13665) );
  INV_X1 U16948 ( .A(n19469), .ZN(n13664) );
  AOI22_X1 U16949 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n13665), .B1(
        n13664), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13666) );
  NAND4_X1 U16950 ( .A1(n13669), .A2(n13668), .A3(n13667), .A4(n13666), .ZN(
        n13670) );
  NAND2_X1 U16951 ( .A1(n13672), .A2(n19282), .ZN(n13673) );
  OAI21_X1 U16952 ( .B1(n13676), .B2(n13675), .A(n13903), .ZN(n19081) );
  INV_X1 U16953 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13682) );
  XNOR2_X1 U16954 ( .A(n13898), .B(n13682), .ZN(n13896) );
  XNOR2_X1 U16955 ( .A(n13897), .B(n13896), .ZN(n13705) );
  INV_X1 U16956 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19234) );
  INV_X1 U16957 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16300) );
  NOR2_X1 U16958 ( .A1(n13677), .A2(n16300), .ZN(n13680) );
  INV_X1 U16959 ( .A(n13681), .ZN(n13683) );
  NAND2_X1 U16960 ( .A1(n13683), .A2(n13682), .ZN(n13891) );
  NAND2_X1 U16961 ( .A1(n13681), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13895) );
  NAND2_X1 U16962 ( .A1(n13891), .A2(n13895), .ZN(n13684) );
  XNOR2_X1 U16963 ( .A(n13892), .B(n13684), .ZN(n13699) );
  NAND2_X1 U16964 ( .A1(n13699), .A2(n19250), .ZN(n13698) );
  NAND2_X1 U16965 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19246) );
  NAND2_X1 U16966 ( .A1(n19265), .A2(n19246), .ZN(n13690) );
  INV_X1 U16967 ( .A(n13690), .ZN(n13685) );
  AND2_X1 U16968 ( .A1(n19245), .A2(n13685), .ZN(n19247) );
  INV_X1 U16969 ( .A(n19246), .ZN(n19252) );
  INV_X1 U16970 ( .A(n19253), .ZN(n13686) );
  AOI21_X1 U16971 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19252), .A(
        n13686), .ZN(n13687) );
  NOR3_X1 U16972 ( .A1(n19244), .A2(n19247), .A3(n13687), .ZN(n16299) );
  OAI21_X1 U16973 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15787), .A(
        n16299), .ZN(n19237) );
  NOR2_X1 U16974 ( .A1(n16277), .A2(n19087), .ZN(n13696) );
  XNOR2_X1 U16975 ( .A(n13689), .B(n13688), .ZN(n19178) );
  NOR2_X1 U16976 ( .A1(n19265), .A2(n19246), .ZN(n13691) );
  OAI211_X1 U16977 ( .C1(n19245), .C2(n13691), .A(n13690), .B(n15579), .ZN(
        n16301) );
  NOR2_X1 U16978 ( .A1(n16300), .A2(n16301), .ZN(n19235) );
  OAI221_X1 U16979 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n13682), .C2(n19234), .A(
        n19235), .ZN(n13694) );
  NOR2_X1 U16980 ( .A1(n19066), .A2(n13692), .ZN(n13701) );
  INV_X1 U16981 ( .A(n13701), .ZN(n13693) );
  OAI211_X1 U16982 ( .C1(n16290), .C2(n19178), .A(n13694), .B(n13693), .ZN(
        n13695) );
  AOI211_X1 U16983 ( .C1(n19237), .C2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13696), .B(n13695), .ZN(n13697) );
  OAI211_X1 U16984 ( .C1(n13705), .C2(n16273), .A(n13698), .B(n13697), .ZN(
        P2_U3041) );
  NAND2_X1 U16985 ( .A1(n13699), .A2(n19227), .ZN(n13704) );
  INV_X1 U16986 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19094) );
  OAI22_X1 U16987 ( .A1(n19231), .A2(n19094), .B1(n16236), .B2(n19086), .ZN(
        n13700) );
  AOI211_X1 U16988 ( .C1(n16239), .C2(n13702), .A(n13701), .B(n13700), .ZN(
        n13703) );
  OAI211_X1 U16989 ( .C1(n13705), .C2(n19224), .A(n13704), .B(n13703), .ZN(
        P2_U3009) );
  XNOR2_X1 U16990 ( .A(n13706), .B(n13707), .ZN(n13716) );
  AOI22_X1 U16991 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n9645), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n13708) );
  OAI21_X1 U16992 ( .B1(n15963), .B2(n20047), .A(n13708), .ZN(n13709) );
  AOI21_X1 U16993 ( .B1(n20056), .B2(n15960), .A(n13709), .ZN(n13710) );
  OAI21_X1 U16994 ( .B1(n20007), .B2(n13716), .A(n13710), .ZN(P1_U2993) );
  INV_X1 U16995 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20754) );
  NOR2_X1 U16996 ( .A1(n20073), .A2(n20754), .ZN(n13714) );
  NOR2_X1 U16997 ( .A1(n13853), .A2(n14935), .ZN(n13712) );
  MUX2_X1 U16998 ( .A(n13712), .B(n13711), .S(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n13713) );
  AOI211_X1 U16999 ( .C1(n16032), .C2(n20052), .A(n13714), .B(n13713), .ZN(
        n13715) );
  OAI21_X1 U17000 ( .B1(n20164), .B2(n13716), .A(n13715), .ZN(P1_U3025) );
  NAND2_X1 U17001 ( .A1(n20087), .A2(n20075), .ZN(n13721) );
  AOI22_X1 U17002 ( .A1(n9664), .A2(n20091), .B1(n20077), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13718) );
  INV_X1 U17003 ( .A(n13796), .ZN(n20041) );
  NAND2_X1 U17004 ( .A1(n15910), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13717) );
  OAI211_X1 U17005 ( .C1(n20084), .C2(n13719), .A(n13718), .B(n13717), .ZN(
        n13720) );
  AOI21_X1 U17006 ( .B1(n13721), .B2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n13720), .ZN(n13722) );
  OAI21_X1 U17007 ( .B1(n13795), .B2(n13723), .A(n13722), .ZN(P1_U2840) );
  NOR2_X1 U17008 ( .A1(n19021), .A2(n13724), .ZN(n13726) );
  XNOR2_X1 U17009 ( .A(n13726), .B(n13725), .ZN(n13735) );
  NOR2_X1 U17010 ( .A1(n19566), .A2(n19108), .ZN(n13734) );
  OAI22_X1 U17011 ( .A1(n13728), .A2(n19099), .B1(n19093), .B2(n13727), .ZN(
        n13731) );
  OAI22_X1 U17012 ( .A1(n19082), .A2(n13729), .B1(n13432), .B2(n19067), .ZN(
        n13730) );
  AOI211_X1 U17013 ( .C1(n16288), .C2(n19076), .A(n13731), .B(n13730), .ZN(
        n13732) );
  OAI21_X1 U17014 ( .B1(n16291), .B2(n19098), .A(n13732), .ZN(n13733) );
  AOI211_X1 U17015 ( .C1(n13735), .C2(n19089), .A(n13734), .B(n13733), .ZN(
        n13736) );
  INV_X1 U17016 ( .A(n13736), .ZN(P2_U2852) );
  AOI21_X1 U17017 ( .B1(n13915), .B2(n13738), .A(n13739), .ZN(n13740) );
  OR2_X1 U17018 ( .A1(n13737), .A2(n13740), .ZN(n20028) );
  INV_X1 U17019 ( .A(n14602), .ZN(n13919) );
  INV_X1 U17020 ( .A(DATAI_8_), .ZN(n13742) );
  NAND2_X1 U17021 ( .A1(n14535), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13741) );
  OAI21_X1 U17022 ( .B1(n14535), .B2(n13742), .A(n13741), .ZN(n20134) );
  AOI22_X1 U17023 ( .A1(n13919), .A2(n20134), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14569), .ZN(n13743) );
  OAI21_X1 U17024 ( .B1(n20028), .B2(n14605), .A(n13743), .ZN(P1_U2896) );
  INV_X1 U17025 ( .A(n13744), .ZN(n13750) );
  INV_X1 U17026 ( .A(n13745), .ZN(n13746) );
  OR2_X1 U17027 ( .A1(n13747), .A2(n13746), .ZN(n13749) );
  INV_X1 U17028 ( .A(n13819), .ZN(n13748) );
  NAND2_X1 U17029 ( .A1(n13749), .A2(n13748), .ZN(n16252) );
  INV_X1 U17030 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19183) );
  OAI222_X1 U17031 ( .A1(n13822), .A2(n13750), .B1(n16252), .B2(n19179), .C1(
        n15130), .C2(n19183), .ZN(P2_U2905) );
  INV_X1 U17032 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13761) );
  INV_X1 U17033 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20102) );
  NAND2_X1 U17034 ( .A1(n14048), .A2(n20102), .ZN(n13753) );
  NAND2_X1 U17035 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13751) );
  OAI211_X1 U17036 ( .C1(n14068), .C2(P1_EBX_REG_7__SCAN_IN), .A(n13751), .B(
        n14066), .ZN(n13752) );
  NAND2_X1 U17037 ( .A1(n13753), .A2(n13752), .ZN(n16030) );
  NOR2_X1 U17038 ( .A1(n16030), .A2(n16024), .ZN(n13754) );
  OAI21_X1 U17039 ( .B1(n10265), .B2(n13755), .A(n14066), .ZN(n13756) );
  OAI21_X1 U17040 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n14068), .A(n13756), .ZN(
        n13758) );
  NAND2_X1 U17041 ( .A1(n10265), .A2(n13761), .ZN(n13757) );
  AND2_X1 U17042 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  NAND2_X1 U17043 ( .A1(n16027), .A2(n13759), .ZN(n13760) );
  NAND2_X1 U17044 ( .A1(n13782), .A2(n13760), .ZN(n20026) );
  OAI222_X1 U17045 ( .A1(n20028), .A2(n14524), .B1(n13761), .B2(n20103), .C1(
        n20026), .C2(n14523), .ZN(P1_U2864) );
  INV_X1 U17046 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13764) );
  NAND2_X1 U17047 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13762) );
  OAI21_X1 U17048 ( .B1(n20041), .B2(n13762), .A(n15910), .ZN(n13788) );
  AOI21_X1 U17049 ( .B1(n13764), .B2(n13763), .A(n13788), .ZN(n13767) );
  NOR2_X1 U17050 ( .A1(n20038), .A2(n13765), .ZN(n13766) );
  AOI211_X1 U17051 ( .C1(n20051), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13767), .B(n13766), .ZN(n13768) );
  OAI21_X1 U17052 ( .B1(n20084), .B2(n20172), .A(n13768), .ZN(n13771) );
  NOR2_X1 U17053 ( .A1(n20087), .A2(n13769), .ZN(n13770) );
  AOI211_X1 U17054 ( .C1(n20091), .C2(n13772), .A(n13771), .B(n13770), .ZN(
        n13773) );
  OAI21_X1 U17055 ( .B1(n13795), .B2(n13774), .A(n13773), .ZN(P1_U2838) );
  OAI21_X1 U17056 ( .B1(n13737), .B2(n13776), .A(n13775), .ZN(n13979) );
  INV_X1 U17057 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13777) );
  NAND2_X1 U17058 ( .A1(n14048), .A2(n13777), .ZN(n13780) );
  NAND2_X1 U17059 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13778) );
  OAI211_X1 U17060 ( .C1(n14068), .C2(P1_EBX_REG_9__SCAN_IN), .A(n13778), .B(
        n14066), .ZN(n13779) );
  NAND2_X1 U17061 ( .A1(n13780), .A2(n13779), .ZN(n13781) );
  AND2_X1 U17062 ( .A1(n13782), .A2(n13781), .ZN(n13783) );
  AOI22_X1 U17063 ( .A1(n9757), .A2(n20098), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14485), .ZN(n13784) );
  OAI21_X1 U17064 ( .B1(n13979), .B2(n14524), .A(n13784), .ZN(P1_U2863) );
  INV_X1 U17065 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20750) );
  AOI22_X1 U17066 ( .A1(n20077), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20051), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13787) );
  NAND2_X1 U17067 ( .A1(n20053), .A2(n13785), .ZN(n13786) );
  OAI211_X1 U17068 ( .C1(n13788), .C2(n20750), .A(n13787), .B(n13786), .ZN(
        n13791) );
  NOR2_X1 U17069 ( .A1(n20087), .A2(n13789), .ZN(n13790) );
  AOI211_X1 U17070 ( .C1(n20091), .C2(n20813), .A(n13791), .B(n13790), .ZN(
        n13793) );
  NAND4_X1 U17071 ( .A1(n20042), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .A4(n20750), .ZN(n13792) );
  OAI211_X1 U17072 ( .C1(n13795), .C2(n13794), .A(n13793), .B(n13792), .ZN(
        P1_U2837) );
  INV_X1 U17073 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20756) );
  NAND4_X1 U17074 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20078)
         );
  NAND3_X1 U17075 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n20024) );
  NOR3_X1 U17076 ( .A1(n20756), .A2(n20078), .A3(n20024), .ZN(n13797) );
  NOR2_X1 U17077 ( .A1(n13999), .A2(n14439), .ZN(n20029) );
  NAND2_X1 U17078 ( .A1(n20042), .A2(n13797), .ZN(n13998) );
  AOI22_X1 U17079 ( .A1(n20077), .A2(P1_EBX_REG_9__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20051), .ZN(n13798) );
  OAI211_X1 U17080 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n13998), .A(n13798), .B(
        n20073), .ZN(n13799) );
  AOI21_X1 U17081 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20029), .A(n13799), .ZN(
        n13802) );
  INV_X1 U17082 ( .A(n13975), .ZN(n13800) );
  AOI22_X1 U17083 ( .A1(n20049), .A2(n13800), .B1(n9757), .B2(n20053), .ZN(
        n13801) );
  OAI211_X1 U17084 ( .C1(n13979), .C2(n15914), .A(n13802), .B(n13801), .ZN(
        P1_U2831) );
  OAI211_X1 U17085 ( .C1(n13807), .C2(n13804), .A(n9634), .B(n13803), .ZN(
        n13823) );
  OAI21_X1 U17086 ( .B1(n9634), .B2(n13805), .A(n13823), .ZN(n13806) );
  INV_X1 U17087 ( .A(n13806), .ZN(n15609) );
  INV_X1 U17088 ( .A(n13807), .ZN(n13942) );
  AOI22_X1 U17089 ( .A1(n19021), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n13942), .B2(n9634), .ZN(n15591) );
  NOR2_X1 U17090 ( .A1(n15591), .A2(n15593), .ZN(n15596) );
  INV_X1 U17091 ( .A(n13808), .ZN(n15607) );
  NAND2_X1 U17092 ( .A1(n12867), .A2(n15607), .ZN(n13815) );
  NAND2_X1 U17093 ( .A1(n13810), .A2(n13809), .ZN(n15588) );
  NOR2_X1 U17094 ( .A1(n13811), .A2(n13134), .ZN(n13813) );
  AOI22_X1 U17095 ( .A1(n15588), .A2(n13813), .B1(n15587), .B2(n13812), .ZN(
        n13814) );
  NAND2_X1 U17096 ( .A1(n13815), .A2(n13814), .ZN(n16304) );
  AOI222_X1 U17097 ( .A1(n15609), .A2(n15596), .B1(n16350), .B2(n19953), .C1(
        n16304), .C2(n19933), .ZN(n13818) );
  NAND2_X1 U17098 ( .A1(n13817), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13816) );
  OAI21_X1 U17099 ( .B1(n13818), .B2(n13817), .A(n13816), .ZN(P2_U3600) );
  OAI21_X1 U17100 ( .B1(n13820), .B2(n13819), .A(n13963), .ZN(n19000) );
  OAI222_X1 U17101 ( .A1(n19000), .A2(n19179), .B1(n13822), .B2(n13821), .C1(
        n15130), .C2(n12732), .ZN(P2_U2904) );
  INV_X1 U17102 ( .A(n19009), .ZN(n13824) );
  OAI22_X1 U17103 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n13824), .B1(
        n13823), .B2(n19851), .ZN(n13825) );
  INV_X1 U17104 ( .A(n13825), .ZN(n13835) );
  INV_X1 U17105 ( .A(n19099), .ZN(n19056) );
  INV_X1 U17106 ( .A(n13826), .ZN(n13829) );
  OAI22_X1 U17107 ( .A1(n13827), .A2(n19093), .B1(n19870), .B2(n19067), .ZN(
        n13828) );
  AOI21_X1 U17108 ( .B1(n19056), .B2(n13829), .A(n13828), .ZN(n13831) );
  NAND2_X1 U17109 ( .A1(n18973), .A2(n19957), .ZN(n13830) );
  OAI211_X1 U17110 ( .C1(n19082), .C2(n13832), .A(n13831), .B(n13830), .ZN(
        n13833) );
  AOI21_X1 U17111 ( .B1(n12867), .B2(n19076), .A(n13833), .ZN(n13834) );
  OAI211_X1 U17112 ( .C1(n19108), .C2(n19275), .A(n13835), .B(n13834), .ZN(
        P2_U2854) );
  INV_X1 U17113 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13836) );
  INV_X1 U17114 ( .A(DATAI_9_), .ZN(n20873) );
  MUX2_X1 U17115 ( .A(n20873), .B(n16455), .S(n14535), .Z(n20136) );
  OAI222_X1 U17116 ( .A1(n13979), .A2(n14605), .B1(n13836), .B2(n14603), .C1(
        n14602), .C2(n20136), .ZN(P1_U2895) );
  OAI21_X1 U17117 ( .B1(n13837), .B2(n13839), .A(n13838), .ZN(n13960) );
  INV_X1 U17118 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n13840) );
  OR2_X1 U17119 ( .A1(n19148), .A2(n13840), .ZN(n13844) );
  OR2_X1 U17120 ( .A1(n15764), .A2(n13841), .ZN(n13842) );
  AND2_X1 U17121 ( .A1(n13842), .A2(n15484), .ZN(n18974) );
  NAND2_X1 U17122 ( .A1(n19148), .A2(n18974), .ZN(n13843) );
  OAI211_X1 U17123 ( .C1(n13960), .C2(n19145), .A(n13844), .B(n13843), .ZN(
        P2_U2870) );
  XNOR2_X1 U17124 ( .A(n13845), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13846) );
  XNOR2_X1 U17125 ( .A(n13847), .B(n13846), .ZN(n13858) );
  AOI22_X1 U17126 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n9645), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13849) );
  NAND2_X1 U17127 ( .A1(n15950), .A2(n20023), .ZN(n13848) );
  OAI211_X1 U17128 ( .C1(n20028), .C2(n15934), .A(n13849), .B(n13848), .ZN(
        n13850) );
  INV_X1 U17129 ( .A(n13850), .ZN(n13851) );
  OAI21_X1 U17130 ( .B1(n13858), .B2(n20007), .A(n13851), .ZN(P1_U2991) );
  OAI21_X1 U17131 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14939), .A(
        n13852), .ZN(n16035) );
  OAI22_X1 U17132 ( .A1(n20173), .A2(n20026), .B1(n20756), .B2(n20073), .ZN(
        n13856) );
  NOR2_X1 U17133 ( .A1(n13592), .A2(n13853), .ZN(n14011) );
  NAND2_X1 U17134 ( .A1(n14011), .A2(n15998), .ZN(n16038) );
  AOI221_X1 U17135 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n13755), .C2(n13854), .A(
        n16038), .ZN(n13855) );
  AOI211_X1 U17136 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n16035), .A(
        n13856), .B(n13855), .ZN(n13857) );
  OAI21_X1 U17137 ( .B1(n20164), .B2(n13858), .A(n13857), .ZN(P1_U3023) );
  INV_X1 U17138 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13860) );
  INV_X1 U17139 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13859) );
  OAI22_X1 U17140 ( .A1(n13860), .A2(n19677), .B1(n13658), .B2(n13859), .ZN(
        n13864) );
  INV_X1 U17141 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13862) );
  INV_X1 U17142 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13861) );
  OAI22_X1 U17143 ( .A1(n19640), .A2(n13862), .B1(n19411), .B2(n13861), .ZN(
        n13863) );
  NOR2_X1 U17144 ( .A1(n13864), .A2(n13863), .ZN(n13887) );
  INV_X1 U17145 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13867) );
  INV_X1 U17146 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13865) );
  OAI22_X1 U17147 ( .A1(n13867), .A2(n13866), .B1(n19380), .B2(n13865), .ZN(
        n13871) );
  INV_X1 U17148 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13869) );
  INV_X1 U17149 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13868) );
  OAI22_X1 U17150 ( .A1(n19785), .A2(n13869), .B1(n19440), .B2(n13868), .ZN(
        n13870) );
  NOR2_X1 U17151 ( .A1(n13871), .A2(n13870), .ZN(n13886) );
  INV_X1 U17152 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13873) );
  INV_X1 U17153 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13872) );
  INV_X1 U17154 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13874) );
  NOR2_X1 U17155 ( .A1(n13876), .A2(n13875), .ZN(n13885) );
  INV_X1 U17156 ( .A(n19606), .ZN(n19611) );
  INV_X1 U17157 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13878) );
  NAND2_X1 U17158 ( .A1(n19576), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13877) );
  OAI21_X1 U17159 ( .B1(n19611), .B2(n13878), .A(n13877), .ZN(n13883) );
  INV_X1 U17160 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13880) );
  INV_X1 U17161 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13879) );
  OAI22_X1 U17162 ( .A1(n13881), .A2(n13880), .B1(n19504), .B2(n13879), .ZN(
        n13882) );
  NOR2_X1 U17163 ( .A1(n13883), .A2(n13882), .ZN(n13884) );
  NAND4_X1 U17164 ( .A1(n13887), .A2(n13886), .A3(n13885), .A4(n13884), .ZN(
        n13890) );
  NAND2_X1 U17165 ( .A1(n13888), .A2(n19282), .ZN(n13889) );
  XNOR2_X2 U17166 ( .A(n14249), .B(n14247), .ZN(n13901) );
  XNOR2_X1 U17167 ( .A(n14250), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16250) );
  NAND2_X1 U17168 ( .A1(n13897), .A2(n13896), .ZN(n13900) );
  NAND2_X1 U17169 ( .A1(n13898), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13899) );
  NAND2_X1 U17170 ( .A1(n13901), .A2(n15158), .ZN(n13905) );
  NAND2_X1 U17171 ( .A1(n13903), .A2(n13902), .ZN(n13904) );
  NAND2_X1 U17172 ( .A1(n10159), .A2(n13904), .ZN(n19069) );
  NAND2_X1 U17173 ( .A1(n13905), .A2(n19069), .ZN(n14102) );
  INV_X1 U17174 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13909) );
  XNOR2_X1 U17175 ( .A(n14101), .B(n14100), .ZN(n16246) );
  NAND3_X1 U17176 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13906) );
  NOR2_X1 U17177 ( .A1(n16301), .A2(n13906), .ZN(n14238) );
  INV_X1 U17178 ( .A(n13906), .ZN(n13907) );
  OAI221_X1 U17179 ( .B1(n15787), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        n15787), .C2(n13907), .A(n16299), .ZN(n16276) );
  INV_X1 U17180 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19877) );
  NOR2_X1 U17181 ( .A1(n19877), .A2(n19066), .ZN(n13908) );
  AOI221_X1 U17182 ( .B1(n14238), .B2(n13909), .C1(n16276), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n13908), .ZN(n13912) );
  INV_X1 U17183 ( .A(n19080), .ZN(n13910) );
  AOI22_X1 U17184 ( .A1(n19262), .A2(n13910), .B1(n19248), .B2(n19075), .ZN(
        n13911) );
  OAI211_X1 U17185 ( .C1(n16246), .C2(n16273), .A(n13912), .B(n13911), .ZN(
        n13913) );
  INV_X1 U17186 ( .A(n13913), .ZN(n13914) );
  OAI21_X1 U17187 ( .B1(n16250), .B2(n16292), .A(n13914), .ZN(P2_U3040) );
  INV_X1 U17188 ( .A(n14555), .ZN(n20228) );
  XOR2_X1 U17189 ( .A(n13738), .B(n13915), .Z(n20100) );
  INV_X1 U17190 ( .A(n20100), .ZN(n13916) );
  INV_X1 U17191 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20117) );
  OAI222_X1 U17192 ( .A1(n14602), .A2(n20228), .B1(n14605), .B2(n13916), .C1(
        n20117), .C2(n14603), .ZN(P1_U2897) );
  AOI21_X1 U17193 ( .B1(n13917), .B2(n13775), .A(n9674), .ZN(n15951) );
  INV_X1 U17194 ( .A(n15951), .ZN(n13927) );
  INV_X1 U17195 ( .A(DATAI_10_), .ZN(n20995) );
  NAND2_X1 U17196 ( .A1(n14535), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13918) );
  OAI21_X1 U17197 ( .B1(n14535), .B2(n20995), .A(n13918), .ZN(n20139) );
  AOI22_X1 U17198 ( .A1(n13919), .A2(n20139), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14569), .ZN(n13920) );
  OAI21_X1 U17199 ( .B1(n13927), .B2(n14605), .A(n13920), .ZN(P1_U2894) );
  INV_X1 U17200 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15921) );
  OAI21_X1 U17201 ( .B1(n10265), .B2(n14930), .A(n14066), .ZN(n13921) );
  OAI21_X1 U17202 ( .B1(P1_EBX_REG_10__SCAN_IN), .B2(n14068), .A(n13921), .ZN(
        n13923) );
  NAND2_X1 U17203 ( .A1(n10265), .A2(n15921), .ZN(n13922) );
  NAND2_X1 U17204 ( .A1(n13923), .A2(n13922), .ZN(n13924) );
  NAND2_X1 U17205 ( .A1(n13925), .A2(n13924), .ZN(n13986) );
  OR2_X1 U17206 ( .A1(n13925), .A2(n13924), .ZN(n13926) );
  NAND2_X1 U17207 ( .A1(n13986), .A2(n13926), .ZN(n15922) );
  OAI222_X1 U17208 ( .A1(n13927), .A2(n14524), .B1(n15921), .B2(n20103), .C1(
        n15922), .C2(n14523), .ZN(P1_U2862) );
  NAND2_X1 U17209 ( .A1(n14206), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13928) );
  MUX2_X1 U17210 ( .A(n14206), .B(n13928), .S(n14142), .Z(n13929) );
  OR2_X1 U17211 ( .A1(n14142), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14175) );
  AND2_X1 U17212 ( .A1(n13929), .A2(n14175), .ZN(n14170) );
  INV_X1 U17213 ( .A(n14170), .ZN(n13941) );
  NAND2_X1 U17214 ( .A1(n9634), .A2(n13930), .ZN(n19010) );
  XOR2_X1 U17215 ( .A(n16186), .B(n19010), .Z(n13931) );
  NAND2_X1 U17216 ( .A1(n13931), .A2(n19089), .ZN(n13940) );
  OAI21_X1 U17217 ( .B1(n13934), .B2(n13933), .A(n13932), .ZN(n19124) );
  INV_X1 U17218 ( .A(n19124), .ZN(n16256) );
  NOR2_X1 U17219 ( .A1(n19098), .A2(n16252), .ZN(n13938) );
  AOI22_X1 U17220 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19095), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19096), .ZN(n13935) );
  OAI211_X1 U17221 ( .C1(n19067), .C2(n13936), .A(n13935), .B(n19066), .ZN(
        n13937) );
  AOI211_X1 U17222 ( .C1(n16256), .C2(n19076), .A(n13938), .B(n13937), .ZN(
        n13939) );
  OAI211_X1 U17223 ( .C1(n13941), .C2(n19099), .A(n13940), .B(n13939), .ZN(
        P2_U2841) );
  NOR2_X1 U17224 ( .A1(n19021), .A2(n19851), .ZN(n18995) );
  NAND2_X1 U17225 ( .A1(n18995), .A2(n13942), .ZN(n13951) );
  NAND2_X1 U17226 ( .A1(n19056), .A2(n13943), .ZN(n13945) );
  OAI21_X1 U17227 ( .B1(n19095), .B2(n19009), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13944) );
  OAI211_X1 U17228 ( .C1(n18922), .C2(n19067), .A(n13945), .B(n13944), .ZN(
        n13946) );
  AOI21_X1 U17229 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19096), .A(n13946), .ZN(
        n13947) );
  OAI21_X1 U17230 ( .B1(n19098), .B2(n13948), .A(n13947), .ZN(n13949) );
  AOI21_X1 U17231 ( .B1(n15590), .B2(n19076), .A(n13949), .ZN(n13950) );
  OAI211_X1 U17232 ( .C1(n19108), .C2(n19961), .A(n13951), .B(n13950), .ZN(
        P2_U2855) );
  OR2_X1 U17233 ( .A1(n13953), .A2(n13952), .ZN(n13954) );
  NAND2_X1 U17234 ( .A1(n13954), .A2(n15487), .ZN(n15784) );
  AOI22_X1 U17235 ( .A1(n19153), .A2(BUF1_REG_17__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U17236 ( .A1(n16127), .A2(n13955), .B1(n19169), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13956) );
  OAI211_X1 U17237 ( .C1(n16119), .C2(n15784), .A(n13957), .B(n13956), .ZN(
        n13958) );
  INV_X1 U17238 ( .A(n13958), .ZN(n13959) );
  OAI21_X1 U17239 ( .B1(n13960), .B2(n16120), .A(n13959), .ZN(P2_U2902) );
  INV_X1 U17240 ( .A(n13961), .ZN(n13962) );
  AOI21_X1 U17241 ( .B1(n13962), .B2(n9734), .A(n13837), .ZN(n19118) );
  INV_X1 U17242 ( .A(n19118), .ZN(n13970) );
  XNOR2_X1 U17243 ( .A(n13964), .B(n13963), .ZN(n18983) );
  INV_X1 U17244 ( .A(n18983), .ZN(n13967) );
  OAI22_X1 U17245 ( .A1(n19274), .A2(n15131), .B1(n15130), .B2(n13965), .ZN(
        n13966) );
  AOI21_X1 U17246 ( .B1(n19150), .B2(n13967), .A(n13966), .ZN(n13969) );
  AOI22_X1 U17247 ( .A1(n19153), .A2(BUF1_REG_16__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n13968) );
  OAI211_X1 U17248 ( .C1(n13970), .C2(n16120), .A(n13969), .B(n13968), .ZN(
        P2_U2903) );
  MUX2_X1 U17249 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n13971), .S(n9971), .Z(n13972) );
  XNOR2_X1 U17250 ( .A(n13973), .B(n13972), .ZN(n16020) );
  NAND2_X1 U17251 ( .A1(n16020), .A2(n15959), .ZN(n13978) );
  INV_X1 U17252 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13974) );
  NOR2_X1 U17253 ( .A1(n20073), .A2(n13974), .ZN(n16018) );
  NOR2_X1 U17254 ( .A1(n15963), .A2(n13975), .ZN(n13976) );
  AOI211_X1 U17255 ( .C1(n15948), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16018), .B(n13976), .ZN(n13977) );
  OAI211_X1 U17256 ( .C1(n15934), .C2(n13979), .A(n13978), .B(n13977), .ZN(
        P1_U2990) );
  OAI21_X1 U17257 ( .B1(n13982), .B2(n13981), .A(n13980), .ZN(n15915) );
  MUX2_X1 U17258 ( .A(n14057), .B(n14293), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13984) );
  NAND2_X1 U17259 ( .A1(n14058), .A2(n14919), .ZN(n13983) );
  NAND2_X1 U17260 ( .A1(n13984), .A2(n13983), .ZN(n13987) );
  OR2_X2 U17261 ( .A1(n13986), .A2(n13987), .ZN(n14520) );
  INV_X1 U17262 ( .A(n14520), .ZN(n13985) );
  AOI21_X1 U17263 ( .B1(n13987), .B2(n13986), .A(n13985), .ZN(n16011) );
  AOI22_X1 U17264 ( .A1(n16011), .A2(n20098), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14485), .ZN(n13988) );
  OAI21_X1 U17265 ( .B1(n15915), .B2(n14524), .A(n13988), .ZN(P1_U2861) );
  INV_X1 U17266 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20110) );
  OAI222_X1 U17267 ( .A1(n15915), .A2(n14605), .B1(n20110), .B2(n14603), .C1(
        n14602), .C2(n14541), .ZN(P1_U2893) );
  AND3_X1 U17268 ( .A1(n13980), .A2(n13991), .A3(n13990), .ZN(n13992) );
  OR2_X1 U17269 ( .A1(n13989), .A2(n13992), .ZN(n14764) );
  NAND2_X1 U17270 ( .A1(n14066), .A2(n13993), .ZN(n13994) );
  OAI211_X1 U17271 ( .C1(n14068), .C2(P1_EBX_REG_12__SCAN_IN), .A(n13994), .B(
        n14293), .ZN(n13996) );
  INV_X1 U17272 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U17273 ( .A1(n10265), .A2(n14002), .ZN(n13995) );
  NAND2_X1 U17274 ( .A1(n13996), .A2(n13995), .ZN(n14517) );
  XNOR2_X1 U17275 ( .A(n14520), .B(n14517), .ZN(n14926) );
  AOI22_X1 U17276 ( .A1(n14926), .A2(n20098), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14485), .ZN(n13997) );
  OAI21_X1 U17277 ( .B1(n14764), .B2(n14524), .A(n13997), .ZN(P1_U2860) );
  INV_X1 U17278 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15920) );
  NOR2_X1 U17279 ( .A1(n13974), .A2(n13998), .ZN(n15925) );
  NAND2_X1 U17280 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n15925), .ZN(n15913) );
  NOR2_X1 U17281 ( .A1(n15920), .A2(n15913), .ZN(n14281) );
  INV_X1 U17282 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n14000) );
  NAND3_X1 U17283 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n13999), .ZN(n15909) );
  NOR3_X1 U17284 ( .A1(n14000), .A2(n15920), .A3(n15909), .ZN(n14276) );
  NOR2_X1 U17285 ( .A1(n14276), .A2(n14439), .ZN(n15904) );
  OAI21_X1 U17286 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n14281), .A(n15904), 
        .ZN(n14006) );
  AOI21_X1 U17287 ( .B1(n20051), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n9645), .ZN(n14001) );
  OAI21_X1 U17288 ( .B1(n20038), .B2(n14002), .A(n14001), .ZN(n14004) );
  NOR2_X1 U17289 ( .A1(n20087), .A2(n14766), .ZN(n14003) );
  AOI211_X1 U17290 ( .C1(n20053), .C2(n14926), .A(n14004), .B(n14003), .ZN(
        n14005) );
  OAI211_X1 U17291 ( .C1(n14764), .C2(n15914), .A(n14006), .B(n14005), .ZN(
        P1_U2828) );
  NAND3_X1 U17292 ( .A1(n17133), .A2(n15726), .A3(n18719), .ZN(n18225) );
  NOR2_X1 U17293 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18225), .ZN(n14007) );
  NAND3_X1 U17294 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18831)
         );
  OAI21_X1 U17295 ( .B1(n14007), .B2(n18831), .A(n18518), .ZN(n18231) );
  INV_X1 U17296 ( .A(n18231), .ZN(n14008) );
  INV_X1 U17297 ( .A(n17805), .ZN(n17862) );
  AOI22_X1 U17298 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n15708), .B2(n17862), .ZN(n15711) );
  NOR2_X1 U17299 ( .A1(n14008), .A2(n15711), .ZN(n14010) );
  INV_X1 U17300 ( .A(n18574), .ZN(n15712) );
  NOR2_X1 U17301 ( .A1(n18833), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18272) );
  INV_X1 U17302 ( .A(n18272), .ZN(n18313) );
  NAND2_X1 U17303 ( .A1(n18313), .A2(n18231), .ZN(n15709) );
  OR2_X1 U17304 ( .A1(n15712), .A2(n15709), .ZN(n14009) );
  MUX2_X1 U17305 ( .A(n14010), .B(n14009), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17306 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15966) );
  INV_X1 U17307 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14888) );
  NAND2_X1 U17308 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15984) );
  NOR2_X1 U17309 ( .A1(n14888), .A2(n15984), .ZN(n15978) );
  NAND2_X1 U17310 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15978), .ZN(
        n14075) );
  NAND3_X1 U17311 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n14011), .ZN(n14936) );
  NOR2_X1 U17312 ( .A1(n14930), .A2(n13971), .ZN(n14013) );
  INV_X1 U17313 ( .A(n14013), .ZN(n14937) );
  NOR2_X1 U17314 ( .A1(n14936), .A2(n14937), .ZN(n15999) );
  NAND3_X1 U17315 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n15999), .ZN(n14914) );
  NOR3_X1 U17316 ( .A1(n14919), .A2(n13993), .A3(n14914), .ZN(n14903) );
  NOR2_X1 U17317 ( .A1(n14012), .A2(n14936), .ZN(n14938) );
  NAND3_X1 U17318 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14013), .A3(
        n14938), .ZN(n14915) );
  NOR2_X1 U17319 ( .A1(n13993), .A2(n14915), .ZN(n14891) );
  AOI21_X1 U17320 ( .B1(n14903), .B2(n14838), .A(n14867), .ZN(n15972) );
  INV_X1 U17321 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16000) );
  INV_X1 U17322 ( .A(n15991), .ZN(n14889) );
  INV_X1 U17323 ( .A(n14862), .ZN(n14079) );
  NAND2_X1 U17324 ( .A1(n15836), .A2(n14079), .ZN(n14856) );
  NOR2_X1 U17325 ( .A1(n14856), .A2(n14082), .ZN(n14831) );
  AND2_X1 U17326 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14088) );
  AND2_X1 U17327 ( .A1(n14831), .A2(n14088), .ZN(n14806) );
  INV_X1 U17328 ( .A(n14058), .ZN(n14071) );
  AOI22_X1 U17329 ( .A1(n14071), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14068), .ZN(n14073) );
  AOI22_X1 U17330 ( .A1(n14071), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14068), .ZN(n14295) );
  MUX2_X1 U17331 ( .A(n14057), .B(n14293), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14015) );
  NAND2_X1 U17332 ( .A1(n14058), .A2(n14907), .ZN(n14014) );
  NAND2_X1 U17333 ( .A1(n14015), .A2(n14014), .ZN(n14518) );
  INV_X1 U17334 ( .A(n14518), .ZN(n14016) );
  NAND2_X1 U17335 ( .A1(n14016), .A2(n14517), .ZN(n14017) );
  NAND2_X1 U17336 ( .A1(n14066), .A2(n16000), .ZN(n14018) );
  OAI211_X1 U17337 ( .C1(n14068), .C2(P1_EBX_REG_14__SCAN_IN), .A(n14018), .B(
        n14293), .ZN(n14020) );
  INV_X1 U17338 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14514) );
  NAND2_X1 U17339 ( .A1(n10265), .A2(n14514), .ZN(n14019) );
  NOR2_X2 U17340 ( .A1(n14521), .A2(n14510), .ZN(n15881) );
  INV_X1 U17341 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15932) );
  NAND2_X1 U17342 ( .A1(n14048), .A2(n15932), .ZN(n14023) );
  NAND2_X1 U17343 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14021) );
  OAI211_X1 U17344 ( .C1(n14068), .C2(P1_EBX_REG_15__SCAN_IN), .A(n14021), .B(
        n14066), .ZN(n14022) );
  AND2_X2 U17345 ( .A1(n15881), .A2(n15880), .ZN(n15883) );
  INV_X1 U17346 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15987) );
  NAND2_X1 U17347 ( .A1(n14066), .A2(n15987), .ZN(n14024) );
  OAI211_X1 U17348 ( .C1(n14068), .C2(P1_EBX_REG_16__SCAN_IN), .A(n14024), .B(
        n14293), .ZN(n14026) );
  INV_X1 U17349 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14504) );
  NAND2_X1 U17350 ( .A1(n10265), .A2(n14504), .ZN(n14025) );
  NAND2_X1 U17351 ( .A1(n14026), .A2(n14025), .ZN(n14463) );
  MUX2_X1 U17352 ( .A(n14057), .B(n14293), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14028) );
  NAND2_X1 U17353 ( .A1(n14058), .A2(n14888), .ZN(n14027) );
  NAND2_X1 U17354 ( .A1(n14028), .A2(n14027), .ZN(n14499) );
  INV_X1 U17355 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15977) );
  NAND2_X1 U17356 ( .A1(n14066), .A2(n15977), .ZN(n14029) );
  OAI211_X1 U17357 ( .C1(n14068), .C2(P1_EBX_REG_18__SCAN_IN), .A(n14029), .B(
        n14293), .ZN(n14031) );
  INV_X1 U17358 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U17359 ( .A1(n10265), .A2(n14493), .ZN(n14030) );
  AND2_X1 U17360 ( .A1(n14031), .A2(n14030), .ZN(n14450) );
  INV_X1 U17361 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14490) );
  NAND2_X1 U17362 ( .A1(n14048), .A2(n14490), .ZN(n14034) );
  NAND2_X1 U17363 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14032) );
  OAI211_X1 U17364 ( .C1(n14068), .C2(P1_EBX_REG_19__SCAN_IN), .A(n14032), .B(
        n14066), .ZN(n14033) );
  OAI21_X1 U17365 ( .B1(n10265), .B2(n14697), .A(n14066), .ZN(n14035) );
  OAI21_X1 U17366 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n14068), .A(n14035), .ZN(
        n14037) );
  INV_X1 U17367 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14489) );
  NAND2_X1 U17368 ( .A1(n10265), .A2(n14489), .ZN(n14036) );
  NAND2_X1 U17369 ( .A1(n14037), .A2(n14036), .ZN(n14420) );
  MUX2_X1 U17370 ( .A(n14057), .B(n14293), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14039) );
  NAND2_X1 U17371 ( .A1(n14058), .A2(n15835), .ZN(n14038) );
  NAND2_X1 U17372 ( .A1(n14039), .A2(n14038), .ZN(n14408) );
  INV_X1 U17373 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14040) );
  NAND2_X1 U17374 ( .A1(n14048), .A2(n14040), .ZN(n14043) );
  NAND2_X1 U17375 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14041) );
  OAI211_X1 U17376 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n14068), .A(n14041), .B(
        n14066), .ZN(n14042) );
  AND2_X1 U17377 ( .A1(n14043), .A2(n14042), .ZN(n14382) );
  INV_X1 U17378 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14679) );
  NAND2_X1 U17379 ( .A1(n14066), .A2(n14679), .ZN(n14044) );
  OAI211_X1 U17380 ( .C1(n14068), .C2(P1_EBX_REG_22__SCAN_IN), .A(n14044), .B(
        n14293), .ZN(n14047) );
  INV_X1 U17381 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14045) );
  NAND2_X1 U17382 ( .A1(n10265), .A2(n14045), .ZN(n14046) );
  NAND2_X1 U17383 ( .A1(n14047), .A2(n14046), .ZN(n14396) );
  INV_X1 U17384 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14481) );
  NAND2_X1 U17385 ( .A1(n14048), .A2(n14481), .ZN(n14051) );
  NAND2_X1 U17386 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14049) );
  OAI211_X1 U17387 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n14068), .A(n14049), .B(
        n14066), .ZN(n14050) );
  AND2_X1 U17388 ( .A1(n14051), .A2(n14050), .ZN(n14357) );
  NAND2_X1 U17389 ( .A1(n14066), .A2(n14835), .ZN(n14052) );
  OAI211_X1 U17390 ( .C1(n14068), .C2(P1_EBX_REG_24__SCAN_IN), .A(n14052), .B(
        n14293), .ZN(n14055) );
  INV_X1 U17391 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14053) );
  NAND2_X1 U17392 ( .A1(n10265), .A2(n14053), .ZN(n14054) );
  NAND2_X1 U17393 ( .A1(n14055), .A2(n14054), .ZN(n14368) );
  NAND2_X1 U17394 ( .A1(n14357), .A2(n14368), .ZN(n14056) );
  MUX2_X1 U17395 ( .A(n14057), .B(n14293), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14060) );
  NAND2_X1 U17396 ( .A1(n14058), .A2(n14812), .ZN(n14059) );
  NAND2_X1 U17397 ( .A1(n14060), .A2(n14059), .ZN(n14334) );
  INV_X1 U17398 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14643) );
  NAND2_X1 U17399 ( .A1(n14066), .A2(n14643), .ZN(n14061) );
  OAI211_X1 U17400 ( .C1(n13171), .C2(P1_EBX_REG_26__SCAN_IN), .A(n14061), .B(
        n14293), .ZN(n14063) );
  INV_X1 U17401 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14480) );
  NAND2_X1 U17402 ( .A1(n10265), .A2(n14480), .ZN(n14062) );
  AND2_X1 U17403 ( .A1(n14063), .A2(n14062), .ZN(n14333) );
  NOR2_X1 U17404 ( .A1(n14334), .A2(n14333), .ZN(n14064) );
  NAND2_X1 U17405 ( .A1(n14066), .A2(n14065), .ZN(n14067) );
  OAI211_X1 U17406 ( .C1(n14068), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14067), .B(
        n14293), .ZN(n14070) );
  INV_X1 U17407 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14478) );
  NAND2_X1 U17408 ( .A1(n10265), .A2(n14478), .ZN(n14069) );
  AND2_X1 U17409 ( .A1(n14070), .A2(n14069), .ZN(n14318) );
  OR2_X2 U17410 ( .A1(n14336), .A2(n14318), .ZN(n14320) );
  OAI22_X1 U17411 ( .A1(n14071), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n13171), .ZN(n14292) );
  MUX2_X1 U17412 ( .A(n14292), .B(P1_EBX_REG_29__SCAN_IN), .S(n10265), .Z(
        n14307) );
  NOR2_X2 U17413 ( .A1(n14320), .A2(n14307), .ZN(n14309) );
  MUX2_X1 U17414 ( .A(n14293), .B(n14295), .S(n14309), .Z(n14072) );
  NOR3_X1 U17415 ( .A1(n14907), .A2(n16000), .A3(n14075), .ZN(n14869) );
  NAND2_X1 U17416 ( .A1(n14903), .A2(n14869), .ZN(n14870) );
  NAND2_X1 U17417 ( .A1(n14869), .A2(n14891), .ZN(n14873) );
  AOI211_X1 U17418 ( .C1(n14870), .C2(n14913), .A(n14076), .B(n14873), .ZN(
        n14077) );
  OR2_X1 U17419 ( .A1(n14077), .A2(n14939), .ZN(n14078) );
  INV_X1 U17420 ( .A(n14894), .ZN(n14918) );
  NAND2_X1 U17421 ( .A1(n14078), .A2(n14918), .ZN(n15834) );
  NOR2_X1 U17422 ( .A1(n14939), .A2(n14079), .ZN(n14080) );
  OR2_X1 U17423 ( .A1(n15834), .A2(n14080), .ZN(n14853) );
  NOR2_X1 U17424 ( .A1(n20168), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14081) );
  NOR2_X1 U17425 ( .A1(n14853), .A2(n14081), .ZN(n14840) );
  INV_X1 U17426 ( .A(n14082), .ZN(n14651) );
  OAI22_X1 U17427 ( .A1(n14651), .A2(n14892), .B1(n20168), .B2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14084) );
  NOR2_X1 U17428 ( .A1(n14890), .A2(n14615), .ZN(n14083) );
  NOR2_X1 U17429 ( .A1(n14084), .A2(n14083), .ZN(n14085) );
  AND2_X1 U17430 ( .A1(n14840), .A2(n14085), .ZN(n14087) );
  NAND2_X1 U17431 ( .A1(n14087), .A2(n14939), .ZN(n14092) );
  INV_X1 U17432 ( .A(n14086), .ZN(n14801) );
  NAND2_X1 U17433 ( .A1(n14092), .A2(n14801), .ZN(n14090) );
  INV_X1 U17434 ( .A(n14087), .ZN(n14829) );
  NOR2_X1 U17435 ( .A1(n14939), .A2(n14088), .ZN(n14089) );
  NOR2_X1 U17436 ( .A1(n14829), .A2(n14089), .ZN(n14813) );
  NAND2_X1 U17437 ( .A1(n14090), .A2(n14813), .ZN(n14792) );
  AOI211_X1 U17438 ( .C1(n14606), .C2(n14895), .A(n14091), .B(n14792), .ZN(
        n14780) );
  INV_X1 U17439 ( .A(n14092), .ZN(n14094) );
  NOR3_X1 U17440 ( .A1(n14780), .A2(n14094), .A3(n14093), .ZN(n14095) );
  OAI21_X1 U17441 ( .B1(n9712), .B2(n20164), .A(n14096), .ZN(P1_U3000) );
  INV_X1 U17442 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n14097) );
  NOR2_X1 U17443 ( .A1(n15154), .A2(n14097), .ZN(n14226) );
  INV_X1 U17444 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n14098) );
  NOR2_X1 U17445 ( .A1(n15154), .A2(n14098), .ZN(n14949) );
  XNOR2_X1 U17446 ( .A(n14950), .B(n14949), .ZN(n16066) );
  INV_X1 U17447 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14258) );
  OAI21_X1 U17448 ( .B1(n16066), .B2(n15158), .A(n14258), .ZN(n15151) );
  INV_X1 U17449 ( .A(n16066), .ZN(n14099) );
  NAND3_X1 U17450 ( .A1(n14099), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13426), .ZN(n15170) );
  NAND2_X1 U17451 ( .A1(n15151), .A2(n15170), .ZN(n14233) );
  NAND2_X1 U17452 ( .A1(n14102), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14103) );
  XNOR2_X1 U17453 ( .A(n14106), .B(n10158), .ZN(n19057) );
  AND2_X1 U17454 ( .A1(n19057), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15574) );
  NOR2_X1 U17455 ( .A1(n14107), .A2(n15158), .ZN(n14113) );
  AND2_X1 U17456 ( .A1(n14113), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16227) );
  INV_X1 U17457 ( .A(n14117), .ZN(n14111) );
  NAND2_X1 U17458 ( .A1(n14206), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14109) );
  MUX2_X1 U17459 ( .A(n14109), .B(n14206), .S(n14108), .Z(n14110) );
  AND2_X1 U17460 ( .A1(n14111), .A2(n14110), .ZN(n14129) );
  NAND2_X1 U17461 ( .A1(n14129), .A2(n13426), .ZN(n14112) );
  NAND2_X1 U17462 ( .A1(n14112), .A2(n15558), .ZN(n15549) );
  INV_X1 U17463 ( .A(n14113), .ZN(n14115) );
  INV_X1 U17464 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14114) );
  NAND2_X1 U17465 ( .A1(n14115), .A2(n14114), .ZN(n16225) );
  INV_X1 U17466 ( .A(n19057), .ZN(n14116) );
  NAND2_X1 U17467 ( .A1(n14116), .A2(n15568), .ZN(n16224) );
  AND2_X1 U17468 ( .A1(n16225), .A2(n16224), .ZN(n15531) );
  NAND2_X1 U17469 ( .A1(n14117), .A2(n19138), .ZN(n14121) );
  NOR2_X1 U17470 ( .A1(n14117), .A2(n19138), .ZN(n14118) );
  NAND2_X1 U17471 ( .A1(n14206), .A2(n14118), .ZN(n14119) );
  AND2_X1 U17472 ( .A1(n14220), .A2(n14119), .ZN(n14120) );
  NAND2_X1 U17473 ( .A1(n14121), .A2(n14120), .ZN(n19035) );
  OR2_X1 U17474 ( .A1(n19035), .A2(n15158), .ZN(n14122) );
  INV_X1 U17475 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16200) );
  NAND2_X1 U17476 ( .A1(n14122), .A2(n16200), .ZN(n16202) );
  NAND2_X1 U17477 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n14121), .ZN(n14124) );
  NOR2_X1 U17478 ( .A1(n15154), .A2(n14124), .ZN(n14125) );
  OR2_X1 U17479 ( .A1(n14126), .A2(n14125), .ZN(n19018) );
  INV_X1 U17480 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14127) );
  OAI21_X1 U17481 ( .B1(n19018), .B2(n15158), .A(n14127), .ZN(n15535) );
  AND4_X1 U17482 ( .A1(n15549), .A2(n15531), .A3(n16202), .A4(n15535), .ZN(
        n14128) );
  INV_X1 U17483 ( .A(n14129), .ZN(n19043) );
  NAND2_X1 U17484 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14130) );
  NAND2_X1 U17485 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14131) );
  OR2_X1 U17486 ( .A1(n19018), .A2(n14131), .ZN(n15534) );
  OR3_X1 U17487 ( .A1(n19035), .A2(n15158), .A3(n16200), .ZN(n16201) );
  AND3_X1 U17488 ( .A1(n16203), .A2(n15534), .A3(n16201), .ZN(n14132) );
  NAND2_X1 U17489 ( .A1(n15521), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14135) );
  NAND3_X1 U17490 ( .A1(n14206), .A2(n14133), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n14134) );
  NAND2_X1 U17491 ( .A1(n14140), .A2(n14134), .ZN(n15028) );
  OR2_X1 U17492 ( .A1(n15028), .A2(n15158), .ZN(n15519) );
  INV_X1 U17493 ( .A(n15521), .ZN(n14136) );
  INV_X1 U17494 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15524) );
  NAND2_X1 U17495 ( .A1(n14140), .A2(n14139), .ZN(n14141) );
  NAND2_X1 U17496 ( .A1(n14142), .A2(n14141), .ZN(n19006) );
  OR2_X1 U17497 ( .A1(n19006), .A2(n15158), .ZN(n14144) );
  INV_X1 U17498 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14143) );
  AND2_X1 U17499 ( .A1(n14144), .A2(n14143), .ZN(n15293) );
  NAND2_X1 U17500 ( .A1(n14206), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14147) );
  MUX2_X1 U17501 ( .A(n14206), .B(n14147), .S(n14146), .Z(n14149) );
  NAND2_X1 U17502 ( .A1(n14149), .A2(n14148), .ZN(n18937) );
  OR2_X1 U17503 ( .A1(n18937), .A2(n15158), .ZN(n14150) );
  INV_X1 U17504 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15452) );
  NAND2_X1 U17505 ( .A1(n14150), .A2(n15452), .ZN(n15256) );
  XNOR2_X1 U17506 ( .A(n9706), .B(n14151), .ZN(n18947) );
  NAND2_X1 U17507 ( .A1(n18947), .A2(n13426), .ZN(n14183) );
  INV_X1 U17508 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U17509 ( .A1(n14183), .A2(n15451), .ZN(n15273) );
  INV_X1 U17510 ( .A(n14152), .ZN(n14153) );
  XNOR2_X1 U17511 ( .A(n14159), .B(n14153), .ZN(n18959) );
  NAND2_X1 U17512 ( .A1(n18959), .A2(n13426), .ZN(n14154) );
  INV_X1 U17513 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15481) );
  NAND2_X1 U17514 ( .A1(n14154), .A2(n15481), .ZN(n15472) );
  AND2_X1 U17515 ( .A1(n15273), .A2(n15472), .ZN(n15253) );
  AND2_X1 U17516 ( .A1(n15256), .A2(n15253), .ZN(n15239) );
  INV_X1 U17517 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14155) );
  OAI21_X1 U17518 ( .B1(n14180), .B2(n15158), .A(n14155), .ZN(n15241) );
  INV_X1 U17519 ( .A(n14156), .ZN(n14158) );
  NAND2_X1 U17520 ( .A1(n14158), .A2(n10154), .ZN(n14160) );
  NAND2_X1 U17521 ( .A1(n14160), .A2(n14159), .ZN(n18969) );
  OR2_X1 U17522 ( .A1(n18969), .A2(n15158), .ZN(n14162) );
  INV_X1 U17523 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14161) );
  NAND2_X1 U17524 ( .A1(n14162), .A2(n14161), .ZN(n15280) );
  NOR2_X1 U17525 ( .A1(n15154), .A2(n14163), .ZN(n14165) );
  INV_X1 U17526 ( .A(n14220), .ZN(n14164) );
  AOI21_X1 U17527 ( .B1(n14176), .B2(n14165), .A(n14164), .ZN(n14166) );
  NAND2_X1 U17528 ( .A1(n14167), .A2(n14166), .ZN(n18979) );
  NAND2_X1 U17529 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14168) );
  INV_X1 U17530 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15770) );
  OAI21_X1 U17531 ( .B1(n18979), .B2(n15158), .A(n15770), .ZN(n14169) );
  INV_X1 U17532 ( .A(n14186), .ZN(n14172) );
  NAND2_X1 U17533 ( .A1(n14172), .A2(n14171), .ZN(n16177) );
  INV_X1 U17534 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14173) );
  NOR2_X1 U17535 ( .A1(n15154), .A2(n14173), .ZN(n14174) );
  NAND2_X1 U17536 ( .A1(n14175), .A2(n14174), .ZN(n14177) );
  NAND2_X1 U17537 ( .A1(n14177), .A2(n14176), .ZN(n18992) );
  INV_X1 U17538 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14178) );
  OAI21_X1 U17539 ( .B1(n18992), .B2(n15158), .A(n14178), .ZN(n15497) );
  AND4_X1 U17540 ( .A1(n15280), .A2(n15762), .A3(n16177), .A4(n15497), .ZN(
        n14179) );
  NAND3_X1 U17541 ( .A1(n15239), .A2(n15241), .A3(n14179), .ZN(n14195) );
  INV_X1 U17542 ( .A(n14180), .ZN(n14182) );
  AND2_X1 U17543 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14181) );
  NAND2_X1 U17544 ( .A1(n14182), .A2(n14181), .ZN(n15240) );
  INV_X1 U17545 ( .A(n14183), .ZN(n14184) );
  NAND2_X1 U17546 ( .A1(n14184), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15274) );
  NAND2_X1 U17547 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14185) );
  OR2_X1 U17548 ( .A1(n18969), .A2(n14185), .ZN(n15279) );
  NAND2_X1 U17549 ( .A1(n15279), .A2(n15281), .ZN(n15234) );
  NAND2_X1 U17550 ( .A1(n14186), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16178) );
  INV_X1 U17551 ( .A(n18992), .ZN(n14188) );
  AND2_X1 U17552 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14187) );
  NAND2_X1 U17553 ( .A1(n14188), .A2(n14187), .ZN(n15496) );
  NAND2_X1 U17554 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14189) );
  OR2_X1 U17555 ( .A1(n19006), .A2(n14189), .ZN(n15291) );
  NAND3_X1 U17556 ( .A1(n16178), .A2(n15496), .A3(n15291), .ZN(n14190) );
  NOR2_X1 U17557 ( .A1(n15234), .A2(n14190), .ZN(n14192) );
  AND2_X1 U17558 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14191) );
  NAND2_X1 U17559 ( .A1(n18959), .A2(n14191), .ZN(n15471) );
  AND3_X1 U17560 ( .A1(n15274), .A2(n14192), .A3(n15471), .ZN(n14193) );
  OR3_X1 U17561 ( .A1(n18937), .A2(n15158), .A3(n15452), .ZN(n15255) );
  AND3_X1 U17562 ( .A1(n15240), .A2(n14193), .A3(n15255), .ZN(n14194) );
  NAND2_X1 U17563 ( .A1(n14197), .A2(n10163), .ZN(n14198) );
  NAND2_X1 U17564 ( .A1(n14202), .A2(n14198), .ZN(n15773) );
  OR2_X1 U17565 ( .A1(n15773), .A2(n15158), .ZN(n14199) );
  INV_X1 U17566 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15409) );
  NAND2_X1 U17567 ( .A1(n14199), .A2(n15409), .ZN(n15404) );
  INV_X1 U17568 ( .A(n14199), .ZN(n14200) );
  NAND2_X1 U17569 ( .A1(n14200), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15405) );
  XNOR2_X1 U17570 ( .A(n14202), .B(n14201), .ZN(n15023) );
  NAND2_X1 U17571 ( .A1(n15023), .A2(n13426), .ZN(n14204) );
  XNOR2_X1 U17572 ( .A(n14204), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15390) );
  INV_X1 U17573 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14203) );
  NOR2_X1 U17574 ( .A1(n14204), .A2(n14203), .ZN(n14205) );
  NAND3_X1 U17575 ( .A1(n14207), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n14206), 
        .ZN(n14208) );
  NAND2_X1 U17576 ( .A1(n14208), .A2(n14220), .ZN(n14209) );
  OR2_X1 U17577 ( .A1(n14209), .A2(n9703), .ZN(n15010) );
  NOR2_X1 U17578 ( .A1(n15010), .A2(n15158), .ZN(n14210) );
  AND2_X1 U17579 ( .A1(n14210), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15376) );
  INV_X1 U17580 ( .A(n14210), .ZN(n14211) );
  INV_X1 U17581 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15380) );
  NAND2_X1 U17582 ( .A1(n14211), .A2(n15380), .ZN(n15375) );
  NAND2_X1 U17583 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n14222), .ZN(n14212) );
  NOR2_X1 U17584 ( .A1(n15154), .A2(n14212), .ZN(n14213) );
  NOR2_X1 U17585 ( .A1(n14951), .A2(n14213), .ZN(n14215) );
  AND2_X1 U17586 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14214) );
  NAND2_X1 U17587 ( .A1(n14215), .A2(n14214), .ZN(n14232) );
  INV_X1 U17588 ( .A(n14215), .ZN(n16078) );
  INV_X1 U17589 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15356) );
  OAI21_X1 U17590 ( .B1(n16078), .B2(n15158), .A(n15356), .ZN(n14216) );
  NAND2_X1 U17591 ( .A1(n14232), .A2(n14216), .ZN(n15215) );
  NOR2_X1 U17592 ( .A1(n14217), .A2(n15158), .ZN(n15193) );
  NOR2_X1 U17593 ( .A1(n9703), .A2(n15070), .ZN(n14218) );
  NAND2_X1 U17594 ( .A1(n14206), .A2(n14218), .ZN(n14219) );
  AND2_X1 U17595 ( .A1(n14220), .A2(n14219), .ZN(n14221) );
  NAND2_X1 U17596 ( .A1(n14222), .A2(n14221), .ZN(n16084) );
  INV_X1 U17597 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15355) );
  NAND2_X1 U17598 ( .A1(n14230), .A2(n15355), .ZN(n15223) );
  INV_X1 U17599 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15197) );
  INV_X1 U17600 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15327) );
  NAND2_X1 U17601 ( .A1(n14227), .A2(n14226), .ZN(n14228) );
  NAND2_X1 U17602 ( .A1(n14950), .A2(n14228), .ZN(n14995) );
  NOR2_X1 U17603 ( .A1(n14995), .A2(n15158), .ZN(n15194) );
  INV_X1 U17604 ( .A(n14230), .ZN(n14231) );
  NAND2_X1 U17605 ( .A1(n14231), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15224) );
  XOR2_X1 U17606 ( .A(n14233), .B(n15152), .Z(n15190) );
  NAND2_X1 U17607 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16281) );
  AOI21_X1 U17608 ( .B1(n15579), .B2(n16281), .A(n16276), .ZN(n15559) );
  NAND3_X1 U17609 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15500) );
  NAND2_X1 U17610 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16259) );
  INV_X1 U17611 ( .A(n16259), .ZN(n15508) );
  NAND2_X1 U17612 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15508), .ZN(
        n15447) );
  NOR2_X1 U17613 ( .A1(n15500), .A2(n15447), .ZN(n15285) );
  NAND4_X1 U17614 ( .A1(n15285), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15440) );
  NAND2_X1 U17615 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15248) );
  NOR3_X1 U17616 ( .A1(n15481), .A2(n15440), .A3(n15248), .ZN(n15426) );
  NAND2_X1 U17617 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15426), .ZN(
        n15393) );
  NAND2_X1 U17618 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15395) );
  NOR2_X1 U17619 ( .A1(n15393), .A2(n15395), .ZN(n14256) );
  NAND2_X1 U17620 ( .A1(n15559), .A2(n14256), .ZN(n14235) );
  INV_X1 U17621 ( .A(n19244), .ZN(n14234) );
  NAND2_X1 U17622 ( .A1(n15787), .A2(n14234), .ZN(n15538) );
  NAND2_X1 U17623 ( .A1(n14235), .A2(n15538), .ZN(n14236) );
  NAND2_X1 U17624 ( .A1(n14236), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15381) );
  NAND2_X1 U17625 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14257) );
  OR2_X1 U17626 ( .A1(n15381), .A2(n14257), .ZN(n14237) );
  NAND2_X1 U17627 ( .A1(n14237), .A2(n15538), .ZN(n15339) );
  NAND2_X1 U17628 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14238), .ZN(
        n15567) );
  INV_X1 U17629 ( .A(n15540), .ZN(n15555) );
  OR2_X1 U17630 ( .A1(n15393), .A2(n15555), .ZN(n15420) );
  NOR2_X1 U17631 ( .A1(n15395), .A2(n15420), .ZN(n15382) );
  NAND2_X1 U17632 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15382), .ZN(
        n15367) );
  NOR2_X1 U17633 ( .A1(n14257), .A2(n15367), .ZN(n15303) );
  NAND2_X1 U17634 ( .A1(n15327), .A2(n15303), .ZN(n15340) );
  NAND2_X1 U17635 ( .A1(n15339), .A2(n15340), .ZN(n15336) );
  AND2_X1 U17636 ( .A1(n14989), .A2(n14239), .ZN(n14240) );
  NOR2_X1 U17637 ( .A1(n19066), .A2(n19915), .ZN(n15183) );
  INV_X1 U17638 ( .A(n15183), .ZN(n14244) );
  INV_X1 U17639 ( .A(n15303), .ZN(n15326) );
  AOI21_X1 U17640 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14258), .A(
        n15197), .ZN(n14241) );
  AOI211_X1 U17641 ( .C1(n14258), .C2(n15197), .A(n15326), .B(n14241), .ZN(
        n14242) );
  INV_X1 U17642 ( .A(n14242), .ZN(n14243) );
  INV_X1 U17643 ( .A(n14245), .ZN(n14246) );
  OAI21_X1 U17644 ( .B1(n16061), .B2(n16277), .A(n14246), .ZN(n14259) );
  NAND2_X1 U17645 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n14254), .ZN(
        n14255) );
  XNOR2_X1 U17646 ( .A(n14252), .B(n15158), .ZN(n15564) );
  INV_X1 U17647 ( .A(n15564), .ZN(n14253) );
  XOR2_X1 U17648 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14254), .Z(
        n16222) );
  INV_X1 U17649 ( .A(n14257), .ZN(n15354) );
  NAND3_X1 U17650 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15301) );
  OAI21_X1 U17651 ( .B1(n15190), .B2(n16273), .A(n14260), .ZN(P2_U3017) );
  INV_X1 U17652 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15178) );
  OAI22_X1 U17653 ( .A1(n14261), .A2(n19918), .B1(n15593), .B2(n15178), .ZN(
        n14262) );
  INV_X1 U17654 ( .A(n14262), .ZN(n14265) );
  NAND2_X1 U17655 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14264) );
  NAND2_X1 U17656 ( .A1(n11962), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14263) );
  AND3_X1 U17657 ( .A1(n14265), .A2(n14264), .A3(n14263), .ZN(n14957) );
  INV_X1 U17658 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n15153) );
  MUX2_X1 U17659 ( .A(n15177), .B(n15153), .S(n12991), .Z(n14266) );
  OAI21_X1 U17660 ( .B1(n14267), .B2(n19145), .A(n14266), .ZN(P2_U2857) );
  NAND2_X1 U17661 ( .A1(n14268), .A2(n19173), .ZN(n14274) );
  OAI22_X1 U17662 ( .A1(n16070), .A2(n16119), .B1(n15130), .B2(n14269), .ZN(
        n14270) );
  AOI21_X1 U17663 ( .B1(n16127), .B2(n14271), .A(n14270), .ZN(n14273) );
  AOI22_X1 U17664 ( .A1(n19153), .A2(BUF1_REG_29__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14272) );
  OAI211_X1 U17665 ( .C1(n12027), .C2(n14274), .A(n14273), .B(n14272), .ZN(
        P2_U2890) );
  INV_X1 U17666 ( .A(n14275), .ZN(n14290) );
  NAND2_X1 U17667 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14285) );
  INV_X1 U17668 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14326) );
  NAND3_X1 U17669 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14277) );
  NAND3_X1 U17670 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n14276), .ZN(n14462) );
  NOR2_X1 U17671 ( .A1(n14277), .A2(n14462), .ZN(n14438) );
  NAND4_X1 U17672 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .A3(P1_REIP_REG_19__SCAN_IN), .A4(n14438), .ZN(n14395) );
  NAND3_X1 U17673 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(P1_REIP_REG_21__SCAN_IN), .ZN(n14284) );
  NOR2_X1 U17674 ( .A1(n14395), .A2(n14284), .ZN(n14356) );
  NAND4_X1 U17675 ( .A1(n14356), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .A4(P1_REIP_REG_26__SCAN_IN), .ZN(n14332) );
  NOR2_X1 U17676 ( .A1(n14326), .A2(n14332), .ZN(n14278) );
  AOI21_X1 U17677 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14278), .A(n14439), 
        .ZN(n14322) );
  AOI21_X1 U17678 ( .B1(n14285), .B2(n15910), .A(n14322), .ZN(n14299) );
  INV_X1 U17679 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14280) );
  AOI22_X1 U17680 ( .A1(n20077), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20051), .ZN(n14279) );
  OAI21_X1 U17681 ( .B1(n14299), .B2(n14280), .A(n14279), .ZN(n14287) );
  NAND2_X1 U17682 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n14281), .ZN(n15908) );
  NAND2_X1 U17683 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14282) );
  NAND4_X1 U17684 ( .A1(n15875), .A2(P1_REIP_REG_17__SCAN_IN), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_15__SCAN_IN), .ZN(n14440) );
  INV_X1 U17685 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20770) );
  NOR2_X1 U17686 ( .A1(n14440), .A2(n20770), .ZN(n14437) );
  AND2_X1 U17687 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14283) );
  NAND2_X1 U17688 ( .A1(n14437), .A2(n14283), .ZN(n14417) );
  NAND3_X1 U17689 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_25__SCAN_IN), .ZN(n14340) );
  INV_X1 U17690 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20943) );
  NOR3_X1 U17691 ( .A1(n14351), .A2(n14340), .A3(n20943), .ZN(n14327) );
  NAND2_X1 U17692 ( .A1(n14327), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14315) );
  NOR3_X1 U17693 ( .A1(n14315), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14285), 
        .ZN(n14286) );
  AOI211_X1 U17694 ( .C1(n14288), .C2(n20053), .A(n14287), .B(n14286), .ZN(
        n14289) );
  OAI21_X1 U17695 ( .B1(n14290), .B2(n15914), .A(n14289), .ZN(P1_U2809) );
  INV_X1 U17696 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14476) );
  OAI22_X1 U17697 ( .A1(n20038), .A2(n14476), .B1(n14291), .B2(n20075), .ZN(
        n14297) );
  OAI22_X1 U17698 ( .A1(n14309), .A2(n14293), .B1(n14292), .B2(n14320), .ZN(
        n14294) );
  XOR2_X1 U17699 ( .A(n14295), .B(n14294), .Z(n14776) );
  NOR2_X1 U17700 ( .A1(n14776), .A2(n20084), .ZN(n14296) );
  AOI211_X1 U17701 ( .C1(n14298), .C2(n20049), .A(n14297), .B(n14296), .ZN(
        n14303) );
  INV_X1 U17702 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20924) );
  NOR2_X1 U17703 ( .A1(n14315), .A2(n20924), .ZN(n14301) );
  INV_X1 U17704 ( .A(n14299), .ZN(n14300) );
  OAI21_X1 U17705 ( .B1(n14301), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14300), 
        .ZN(n14302) );
  OAI211_X1 U17706 ( .C1(n14529), .C2(n15914), .A(n14303), .B(n14302), .ZN(
        P1_U2810) );
  AOI21_X1 U17707 ( .B1(n14306), .B2(n14304), .A(n14305), .ZN(n14530) );
  NAND2_X1 U17708 ( .A1(n14530), .A2(n20055), .ZN(n14314) );
  AND2_X1 U17709 ( .A1(n14320), .A2(n14307), .ZN(n14308) );
  NOR2_X1 U17710 ( .A1(n14309), .A2(n14308), .ZN(n14788) );
  AOI22_X1 U17711 ( .A1(n20077), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20051), .ZN(n14311) );
  NAND2_X1 U17712 ( .A1(n14322), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14310) );
  OAI211_X1 U17713 ( .C1(n20087), .C2(n14610), .A(n14311), .B(n14310), .ZN(
        n14312) );
  AOI21_X1 U17714 ( .B1(n14788), .B2(n20053), .A(n14312), .ZN(n14313) );
  OAI211_X1 U17715 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14315), .A(n14314), 
        .B(n14313), .ZN(P1_U2811) );
  OAI21_X1 U17716 ( .B1(n14316), .B2(n14317), .A(n14304), .ZN(n14627) );
  NAND2_X1 U17717 ( .A1(n14336), .A2(n14318), .ZN(n14319) );
  NAND2_X1 U17718 ( .A1(n14320), .A2(n14319), .ZN(n14798) );
  INV_X1 U17719 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14624) );
  OAI22_X1 U17720 ( .A1(n20038), .A2(n14478), .B1(n14624), .B2(n20075), .ZN(
        n14321) );
  AOI21_X1 U17721 ( .B1(n14322), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14321), 
        .ZN(n14324) );
  NAND2_X1 U17722 ( .A1(n20049), .A2(n14622), .ZN(n14323) );
  OAI211_X1 U17723 ( .C1(n14798), .C2(n20084), .A(n14324), .B(n14323), .ZN(
        n14325) );
  AOI21_X1 U17724 ( .B1(n14327), .B2(n14326), .A(n14325), .ZN(n14328) );
  OAI21_X1 U17725 ( .B1(n14627), .B2(n15914), .A(n14328), .ZN(P1_U2812) );
  AOI21_X1 U17726 ( .B1(n14330), .B2(n14329), .A(n14316), .ZN(n14331) );
  INV_X1 U17727 ( .A(n14331), .ZN(n14638) );
  AND2_X1 U17728 ( .A1(n14332), .A2(n15910), .ZN(n14350) );
  INV_X1 U17729 ( .A(n14333), .ZN(n14346) );
  NAND2_X1 U17730 ( .A1(n14358), .A2(n14346), .ZN(n14335) );
  NAND2_X1 U17731 ( .A1(n14335), .A2(n14334), .ZN(n14337) );
  AND2_X1 U17732 ( .A1(n14337), .A2(n14336), .ZN(n14809) );
  NAND2_X1 U17733 ( .A1(n14809), .A2(n20053), .ZN(n14339) );
  AOI22_X1 U17734 ( .A1(n20077), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20051), .ZN(n14338) );
  OAI211_X1 U17735 ( .C1(n20087), .C2(n14635), .A(n14339), .B(n14338), .ZN(
        n14342) );
  NOR3_X1 U17736 ( .A1(n14351), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14340), 
        .ZN(n14341) );
  AOI211_X1 U17737 ( .C1(n14350), .C2(P1_REIP_REG_27__SCAN_IN), .A(n14342), 
        .B(n14341), .ZN(n14343) );
  OAI21_X1 U17738 ( .B1(n14638), .B2(n15914), .A(n14343), .ZN(P1_U2813) );
  XNOR2_X1 U17739 ( .A(n14344), .B(n14345), .ZN(n14650) );
  XNOR2_X1 U17740 ( .A(n14358), .B(n14346), .ZN(n14819) );
  AOI22_X1 U17741 ( .A1(n20077), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20051), .ZN(n14348) );
  NAND2_X1 U17742 ( .A1(n20049), .A2(n14645), .ZN(n14347) );
  OAI211_X1 U17743 ( .C1(n14819), .C2(n20084), .A(n14348), .B(n14347), .ZN(
        n14349) );
  AOI21_X1 U17744 ( .B1(n14350), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14349), 
        .ZN(n14353) );
  INV_X1 U17745 ( .A(n14351), .ZN(n14376) );
  INV_X1 U17746 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20905) );
  NAND4_X1 U17747 ( .A1(n14376), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .A4(n20905), .ZN(n14352) );
  OAI211_X1 U17748 ( .C1(n14650), .C2(n15914), .A(n14353), .B(n14352), .ZN(
        P1_U2814) );
  OAI21_X1 U17749 ( .B1(n14355), .B2(n14354), .A(n14344), .ZN(n14656) );
  XOR2_X1 U17750 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .Z(n14365) );
  OR2_X1 U17751 ( .A1(n14356), .A2(n14439), .ZN(n14387) );
  INV_X1 U17752 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20882) );
  NOR2_X1 U17753 ( .A1(n14387), .A2(n20882), .ZN(n14364) );
  INV_X1 U17754 ( .A(n14369), .ZN(n14383) );
  AOI21_X1 U17755 ( .B1(n14383), .B2(n14368), .A(n14357), .ZN(n14359) );
  OR2_X1 U17756 ( .A1(n14359), .A2(n14358), .ZN(n14827) );
  AOI22_X1 U17757 ( .A1(n20077), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20051), .ZN(n14362) );
  NAND2_X1 U17758 ( .A1(n20049), .A2(n14360), .ZN(n14361) );
  OAI211_X1 U17759 ( .C1(n14827), .C2(n20084), .A(n14362), .B(n14361), .ZN(
        n14363) );
  AOI211_X1 U17760 ( .C1(n14376), .C2(n14365), .A(n14364), .B(n14363), .ZN(
        n14366) );
  OAI21_X1 U17761 ( .B1(n14656), .B2(n15914), .A(n14366), .ZN(P1_U2815) );
  XNOR2_X1 U17762 ( .A(n14381), .B(n14367), .ZN(n14670) );
  INV_X1 U17763 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14375) );
  XNOR2_X1 U17764 ( .A(n14369), .B(n14368), .ZN(n14841) );
  INV_X1 U17765 ( .A(n14665), .ZN(n14371) );
  AOI22_X1 U17766 ( .A1(n20077), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20051), .ZN(n14370) );
  OAI21_X1 U17767 ( .B1(n20087), .B2(n14371), .A(n14370), .ZN(n14372) );
  AOI21_X1 U17768 ( .B1(n20053), .B2(n14841), .A(n14372), .ZN(n14373) );
  OAI21_X1 U17769 ( .B1(n14387), .B2(n14375), .A(n14373), .ZN(n14374) );
  AOI21_X1 U17770 ( .B1(n14376), .B2(n14375), .A(n14374), .ZN(n14377) );
  OAI21_X1 U17771 ( .B1(n14670), .B2(n15914), .A(n14377), .ZN(P1_U2816) );
  NAND2_X1 U17772 ( .A1(n14379), .A2(n14378), .ZN(n14380) );
  NAND2_X1 U17773 ( .A1(n14381), .A2(n14380), .ZN(n14676) );
  INV_X1 U17774 ( .A(n14673), .ZN(n14391) );
  AOI21_X1 U17775 ( .B1(n10015), .B2(n14396), .A(n14382), .ZN(n14384) );
  NOR2_X1 U17776 ( .A1(n14384), .A2(n14383), .ZN(n14483) );
  INV_X1 U17777 ( .A(n14483), .ZN(n14850) );
  AOI22_X1 U17778 ( .A1(n20077), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20051), .ZN(n14385) );
  OAI21_X1 U17779 ( .B1(n14850), .B2(n20084), .A(n14385), .ZN(n14390) );
  INV_X1 U17780 ( .A(n14417), .ZN(n14386) );
  NAND3_X1 U17781 ( .A1(n14386), .A2(P1_REIP_REG_22__SCAN_IN), .A3(
        P1_REIP_REG_21__SCAN_IN), .ZN(n14388) );
  INV_X1 U17782 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20960) );
  AOI21_X1 U17783 ( .B1(n14388), .B2(n20960), .A(n14387), .ZN(n14389) );
  AOI211_X1 U17784 ( .C1(n20049), .C2(n14391), .A(n14390), .B(n14389), .ZN(
        n14392) );
  OAI21_X1 U17785 ( .B1(n14676), .B2(n15914), .A(n14392), .ZN(P1_U2817) );
  XNOR2_X1 U17786 ( .A(P1_REIP_REG_22__SCAN_IN), .B(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14403) );
  XNOR2_X1 U17787 ( .A(n14406), .B(n14393), .ZN(n14686) );
  INV_X1 U17788 ( .A(n14686), .ZN(n14394) );
  NAND2_X1 U17789 ( .A1(n14394), .A2(n20055), .ZN(n14402) );
  AND2_X1 U17790 ( .A1(n14395), .A2(n15910), .ZN(n14424) );
  XNOR2_X1 U17791 ( .A(n14410), .B(n14396), .ZN(n14858) );
  NAND2_X1 U17792 ( .A1(n14858), .A2(n20053), .ZN(n14399) );
  AOI22_X1 U17793 ( .A1(n20077), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20051), .ZN(n14398) );
  NAND2_X1 U17794 ( .A1(n20049), .A2(n14681), .ZN(n14397) );
  NAND3_X1 U17795 ( .A1(n14399), .A2(n14398), .A3(n14397), .ZN(n14400) );
  AOI21_X1 U17796 ( .B1(n14424), .B2(P1_REIP_REG_22__SCAN_IN), .A(n14400), 
        .ZN(n14401) );
  OAI211_X1 U17797 ( .C1(n14417), .C2(n14403), .A(n14402), .B(n14401), .ZN(
        P1_U2818) );
  NOR2_X1 U17798 ( .A1(n14405), .A2(n14404), .ZN(n14407) );
  NOR2_X1 U17799 ( .A1(n14407), .A2(n14406), .ZN(n14693) );
  NAND2_X1 U17800 ( .A1(n14693), .A2(n20055), .ZN(n14416) );
  NAND2_X1 U17801 ( .A1(n14422), .A2(n14408), .ZN(n14409) );
  NAND2_X1 U17802 ( .A1(n14410), .A2(n14409), .ZN(n15838) );
  INV_X1 U17803 ( .A(n14691), .ZN(n14411) );
  NAND2_X1 U17804 ( .A1(n20049), .A2(n14411), .ZN(n14413) );
  AOI22_X1 U17805 ( .A1(n20077), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20051), .ZN(n14412) );
  OAI211_X1 U17806 ( .C1(n15838), .C2(n20084), .A(n14413), .B(n14412), .ZN(
        n14414) );
  AOI21_X1 U17807 ( .B1(n14424), .B2(P1_REIP_REG_21__SCAN_IN), .A(n14414), 
        .ZN(n14415) );
  OAI211_X1 U17808 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n14417), .A(n14416), 
        .B(n14415), .ZN(P1_U2819) );
  XNOR2_X1 U17809 ( .A(n14419), .B(n14418), .ZN(n14704) );
  OR2_X1 U17810 ( .A1(n14434), .A2(n14420), .ZN(n14421) );
  NAND2_X1 U17811 ( .A1(n14422), .A2(n14421), .ZN(n14874) );
  AOI22_X1 U17812 ( .A1(n20077), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20051), .ZN(n14423) );
  OAI21_X1 U17813 ( .B1(n14874), .B2(n20084), .A(n14423), .ZN(n14428) );
  AOI21_X1 U17814 ( .B1(n14437), .B2(P1_REIP_REG_19__SCAN_IN), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n14426) );
  INV_X1 U17815 ( .A(n14424), .ZN(n14425) );
  NOR2_X1 U17816 ( .A1(n14426), .A2(n14425), .ZN(n14427) );
  AOI211_X1 U17817 ( .C1(n20049), .C2(n14699), .A(n14428), .B(n14427), .ZN(
        n14429) );
  OAI21_X1 U17818 ( .B1(n14704), .B2(n15914), .A(n14429), .ZN(P1_U2820) );
  XNOR2_X1 U17819 ( .A(n14430), .B(n14431), .ZN(n14708) );
  INV_X1 U17820 ( .A(n14710), .ZN(n14446) );
  NOR2_X1 U17821 ( .A1(n9735), .A2(n14432), .ZN(n14433) );
  OR2_X1 U17822 ( .A1(n14434), .A2(n14433), .ZN(n15967) );
  NOR2_X1 U17823 ( .A1(n20038), .A2(n14490), .ZN(n14435) );
  AOI211_X1 U17824 ( .C1(n20051), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n9645), .B(n14435), .ZN(n14436) );
  OAI21_X1 U17825 ( .B1(n15967), .B2(n20084), .A(n14436), .ZN(n14445) );
  INV_X1 U17826 ( .A(n14437), .ZN(n14443) );
  INV_X1 U17827 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14442) );
  NOR2_X1 U17828 ( .A1(n14439), .A2(n14438), .ZN(n15873) );
  NOR2_X1 U17829 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14440), .ZN(n14452) );
  NOR3_X1 U17830 ( .A1(n15873), .A2(n14452), .A3(n14442), .ZN(n14441) );
  AOI21_X1 U17831 ( .B1(n14443), .B2(n14442), .A(n14441), .ZN(n14444) );
  AOI211_X1 U17832 ( .C1(n20049), .C2(n14446), .A(n14445), .B(n14444), .ZN(
        n14447) );
  OAI21_X1 U17833 ( .B1(n14708), .B2(n15914), .A(n14447), .ZN(P1_U2821) );
  AND2_X1 U17834 ( .A1(n14458), .A2(n14448), .ZN(n14498) );
  OAI21_X1 U17835 ( .B1(n14498), .B2(n14449), .A(n14430), .ZN(n14721) );
  AND2_X1 U17836 ( .A1(n14502), .A2(n14450), .ZN(n14451) );
  OR2_X1 U17837 ( .A1(n14451), .A2(n9735), .ZN(n15973) );
  NOR2_X1 U17838 ( .A1(n15973), .A2(n20084), .ZN(n14455) );
  AOI211_X1 U17839 ( .C1(n20051), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14452), .B(n9645), .ZN(n14453) );
  OAI21_X1 U17840 ( .B1(n14493), .B2(n20038), .A(n14453), .ZN(n14454) );
  AOI211_X1 U17841 ( .C1(n20049), .C2(n14719), .A(n14455), .B(n14454), .ZN(
        n14457) );
  NAND2_X1 U17842 ( .A1(n15873), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14456) );
  OAI211_X1 U17843 ( .C1(n14721), .C2(n15914), .A(n14457), .B(n14456), .ZN(
        P1_U2822) );
  INV_X1 U17844 ( .A(n14458), .ZN(n14595) );
  INV_X1 U17845 ( .A(n14497), .ZN(n14460) );
  NAND2_X1 U17846 ( .A1(n15910), .A2(n14462), .ZN(n15893) );
  INV_X1 U17847 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15988) );
  NAND2_X1 U17848 ( .A1(n15875), .A2(n15988), .ZN(n15887) );
  INV_X1 U17849 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20767) );
  AOI21_X1 U17850 ( .B1(n15893), .B2(n15887), .A(n20767), .ZN(n14472) );
  NAND3_X1 U17851 ( .A1(n15875), .A2(P1_REIP_REG_15__SCAN_IN), .A3(n20767), 
        .ZN(n14470) );
  OR2_X1 U17852 ( .A1(n15883), .A2(n14463), .ZN(n14464) );
  NAND2_X1 U17853 ( .A1(n14500), .A2(n14464), .ZN(n15982) );
  INV_X1 U17854 ( .A(n15982), .ZN(n14465) );
  AOI22_X1 U17855 ( .A1(n20053), .A2(n14465), .B1(n20077), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14466) );
  OAI211_X1 U17856 ( .C1(n20075), .C2(n14467), .A(n14466), .B(n20073), .ZN(
        n14468) );
  AOI21_X1 U17857 ( .B1(n20049), .B2(n14733), .A(n14468), .ZN(n14469) );
  NAND2_X1 U17858 ( .A1(n14470), .A2(n14469), .ZN(n14471) );
  AOI211_X1 U17859 ( .C1(n14737), .C2(n20055), .A(n14472), .B(n14471), .ZN(
        n14473) );
  INV_X1 U17860 ( .A(n14473), .ZN(P1_U2824) );
  OAI22_X1 U17861 ( .A1(n14475), .A2(n14523), .B1(n20103), .B2(n14474), .ZN(
        P1_U2841) );
  OAI222_X1 U17862 ( .A1(n14523), .A2(n14776), .B1(n14476), .B2(n20103), .C1(
        n14529), .C2(n14524), .ZN(P1_U2842) );
  INV_X1 U17863 ( .A(n14530), .ZN(n14613) );
  AOI22_X1 U17864 ( .A1(n14788), .A2(n20098), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14485), .ZN(n14477) );
  OAI21_X1 U17865 ( .B1(n14613), .B2(n14524), .A(n14477), .ZN(P1_U2843) );
  OAI222_X1 U17866 ( .A1(n14798), .A2(n14523), .B1(n14478), .B2(n20103), .C1(
        n14627), .C2(n14524), .ZN(P1_U2844) );
  AOI22_X1 U17867 ( .A1(n14809), .A2(n20098), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14485), .ZN(n14479) );
  OAI21_X1 U17868 ( .B1(n14638), .B2(n14524), .A(n14479), .ZN(P1_U2845) );
  OAI222_X1 U17869 ( .A1(n14524), .A2(n14650), .B1(n14480), .B2(n20103), .C1(
        n14523), .C2(n14819), .ZN(P1_U2846) );
  OAI222_X1 U17870 ( .A1(n14827), .A2(n14523), .B1(n14481), .B2(n20103), .C1(
        n14656), .C2(n14524), .ZN(P1_U2847) );
  AOI22_X1 U17871 ( .A1(n14841), .A2(n20098), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14485), .ZN(n14482) );
  OAI21_X1 U17872 ( .B1(n14670), .B2(n14524), .A(n14482), .ZN(P1_U2848) );
  AOI22_X1 U17873 ( .A1(n14483), .A2(n20098), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14485), .ZN(n14484) );
  OAI21_X1 U17874 ( .B1(n14676), .B2(n14524), .A(n14484), .ZN(P1_U2849) );
  AOI22_X1 U17875 ( .A1(n14858), .A2(n20098), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14485), .ZN(n14486) );
  OAI21_X1 U17876 ( .B1(n14686), .B2(n14524), .A(n14486), .ZN(P1_U2850) );
  INV_X1 U17877 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14488) );
  INV_X1 U17878 ( .A(n14693), .ZN(n14487) );
  OAI222_X1 U17879 ( .A1(n15838), .A2(n14523), .B1(n14488), .B2(n20103), .C1(
        n14487), .C2(n14524), .ZN(P1_U2851) );
  OAI222_X1 U17880 ( .A1(n14874), .A2(n14523), .B1(n14489), .B2(n20103), .C1(
        n14704), .C2(n14524), .ZN(P1_U2852) );
  OAI22_X1 U17881 ( .A1(n15967), .A2(n14523), .B1(n14490), .B2(n20103), .ZN(
        n14491) );
  INV_X1 U17882 ( .A(n14491), .ZN(n14492) );
  OAI21_X1 U17883 ( .B1(n14708), .B2(n14524), .A(n14492), .ZN(P1_U2853) );
  OAI22_X1 U17884 ( .A1(n15973), .A2(n14523), .B1(n14493), .B2(n20103), .ZN(
        n14494) );
  INV_X1 U17885 ( .A(n14494), .ZN(n14495) );
  OAI21_X1 U17886 ( .B1(n14721), .B2(n14524), .A(n14495), .ZN(P1_U2854) );
  INV_X1 U17887 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14503) );
  NAND2_X1 U17888 ( .A1(n14500), .A2(n14499), .ZN(n14501) );
  NAND2_X1 U17889 ( .A1(n14502), .A2(n14501), .ZN(n15871) );
  OAI222_X1 U17890 ( .A1(n15935), .A2(n14524), .B1(n14503), .B2(n20103), .C1(
        n15871), .C2(n14523), .ZN(P1_U2855) );
  INV_X1 U17891 ( .A(n14524), .ZN(n20099) );
  OAI22_X1 U17892 ( .A1(n15982), .A2(n14523), .B1(n14504), .B2(n20103), .ZN(
        n14505) );
  AOI21_X1 U17893 ( .B1(n14737), .B2(n20099), .A(n14505), .ZN(n14506) );
  INV_X1 U17894 ( .A(n14506), .ZN(P1_U2856) );
  OR2_X1 U17895 ( .A1(n14507), .A2(n14508), .ZN(n14509) );
  NAND2_X1 U17896 ( .A1(n15896), .A2(n20099), .ZN(n14513) );
  AND2_X1 U17897 ( .A1(n14521), .A2(n14510), .ZN(n14511) );
  NOR2_X1 U17898 ( .A1(n15881), .A2(n14511), .ZN(n16002) );
  NAND2_X1 U17899 ( .A1(n16002), .A2(n20098), .ZN(n14512) );
  OAI211_X1 U17900 ( .C1(n14514), .C2(n20103), .A(n14513), .B(n14512), .ZN(
        P1_U2858) );
  NOR2_X1 U17901 ( .A1(n13989), .A2(n14515), .ZN(n14516) );
  INV_X1 U17902 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15900) );
  INV_X1 U17903 ( .A(n14517), .ZN(n14519) );
  OAI21_X1 U17904 ( .B1(n14520), .B2(n14519), .A(n14518), .ZN(n14522) );
  NAND2_X1 U17905 ( .A1(n14522), .A2(n14521), .ZN(n15901) );
  OAI222_X1 U17906 ( .A1(n14752), .A2(n14524), .B1(n15900), .B2(n20103), .C1(
        n15901), .C2(n14523), .ZN(P1_U2859) );
  NAND3_X1 U17907 ( .A1(n14603), .A2(n20213), .A3(n14525), .ZN(n14586) );
  INV_X1 U17908 ( .A(DATAI_14_), .ZN(n20927) );
  MUX2_X1 U17909 ( .A(n20927), .B(n16446), .S(n14535), .Z(n20147) );
  OAI22_X1 U17910 ( .A1(n14586), .A2(n20147), .B1(n14603), .B2(n13275), .ZN(
        n14526) );
  AOI21_X1 U17911 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14588), .A(n14526), .ZN(
        n14528) );
  NAND2_X1 U17912 ( .A1(n14589), .A2(DATAI_30_), .ZN(n14527) );
  OAI211_X1 U17913 ( .C1(n14529), .C2(n14605), .A(n14528), .B(n14527), .ZN(
        P1_U2874) );
  INV_X1 U17914 ( .A(DATAI_29_), .ZN(n14534) );
  NAND2_X1 U17915 ( .A1(n14530), .A2(n14563), .ZN(n14533) );
  INV_X1 U17916 ( .A(DATAI_13_), .ZN(n20970) );
  MUX2_X1 U17917 ( .A(n20970), .B(n16448), .S(n14535), .Z(n20144) );
  OAI22_X1 U17918 ( .A1(n14586), .A2(n20144), .B1(n14603), .B2(n13270), .ZN(
        n14531) );
  AOI21_X1 U17919 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14588), .A(n14531), .ZN(
        n14532) );
  OAI211_X1 U17920 ( .C1(n14568), .C2(n14534), .A(n14533), .B(n14532), .ZN(
        P1_U2875) );
  INV_X1 U17921 ( .A(DATAI_12_), .ZN(n14536) );
  MUX2_X1 U17922 ( .A(n14536), .B(n16450), .S(n14535), .Z(n20141) );
  OAI22_X1 U17923 ( .A1(n14586), .A2(n20141), .B1(n14603), .B2(n14537), .ZN(
        n14538) );
  AOI21_X1 U17924 ( .B1(n14588), .B2(BUF1_REG_28__SCAN_IN), .A(n14538), .ZN(
        n14540) );
  NAND2_X1 U17925 ( .A1(n14589), .A2(DATAI_28_), .ZN(n14539) );
  OAI211_X1 U17926 ( .C1(n14627), .C2(n14605), .A(n14540), .B(n14539), .ZN(
        P1_U2876) );
  OAI22_X1 U17927 ( .A1(n14586), .A2(n14541), .B1(n14603), .B2(n12979), .ZN(
        n14542) );
  AOI21_X1 U17928 ( .B1(n14588), .B2(BUF1_REG_27__SCAN_IN), .A(n14542), .ZN(
        n14544) );
  NAND2_X1 U17929 ( .A1(n14589), .A2(DATAI_27_), .ZN(n14543) );
  OAI211_X1 U17930 ( .C1(n14638), .C2(n14605), .A(n14544), .B(n14543), .ZN(
        P1_U2877) );
  INV_X1 U17931 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20198) );
  INV_X1 U17932 ( .A(n14586), .ZN(n14571) );
  AOI22_X1 U17933 ( .A1(n14571), .A2(n20139), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n14569), .ZN(n14545) );
  OAI21_X1 U17934 ( .B1(n14573), .B2(n20198), .A(n14545), .ZN(n14546) );
  AOI21_X1 U17935 ( .B1(n14589), .B2(DATAI_26_), .A(n14546), .ZN(n14547) );
  OAI21_X1 U17936 ( .B1(n14650), .B2(n14605), .A(n14547), .ZN(P1_U2878) );
  INV_X1 U17937 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20190) );
  NOR2_X1 U17938 ( .A1(n14573), .A2(n20190), .ZN(n14550) );
  OAI22_X1 U17939 ( .A1(n14586), .A2(n20136), .B1(n14603), .B2(n14548), .ZN(
        n14549) );
  AOI211_X1 U17940 ( .C1(DATAI_25_), .C2(n14589), .A(n14550), .B(n14549), .ZN(
        n14551) );
  OAI21_X1 U17941 ( .B1(n14656), .B2(n14605), .A(n14551), .ZN(P1_U2879) );
  INV_X1 U17942 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20183) );
  AOI22_X1 U17943 ( .A1(n14571), .A2(n20134), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n14569), .ZN(n14552) );
  OAI21_X1 U17944 ( .B1(n14573), .B2(n20183), .A(n14552), .ZN(n14553) );
  AOI21_X1 U17945 ( .B1(n14589), .B2(DATAI_24_), .A(n14553), .ZN(n14554) );
  OAI21_X1 U17946 ( .B1(n14670), .B2(n14605), .A(n14554), .ZN(P1_U2880) );
  INV_X1 U17947 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20219) );
  AOI22_X1 U17948 ( .A1(n14571), .A2(n14555), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n14569), .ZN(n14556) );
  OAI21_X1 U17949 ( .B1(n14573), .B2(n20219), .A(n14556), .ZN(n14557) );
  AOI21_X1 U17950 ( .B1(n14589), .B2(DATAI_23_), .A(n14557), .ZN(n14558) );
  OAI21_X1 U17951 ( .B1(n14676), .B2(n14605), .A(n14558), .ZN(P1_U2881) );
  AOI22_X1 U17952 ( .A1(n14571), .A2(n14559), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n14569), .ZN(n14560) );
  OAI21_X1 U17953 ( .B1(n14573), .B2(n16435), .A(n14560), .ZN(n14561) );
  AOI21_X1 U17954 ( .B1(n14589), .B2(DATAI_22_), .A(n14561), .ZN(n14562) );
  OAI21_X1 U17955 ( .B1(n14686), .B2(n14605), .A(n14562), .ZN(P1_U2882) );
  INV_X1 U17956 ( .A(DATAI_21_), .ZN(n14567) );
  NAND2_X1 U17957 ( .A1(n14693), .A2(n14563), .ZN(n14566) );
  OAI22_X1 U17958 ( .A1(n14586), .A2(n20214), .B1(n14603), .B2(n12981), .ZN(
        n14564) );
  AOI21_X1 U17959 ( .B1(n14588), .B2(BUF1_REG_21__SCAN_IN), .A(n14564), .ZN(
        n14565) );
  OAI211_X1 U17960 ( .C1(n14568), .C2(n14567), .A(n14566), .B(n14565), .ZN(
        P1_U2883) );
  AOI22_X1 U17961 ( .A1(n14571), .A2(n14570), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n14569), .ZN(n14572) );
  OAI21_X1 U17962 ( .B1(n14573), .B2(n16438), .A(n14572), .ZN(n14574) );
  AOI21_X1 U17963 ( .B1(n14589), .B2(DATAI_20_), .A(n14574), .ZN(n14575) );
  OAI21_X1 U17964 ( .B1(n14704), .B2(n14605), .A(n14575), .ZN(P1_U2884) );
  OAI22_X1 U17965 ( .A1(n14586), .A2(n20206), .B1(n14603), .B2(n14576), .ZN(
        n14577) );
  AOI21_X1 U17966 ( .B1(n14588), .B2(BUF1_REG_19__SCAN_IN), .A(n14577), .ZN(
        n14579) );
  NAND2_X1 U17967 ( .A1(n14589), .A2(DATAI_19_), .ZN(n14578) );
  OAI211_X1 U17968 ( .C1(n14708), .C2(n14605), .A(n14579), .B(n14578), .ZN(
        P1_U2885) );
  OAI22_X1 U17969 ( .A1(n14586), .A2(n20199), .B1(n14603), .B2(n12969), .ZN(
        n14580) );
  AOI21_X1 U17970 ( .B1(n14588), .B2(BUF1_REG_18__SCAN_IN), .A(n14580), .ZN(
        n14582) );
  NAND2_X1 U17971 ( .A1(n14589), .A2(DATAI_18_), .ZN(n14581) );
  OAI211_X1 U17972 ( .C1(n14721), .C2(n14605), .A(n14582), .B(n14581), .ZN(
        P1_U2886) );
  OAI22_X1 U17973 ( .A1(n14586), .A2(n20193), .B1(n14603), .B2(n12972), .ZN(
        n14583) );
  AOI21_X1 U17974 ( .B1(n14588), .B2(BUF1_REG_17__SCAN_IN), .A(n14583), .ZN(
        n14585) );
  NAND2_X1 U17975 ( .A1(n14589), .A2(DATAI_17_), .ZN(n14584) );
  OAI211_X1 U17976 ( .C1(n15935), .C2(n14605), .A(n14585), .B(n14584), .ZN(
        P1_U2887) );
  INV_X1 U17977 ( .A(n14737), .ZN(n14592) );
  OAI22_X1 U17978 ( .A1(n14586), .A2(n20185), .B1(n14603), .B2(n12974), .ZN(
        n14587) );
  AOI21_X1 U17979 ( .B1(n14588), .B2(BUF1_REG_16__SCAN_IN), .A(n14587), .ZN(
        n14591) );
  NAND2_X1 U17980 ( .A1(n14589), .A2(DATAI_16_), .ZN(n14590) );
  OAI211_X1 U17981 ( .C1(n14592), .C2(n14605), .A(n14591), .B(n14590), .ZN(
        P1_U2888) );
  INV_X1 U17982 ( .A(n14593), .ZN(n14594) );
  INV_X1 U17983 ( .A(n15945), .ZN(n14598) );
  OAI222_X1 U17984 ( .A1(n14605), .A2(n14598), .B1(n14603), .B2(n13040), .C1(
        n14602), .C2(n14597), .ZN(P1_U2889) );
  INV_X1 U17985 ( .A(n15896), .ZN(n14600) );
  INV_X1 U17986 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14599) );
  OAI222_X1 U17987 ( .A1(n14600), .A2(n14605), .B1(n14599), .B2(n14603), .C1(
        n14602), .C2(n20147), .ZN(P1_U2890) );
  INV_X1 U17988 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14601) );
  OAI222_X1 U17989 ( .A1(n14752), .A2(n14605), .B1(n14601), .B2(n14603), .C1(
        n14602), .C2(n20144), .ZN(P1_U2891) );
  INV_X1 U17990 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14604) );
  OAI222_X1 U17991 ( .A1(n14764), .A2(n14605), .B1(n14604), .B2(n14603), .C1(
        n14602), .C2(n20141), .ZN(P1_U2892) );
  XNOR2_X1 U17992 ( .A(n9971), .B(n14606), .ZN(n14607) );
  XNOR2_X1 U17993 ( .A(n14608), .B(n14607), .ZN(n14787) );
  NAND2_X1 U17994 ( .A1(n9645), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14789) );
  NAND2_X1 U17995 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14609) );
  OAI211_X1 U17996 ( .C1(n14610), .C2(n15963), .A(n14789), .B(n14609), .ZN(
        n14611) );
  AOI21_X1 U17997 ( .B1(n14787), .B2(n15959), .A(n14611), .ZN(n14612) );
  OAI21_X1 U17998 ( .B1(n14613), .B2(n15934), .A(n14612), .ZN(P1_U2970) );
  NAND2_X1 U17999 ( .A1(n9971), .A2(n11252), .ZN(n14639) );
  NAND2_X1 U18000 ( .A1(n14614), .A2(n14639), .ZN(n14620) );
  INV_X1 U18001 ( .A(n14616), .ZN(n14617) );
  OAI21_X1 U18002 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14617), .A(
        n14620), .ZN(n14619) );
  MUX2_X1 U18003 ( .A(n14812), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9971), .Z(n14618) );
  OAI211_X1 U18004 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14620), .A(
        n14619), .B(n14618), .ZN(n14621) );
  XNOR2_X1 U18005 ( .A(n14621), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14796) );
  NAND2_X1 U18006 ( .A1(n14622), .A2(n15950), .ZN(n14623) );
  NAND2_X1 U18007 ( .A1(n9645), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14797) );
  OAI211_X1 U18008 ( .C1(n14772), .C2(n14624), .A(n14623), .B(n14797), .ZN(
        n14625) );
  AOI21_X1 U18009 ( .B1(n14796), .B2(n15959), .A(n14625), .ZN(n14626) );
  OAI21_X1 U18010 ( .B1(n14627), .B2(n15934), .A(n14626), .ZN(P1_U2971) );
  NAND3_X1 U18011 ( .A1(n14628), .A2(n9648), .A3(n14837), .ZN(n14663) );
  NOR2_X1 U18012 ( .A1(n14663), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14652) );
  NAND2_X1 U18013 ( .A1(n14652), .A2(n14830), .ZN(n14631) );
  NAND2_X1 U18014 ( .A1(n14653), .A2(n9971), .ZN(n14629) );
  OAI22_X1 U18015 ( .A1(n14632), .A2(n14631), .B1(n14630), .B2(n14629), .ZN(
        n14633) );
  XNOR2_X1 U18016 ( .A(n14633), .B(n14812), .ZN(n14815) );
  NAND2_X1 U18017 ( .A1(n9645), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14807) );
  NAND2_X1 U18018 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14634) );
  OAI211_X1 U18019 ( .C1(n14635), .C2(n15963), .A(n14807), .B(n14634), .ZN(
        n14636) );
  AOI21_X1 U18020 ( .B1(n14815), .B2(n15959), .A(n14636), .ZN(n14637) );
  OAI21_X1 U18021 ( .B1(n14638), .B2(n15934), .A(n14637), .ZN(P1_U2972) );
  INV_X1 U18022 ( .A(n14639), .ZN(n14641) );
  AOI211_X1 U18023 ( .C1(n9648), .C2(n14642), .A(n14641), .B(n14640), .ZN(
        n14644) );
  XNOR2_X1 U18024 ( .A(n14644), .B(n14643), .ZN(n14817) );
  NAND2_X1 U18025 ( .A1(n14645), .A2(n15950), .ZN(n14646) );
  NAND2_X1 U18026 ( .A1(n9645), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14818) );
  OAI211_X1 U18027 ( .C1(n14772), .C2(n14647), .A(n14646), .B(n14818), .ZN(
        n14648) );
  AOI21_X1 U18028 ( .B1(n14817), .B2(n15959), .A(n14648), .ZN(n14649) );
  OAI21_X1 U18029 ( .B1(n14650), .B2(n15934), .A(n14649), .ZN(P1_U2973) );
  AND2_X1 U18030 ( .A1(n9971), .A2(n14651), .ZN(n14654) );
  AOI21_X1 U18031 ( .B1(n14654), .B2(n14653), .A(n14652), .ZN(n14655) );
  XNOR2_X1 U18032 ( .A(n14655), .B(n14830), .ZN(n14834) );
  INV_X1 U18033 ( .A(n14656), .ZN(n14660) );
  AND2_X1 U18034 ( .A1(n9645), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14825) );
  AOI21_X1 U18035 ( .B1(n15948), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14825), .ZN(n14657) );
  OAI21_X1 U18036 ( .B1(n14658), .B2(n15963), .A(n14657), .ZN(n14659) );
  AOI21_X1 U18037 ( .B1(n14660), .B2(n15960), .A(n14659), .ZN(n14661) );
  OAI21_X1 U18038 ( .B1(n14834), .B2(n20007), .A(n14661), .ZN(P1_U2974) );
  NAND3_X1 U18039 ( .A1(n14614), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n9971), .ZN(n14662) );
  NAND2_X1 U18040 ( .A1(n14663), .A2(n14662), .ZN(n14664) );
  XNOR2_X1 U18041 ( .A(n14664), .B(n14835), .ZN(n14836) );
  NAND2_X1 U18042 ( .A1(n14665), .A2(n15950), .ZN(n14666) );
  NAND2_X1 U18043 ( .A1(n9645), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14842) );
  OAI211_X1 U18044 ( .C1(n14772), .C2(n14667), .A(n14666), .B(n14842), .ZN(
        n14668) );
  AOI21_X1 U18045 ( .B1(n14836), .B2(n15959), .A(n14668), .ZN(n14669) );
  OAI21_X1 U18046 ( .B1(n14670), .B2(n15934), .A(n14669), .ZN(P1_U2975) );
  XNOR2_X1 U18047 ( .A(n9971), .B(n14837), .ZN(n14671) );
  XNOR2_X1 U18048 ( .A(n14614), .B(n14671), .ZN(n14849) );
  NOR2_X1 U18049 ( .A1(n20073), .A2(n20960), .ZN(n14852) );
  AOI21_X1 U18050 ( .B1(n15948), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14852), .ZN(n14672) );
  OAI21_X1 U18051 ( .B1(n14673), .B2(n15963), .A(n14672), .ZN(n14674) );
  AOI21_X1 U18052 ( .B1(n14849), .B2(n15959), .A(n14674), .ZN(n14675) );
  OAI21_X1 U18053 ( .B1(n14676), .B2(n15934), .A(n14675), .ZN(P1_U2976) );
  INV_X1 U18054 ( .A(n14688), .ZN(n14677) );
  AOI21_X1 U18055 ( .B1(n14677), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n9972), .ZN(n14678) );
  NOR2_X1 U18056 ( .A1(n14678), .A2(n9969), .ZN(n14680) );
  XNOR2_X1 U18057 ( .A(n14680), .B(n14679), .ZN(n14857) );
  INV_X1 U18058 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14683) );
  NAND2_X1 U18059 ( .A1(n15950), .A2(n14681), .ZN(n14682) );
  NAND2_X1 U18060 ( .A1(n9645), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14859) );
  OAI211_X1 U18061 ( .C1(n14772), .C2(n14683), .A(n14682), .B(n14859), .ZN(
        n14684) );
  AOI21_X1 U18062 ( .B1(n14857), .B2(n15959), .A(n14684), .ZN(n14685) );
  OAI21_X1 U18063 ( .B1(n14686), .B2(n15934), .A(n14685), .ZN(P1_U2977) );
  NAND3_X1 U18064 ( .A1(n11251), .A2(n9648), .A3(n14687), .ZN(n14695) );
  OAI22_X1 U18065 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14695), .B1(
        n14688), .B2(n9648), .ZN(n14689) );
  XNOR2_X1 U18066 ( .A(n14689), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15837) );
  AOI22_X1 U18067 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n9645), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n14690) );
  OAI21_X1 U18068 ( .B1(n15963), .B2(n14691), .A(n14690), .ZN(n14692) );
  AOI21_X1 U18069 ( .B1(n14693), .B2(n15960), .A(n14692), .ZN(n14694) );
  OAI21_X1 U18070 ( .B1(n15837), .B2(n20007), .A(n14694), .ZN(P1_U2978) );
  NAND2_X1 U18071 ( .A1(n9971), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14696) );
  OAI21_X1 U18072 ( .B1(n14715), .B2(n14696), .A(n14695), .ZN(n14698) );
  XNOR2_X1 U18073 ( .A(n14698), .B(n14697), .ZN(n14866) );
  INV_X1 U18074 ( .A(n14699), .ZN(n14701) );
  AOI22_X1 U18075 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n9645), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n14700) );
  OAI21_X1 U18076 ( .B1(n15963), .B2(n14701), .A(n14700), .ZN(n14702) );
  AOI21_X1 U18077 ( .B1(n14866), .B2(n15959), .A(n14702), .ZN(n14703) );
  OAI21_X1 U18078 ( .B1(n14704), .B2(n15934), .A(n14703), .ZN(P1_U2979) );
  NOR2_X1 U18079 ( .A1(n9971), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14706) );
  MUX2_X1 U18080 ( .A(n9971), .B(n14706), .S(n14715), .Z(n14707) );
  XNOR2_X1 U18081 ( .A(n14707), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15964) );
  INV_X1 U18082 ( .A(n14708), .ZN(n14712) );
  AOI22_X1 U18083 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n9645), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14709) );
  OAI21_X1 U18084 ( .B1(n15963), .B2(n14710), .A(n14709), .ZN(n14711) );
  AOI21_X1 U18085 ( .B1(n14712), .B2(n15960), .A(n14711), .ZN(n14713) );
  OAI21_X1 U18086 ( .B1(n20007), .B2(n15964), .A(n14713), .ZN(P1_U2980) );
  OAI22_X1 U18087 ( .A1(n14772), .A2(n14714), .B1(n20073), .B2(n20770), .ZN(
        n14718) );
  OAI21_X1 U18088 ( .B1(n11250), .B2(n14716), .A(n14715), .ZN(n15974) );
  NOR2_X1 U18089 ( .A1(n15974), .A2(n20007), .ZN(n14717) );
  AOI211_X1 U18090 ( .C1(n15950), .C2(n14719), .A(n14718), .B(n14717), .ZN(
        n14720) );
  OAI21_X1 U18091 ( .B1(n14721), .B2(n15934), .A(n14720), .ZN(P1_U2981) );
  OR2_X1 U18092 ( .A1(n14722), .A2(n14723), .ZN(n14727) );
  INV_X1 U18093 ( .A(n14724), .ZN(n14725) );
  AND2_X1 U18094 ( .A1(n14725), .A2(n14739), .ZN(n14726) );
  NAND2_X1 U18095 ( .A1(n14727), .A2(n14726), .ZN(n15941) );
  INV_X1 U18096 ( .A(n14730), .ZN(n14729) );
  OR2_X1 U18097 ( .A1(n14729), .A2(n14728), .ZN(n15940) );
  NAND2_X1 U18098 ( .A1(n15943), .A2(n14730), .ZN(n14731) );
  XOR2_X1 U18099 ( .A(n14732), .B(n14731), .Z(n15981) );
  INV_X1 U18100 ( .A(n14733), .ZN(n14735) );
  AOI22_X1 U18101 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n9645), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14734) );
  OAI21_X1 U18102 ( .B1(n15963), .B2(n14735), .A(n14734), .ZN(n14736) );
  AOI21_X1 U18103 ( .B1(n14737), .B2(n15960), .A(n14736), .ZN(n14738) );
  OAI21_X1 U18104 ( .B1(n20007), .B2(n15981), .A(n14738), .ZN(P1_U2983) );
  MUX2_X1 U18105 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n16000), .S(
        n9971), .Z(n14744) );
  INV_X1 U18106 ( .A(n14739), .ZN(n14749) );
  OAI21_X1 U18107 ( .B1(n14883), .B2(n14749), .A(n14740), .ZN(n14742) );
  NAND2_X1 U18108 ( .A1(n14742), .A2(n14741), .ZN(n14743) );
  XOR2_X1 U18109 ( .A(n14744), .B(n14743), .Z(n16003) );
  AND2_X1 U18110 ( .A1(n9645), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16001) );
  AOI21_X1 U18111 ( .B1(n15948), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16001), .ZN(n14745) );
  OAI21_X1 U18112 ( .B1(n15963), .B2(n15890), .A(n14745), .ZN(n14746) );
  AOI21_X1 U18113 ( .B1(n15896), .B2(n15960), .A(n14746), .ZN(n14747) );
  OAI21_X1 U18114 ( .B1(n16003), .B2(n20007), .A(n14747), .ZN(P1_U2985) );
  AND2_X1 U18115 ( .A1(n14883), .A2(n14748), .ZN(n14759) );
  OAI21_X1 U18116 ( .B1(n14759), .B2(n14749), .A(n14760), .ZN(n14751) );
  XNOR2_X1 U18117 ( .A(n14751), .B(n14750), .ZN(n14911) );
  INV_X1 U18118 ( .A(n14752), .ZN(n15905) );
  INV_X1 U18119 ( .A(n14753), .ZN(n15902) );
  AOI22_X1 U18120 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n9645), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14754) );
  OAI21_X1 U18121 ( .B1(n15963), .B2(n15902), .A(n14754), .ZN(n14755) );
  AOI21_X1 U18122 ( .B1(n15905), .B2(n15960), .A(n14755), .ZN(n14756) );
  OAI21_X1 U18123 ( .B1(n14911), .B2(n20007), .A(n14756), .ZN(P1_U2986) );
  INV_X1 U18124 ( .A(n14757), .ZN(n14758) );
  NOR2_X1 U18125 ( .A1(n14759), .A2(n14758), .ZN(n14763) );
  NAND2_X1 U18126 ( .A1(n14761), .A2(n14760), .ZN(n14762) );
  XNOR2_X1 U18127 ( .A(n14763), .B(n14762), .ZN(n14928) );
  INV_X1 U18128 ( .A(n14764), .ZN(n14768) );
  AND2_X1 U18129 ( .A1(n9645), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14925) );
  AOI21_X1 U18130 ( .B1(n15948), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n14925), .ZN(n14765) );
  OAI21_X1 U18131 ( .B1(n15963), .B2(n14766), .A(n14765), .ZN(n14767) );
  AOI21_X1 U18132 ( .B1(n14768), .B2(n15960), .A(n14767), .ZN(n14769) );
  OAI21_X1 U18133 ( .B1(n14928), .B2(n20007), .A(n14769), .ZN(P1_U2987) );
  NAND2_X1 U18134 ( .A1(n9648), .A2(n14930), .ZN(n14770) );
  NAND3_X1 U18135 ( .A1(n14883), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9971), .ZN(n14933) );
  OAI21_X1 U18136 ( .B1(n14929), .B2(n14770), .A(n14933), .ZN(n14771) );
  XNOR2_X1 U18137 ( .A(n14771), .B(n14919), .ZN(n16013) );
  NAND2_X1 U18138 ( .A1(n16013), .A2(n15959), .ZN(n14775) );
  NAND2_X1 U18139 ( .A1(n9645), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n16009) );
  OAI21_X1 U18140 ( .B1(n14772), .B2(n15912), .A(n16009), .ZN(n14773) );
  AOI21_X1 U18141 ( .B1(n15950), .B2(n15918), .A(n14773), .ZN(n14774) );
  OAI211_X1 U18142 ( .C1(n15934), .C2(n15915), .A(n14775), .B(n14774), .ZN(
        P1_U2988) );
  INV_X1 U18143 ( .A(n14776), .ZN(n14779) );
  INV_X1 U18144 ( .A(n14777), .ZN(n14778) );
  AOI21_X1 U18145 ( .B1(n14779), .B2(n16032), .A(n14778), .ZN(n14784) );
  INV_X1 U18146 ( .A(n14780), .ZN(n14782) );
  OAI211_X1 U18147 ( .C1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n14786), .A(
        n14782), .B(n14781), .ZN(n14783) );
  OAI211_X1 U18148 ( .C1(n14785), .C2(n20164), .A(n14784), .B(n14783), .ZN(
        P1_U3001) );
  INV_X1 U18149 ( .A(n14786), .ZN(n14795) );
  NAND2_X1 U18150 ( .A1(n14787), .A2(n16033), .ZN(n14794) );
  NAND2_X1 U18151 ( .A1(n14788), .A2(n16032), .ZN(n14790) );
  NAND2_X1 U18152 ( .A1(n14790), .A2(n14789), .ZN(n14791) );
  AOI21_X1 U18153 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14792), .A(
        n14791), .ZN(n14793) );
  OAI211_X1 U18154 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14795), .A(
        n14794), .B(n14793), .ZN(P1_U3002) );
  INV_X1 U18155 ( .A(n14796), .ZN(n14805) );
  INV_X1 U18156 ( .A(n14813), .ZN(n14800) );
  OAI21_X1 U18157 ( .B1(n14798), .B2(n20173), .A(n14797), .ZN(n14799) );
  AOI21_X1 U18158 ( .B1(n14800), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14799), .ZN(n14804) );
  NAND3_X1 U18159 ( .A1(n14806), .A2(n14802), .A3(n14801), .ZN(n14803) );
  OAI211_X1 U18160 ( .C1(n14805), .C2(n20164), .A(n14804), .B(n14803), .ZN(
        P1_U3003) );
  NAND2_X1 U18161 ( .A1(n14806), .A2(n14812), .ZN(n14811) );
  INV_X1 U18162 ( .A(n14807), .ZN(n14808) );
  AOI21_X1 U18163 ( .B1(n14809), .B2(n16032), .A(n14808), .ZN(n14810) );
  OAI211_X1 U18164 ( .C1(n14813), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        n14814) );
  AOI21_X1 U18165 ( .B1(n14815), .B2(n16033), .A(n14814), .ZN(n14816) );
  INV_X1 U18166 ( .A(n14816), .ZN(P1_U3004) );
  INV_X1 U18167 ( .A(n14831), .ZN(n14824) );
  XNOR2_X1 U18168 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14823) );
  NAND2_X1 U18169 ( .A1(n14817), .A2(n16033), .ZN(n14822) );
  OAI21_X1 U18170 ( .B1(n14819), .B2(n20173), .A(n14818), .ZN(n14820) );
  AOI21_X1 U18171 ( .B1(n14829), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14820), .ZN(n14821) );
  OAI211_X1 U18172 ( .C1(n14824), .C2(n14823), .A(n14822), .B(n14821), .ZN(
        P1_U3005) );
  INV_X1 U18173 ( .A(n14825), .ZN(n14826) );
  OAI21_X1 U18174 ( .B1(n14827), .B2(n20173), .A(n14826), .ZN(n14828) );
  AOI21_X1 U18175 ( .B1(n14829), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14828), .ZN(n14833) );
  NAND2_X1 U18176 ( .A1(n14831), .A2(n14830), .ZN(n14832) );
  OAI211_X1 U18177 ( .C1(n14834), .C2(n20164), .A(n14833), .B(n14832), .ZN(
        P1_U3006) );
  NAND2_X1 U18178 ( .A1(n14835), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14848) );
  NAND2_X1 U18179 ( .A1(n14836), .A2(n16033), .ZN(n14847) );
  NAND2_X1 U18180 ( .A1(n14838), .A2(n14837), .ZN(n14839) );
  NAND2_X1 U18181 ( .A1(n14840), .A2(n14839), .ZN(n14845) );
  NAND2_X1 U18182 ( .A1(n14841), .A2(n16032), .ZN(n14843) );
  NAND2_X1 U18183 ( .A1(n14843), .A2(n14842), .ZN(n14844) );
  AOI21_X1 U18184 ( .B1(n14845), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14844), .ZN(n14846) );
  OAI211_X1 U18185 ( .C1(n14856), .C2(n14848), .A(n14847), .B(n14846), .ZN(
        P1_U3007) );
  NAND2_X1 U18186 ( .A1(n14849), .A2(n16033), .ZN(n14855) );
  NOR2_X1 U18187 ( .A1(n14850), .A2(n20173), .ZN(n14851) );
  AOI211_X1 U18188 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14853), .A(
        n14852), .B(n14851), .ZN(n14854) );
  OAI211_X1 U18189 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14856), .A(
        n14855), .B(n14854), .ZN(P1_U3008) );
  INV_X1 U18190 ( .A(n14857), .ZN(n14865) );
  INV_X1 U18191 ( .A(n14858), .ZN(n14860) );
  OAI21_X1 U18192 ( .B1(n14860), .B2(n20173), .A(n14859), .ZN(n14861) );
  AOI21_X1 U18193 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15834), .A(
        n14861), .ZN(n14864) );
  OAI211_X1 U18194 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15836), .B(n14862), .ZN(
        n14863) );
  OAI211_X1 U18195 ( .C1(n14865), .C2(n20164), .A(n14864), .B(n14863), .ZN(
        P1_U3009) );
  NAND2_X1 U18196 ( .A1(n14866), .A2(n16033), .ZN(n14879) );
  NOR2_X1 U18197 ( .A1(n20166), .A2(n14892), .ZN(n14868) );
  AOI21_X1 U18198 ( .B1(n14903), .B2(n14868), .A(n14867), .ZN(n14900) );
  NAND2_X1 U18199 ( .A1(n14869), .A2(n15966), .ZN(n15971) );
  OAI21_X1 U18200 ( .B1(n14870), .B2(n15966), .A(n14913), .ZN(n14871) );
  INV_X1 U18201 ( .A(n14871), .ZN(n14872) );
  AOI211_X1 U18202 ( .C1(n14916), .C2(n14873), .A(n14894), .B(n14872), .ZN(
        n15965) );
  OAI21_X1 U18203 ( .B1(n14900), .B2(n15971), .A(n15965), .ZN(n14877) );
  INV_X1 U18204 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20884) );
  NOR2_X1 U18205 ( .A1(n20073), .A2(n20884), .ZN(n14876) );
  NOR2_X1 U18206 ( .A1(n14874), .A2(n20173), .ZN(n14875) );
  AOI211_X1 U18207 ( .C1(n14877), .C2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14876), .B(n14875), .ZN(n14878) );
  OAI211_X1 U18208 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n14880), .A(
        n14879), .B(n14878), .ZN(P1_U3011) );
  OAI21_X1 U18209 ( .B1(n14883), .B2(n14882), .A(n14881), .ZN(n14886) );
  NAND2_X1 U18210 ( .A1(n14886), .A2(n15987), .ZN(n14885) );
  MUX2_X1 U18211 ( .A(n14886), .B(n14885), .S(n9648), .Z(n14887) );
  XNOR2_X1 U18212 ( .A(n14887), .B(n14888), .ZN(n15939) );
  OAI21_X1 U18213 ( .B1(n15984), .B2(n14889), .A(n14888), .ZN(n14898) );
  AOI21_X1 U18214 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14903), .A(
        n14890), .ZN(n14902) );
  OAI22_X1 U18215 ( .A1(n14903), .A2(n14892), .B1(n14891), .B2(n20168), .ZN(
        n14893) );
  NOR3_X1 U18216 ( .A1(n14902), .A2(n14894), .A3(n14893), .ZN(n14908) );
  OAI21_X1 U18217 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14900), .A(
        n14908), .ZN(n16004) );
  AOI21_X1 U18218 ( .B1(n16000), .B2(n14895), .A(n16004), .ZN(n15997) );
  OAI21_X1 U18219 ( .B1(n14939), .B2(n15978), .A(n15997), .ZN(n15976) );
  INV_X1 U18220 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14896) );
  OAI22_X1 U18221 ( .A1(n15871), .A2(n20173), .B1(n20073), .B2(n14896), .ZN(
        n14897) );
  AOI21_X1 U18222 ( .B1(n14898), .B2(n15976), .A(n14897), .ZN(n14899) );
  OAI21_X1 U18223 ( .B1(n15939), .B2(n20164), .A(n14899), .ZN(P1_U3014) );
  NOR2_X1 U18224 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14900), .ZN(
        n14906) );
  AND2_X1 U18225 ( .A1(n9645), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n14901) );
  AOI21_X1 U18226 ( .B1(n14903), .B2(n14902), .A(n14901), .ZN(n14904) );
  OAI21_X1 U18227 ( .B1(n15901), .B2(n20173), .A(n14904), .ZN(n14905) );
  NOR2_X1 U18228 ( .A1(n14906), .A2(n14905), .ZN(n14910) );
  OR2_X1 U18229 ( .A1(n14908), .A2(n14907), .ZN(n14909) );
  OAI211_X1 U18230 ( .C1(n14911), .C2(n20164), .A(n14910), .B(n14909), .ZN(
        P1_U3018) );
  NOR2_X1 U18231 ( .A1(n14912), .A2(n14915), .ZN(n14923) );
  AOI22_X1 U18232 ( .A1(n14916), .A2(n14915), .B1(n14914), .B2(n14913), .ZN(
        n14917) );
  NAND2_X1 U18233 ( .A1(n14918), .A2(n14917), .ZN(n16012) );
  AOI21_X1 U18234 ( .B1(n14920), .B2(n14919), .A(n16012), .ZN(n14921) );
  INV_X1 U18235 ( .A(n14921), .ZN(n14922) );
  MUX2_X1 U18236 ( .A(n14923), .B(n14922), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n14924) );
  AOI211_X1 U18237 ( .C1(n16032), .C2(n14926), .A(n14925), .B(n14924), .ZN(
        n14927) );
  OAI21_X1 U18238 ( .B1(n14928), .B2(n20164), .A(n14927), .ZN(P1_U3019) );
  XNOR2_X1 U18239 ( .A(n14929), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14932) );
  NAND2_X1 U18240 ( .A1(n14722), .A2(n14930), .ZN(n14931) );
  MUX2_X1 U18241 ( .A(n14932), .B(n14931), .S(n9971), .Z(n14934) );
  NAND2_X1 U18242 ( .A1(n14934), .A2(n14933), .ZN(n15954) );
  NOR2_X1 U18243 ( .A1(n14936), .A2(n14935), .ZN(n16019) );
  OAI211_X1 U18244 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16019), .B(n14937), .ZN(n14942) );
  OAI21_X1 U18245 ( .B1(n14939), .B2(n14938), .A(n20179), .ZN(n16017) );
  INV_X1 U18246 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15929) );
  OAI22_X1 U18247 ( .A1(n15922), .A2(n20173), .B1(n15929), .B2(n20073), .ZN(
        n14940) );
  AOI21_X1 U18248 ( .B1(n16017), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n14940), .ZN(n14941) );
  OAI211_X1 U18249 ( .C1(n15954), .C2(n20164), .A(n14942), .B(n14941), .ZN(
        P1_U3021) );
  INV_X1 U18250 ( .A(n14943), .ZN(n20820) );
  NAND2_X1 U18251 ( .A1(n20974), .A2(n20671), .ZN(n20484) );
  MUX2_X1 U18252 ( .A(n20820), .B(n20484), .S(n9656), .Z(n14944) );
  OAI21_X1 U18253 ( .B1(n14947), .B2(n9637), .A(n14944), .ZN(n14945) );
  MUX2_X1 U18254 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14945), .S(
        n20823), .Z(P1_U3477) );
  AND2_X1 U18255 ( .A1(n9656), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20523) );
  AOI21_X1 U18256 ( .B1(n13507), .B2(n20523), .A(n20664), .ZN(n20668) );
  OAI21_X1 U18257 ( .B1(n11172), .B2(n20523), .A(n20668), .ZN(n14946) );
  OAI21_X1 U18258 ( .B1(n14947), .B2(n13095), .A(n14946), .ZN(n14948) );
  MUX2_X1 U18259 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14948), .S(
        n20823), .Z(P1_U3476) );
  OAI21_X1 U18260 ( .B1(n9771), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14953), .ZN(n14954) );
  INV_X1 U18261 ( .A(n14954), .ZN(n16059) );
  AOI21_X1 U18262 ( .B1(n15198), .B2(n14955), .A(n9771), .ZN(n15205) );
  NOR2_X1 U18263 ( .A1(n15205), .A2(n14980), .ZN(n14979) );
  NOR2_X1 U18264 ( .A1(n19021), .A2(n14979), .ZN(n16060) );
  XNOR2_X1 U18265 ( .A(n14953), .B(n15178), .ZN(n16050) );
  NAND4_X1 U18266 ( .A1(n16058), .A2(n9634), .A3(n19089), .A4(n16050), .ZN(
        n14978) );
  NAND2_X1 U18267 ( .A1(n11966), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14963) );
  NAND2_X1 U18268 ( .A1(n12008), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14962) );
  NAND2_X1 U18269 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14961) );
  NAND2_X1 U18270 ( .A1(n14959), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14960) );
  NAND4_X1 U18271 ( .A1(n14963), .A2(n14962), .A3(n14961), .A4(n14960), .ZN(
        n14964) );
  INV_X1 U18272 ( .A(n16098), .ZN(n14976) );
  INV_X1 U18273 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19921) );
  OAI22_X1 U18274 ( .A1(n12594), .A2(n19093), .B1(n19921), .B2(n19067), .ZN(
        n14975) );
  NAND2_X1 U18275 ( .A1(n14967), .A2(n14966), .ZN(n14972) );
  NAND2_X1 U18276 ( .A1(n14968), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14970) );
  AOI22_X1 U18277 ( .A1(n12211), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12115), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14969) );
  AND2_X1 U18278 ( .A1(n14970), .A2(n14969), .ZN(n14971) );
  OAI22_X1 U18279 ( .A1(n19149), .A2(n19098), .B1(n12661), .B2(n14973), .ZN(
        n14974) );
  AOI211_X1 U18280 ( .C1(n14976), .C2(n19076), .A(n14975), .B(n14974), .ZN(
        n14977) );
  OAI211_X1 U18281 ( .C1(n15159), .C2(n19099), .A(n14978), .B(n14977), .ZN(
        P2_U2824) );
  AOI21_X1 U18282 ( .B1(n14980), .B2(n15205), .A(n14979), .ZN(n14981) );
  NAND2_X1 U18283 ( .A1(n14981), .A2(n19089), .ZN(n14994) );
  NAND2_X1 U18284 ( .A1(n14983), .A2(n14982), .ZN(n14984) );
  NAND2_X1 U18285 ( .A1(n14987), .A2(n14986), .ZN(n14988) );
  NAND2_X1 U18286 ( .A1(n14989), .A2(n14988), .ZN(n15090) );
  AOI22_X1 U18287 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19095), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19102), .ZN(n14991) );
  NAND2_X1 U18288 ( .A1(n19096), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14990) );
  OAI211_X1 U18289 ( .C1(n15090), .C2(n19098), .A(n14991), .B(n14990), .ZN(
        n14992) );
  AOI21_X1 U18290 ( .B1(n15325), .B2(n19076), .A(n14992), .ZN(n14993) );
  OAI211_X1 U18291 ( .C1(n14995), .C2(n19099), .A(n14994), .B(n14993), .ZN(
        P2_U2827) );
  AOI211_X1 U18292 ( .C1(n14998), .C2(n14996), .A(n14997), .B(n19851), .ZN(
        n14999) );
  INV_X1 U18293 ( .A(n14999), .ZN(n15009) );
  OR2_X1 U18294 ( .A1(n15011), .A2(n15000), .ZN(n15001) );
  AND2_X1 U18295 ( .A1(n9711), .A2(n15001), .ZN(n15383) );
  NAND2_X1 U18296 ( .A1(n15002), .A2(n15003), .ZN(n15004) );
  NAND2_X1 U18297 ( .A1(n15112), .A2(n15004), .ZN(n15386) );
  NAND2_X1 U18298 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19096), .ZN(n15006) );
  AOI22_X1 U18299 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19095), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19102), .ZN(n15005) );
  OAI211_X1 U18300 ( .C1(n19098), .C2(n15386), .A(n15006), .B(n15005), .ZN(
        n15007) );
  AOI21_X1 U18301 ( .B1(n15383), .B2(n19076), .A(n15007), .ZN(n15008) );
  OAI211_X1 U18302 ( .C1(n15010), .C2(n19099), .A(n15009), .B(n15008), .ZN(
        P2_U2831) );
  INV_X1 U18303 ( .A(n15413), .ZN(n15012) );
  AOI21_X1 U18304 ( .B1(n9773), .B2(n15012), .A(n15011), .ZN(n16143) );
  INV_X1 U18305 ( .A(n16143), .ZN(n15018) );
  OR2_X1 U18306 ( .A1(n15418), .A2(n15013), .ZN(n15014) );
  NAND2_X1 U18307 ( .A1(n15002), .A2(n15014), .ZN(n15401) );
  AOI22_X1 U18308 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19095), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19102), .ZN(n15015) );
  OAI21_X1 U18309 ( .B1(n19098), .B2(n15401), .A(n15015), .ZN(n15016) );
  AOI21_X1 U18310 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n19096), .A(n15016), .ZN(
        n15017) );
  OAI21_X1 U18311 ( .B1(n15018), .B2(n19107), .A(n15017), .ZN(n15022) );
  AOI211_X1 U18312 ( .C1(n16142), .C2(n15020), .A(n15019), .B(n19851), .ZN(
        n15021) );
  AOI211_X1 U18313 ( .C1(n19056), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        n15024) );
  INV_X1 U18314 ( .A(n15024), .ZN(P2_U2832) );
  NAND2_X1 U18315 ( .A1(n9634), .A2(n15025), .ZN(n15026) );
  XOR2_X1 U18316 ( .A(n16192), .B(n15026), .Z(n15027) );
  NAND2_X1 U18317 ( .A1(n15027), .A2(n19089), .ZN(n15045) );
  INV_X1 U18318 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n19130) );
  INV_X1 U18319 ( .A(n15028), .ZN(n15029) );
  AOI22_X1 U18320 ( .A1(n19056), .A2(n15029), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19095), .ZN(n15030) );
  OAI21_X1 U18321 ( .B1(n19082), .B2(n19130), .A(n15030), .ZN(n15031) );
  AOI211_X1 U18322 ( .C1(n19102), .C2(P2_REIP_REG_12__SCAN_IN), .A(n15785), 
        .B(n15031), .ZN(n15044) );
  NAND2_X1 U18323 ( .A1(n15033), .A2(n15032), .ZN(n15034) );
  AND2_X1 U18324 ( .A1(n15035), .A2(n15034), .ZN(n19126) );
  NAND2_X1 U18325 ( .A1(n19126), .A2(n19076), .ZN(n15043) );
  INV_X1 U18326 ( .A(n15036), .ZN(n15037) );
  OR2_X1 U18327 ( .A1(n15038), .A2(n15037), .ZN(n15041) );
  INV_X1 U18328 ( .A(n15039), .ZN(n15040) );
  NAND2_X1 U18329 ( .A1(n18973), .A2(n19156), .ZN(n15042) );
  NAND4_X1 U18330 ( .A1(n15045), .A2(n15044), .A3(n15043), .A4(n15042), .ZN(
        P2_U2843) );
  NAND2_X1 U18331 ( .A1(n15047), .A2(n15046), .ZN(n15049) );
  XNOR2_X1 U18332 ( .A(n15049), .B(n15048), .ZN(n15095) );
  NAND2_X1 U18333 ( .A1(n12991), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15051) );
  NAND2_X1 U18334 ( .A1(n15325), .A2(n19148), .ZN(n15050) );
  OAI211_X1 U18335 ( .C1(n15095), .C2(n19145), .A(n15051), .B(n15050), .ZN(
        P2_U2859) );
  AOI21_X1 U18336 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(n15096) );
  NAND2_X1 U18337 ( .A1(n15096), .A2(n19127), .ZN(n15056) );
  NAND2_X1 U18338 ( .A1(n12991), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15055) );
  OAI211_X1 U18339 ( .C1(n15345), .C2(n12991), .A(n15056), .B(n15055), .ZN(
        P2_U2860) );
  AND2_X1 U18340 ( .A1(n9672), .A2(n15057), .ZN(n15059) );
  OR2_X1 U18341 ( .A1(n15059), .A2(n15058), .ZN(n15361) );
  AOI21_X1 U18342 ( .B1(n15060), .B2(n15062), .A(n15061), .ZN(n15102) );
  NAND2_X1 U18343 ( .A1(n15102), .A2(n19127), .ZN(n15064) );
  NAND2_X1 U18344 ( .A1(n12991), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15063) );
  OAI211_X1 U18345 ( .C1(n15361), .C2(n12991), .A(n15064), .B(n15063), .ZN(
        P2_U2861) );
  OAI21_X1 U18346 ( .B1(n15065), .B2(n15067), .A(n15066), .ZN(n15118) );
  NAND2_X1 U18347 ( .A1(n9711), .A2(n15068), .ZN(n15069) );
  NAND2_X1 U18348 ( .A1(n9672), .A2(n15069), .ZN(n16088) );
  MUX2_X1 U18349 ( .A(n16088), .B(n15070), .S(n12991), .Z(n15071) );
  OAI21_X1 U18350 ( .B1(n15118), .B2(n19145), .A(n15071), .ZN(P2_U2862) );
  AOI21_X1 U18351 ( .B1(n9743), .B2(n15073), .A(n15072), .ZN(n15074) );
  XOR2_X1 U18352 ( .A(n15075), .B(n15074), .Z(n15124) );
  INV_X1 U18353 ( .A(n15383), .ZN(n16133) );
  NOR2_X1 U18354 ( .A1(n16133), .A2(n12991), .ZN(n15076) );
  AOI21_X1 U18355 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n12991), .A(n15076), .ZN(
        n15077) );
  OAI21_X1 U18356 ( .B1(n15124), .B2(n19145), .A(n15077), .ZN(P2_U2863) );
  OAI21_X1 U18357 ( .B1(n15078), .B2(n15080), .A(n15079), .ZN(n15142) );
  NOR2_X1 U18358 ( .A1(n15432), .A2(n12991), .ZN(n15081) );
  AOI21_X1 U18359 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n12991), .A(n15081), .ZN(
        n15082) );
  OAI21_X1 U18360 ( .B1(n15142), .B2(n19145), .A(n15082), .ZN(P2_U2866) );
  AND2_X1 U18361 ( .A1(n15486), .A2(n15083), .ZN(n15084) );
  OR2_X1 U18362 ( .A1(n15084), .A2(n9736), .ZN(n18943) );
  AOI21_X1 U18363 ( .B1(n15087), .B2(n15085), .A(n15086), .ZN(n15149) );
  NAND2_X1 U18364 ( .A1(n15149), .A2(n19127), .ZN(n15089) );
  NAND2_X1 U18365 ( .A1(n12991), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15088) );
  OAI211_X1 U18366 ( .C1(n18943), .C2(n12991), .A(n15089), .B(n15088), .ZN(
        P2_U2868) );
  INV_X1 U18367 ( .A(n15090), .ZN(n15330) );
  OAI22_X1 U18368 ( .A1(n15091), .A2(n15131), .B1(n15130), .B2(n12781), .ZN(
        n15092) );
  AOI21_X1 U18369 ( .B1(n19150), .B2(n15330), .A(n15092), .ZN(n15094) );
  AOI22_X1 U18370 ( .A1(n19153), .A2(BUF1_REG_28__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15093) );
  OAI211_X1 U18371 ( .C1(n15095), .C2(n16120), .A(n15094), .B(n15093), .ZN(
        P2_U2891) );
  NAND2_X1 U18372 ( .A1(n15096), .A2(n19173), .ZN(n15101) );
  AOI22_X1 U18373 ( .A1(n19150), .A2(n15343), .B1(n19169), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U18374 ( .A1(n19153), .A2(BUF1_REG_27__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15099) );
  NAND2_X1 U18375 ( .A1(n16127), .A2(n15097), .ZN(n15098) );
  NAND4_X1 U18376 ( .A1(n15101), .A2(n15100), .A3(n15099), .A4(n15098), .ZN(
        P2_U2892) );
  NAND2_X1 U18377 ( .A1(n15102), .A2(n19173), .ZN(n15109) );
  OR2_X1 U18378 ( .A1(n15104), .A2(n15103), .ZN(n15105) );
  AND2_X1 U18379 ( .A1(n12670), .A2(n15105), .ZN(n16081) );
  AOI22_X1 U18380 ( .A1(n19150), .A2(n16081), .B1(n19169), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15108) );
  AOI22_X1 U18381 ( .A1(n19153), .A2(BUF1_REG_26__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15107) );
  NAND2_X1 U18382 ( .A1(n16127), .A2(n19160), .ZN(n15106) );
  NAND4_X1 U18383 ( .A1(n15109), .A2(n15108), .A3(n15107), .A4(n15106), .ZN(
        P2_U2893) );
  AOI22_X1 U18384 ( .A1(n19153), .A2(BUF1_REG_25__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15114) );
  INV_X1 U18385 ( .A(n15110), .ZN(n15111) );
  XNOR2_X1 U18386 ( .A(n15112), .B(n15111), .ZN(n16086) );
  AOI22_X1 U18387 ( .A1(n19150), .A2(n16086), .B1(n19169), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15113) );
  OAI211_X1 U18388 ( .C1(n15115), .C2(n15131), .A(n15114), .B(n15113), .ZN(
        n15116) );
  INV_X1 U18389 ( .A(n15116), .ZN(n15117) );
  OAI21_X1 U18390 ( .B1(n15118), .B2(n16120), .A(n15117), .ZN(P2_U2894) );
  INV_X1 U18391 ( .A(n15386), .ZN(n15121) );
  OAI22_X1 U18392 ( .A1(n15119), .A2(n15131), .B1(n15130), .B2(n13000), .ZN(
        n15120) );
  AOI21_X1 U18393 ( .B1(n19150), .B2(n15121), .A(n15120), .ZN(n15123) );
  AOI22_X1 U18394 ( .A1(n19153), .A2(BUF1_REG_24__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15122) );
  OAI211_X1 U18395 ( .C1(n15124), .C2(n16120), .A(n15123), .B(n15122), .ZN(
        P2_U2895) );
  INV_X1 U18396 ( .A(n15126), .ZN(n15127) );
  AOI21_X1 U18397 ( .B1(n15125), .B2(n15128), .A(n15127), .ZN(n16099) );
  INV_X1 U18398 ( .A(n16099), .ZN(n15136) );
  INV_X1 U18399 ( .A(n15401), .ZN(n15133) );
  OAI22_X1 U18400 ( .A1(n19308), .A2(n15131), .B1(n15130), .B2(n15129), .ZN(
        n15132) );
  AOI21_X1 U18401 ( .B1(n19150), .B2(n15133), .A(n15132), .ZN(n15135) );
  AOI22_X1 U18402 ( .A1(n19153), .A2(BUF1_REG_23__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15134) );
  OAI211_X1 U18403 ( .C1(n15136), .C2(n16120), .A(n15135), .B(n15134), .ZN(
        P2_U2896) );
  AOI22_X1 U18404 ( .A1(n19153), .A2(BUF1_REG_21__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U18405 ( .A1(n16127), .A2(n19170), .B1(n19169), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15137) );
  OAI211_X1 U18406 ( .C1(n16119), .C2(n15139), .A(n15138), .B(n15137), .ZN(
        n15140) );
  INV_X1 U18407 ( .A(n15140), .ZN(n15141) );
  OAI21_X1 U18408 ( .B1(n15142), .B2(n16120), .A(n15141), .ZN(P2_U2898) );
  NOR2_X1 U18409 ( .A1(n15143), .A2(n15489), .ZN(n15144) );
  OR2_X1 U18410 ( .A1(n15442), .A2(n15144), .ZN(n18942) );
  AOI22_X1 U18411 ( .A1(n19153), .A2(BUF1_REG_19__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15147) );
  AOI22_X1 U18412 ( .A1(n16127), .A2(n15145), .B1(n19169), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15146) );
  OAI211_X1 U18413 ( .C1(n16119), .C2(n18942), .A(n15147), .B(n15146), .ZN(
        n15148) );
  AOI21_X1 U18414 ( .B1(n15149), .B2(n19173), .A(n15148), .ZN(n15150) );
  INV_X1 U18415 ( .A(n15150), .ZN(P2_U2900) );
  NOR2_X1 U18416 ( .A1(n15154), .A2(n15153), .ZN(n15155) );
  XNOR2_X1 U18417 ( .A(n15156), .B(n15155), .ZN(n16046) );
  AOI21_X1 U18418 ( .B1(n16046), .B2(n13426), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15174) );
  AND2_X1 U18419 ( .A1(n13426), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15157) );
  NAND2_X1 U18420 ( .A1(n16046), .A2(n15157), .ZN(n15172) );
  NOR2_X1 U18421 ( .A1(n15159), .A2(n15158), .ZN(n15160) );
  XOR2_X1 U18422 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n15160), .Z(
        n15161) );
  NAND2_X1 U18423 ( .A1(n15186), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15162) );
  XNOR2_X1 U18424 ( .A(n15162), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15308) );
  INV_X1 U18425 ( .A(n15308), .ZN(n15167) );
  NAND2_X1 U18426 ( .A1(n16187), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15164) );
  NAND2_X1 U18427 ( .A1(n15785), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15304) );
  OAI211_X1 U18428 ( .C1(n16098), .C2(n19223), .A(n15164), .B(n15304), .ZN(
        n15165) );
  INV_X1 U18429 ( .A(n15165), .ZN(n15166) );
  INV_X1 U18430 ( .A(n15168), .ZN(n15169) );
  OAI21_X1 U18431 ( .B1(n15310), .B2(n19224), .A(n15169), .ZN(P2_U2983) );
  NAND2_X1 U18432 ( .A1(n15171), .A2(n15170), .ZN(n15176) );
  INV_X1 U18433 ( .A(n15172), .ZN(n15173) );
  NOR2_X1 U18434 ( .A1(n15174), .A2(n15173), .ZN(n15175) );
  XNOR2_X1 U18435 ( .A(n15176), .B(n15175), .ZN(n15324) );
  XOR2_X1 U18436 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15186), .Z(
        n15322) );
  INV_X1 U18437 ( .A(n15177), .ZN(n16052) );
  NAND2_X1 U18438 ( .A1(n15785), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15312) );
  OAI21_X1 U18439 ( .B1(n19231), .B2(n15178), .A(n15312), .ZN(n15179) );
  AOI21_X1 U18440 ( .B1(n16052), .B2(n16239), .A(n15179), .ZN(n15180) );
  OAI21_X1 U18441 ( .B1(n16050), .B2(n16236), .A(n15180), .ZN(n15181) );
  AOI21_X1 U18442 ( .B1(n15322), .B2(n19227), .A(n15181), .ZN(n15182) );
  OAI21_X1 U18443 ( .B1(n15324), .B2(n19224), .A(n15182), .ZN(P2_U2984) );
  AOI21_X1 U18444 ( .B1(n16187), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15183), .ZN(n15184) );
  OAI21_X1 U18445 ( .B1(n16061), .B2(n19223), .A(n15184), .ZN(n15188) );
  NOR3_X1 U18446 ( .A1(n15186), .A2(n15185), .A3(n16251), .ZN(n15187) );
  AOI211_X1 U18447 ( .C1(n19216), .C2(n16059), .A(n15188), .B(n15187), .ZN(
        n15189) );
  OAI21_X1 U18448 ( .B1(n15190), .B2(n19224), .A(n15189), .ZN(P2_U2985) );
  XNOR2_X1 U18449 ( .A(n15191), .B(n15193), .ZN(n15207) );
  INV_X1 U18450 ( .A(n15191), .ZN(n15192) );
  AOI22_X1 U18451 ( .A1(n15207), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n15193), .B2(n15192), .ZN(n15196) );
  XNOR2_X1 U18452 ( .A(n15194), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15195) );
  XNOR2_X1 U18453 ( .A(n15196), .B(n15195), .ZN(n15338) );
  XNOR2_X1 U18454 ( .A(n15197), .B(n15346), .ZN(n15331) );
  NAND2_X1 U18455 ( .A1(n15331), .A2(n19227), .ZN(n15203) );
  NAND2_X1 U18456 ( .A1(n15325), .A2(n16239), .ZN(n15201) );
  NOR2_X1 U18457 ( .A1(n19066), .A2(n15199), .ZN(n15329) );
  NAND2_X1 U18458 ( .A1(n15203), .A2(n15202), .ZN(n15204) );
  AOI21_X1 U18459 ( .B1(n15205), .B2(n19216), .A(n15204), .ZN(n15206) );
  OAI21_X1 U18460 ( .B1(n15338), .B2(n19224), .A(n15206), .ZN(P2_U2986) );
  XNOR2_X1 U18461 ( .A(n15207), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15352) );
  NOR2_X1 U18462 ( .A1(n19066), .A2(n19913), .ZN(n15341) );
  AOI21_X1 U18463 ( .B1(n16187), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15341), .ZN(n15208) );
  OAI21_X1 U18464 ( .B1(n15345), .B2(n19223), .A(n15208), .ZN(n15210) );
  AND2_X1 U18465 ( .A1(n15216), .A2(n15327), .ZN(n15347) );
  NOR3_X1 U18466 ( .A1(n15347), .A2(n15346), .A3(n16251), .ZN(n15209) );
  AOI211_X1 U18467 ( .C1(n19216), .C2(n15211), .A(n15210), .B(n15209), .ZN(
        n15212) );
  OAI21_X1 U18468 ( .B1(n15352), .B2(n19224), .A(n15212), .ZN(P2_U2987) );
  OAI21_X1 U18469 ( .B1(n15213), .B2(n14223), .A(n15224), .ZN(n15214) );
  XOR2_X1 U18470 ( .A(n15215), .B(n15214), .Z(n15365) );
  INV_X1 U18471 ( .A(n15379), .ZN(n15227) );
  NOR2_X1 U18472 ( .A1(n15227), .A2(n15355), .ZN(n15226) );
  OAI21_X1 U18473 ( .B1(n15226), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15216), .ZN(n15217) );
  INV_X1 U18474 ( .A(n15217), .ZN(n15363) );
  INV_X1 U18475 ( .A(n15361), .ZN(n16076) );
  NAND2_X1 U18476 ( .A1(n15785), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15353) );
  OAI21_X1 U18477 ( .B1(n19231), .B2(n10124), .A(n15353), .ZN(n15218) );
  AOI21_X1 U18478 ( .B1(n16076), .B2(n16239), .A(n15218), .ZN(n15219) );
  OAI21_X1 U18479 ( .B1(n15220), .B2(n16236), .A(n15219), .ZN(n15221) );
  AOI21_X1 U18480 ( .B1(n15363), .B2(n19227), .A(n15221), .ZN(n15222) );
  OAI21_X1 U18481 ( .B1(n15365), .B2(n19224), .A(n15222), .ZN(P2_U2988) );
  NAND2_X1 U18482 ( .A1(n15224), .A2(n15223), .ZN(n15225) );
  XNOR2_X1 U18483 ( .A(n15213), .B(n15225), .ZN(n15374) );
  AOI21_X1 U18484 ( .B1(n15227), .B2(n15355), .A(n15226), .ZN(n15372) );
  OAI22_X1 U18485 ( .A1(n19231), .A2(n16083), .B1(n19908), .B2(n19066), .ZN(
        n15228) );
  AOI21_X1 U18486 ( .B1(n19216), .B2(n16092), .A(n15228), .ZN(n15229) );
  OAI21_X1 U18487 ( .B1(n16088), .B2(n19223), .A(n15229), .ZN(n15230) );
  AOI21_X1 U18488 ( .B1(n15372), .B2(n19227), .A(n15230), .ZN(n15231) );
  OAI21_X1 U18489 ( .B1(n19224), .B2(n15374), .A(n15231), .ZN(P2_U2989) );
  NAND2_X1 U18490 ( .A1(n15232), .A2(n15497), .ZN(n15763) );
  INV_X1 U18491 ( .A(n15762), .ZN(n15233) );
  INV_X1 U18492 ( .A(n15234), .ZN(n15236) );
  INV_X1 U18493 ( .A(n15280), .ZN(n15235) );
  INV_X1 U18494 ( .A(n15471), .ZN(n15237) );
  NAND2_X1 U18495 ( .A1(n15272), .A2(n15274), .ZN(n15254) );
  INV_X1 U18496 ( .A(n15255), .ZN(n15238) );
  AOI21_X1 U18497 ( .B1(n15254), .B2(n15239), .A(n15238), .ZN(n15243) );
  NAND2_X1 U18498 ( .A1(n15241), .A2(n15240), .ZN(n15242) );
  XNOR2_X1 U18499 ( .A(n15243), .B(n15242), .ZN(n15438) );
  NAND2_X1 U18500 ( .A1(n19216), .A2(n15244), .ZN(n15245) );
  NAND2_X1 U18501 ( .A1(n15785), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15427) );
  OAI211_X1 U18502 ( .C1(n19231), .C2(n15246), .A(n15245), .B(n15427), .ZN(
        n15250) );
  INV_X1 U18503 ( .A(n15440), .ZN(n15478) );
  NAND2_X1 U18504 ( .A1(n15548), .A2(n15478), .ZN(n15475) );
  INV_X1 U18505 ( .A(n15475), .ZN(n15247) );
  NOR2_X2 U18506 ( .A1(n15477), .A2(n15248), .ZN(n15259) );
  NAND2_X1 U18507 ( .A1(n15259), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15410) );
  OAI21_X1 U18508 ( .B1(n15259), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15410), .ZN(n15433) );
  NOR2_X1 U18509 ( .A1(n15433), .A2(n16251), .ZN(n15249) );
  AOI211_X1 U18510 ( .C1(n16239), .C2(n15251), .A(n15250), .B(n15249), .ZN(
        n15252) );
  OAI21_X1 U18511 ( .B1(n15438), .B2(n19224), .A(n15252), .ZN(P2_U2993) );
  NAND2_X1 U18512 ( .A1(n15254), .A2(n15253), .ZN(n15258) );
  NAND2_X1 U18513 ( .A1(n15256), .A2(n15255), .ZN(n15257) );
  XNOR2_X1 U18514 ( .A(n15258), .B(n15257), .ZN(n15458) );
  INV_X1 U18515 ( .A(n15477), .ZN(n15268) );
  NAND2_X1 U18516 ( .A1(n15268), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15267) );
  AOI21_X1 U18517 ( .B1(n15452), .B2(n15267), .A(n15259), .ZN(n15439) );
  NAND2_X1 U18518 ( .A1(n15785), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15445) );
  OAI21_X1 U18519 ( .B1(n16236), .B2(n15260), .A(n15445), .ZN(n15265) );
  OR2_X1 U18520 ( .A1(n9736), .A2(n15261), .ZN(n15262) );
  NAND2_X1 U18521 ( .A1(n12683), .A2(n15262), .ZN(n18931) );
  INV_X1 U18522 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15263) );
  OAI22_X1 U18523 ( .A1(n18931), .A2(n19223), .B1(n15263), .B2(n19231), .ZN(
        n15264) );
  AOI211_X1 U18524 ( .C1(n15439), .C2(n19227), .A(n15265), .B(n15264), .ZN(
        n15266) );
  OAI21_X1 U18525 ( .B1(n19224), .B2(n15458), .A(n15266), .ZN(P2_U2994) );
  OAI21_X1 U18526 ( .B1(n15268), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15267), .ZN(n15470) );
  NOR2_X1 U18527 ( .A1(n18943), .A2(n19223), .ZN(n15271) );
  NAND2_X1 U18528 ( .A1(n15785), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15460) );
  OAI21_X1 U18529 ( .B1(n19231), .B2(n15269), .A(n15460), .ZN(n15270) );
  AOI211_X1 U18530 ( .C1(n18946), .C2(n19216), .A(n15271), .B(n15270), .ZN(
        n15278) );
  NAND2_X1 U18531 ( .A1(n15274), .A2(n15273), .ZN(n15275) );
  XNOR2_X1 U18532 ( .A(n15276), .B(n15275), .ZN(n15467) );
  NAND2_X1 U18533 ( .A1(n15467), .A2(n16240), .ZN(n15277) );
  OAI211_X1 U18534 ( .C1(n15470), .C2(n16251), .A(n15278), .B(n15277), .ZN(
        P2_U2995) );
  NAND2_X1 U18535 ( .A1(n15280), .A2(n15279), .ZN(n15284) );
  NAND2_X1 U18536 ( .A1(n15282), .A2(n15281), .ZN(n15283) );
  XOR2_X1 U18537 ( .A(n15284), .B(n15283), .Z(n15792) );
  OAI211_X1 U18538 ( .C1(n15759), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19227), .B(n15475), .ZN(n15289) );
  NOR2_X1 U18539 ( .A1(n19896), .A2(n19066), .ZN(n15287) );
  OAI22_X1 U18540 ( .A1(n19231), .A2(n18968), .B1(n16236), .B2(n18966), .ZN(
        n15286) );
  AOI211_X1 U18541 ( .C1(n16239), .C2(n18974), .A(n15287), .B(n15286), .ZN(
        n15288) );
  OAI211_X1 U18542 ( .C1(n15792), .C2(n19224), .A(n15289), .B(n15288), .ZN(
        P2_U2997) );
  NAND2_X1 U18543 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15517), .ZN(
        n15516) );
  NOR2_X1 U18544 ( .A1(n16259), .A2(n15530), .ZN(n16182) );
  AOI21_X1 U18545 ( .B1(n14143), .B2(n15516), .A(n16182), .ZN(n15290) );
  INV_X1 U18546 ( .A(n15290), .ZN(n15515) );
  INV_X1 U18547 ( .A(n15291), .ZN(n15292) );
  NOR2_X1 U18548 ( .A1(n15293), .A2(n15292), .ZN(n15294) );
  XNOR2_X1 U18549 ( .A(n15295), .B(n15294), .ZN(n15512) );
  OAI22_X1 U18550 ( .A1(n19231), .A2(n15296), .B1(n16236), .B2(n19012), .ZN(
        n15299) );
  INV_X1 U18551 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15297) );
  OAI22_X1 U18552 ( .A1(n19001), .A2(n19223), .B1(n19066), .B2(n15297), .ZN(
        n15298) );
  AOI211_X1 U18553 ( .C1(n15512), .C2(n16240), .A(n15299), .B(n15298), .ZN(
        n15300) );
  OAI21_X1 U18554 ( .B1(n15515), .B2(n16251), .A(n15300), .ZN(P2_U3001) );
  NAND2_X1 U18555 ( .A1(n15579), .A2(n15301), .ZN(n15302) );
  AND2_X1 U18556 ( .A1(n15339), .A2(n15302), .ZN(n15316) );
  OAI21_X1 U18557 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15787), .A(
        n15316), .ZN(n15307) );
  AND4_X1 U18558 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A4(n15303), .ZN(n15311) );
  NAND3_X1 U18559 ( .A1(n15311), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12596), .ZN(n15305) );
  OAI211_X1 U18560 ( .C1(n19149), .C2(n16290), .A(n15305), .B(n15304), .ZN(
        n15306) );
  NAND2_X1 U18561 ( .A1(n15308), .A2(n19250), .ZN(n15309) );
  INV_X1 U18562 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15315) );
  NAND2_X1 U18563 ( .A1(n15311), .A2(n15315), .ZN(n15313) );
  NAND2_X1 U18564 ( .A1(n15313), .A2(n15312), .ZN(n15314) );
  AOI21_X1 U18565 ( .B1(n15322), .B2(n19250), .A(n15321), .ZN(n15323) );
  OAI21_X1 U18566 ( .B1(n15324), .B2(n16273), .A(n15323), .ZN(P2_U3016) );
  INV_X1 U18567 ( .A(n15325), .ZN(n15334) );
  NOR3_X1 U18568 ( .A1(n15327), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15326), .ZN(n15328) );
  AOI211_X1 U18569 ( .C1(n19262), .C2(n15330), .A(n15329), .B(n15328), .ZN(
        n15333) );
  NAND2_X1 U18570 ( .A1(n19250), .A2(n15331), .ZN(n15332) );
  OAI211_X1 U18571 ( .C1(n15334), .C2(n16277), .A(n15333), .B(n15332), .ZN(
        n15335) );
  AOI21_X1 U18572 ( .B1(n15336), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15335), .ZN(n15337) );
  OAI21_X1 U18573 ( .B1(n15338), .B2(n16273), .A(n15337), .ZN(P2_U3018) );
  INV_X1 U18574 ( .A(n15339), .ZN(n15350) );
  INV_X1 U18575 ( .A(n15340), .ZN(n15342) );
  AOI211_X1 U18576 ( .C1(n19262), .C2(n15343), .A(n15342), .B(n15341), .ZN(
        n15344) );
  OAI21_X1 U18577 ( .B1(n15345), .B2(n16277), .A(n15344), .ZN(n15349) );
  NOR3_X1 U18578 ( .A1(n15347), .A2(n15346), .A3(n16292), .ZN(n15348) );
  AOI211_X1 U18579 ( .C1(n15350), .C2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15349), .B(n15348), .ZN(n15351) );
  OAI21_X1 U18580 ( .B1(n15352), .B2(n16273), .A(n15351), .ZN(P2_U3019) );
  NAND3_X1 U18581 ( .A1(n15381), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15538), .ZN(n15360) );
  INV_X1 U18582 ( .A(n15353), .ZN(n15358) );
  AOI211_X1 U18583 ( .C1(n15356), .C2(n15355), .A(n15367), .B(n15354), .ZN(
        n15357) );
  AOI211_X1 U18584 ( .C1(n19262), .C2(n16081), .A(n15358), .B(n15357), .ZN(
        n15359) );
  OAI211_X1 U18585 ( .C1(n15361), .C2(n16277), .A(n15360), .B(n15359), .ZN(
        n15362) );
  AOI21_X1 U18586 ( .B1(n15363), .B2(n19250), .A(n15362), .ZN(n15364) );
  OAI21_X1 U18587 ( .B1(n15365), .B2(n16273), .A(n15364), .ZN(P2_U3020) );
  NAND3_X1 U18588 ( .A1(n15381), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15538), .ZN(n15370) );
  NAND2_X1 U18589 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n12657), .ZN(n15366) );
  OAI21_X1 U18590 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15367), .A(
        n15366), .ZN(n15368) );
  AOI21_X1 U18591 ( .B1(n19262), .B2(n16086), .A(n15368), .ZN(n15369) );
  OAI211_X1 U18592 ( .C1(n16088), .C2(n16277), .A(n15370), .B(n15369), .ZN(
        n15371) );
  AOI21_X1 U18593 ( .B1(n15372), .B2(n19250), .A(n15371), .ZN(n15373) );
  OAI21_X1 U18594 ( .B1(n16273), .B2(n15374), .A(n15373), .ZN(P2_U3021) );
  NOR2_X1 U18595 ( .A1(n10219), .A2(n15376), .ZN(n15377) );
  XNOR2_X1 U18596 ( .A(n15378), .B(n15377), .ZN(n16134) );
  AOI21_X1 U18597 ( .B1(n15380), .B2(n15389), .A(n15379), .ZN(n16136) );
  OAI21_X1 U18598 ( .B1(n15382), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15381), .ZN(n15385) );
  AOI22_X1 U18599 ( .A1(n15383), .A2(n19248), .B1(P2_REIP_REG_24__SCAN_IN), 
        .B2(n15785), .ZN(n15384) );
  OAI211_X1 U18600 ( .C1(n16290), .C2(n15386), .A(n15385), .B(n15384), .ZN(
        n15387) );
  AOI21_X1 U18601 ( .B1(n16136), .B2(n19250), .A(n15387), .ZN(n15388) );
  OAI21_X1 U18602 ( .B1(n16134), .B2(n16273), .A(n15388), .ZN(P2_U3022) );
  NOR2_X1 U18603 ( .A1(n15409), .A2(n15410), .ZN(n15408) );
  OAI21_X1 U18604 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15408), .A(
        n15389), .ZN(n16147) );
  INV_X1 U18605 ( .A(n15390), .ZN(n15392) );
  AOI21_X1 U18606 ( .B1(n9708), .B2(n15392), .A(n15391), .ZN(n16144) );
  INV_X1 U18607 ( .A(n15393), .ZN(n15394) );
  OAI21_X1 U18608 ( .B1(n15787), .B2(n15394), .A(n15559), .ZN(n15436) );
  NAND2_X1 U18609 ( .A1(n15436), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15400) );
  NOR2_X1 U18610 ( .A1(n19904), .A2(n19066), .ZN(n15398) );
  OAI21_X1 U18611 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15395), .ZN(n15396) );
  NOR2_X1 U18612 ( .A1(n15396), .A2(n15420), .ZN(n15397) );
  AOI211_X1 U18613 ( .C1(n16143), .C2(n19248), .A(n15398), .B(n15397), .ZN(
        n15399) );
  OAI211_X1 U18614 ( .C1(n16290), .C2(n15401), .A(n15400), .B(n15399), .ZN(
        n15402) );
  AOI21_X1 U18615 ( .B1(n16144), .B2(n19255), .A(n15402), .ZN(n15403) );
  OAI21_X1 U18616 ( .B1(n16147), .B2(n16292), .A(n15403), .ZN(P2_U3023) );
  NAND2_X1 U18617 ( .A1(n15405), .A2(n15404), .ZN(n15407) );
  XOR2_X1 U18618 ( .A(n15407), .B(n15406), .Z(n16149) );
  AOI21_X1 U18619 ( .B1(n15410), .B2(n15409), .A(n15408), .ZN(n16151) );
  NAND2_X1 U18620 ( .A1(n16151), .A2(n19250), .ZN(n15425) );
  AND2_X1 U18621 ( .A1(n15412), .A2(n15411), .ZN(n15414) );
  OR2_X1 U18622 ( .A1(n15414), .A2(n15413), .ZN(n16148) );
  NOR2_X1 U18623 ( .A1(n15416), .A2(n15415), .ZN(n15417) );
  OR2_X1 U18624 ( .A1(n15418), .A2(n15417), .ZN(n15775) );
  INV_X1 U18625 ( .A(n15775), .ZN(n16112) );
  NAND2_X1 U18626 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n12657), .ZN(n15419) );
  OAI21_X1 U18627 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15420), .A(
        n15419), .ZN(n15421) );
  AOI21_X1 U18628 ( .B1(n19262), .B2(n16112), .A(n15421), .ZN(n15422) );
  OAI21_X1 U18629 ( .B1(n16148), .B2(n16277), .A(n15422), .ZN(n15423) );
  AOI21_X1 U18630 ( .B1(n15436), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15423), .ZN(n15424) );
  OAI211_X1 U18631 ( .C1(n16149), .C2(n16273), .A(n15425), .B(n15424), .ZN(
        P2_U3024) );
  NAND3_X1 U18632 ( .A1(n15426), .A2(n15540), .A3(n14155), .ZN(n15431) );
  INV_X1 U18633 ( .A(n15427), .ZN(n15428) );
  AOI21_X1 U18634 ( .B1(n19262), .B2(n15429), .A(n15428), .ZN(n15430) );
  OAI211_X1 U18635 ( .C1(n16277), .C2(n15432), .A(n15431), .B(n15430), .ZN(
        n15435) );
  NOR2_X1 U18636 ( .A1(n15433), .A2(n16292), .ZN(n15434) );
  AOI211_X1 U18637 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15436), .A(
        n15435), .B(n15434), .ZN(n15437) );
  OAI21_X1 U18638 ( .B1(n15438), .B2(n16273), .A(n15437), .ZN(P2_U3025) );
  NAND2_X1 U18639 ( .A1(n15439), .A2(n19250), .ZN(n15457) );
  NOR4_X1 U18640 ( .A1(n15440), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15451), .A4(n15481), .ZN(n15455) );
  NOR2_X1 U18641 ( .A1(n15442), .A2(n15441), .ZN(n15443) );
  NOR2_X1 U18642 ( .A1(n15444), .A2(n15443), .ZN(n16118) );
  NAND2_X1 U18643 ( .A1(n19262), .A2(n16118), .ZN(n15446) );
  OAI211_X1 U18644 ( .C1(n16277), .C2(n18931), .A(n15446), .B(n15445), .ZN(
        n15454) );
  NAND3_X1 U18645 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15449) );
  INV_X1 U18646 ( .A(n15447), .ZN(n15501) );
  INV_X1 U18647 ( .A(n15559), .ZN(n15448) );
  OAI21_X1 U18648 ( .B1(n15500), .B2(n15448), .A(n15538), .ZN(n15523) );
  OAI21_X1 U18649 ( .B1(n15501), .B2(n15787), .A(n15523), .ZN(n15761) );
  AOI21_X1 U18650 ( .B1(n15449), .B2(n15579), .A(n15761), .ZN(n15480) );
  INV_X1 U18651 ( .A(n15480), .ZN(n15450) );
  AOI21_X1 U18652 ( .B1(n15481), .B2(n15579), .A(n15450), .ZN(n15459) );
  NAND4_X1 U18653 ( .A1(n15540), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15451), .A4(n15478), .ZN(n15464) );
  AOI21_X1 U18654 ( .B1(n15459), .B2(n15464), .A(n15452), .ZN(n15453) );
  AOI211_X1 U18655 ( .C1(n15540), .C2(n15455), .A(n15454), .B(n15453), .ZN(
        n15456) );
  OAI211_X1 U18656 ( .C1(n15458), .C2(n16273), .A(n15457), .B(n15456), .ZN(
        P2_U3026) );
  INV_X1 U18657 ( .A(n15459), .ZN(n15466) );
  INV_X1 U18658 ( .A(n18943), .ZN(n15462) );
  INV_X1 U18659 ( .A(n15460), .ZN(n15461) );
  AOI21_X1 U18660 ( .B1(n15462), .B2(n19248), .A(n15461), .ZN(n15463) );
  OAI211_X1 U18661 ( .C1(n16290), .C2(n18942), .A(n15464), .B(n15463), .ZN(
        n15465) );
  AOI21_X1 U18662 ( .B1(n15466), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15465), .ZN(n15469) );
  NAND2_X1 U18663 ( .A1(n15467), .A2(n19255), .ZN(n15468) );
  OAI211_X1 U18664 ( .C1(n15470), .C2(n16292), .A(n15469), .B(n15468), .ZN(
        P2_U3027) );
  AND2_X1 U18665 ( .A1(n15472), .A2(n15471), .ZN(n15473) );
  XNOR2_X1 U18666 ( .A(n15474), .B(n15473), .ZN(n16155) );
  NAND2_X1 U18667 ( .A1(n15475), .A2(n15481), .ZN(n15476) );
  NAND2_X1 U18668 ( .A1(n15477), .A2(n15476), .ZN(n16156) );
  INV_X1 U18669 ( .A(n16156), .ZN(n15494) );
  NAND2_X1 U18670 ( .A1(n15478), .A2(n15540), .ZN(n15482) );
  NAND2_X1 U18671 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n12657), .ZN(n15479) );
  OAI221_X1 U18672 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15482), 
        .C1(n15481), .C2(n15480), .A(n15479), .ZN(n15493) );
  NAND2_X1 U18673 ( .A1(n15484), .A2(n15483), .ZN(n15485) );
  NAND2_X1 U18674 ( .A1(n15486), .A2(n15485), .ZN(n18954) );
  NAND2_X1 U18675 ( .A1(n15488), .A2(n15487), .ZN(n15491) );
  INV_X1 U18676 ( .A(n15489), .ZN(n15490) );
  NAND2_X1 U18677 ( .A1(n15491), .A2(n15490), .ZN(n18953) );
  OAI22_X1 U18678 ( .A1(n16277), .A2(n18954), .B1(n16290), .B2(n18953), .ZN(
        n15492) );
  AOI211_X1 U18679 ( .C1(n15494), .C2(n19250), .A(n15493), .B(n15492), .ZN(
        n15495) );
  OAI21_X1 U18680 ( .B1(n16273), .B2(n16155), .A(n15495), .ZN(P2_U3028) );
  NAND2_X1 U18681 ( .A1(n15497), .A2(n15496), .ZN(n15498) );
  XNOR2_X1 U18682 ( .A(n15499), .B(n15498), .ZN(n16171) );
  NOR2_X1 U18683 ( .A1(n15500), .A2(n15555), .ZN(n15507) );
  NAND2_X1 U18684 ( .A1(n15501), .A2(n15507), .ZN(n15757) );
  OAI22_X1 U18685 ( .A1(n16277), .A2(n15502), .B1(n16290), .B2(n19000), .ZN(
        n15504) );
  AOI21_X1 U18686 ( .B1(n14178), .B2(n16181), .A(n16166), .ZN(n16170) );
  INV_X1 U18687 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19892) );
  NOR2_X1 U18688 ( .A1(n19892), .A2(n19066), .ZN(n15503) );
  AOI21_X1 U18689 ( .B1(n15761), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15505), .ZN(n15506) );
  OAI21_X1 U18690 ( .B1(n16171), .B2(n16273), .A(n15506), .ZN(P2_U3031) );
  INV_X1 U18691 ( .A(n15507), .ZN(n16258) );
  OAI21_X1 U18692 ( .B1(n15524), .B2(n16258), .A(n14143), .ZN(n15511) );
  OAI21_X1 U18693 ( .B1(n15508), .B2(n16258), .A(n15523), .ZN(n16254) );
  NOR2_X1 U18694 ( .A1(n16277), .A2(n19001), .ZN(n15510) );
  OAI22_X1 U18695 ( .A1(n16290), .A2(n19016), .B1(n15297), .B2(n19066), .ZN(
        n15509) );
  AOI211_X1 U18696 ( .C1(n15511), .C2(n16254), .A(n15510), .B(n15509), .ZN(
        n15514) );
  NAND2_X1 U18697 ( .A1(n15512), .A2(n19255), .ZN(n15513) );
  OAI211_X1 U18698 ( .C1(n15515), .C2(n16292), .A(n15514), .B(n15513), .ZN(
        P2_U3033) );
  OAI21_X1 U18699 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15517), .A(
        n15516), .ZN(n15518) );
  INV_X1 U18700 ( .A(n15518), .ZN(n16188) );
  NAND2_X1 U18701 ( .A1(n16188), .A2(n19250), .ZN(n15529) );
  AOI22_X1 U18702 ( .A1(n19262), .A2(n19156), .B1(n19248), .B2(n19126), .ZN(
        n15528) );
  XNOR2_X1 U18703 ( .A(n15519), .B(n15524), .ZN(n15520) );
  XNOR2_X1 U18704 ( .A(n15521), .B(n15520), .ZN(n16189) );
  NAND2_X1 U18705 ( .A1(n16189), .A2(n19255), .ZN(n15527) );
  NAND2_X1 U18706 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n12657), .ZN(n15522) );
  OAI221_X1 U18707 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16258), 
        .C1(n15524), .C2(n15523), .A(n15522), .ZN(n15525) );
  INV_X1 U18708 ( .A(n15525), .ZN(n15526) );
  NAND4_X1 U18709 ( .A1(n15529), .A2(n15528), .A3(n15527), .A4(n15526), .ZN(
        P2_U3034) );
  NOR2_X1 U18710 ( .A1(n16200), .A2(n16199), .ZN(n16198) );
  OAI21_X1 U18711 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16198), .A(
        n15530), .ZN(n16194) );
  NAND2_X1 U18712 ( .A1(n15551), .A2(n15549), .ZN(n16204) );
  INV_X1 U18713 ( .A(n16202), .ZN(n15533) );
  OAI211_X1 U18714 ( .C1(n16204), .C2(n15533), .A(n16201), .B(n16203), .ZN(
        n15537) );
  AND2_X1 U18715 ( .A1(n15535), .A2(n15534), .ZN(n15536) );
  XNOR2_X1 U18716 ( .A(n15537), .B(n15536), .ZN(n16193) );
  INV_X1 U18717 ( .A(n15538), .ZN(n15539) );
  AOI21_X1 U18718 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15559), .A(
        n15539), .ZN(n16269) );
  NAND2_X1 U18719 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15540), .ZN(
        n16266) );
  AOI221_X1 U18720 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n16200), .C2(n14127), .A(
        n16266), .ZN(n15542) );
  NOR2_X1 U18721 ( .A1(n12219), .A2(n19066), .ZN(n15541) );
  AOI211_X1 U18722 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16269), .A(
        n15542), .B(n15541), .ZN(n15545) );
  INV_X1 U18723 ( .A(n19025), .ZN(n15543) );
  AOI22_X1 U18724 ( .A1(n19262), .A2(n15543), .B1(n19248), .B2(n19024), .ZN(
        n15544) );
  OAI211_X1 U18725 ( .C1(n16193), .C2(n16273), .A(n15545), .B(n15544), .ZN(
        n15546) );
  INV_X1 U18726 ( .A(n15546), .ZN(n15547) );
  OAI21_X1 U18727 ( .B1(n16194), .B2(n16292), .A(n15547), .ZN(P2_U3035) );
  OAI21_X1 U18728 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15548), .A(
        n16199), .ZN(n16219) );
  INV_X1 U18729 ( .A(n15551), .ZN(n15553) );
  AND2_X1 U18730 ( .A1(n15549), .A2(n16203), .ZN(n15550) );
  OAI21_X1 U18731 ( .B1(n15551), .B2(n15550), .A(n16204), .ZN(n15552) );
  OAI21_X1 U18732 ( .B1(n15553), .B2(n16203), .A(n15552), .ZN(n16216) );
  AOI22_X1 U18733 ( .A1(n19248), .A2(n16215), .B1(n12657), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n15554) );
  OAI21_X1 U18734 ( .B1(n15555), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15554), .ZN(n15561) );
  OAI21_X1 U18735 ( .B1(n15557), .B2(n15556), .A(n16265), .ZN(n19165) );
  OAI22_X1 U18736 ( .A1(n15559), .A2(n15558), .B1(n19165), .B2(n16290), .ZN(
        n15560) );
  AOI211_X1 U18737 ( .C1(n16216), .C2(n19255), .A(n15561), .B(n15560), .ZN(
        n15562) );
  OAI21_X1 U18738 ( .B1(n16219), .B2(n16292), .A(n15562), .ZN(P2_U3037) );
  OAI21_X1 U18739 ( .B1(n15565), .B2(n15564), .A(n15563), .ZN(n15566) );
  XOR2_X1 U18740 ( .A(n15566), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n16244) );
  INV_X1 U18741 ( .A(n15567), .ZN(n16282) );
  NAND2_X1 U18742 ( .A1(n16282), .A2(n15568), .ZN(n15570) );
  AOI22_X1 U18743 ( .A1(n19248), .A2(n19059), .B1(n15785), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n15569) );
  OAI211_X1 U18744 ( .C1(n16290), .C2(n19060), .A(n15570), .B(n15569), .ZN(
        n15571) );
  AOI21_X1 U18745 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16276), .A(
        n15571), .ZN(n15578) );
  INV_X1 U18746 ( .A(n16224), .ZN(n15576) );
  OAI21_X1 U18747 ( .B1(n15574), .B2(n15576), .A(n15573), .ZN(n15575) );
  OAI21_X1 U18748 ( .B1(n15572), .B2(n15576), .A(n15575), .ZN(n16241) );
  NAND2_X1 U18749 ( .A1(n16241), .A2(n19255), .ZN(n15577) );
  OAI211_X1 U18750 ( .C1(n16244), .C2(n16292), .A(n15578), .B(n15577), .ZN(
        P2_U3039) );
  OAI211_X1 U18751 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n19246), .B(n15579), .ZN(n15586) );
  AOI22_X1 U18752 ( .A1(n19244), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19255), .B2(n15580), .ZN(n15585) );
  AOI21_X1 U18753 ( .B1(n19248), .B2(n12867), .A(n15581), .ZN(n15584) );
  AOI22_X1 U18754 ( .A1(n19262), .A2(n19957), .B1(n19250), .B2(n15582), .ZN(
        n15583) );
  NAND4_X1 U18755 ( .A1(n15586), .A2(n15585), .A3(n15584), .A4(n15583), .ZN(
        P2_U3045) );
  MUX2_X1 U18756 ( .A(n15588), .B(n15587), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15589) );
  AOI21_X1 U18757 ( .B1(n15590), .B2(n15607), .A(n15589), .ZN(n16302) );
  INV_X1 U18758 ( .A(n15591), .ZN(n15592) );
  OAI222_X1 U18759 ( .A1(n15860), .A2(n15594), .B1(n15608), .B2(n16302), .C1(
        n15593), .C2(n15592), .ZN(n15595) );
  MUX2_X1 U18760 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15595), .S(
        n15611), .Z(P2_U3601) );
  INV_X1 U18761 ( .A(n15596), .ZN(n15610) );
  NOR2_X1 U18762 ( .A1(n16308), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15605) );
  OAI21_X1 U18763 ( .B1(n15598), .B2(n15600), .A(n15597), .ZN(n15602) );
  NAND3_X1 U18764 ( .A1(n15600), .A2(n11319), .A3(n15599), .ZN(n15601) );
  NAND2_X1 U18765 ( .A1(n15602), .A2(n15601), .ZN(n15603) );
  OAI21_X1 U18766 ( .B1(n15605), .B2(n15604), .A(n15603), .ZN(n15606) );
  AOI21_X1 U18767 ( .B1(n12843), .B2(n15607), .A(n15606), .ZN(n16310) );
  OAI222_X1 U18768 ( .A1(n15610), .A2(n15609), .B1(n15608), .B2(n16310), .C1(
        n15860), .C2(n19412), .ZN(n15612) );
  MUX2_X1 U18769 ( .A(n16308), .B(n15612), .S(n15611), .Z(P2_U3599) );
  INV_X1 U18770 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U18771 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15613) );
  OAI21_X1 U18772 ( .B1(n17181), .B2(n17247), .A(n15613), .ZN(n15622) );
  INV_X1 U18773 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U18774 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15620) );
  INV_X1 U18775 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17130) );
  OAI22_X1 U18776 ( .A1(n17133), .A2(n17130), .B1(n15668), .B2(n17025), .ZN(
        n15618) );
  AOI22_X1 U18777 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15616) );
  AOI22_X1 U18778 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15615) );
  AOI22_X1 U18779 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15614) );
  NAND3_X1 U18780 ( .A1(n15616), .A2(n15615), .A3(n15614), .ZN(n15617) );
  AOI211_X1 U18781 ( .C1(n17030), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n15618), .B(n15617), .ZN(n15619) );
  OAI211_X1 U18782 ( .C1(n16984), .C2(n17141), .A(n15620), .B(n15619), .ZN(
        n15621) );
  AOI211_X1 U18783 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n15622), .B(n15621), .ZN(n16958) );
  AOI22_X1 U18784 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15624) );
  OAI21_X1 U18785 ( .B1(n21028), .B2(n15625), .A(n15624), .ZN(n15636) );
  INV_X1 U18786 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15634) );
  AOI22_X1 U18787 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15633) );
  INV_X1 U18788 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17167) );
  OAI22_X1 U18789 ( .A1(n12308), .A2(n17180), .B1(n17133), .B2(n17167), .ZN(
        n15631) );
  AOI22_X1 U18790 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15629) );
  AOI22_X1 U18791 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15628) );
  AOI22_X1 U18792 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15627) );
  NAND3_X1 U18793 ( .A1(n15629), .A2(n15628), .A3(n15627), .ZN(n15630) );
  AOI211_X1 U18794 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n15631), .B(n15630), .ZN(n15632) );
  OAI211_X1 U18795 ( .C1(n12307), .C2(n15634), .A(n15633), .B(n15632), .ZN(
        n15635) );
  AOI211_X1 U18796 ( .C1(n17187), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n15636), .B(n15635), .ZN(n16968) );
  AOI22_X1 U18797 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15637) );
  OAI21_X1 U18798 ( .B1(n16984), .B2(n17226), .A(n15637), .ZN(n15647) );
  AOI22_X1 U18799 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15645) );
  OAI22_X1 U18800 ( .A1(n12307), .A2(n17079), .B1(n12308), .B2(n15638), .ZN(
        n15643) );
  AOI22_X1 U18801 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15641) );
  AOI22_X1 U18802 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15640) );
  AOI22_X1 U18803 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15639) );
  NAND3_X1 U18804 ( .A1(n15641), .A2(n15640), .A3(n15639), .ZN(n15642) );
  AOI211_X1 U18805 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n15643), .B(n15642), .ZN(n15644) );
  OAI211_X1 U18806 ( .C1(n17080), .C2(n17078), .A(n15645), .B(n15644), .ZN(
        n15646) );
  AOI211_X1 U18807 ( .C1(n17187), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n15647), .B(n15646), .ZN(n16978) );
  AOI22_X1 U18808 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15648) );
  OAI21_X1 U18809 ( .B1(n17190), .B2(n17098), .A(n15648), .ZN(n15657) );
  AOI22_X1 U18810 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17030), .B1(
        n17169), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15655) );
  AOI22_X1 U18811 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17151), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17194), .ZN(n15649) );
  OAI21_X1 U18812 ( .B1(n17133), .B2(n17235), .A(n15649), .ZN(n15653) );
  AOI22_X1 U18813 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17147), .ZN(n15651) );
  AOI22_X1 U18814 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n15698), .ZN(n15650) );
  OAI211_X1 U18815 ( .C1(n15668), .C2(n17104), .A(n15651), .B(n15650), .ZN(
        n15652) );
  AOI211_X1 U18816 ( .C1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .C2(n17195), .A(
        n15653), .B(n15652), .ZN(n15654) );
  OAI211_X1 U18817 ( .C1(n17097), .C2(n17181), .A(n15655), .B(n15654), .ZN(
        n15656) );
  AOI211_X1 U18818 ( .C1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .C2(n9646), .A(
        n15657), .B(n15656), .ZN(n16979) );
  NOR2_X1 U18819 ( .A1(n16978), .A2(n16979), .ZN(n16977) );
  AOI22_X1 U18820 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15667) );
  AOI22_X1 U18821 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15666) );
  AOI22_X1 U18822 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9658), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15665) );
  OAI22_X1 U18823 ( .A1(n17133), .A2(n17063), .B1(n17215), .B2(n17189), .ZN(
        n15663) );
  AOI22_X1 U18824 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9657), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15661) );
  AOI22_X1 U18825 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15660) );
  AOI22_X1 U18826 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15659) );
  NAND2_X1 U18827 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n15658) );
  NAND4_X1 U18828 ( .A1(n15661), .A2(n15660), .A3(n15659), .A4(n15658), .ZN(
        n15662) );
  AOI211_X1 U18829 ( .C1(n9646), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n15663), .B(n15662), .ZN(n15664) );
  NAND4_X1 U18830 ( .A1(n15667), .A2(n15666), .A3(n15665), .A4(n15664), .ZN(
        n16973) );
  NAND2_X1 U18831 ( .A1(n16977), .A2(n16973), .ZN(n16972) );
  NOR2_X1 U18832 ( .A1(n16968), .A2(n16972), .ZN(n16967) );
  AOI22_X1 U18833 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9657), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15678) );
  AOI22_X1 U18834 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15677) );
  AOI22_X1 U18835 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15676) );
  OAI22_X1 U18836 ( .A1(n12307), .A2(n17160), .B1(n15668), .B2(n17034), .ZN(
        n15674) );
  AOI22_X1 U18837 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15672) );
  AOI22_X1 U18838 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15671) );
  AOI22_X1 U18839 ( .A1(n17194), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15670) );
  NAND2_X1 U18840 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n15669) );
  NAND4_X1 U18841 ( .A1(n15672), .A2(n15671), .A3(n15670), .A4(n15669), .ZN(
        n15673) );
  AOI211_X1 U18842 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n15674), .B(n15673), .ZN(n15675) );
  NAND4_X1 U18843 ( .A1(n15678), .A2(n15677), .A3(n15676), .A4(n15675), .ZN(
        n16963) );
  NAND2_X1 U18844 ( .A1(n16967), .A2(n16963), .ZN(n16962) );
  NOR2_X1 U18845 ( .A1(n16958), .A2(n16962), .ZN(n16957) );
  INV_X1 U18846 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15697) );
  AOI22_X1 U18847 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15688) );
  AOI22_X1 U18848 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U18849 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15679) );
  OAI211_X1 U18850 ( .C1(n17172), .C2(n17008), .A(n15680), .B(n15679), .ZN(
        n15686) );
  AOI22_X1 U18851 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9657), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15684) );
  AOI22_X1 U18852 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15683) );
  AOI22_X1 U18853 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15682) );
  NAND2_X1 U18854 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n15681) );
  NAND4_X1 U18855 ( .A1(n15684), .A2(n15683), .A3(n15682), .A4(n15681), .ZN(
        n15685) );
  AOI211_X1 U18856 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n15686), .B(n15685), .ZN(n15687) );
  OAI211_X1 U18857 ( .C1(n12307), .C2(n15697), .A(n15688), .B(n15687), .ZN(
        n15689) );
  NAND2_X1 U18858 ( .A1(n16957), .A2(n15689), .ZN(n16950) );
  OAI21_X1 U18859 ( .B1(n16957), .B2(n15689), .A(n16950), .ZN(n17290) );
  NOR3_X1 U18860 ( .A1(n17365), .A2(n15735), .A3(n15690), .ZN(n15691) );
  INV_X1 U18861 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16913) );
  INV_X1 U18862 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16912) );
  INV_X1 U18863 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16623) );
  INV_X1 U18864 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16641) );
  INV_X1 U18865 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17011) );
  INV_X1 U18866 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17059) );
  INV_X1 U18867 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17076) );
  INV_X1 U18868 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17268) );
  INV_X1 U18869 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17262) );
  NOR2_X1 U18870 ( .A1(n17268), .A2(n17262), .ZN(n17245) );
  AND4_X1 U18871 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .A4(n17245), .ZN(n15693) );
  INV_X1 U18872 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16821) );
  INV_X1 U18873 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17231) );
  NAND4_X1 U18874 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n17091) );
  NOR4_X1 U18875 ( .A1(n16821), .A2(n17231), .A3(n17240), .A4(n17091), .ZN(
        n15694) );
  AND4_X1 U18876 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(P3_EBX_REG_12__SCAN_IN), .ZN(n17092)
         );
  NAND4_X1 U18877 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n15693), .A3(n15694), 
        .A4(n17092), .ZN(n17073) );
  NOR2_X1 U18878 ( .A1(n17076), .A2(n17073), .ZN(n17072) );
  NAND2_X1 U18879 ( .A1(n17269), .A2(n17072), .ZN(n17058) );
  NAND2_X1 U18880 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17057), .ZN(n17045) );
  NOR2_X1 U18881 ( .A1(n17365), .A2(n17045), .ZN(n17016) );
  NAND2_X1 U18882 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17016), .ZN(n17015) );
  NAND2_X1 U18883 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16983), .ZN(n16976) );
  NAND2_X1 U18884 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16982), .ZN(n16966) );
  NAND2_X1 U18885 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16971), .ZN(n16956) );
  NOR3_X1 U18886 ( .A1(n16913), .A2(n16912), .A3(n16956), .ZN(n16952) );
  NOR2_X1 U18887 ( .A1(n17266), .A2(n16952), .ZN(n16948) );
  NOR2_X1 U18888 ( .A1(n16912), .A2(n16956), .ZN(n16961) );
  AOI22_X1 U18889 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16948), .B1(n16961), 
        .B2(n16913), .ZN(n15692) );
  OAI21_X1 U18890 ( .B1(n17290), .B2(n17256), .A(n15692), .ZN(P3_U2675) );
  NAND2_X1 U18891 ( .A1(n17269), .A2(n15693), .ZN(n17239) );
  NOR2_X1 U18892 ( .A1(n17365), .A2(n17239), .ZN(n17249) );
  NAND3_X1 U18893 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n15694), .A3(n17249), 
        .ZN(n17144) );
  AOI22_X1 U18894 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15695) );
  OAI21_X1 U18895 ( .B1(n21028), .B2(n17003), .A(n15695), .ZN(n15706) );
  AOI22_X1 U18896 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15704) );
  AOI22_X1 U18897 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9659), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15696) );
  OAI21_X1 U18898 ( .B1(n10260), .B2(n15697), .A(n15696), .ZN(n15702) );
  AOI22_X1 U18899 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15700) );
  AOI22_X1 U18900 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15699) );
  OAI211_X1 U18901 ( .C1(n17215), .C2(n17242), .A(n15700), .B(n15699), .ZN(
        n15701) );
  AOI211_X1 U18902 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n15702), .B(n15701), .ZN(n15703) );
  OAI211_X1 U18903 ( .C1(n16984), .C2(n17008), .A(n15704), .B(n15703), .ZN(
        n15705) );
  AOI211_X1 U18904 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n15706), .B(n15705), .ZN(n17366) );
  NAND3_X1 U18905 ( .A1(n17144), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n17260), 
        .ZN(n15707) );
  OAI221_X1 U18906 ( .B1(n17144), .B2(P3_EBX_REG_13__SCAN_IN), .C1(n17256), 
        .C2(n17366), .A(n15707), .ZN(P3_U2690) );
  NAND2_X1 U18907 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18446) );
  INV_X1 U18908 ( .A(n15708), .ZN(n18879) );
  NOR2_X1 U18909 ( .A1(n18879), .A2(n17805), .ZN(n15710) );
  AOI221_X1 U18910 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18446), .C1(n15710), 
        .C2(n18446), .A(n15709), .ZN(n18230) );
  NOR2_X1 U18911 ( .A1(n15711), .A2(n18693), .ZN(n15713) );
  OAI21_X1 U18912 ( .B1(n15713), .B2(n15712), .A(n18231), .ZN(n18228) );
  AOI22_X1 U18913 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18230), .B1(
        n18228), .B2(n18698), .ZN(P3_U2865) );
  NOR2_X1 U18914 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18833), .ZN(n18236) );
  AND2_X1 U18915 ( .A1(n18708), .A2(n15714), .ZN(n15723) );
  NAND2_X1 U18916 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18885) );
  INV_X1 U18917 ( .A(n18885), .ZN(n18751) );
  INV_X2 U18918 ( .A(n18894), .ZN(n18893) );
  OAI211_X1 U18919 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18758), .B(n18822), .ZN(n18882) );
  NOR4_X1 U18920 ( .A1(n18751), .A2(n16517), .A3(n17427), .A4(n18882), .ZN(
        n15722) );
  OAI21_X1 U18921 ( .B1(n15719), .B2(n15718), .A(n15717), .ZN(n15721) );
  NAND2_X1 U18922 ( .A1(n15721), .A2(n15720), .ZN(n15732) );
  NOR4_X2 U18923 ( .A1(n15723), .A2(n15865), .A3(n15722), .A4(n15732), .ZN(
        n18696) );
  INV_X1 U18924 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18226) );
  OAI22_X1 U18925 ( .A1(n18696), .A2(n18732), .B1(n18226), .B2(n18831), .ZN(
        n15724) );
  AOI21_X1 U18926 ( .B1(n15726), .B2(n18719), .A(n15725), .ZN(n18714) );
  NAND3_X1 U18927 ( .A1(n18864), .A2(n18862), .A3(n18714), .ZN(n15727) );
  OAI21_X1 U18928 ( .B1(n18864), .B2(n18719), .A(n15727), .ZN(P3_U3284) );
  INV_X1 U18929 ( .A(n15728), .ZN(n15734) );
  OAI21_X1 U18930 ( .B1(n18244), .B2(n16544), .A(n18882), .ZN(n15729) );
  OAI21_X1 U18931 ( .B1(n15730), .B2(n15729), .A(n18885), .ZN(n16521) );
  NOR3_X1 U18932 ( .A1(n15731), .A2(n16517), .A3(n16521), .ZN(n15733) );
  OAI21_X1 U18933 ( .B1(n15736), .B2(n15735), .A(n18708), .ZN(n15737) );
  NOR2_X2 U18934 ( .A1(n17394), .A2(n18221), .ZN(n18133) );
  INV_X1 U18935 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16394) );
  NOR2_X1 U18936 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n10010), .ZN(
        n15739) );
  AOI21_X1 U18937 ( .B1(n15740), .B2(n16413), .A(n15739), .ZN(n15741) );
  XOR2_X1 U18938 ( .A(n16394), .B(n15741), .Z(n16390) );
  NOR2_X1 U18939 ( .A1(n18664), .A2(n18707), .ZN(n18072) );
  INV_X1 U18940 ( .A(n18072), .ZN(n18102) );
  INV_X1 U18941 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17921) );
  NAND2_X1 U18942 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18146) );
  NOR2_X1 U18943 ( .A1(n18177), .A2(n18146), .ZN(n18009) );
  AOI21_X1 U18944 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18188) );
  INV_X1 U18945 ( .A(n18188), .ZN(n18163) );
  NAND2_X1 U18946 ( .A1(n18009), .A2(n18163), .ZN(n18125) );
  NAND3_X1 U18947 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15743) );
  NOR2_X1 U18948 ( .A1(n18125), .A2(n15743), .ZN(n18025) );
  NAND2_X1 U18949 ( .A1(n16406), .A2(n18025), .ZN(n18004) );
  INV_X1 U18950 ( .A(n18004), .ZN(n17964) );
  NAND2_X1 U18951 ( .A1(n15742), .A2(n17964), .ZN(n15752) );
  INV_X1 U18952 ( .A(n15752), .ZN(n17946) );
  NAND2_X1 U18953 ( .A1(n17905), .A2(n17946), .ZN(n17926) );
  OAI21_X1 U18954 ( .B1(n17921), .B2(n17926), .A(n18707), .ZN(n17909) );
  INV_X1 U18955 ( .A(n15742), .ZN(n16408) );
  NAND3_X1 U18956 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18009), .ZN(n18123) );
  NOR2_X1 U18957 ( .A1(n15743), .A2(n18123), .ZN(n18023) );
  NAND2_X1 U18958 ( .A1(n16406), .A2(n18023), .ZN(n18003) );
  NOR2_X1 U18959 ( .A1(n16408), .A2(n18003), .ZN(n17907) );
  NAND2_X1 U18960 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17907), .ZN(
        n15744) );
  NAND2_X1 U18961 ( .A1(n9777), .A2(n17929), .ZN(n16370) );
  INV_X1 U18962 ( .A(n16370), .ZN(n15753) );
  NAND2_X1 U18963 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15753), .ZN(
        n16407) );
  OAI21_X1 U18964 ( .B1(n15744), .B2(n16407), .A(n18687), .ZN(n15747) );
  AOI21_X1 U18965 ( .B1(n17907), .B2(n15753), .A(n18689), .ZN(n15745) );
  INV_X1 U18966 ( .A(n15745), .ZN(n15746) );
  NAND3_X1 U18967 ( .A1(n17909), .A2(n15747), .A3(n15746), .ZN(n15847) );
  AOI21_X1 U18968 ( .B1(n9880), .B2(n18102), .A(n15847), .ZN(n16409) );
  INV_X1 U18969 ( .A(n18167), .ZN(n18122) );
  NAND2_X1 U18970 ( .A1(n18122), .A2(n16416), .ZN(n15749) );
  INV_X2 U18971 ( .A(n18108), .ZN(n18210) );
  NOR2_X1 U18972 ( .A1(n18187), .A2(n18126), .ZN(n18209) );
  INV_X1 U18973 ( .A(n16415), .ZN(n18713) );
  NAND2_X1 U18974 ( .A1(n18215), .A2(n17940), .ZN(n18059) );
  OAI22_X1 U18975 ( .A1(n16377), .A2(n18223), .B1(n16386), .B2(n18059), .ZN(
        n15748) );
  NOR2_X1 U18976 ( .A1(n18084), .A2(n15748), .ZN(n15848) );
  OAI221_X1 U18977 ( .B1(n18126), .B2(n16409), .C1(n18126), .C2(n15749), .A(
        n15848), .ZN(n15755) );
  INV_X1 U18978 ( .A(n17545), .ZN(n17906) );
  NAND2_X1 U18979 ( .A1(n16372), .A2(n17906), .ZN(n16412) );
  INV_X1 U18980 ( .A(n18059), .ZN(n18134) );
  NOR2_X1 U18981 ( .A1(n17912), .A2(n15750), .ZN(n16410) );
  NAND2_X1 U18982 ( .A1(n18134), .A2(n16410), .ZN(n15754) );
  OAI221_X1 U18983 ( .B1(n18664), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n18664), .C2(n18687), .A(n17907), .ZN(n15751) );
  OAI21_X1 U18984 ( .B1(n18190), .B2(n15752), .A(n15751), .ZN(n17928) );
  NAND4_X1 U18985 ( .A1(n18215), .A2(n16372), .A3(n15753), .A4(n17928), .ZN(
        n16392) );
  OAI211_X1 U18986 ( .C1(n18223), .C2(n16412), .A(n15754), .B(n16392), .ZN(
        n15849) );
  AOI22_X1 U18987 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15755), .B1(
        n15849), .B2(n16394), .ZN(n15756) );
  NAND2_X1 U18988 ( .A1(n18210), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16380) );
  OAI211_X1 U18989 ( .C1(n18111), .C2(n16390), .A(n15756), .B(n16380), .ZN(
        P3_U2833) );
  OAI21_X1 U18990 ( .B1(n16181), .B2(n16292), .A(n15757), .ZN(n15758) );
  AND2_X1 U18991 ( .A1(n15758), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15789) );
  INV_X1 U18992 ( .A(n15789), .ZN(n15771) );
  INV_X1 U18993 ( .A(n19245), .ZN(n15760) );
  XNOR2_X1 U18994 ( .A(n15763), .B(n15762), .ZN(n16164) );
  NOR2_X1 U18995 ( .A1(n16290), .A2(n18983), .ZN(n15768) );
  INV_X1 U18996 ( .A(n15764), .ZN(n15765) );
  OAI21_X1 U18997 ( .B1(n13628), .B2(n15766), .A(n15765), .ZN(n19120) );
  NAND2_X1 U18998 ( .A1(n15785), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16161) );
  OAI21_X1 U18999 ( .B1(n16277), .B2(n19120), .A(n16161), .ZN(n15767) );
  AOI211_X1 U19000 ( .C1(n16164), .C2(n19255), .A(n15768), .B(n15767), .ZN(
        n15769) );
  OAI221_X1 U19001 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15771), 
        .C1(n15770), .C2(n15786), .A(n15769), .ZN(P2_U3030) );
  AOI22_X1 U19002 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19095), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19102), .ZN(n15783) );
  INV_X1 U19003 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15772) );
  OAI22_X1 U19004 ( .A1(n15773), .A2(n19099), .B1(n19082), .B2(n15772), .ZN(
        n15774) );
  INV_X1 U19005 ( .A(n15774), .ZN(n15782) );
  OAI22_X1 U19006 ( .A1(n16148), .A2(n19107), .B1(n19098), .B2(n15775), .ZN(
        n15776) );
  INV_X1 U19007 ( .A(n15776), .ZN(n15781) );
  AOI21_X1 U19008 ( .B1(n15778), .B2(n9766), .A(n15777), .ZN(n15779) );
  NAND2_X1 U19009 ( .A1(n19089), .A2(n15779), .ZN(n15780) );
  NAND4_X1 U19010 ( .A1(n15783), .A2(n15782), .A3(n15781), .A4(n15780), .ZN(
        P2_U2833) );
  INV_X1 U19011 ( .A(n15784), .ZN(n18972) );
  AOI222_X1 U19012 ( .A1(P2_REIP_REG_17__SCAN_IN), .A2(n15785), .B1(n19262), 
        .B2(n18972), .C1(n19248), .C2(n18974), .ZN(n15791) );
  OAI211_X1 U19013 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15787), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n15786), .ZN(n15788) );
  OAI221_X1 U19014 ( .B1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n15789), .A(n15788), .ZN(
        n15790) );
  OAI211_X1 U19015 ( .C1(n15792), .C2(n16273), .A(n15791), .B(n15790), .ZN(
        P2_U3029) );
  AOI22_X1 U19016 ( .A1(n9664), .A2(n15794), .B1(n15793), .B2(n10275), .ZN(
        n20799) );
  INV_X1 U19017 ( .A(n15795), .ZN(n15796) );
  NAND2_X1 U19018 ( .A1(n15796), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n20808) );
  AND3_X1 U19019 ( .A1(n20799), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        n20808), .ZN(n15801) );
  AOI211_X1 U19020 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n15801), .A(
        n15798), .B(n15797), .ZN(n15799) );
  INV_X1 U19021 ( .A(n15799), .ZN(n15800) );
  OAI21_X1 U19022 ( .B1(n15801), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15800), .ZN(n15802) );
  AOI222_X1 U19023 ( .A1(n11119), .A2(n15803), .B1(n11119), .B2(n15802), .C1(
        n15803), .C2(n15802), .ZN(n15805) );
  AOI21_X1 U19024 ( .B1(n15805), .B2(n15804), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15807) );
  NOR2_X1 U19025 ( .A1(n15805), .A2(n15804), .ZN(n15806) );
  OAI21_X1 U19026 ( .B1(n15807), .B2(n15806), .A(n20182), .ZN(n15817) );
  NAND2_X1 U19027 ( .A1(n20968), .A2(n20944), .ZN(n15812) );
  INV_X1 U19028 ( .A(n15808), .ZN(n15809) );
  OR3_X1 U19029 ( .A1(n15810), .A2(n15809), .A3(n16039), .ZN(n15811) );
  AOI21_X1 U19030 ( .B1(n15813), .B2(n15812), .A(n15811), .ZN(n15815) );
  NAND4_X1 U19031 ( .A1(n15817), .A2(n15816), .A3(n15815), .A4(n15814), .ZN(
        n15826) );
  NAND2_X1 U19032 ( .A1(n15818), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n15825) );
  NOR3_X1 U19033 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20728), .A3(n20738), 
        .ZN(n15821) );
  OAI22_X1 U19034 ( .A1(n15822), .A2(n15821), .B1(n15820), .B2(n15819), .ZN(
        n16044) );
  AOI21_X1 U19035 ( .B1(n15826), .B2(n15823), .A(n16044), .ZN(n16040) );
  AOI211_X1 U19036 ( .C1(n15826), .C2(n15825), .A(n15824), .B(n16040), .ZN(
        n15832) );
  AOI21_X1 U19037 ( .B1(n20731), .B2(n20728), .A(n15827), .ZN(n16041) );
  AOI21_X1 U19038 ( .B1(n15829), .B2(n15828), .A(n16040), .ZN(n15830) );
  INV_X1 U19039 ( .A(n15830), .ZN(n15831) );
  AOI22_X1 U19040 ( .A1(n15832), .A2(n16041), .B1(n16039), .B2(n15831), .ZN(
        P1_U3161) );
  INV_X1 U19041 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20899) );
  NOR2_X1 U19042 ( .A1(n20073), .A2(n20899), .ZN(n15833) );
  AOI221_X1 U19043 ( .B1(n15836), .B2(n15835), .C1(n15834), .C2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(n15833), .ZN(n15842) );
  INV_X1 U19044 ( .A(n15837), .ZN(n15840) );
  INV_X1 U19045 ( .A(n15838), .ZN(n15839) );
  AOI22_X1 U19046 ( .A1(n15840), .A2(n16033), .B1(n16032), .B2(n15839), .ZN(
        n15841) );
  NAND2_X1 U19047 ( .A1(n15842), .A2(n15841), .ZN(P1_U3010) );
  XNOR2_X1 U19048 ( .A(n15844), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16375) );
  NAND2_X1 U19049 ( .A1(n18679), .A2(n18190), .ZN(n18204) );
  OAI21_X1 U19050 ( .B1(n18664), .B2(n18204), .A(n18215), .ZN(n18203) );
  INV_X1 U19051 ( .A(n18203), .ZN(n15845) );
  AOI22_X1 U19052 ( .A1(n18215), .A2(n15847), .B1(n15846), .B2(n15845), .ZN(
        n16391) );
  NAND2_X1 U19053 ( .A1(n16391), .A2(n15848), .ZN(n15850) );
  NOR2_X1 U19054 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16394), .ZN(
        n16371) );
  AOI22_X1 U19055 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15850), .B1(
        n16371), .B2(n15849), .ZN(n15851) );
  NAND2_X1 U19056 ( .A1(n18210), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16362) );
  OAI211_X1 U19057 ( .C1(n16375), .C2(n18111), .A(n15851), .B(n16362), .ZN(
        P3_U2832) );
  INV_X1 U19058 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20745) );
  OAI221_X1 U19059 ( .B1(n20731), .B2(HOLD), .C1(n20731), .C2(n20745), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n15854) );
  INV_X1 U19060 ( .A(HOLD), .ZN(n20976) );
  OAI211_X1 U19061 ( .C1(n20745), .C2(n20976), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15852) );
  NAND3_X1 U19062 ( .A1(n15854), .A2(n15853), .A3(n15852), .ZN(P1_U3195) );
  AND2_X1 U19063 ( .A1(n15855), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19064 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15856) );
  NOR2_X1 U19065 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16349) );
  NOR2_X1 U19066 ( .A1(n19986), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19849) );
  AND2_X1 U19067 ( .A1(n19985), .A2(n19849), .ZN(n16343) );
  NOR4_X1 U19068 ( .A1(n15856), .A2(n16349), .A3(n16358), .A4(n16343), .ZN(
        P2_U3178) );
  INV_X1 U19069 ( .A(n16349), .ZN(n15858) );
  NAND2_X1 U19070 ( .A1(n15858), .A2(n15857), .ZN(n15859) );
  AOI221_X1 U19071 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16358), .C1(n19970), .C2(
        n16358), .A(n19781), .ZN(n19967) );
  INV_X1 U19072 ( .A(n19967), .ZN(n19964) );
  NOR2_X1 U19073 ( .A1(n15862), .A2(n19964), .ZN(P2_U3047) );
  NOR3_X1 U19074 ( .A1(n15863), .A2(n17428), .A3(n16544), .ZN(n15864) );
  NAND2_X1 U19075 ( .A1(n18268), .A2(n17270), .ZN(n17421) );
  INV_X1 U19076 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17500) );
  NOR2_X2 U19077 ( .A1(n15867), .A2(n15866), .ZN(n17419) );
  AOI22_X1 U19078 ( .A1(n17420), .A2(BUF2_REG_0__SCAN_IN), .B1(n17419), .B2(
        n15868), .ZN(n15869) );
  OAI221_X1 U19079 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17421), .C1(n17500), 
        .C2(n17270), .A(n15869), .ZN(P3_U2735) );
  AOI22_X1 U19080 ( .A1(n20077), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20051), .ZN(n15879) );
  AOI21_X1 U19081 ( .B1(n20049), .B2(n15870), .A(n9645), .ZN(n15878) );
  OAI22_X1 U19082 ( .A1(n15935), .A2(n15914), .B1(n20084), .B2(n15871), .ZN(
        n15872) );
  INV_X1 U19083 ( .A(n15872), .ZN(n15877) );
  NOR2_X1 U19084 ( .A1(n20767), .A2(n15988), .ZN(n15874) );
  OAI221_X1 U19085 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15875), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(n15874), .A(n15873), .ZN(n15876) );
  NAND4_X1 U19086 ( .A1(n15879), .A2(n15878), .A3(n15877), .A4(n15876), .ZN(
        P1_U2823) );
  NOR2_X1 U19087 ( .A1(n15881), .A2(n15880), .ZN(n15882) );
  OR2_X1 U19088 ( .A1(n15883), .A2(n15882), .ZN(n15989) );
  INV_X1 U19089 ( .A(n15989), .ZN(n15930) );
  AOI22_X1 U19090 ( .A1(n20049), .A2(n15944), .B1(n20053), .B2(n15930), .ZN(
        n15889) );
  AOI21_X1 U19091 ( .B1(n20051), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n9645), .ZN(n15885) );
  NAND2_X1 U19092 ( .A1(n20077), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n15884) );
  OAI211_X1 U19093 ( .C1(n15893), .C2(n15988), .A(n15885), .B(n15884), .ZN(
        n15886) );
  AOI21_X1 U19094 ( .B1(n15945), .B2(n20055), .A(n15886), .ZN(n15888) );
  NAND3_X1 U19095 ( .A1(n15889), .A2(n15888), .A3(n15887), .ZN(P1_U2825) );
  INV_X1 U19096 ( .A(n15890), .ZN(n15891) );
  AOI22_X1 U19097 ( .A1(n20049), .A2(n15891), .B1(n20077), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n15899) );
  AOI22_X1 U19098 ( .A1(n16002), .A2(n20053), .B1(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n20051), .ZN(n15898) );
  INV_X1 U19099 ( .A(n15908), .ZN(n15892) );
  AOI21_X1 U19100 ( .B1(n15892), .B2(P1_REIP_REG_13__SCAN_IN), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15894) );
  NOR2_X1 U19101 ( .A1(n15894), .A2(n15893), .ZN(n15895) );
  AOI21_X1 U19102 ( .B1(n15896), .B2(n20055), .A(n15895), .ZN(n15897) );
  NAND4_X1 U19103 ( .A1(n15899), .A2(n15898), .A3(n15897), .A4(n20073), .ZN(
        P1_U2826) );
  OAI222_X1 U19104 ( .A1(n15902), .A2(n20087), .B1(n15901), .B2(n20084), .C1(
        n20038), .C2(n15900), .ZN(n15903) );
  AOI211_X1 U19105 ( .C1(n20051), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n9645), .B(n15903), .ZN(n15907) );
  AOI22_X1 U19106 ( .A1(n15905), .A2(n20055), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n15904), .ZN(n15906) );
  OAI211_X1 U19107 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n15908), .A(n15907), 
        .B(n15906), .ZN(P1_U2827) );
  NAND2_X1 U19108 ( .A1(n15910), .A2(n15909), .ZN(n15928) );
  AOI22_X1 U19109 ( .A1(n16011), .A2(n20053), .B1(n20077), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15911) );
  OAI211_X1 U19110 ( .C1(n20075), .C2(n15912), .A(n15911), .B(n20073), .ZN(
        n15917) );
  OAI22_X1 U19111 ( .A1(n15915), .A2(n15914), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n15913), .ZN(n15916) );
  AOI211_X1 U19112 ( .C1(n15918), .C2(n20049), .A(n15917), .B(n15916), .ZN(
        n15919) );
  OAI21_X1 U19113 ( .B1(n15920), .B2(n15928), .A(n15919), .ZN(P1_U2829) );
  OAI222_X1 U19114 ( .A1(n15923), .A2(n20087), .B1(n15922), .B2(n20084), .C1(
        n20038), .C2(n15921), .ZN(n15924) );
  AOI211_X1 U19115 ( .C1(n20051), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n9645), .B(n15924), .ZN(n15927) );
  AOI22_X1 U19116 ( .A1(n15951), .A2(n20055), .B1(n15929), .B2(n15925), .ZN(
        n15926) );
  OAI211_X1 U19117 ( .C1(n15929), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        P1_U2830) );
  AOI22_X1 U19118 ( .A1(n15945), .A2(n20099), .B1(n20098), .B2(n15930), .ZN(
        n15931) );
  OAI21_X1 U19119 ( .B1(n20103), .B2(n15932), .A(n15931), .ZN(P1_U2857) );
  AOI22_X1 U19120 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16031), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15938) );
  OAI22_X1 U19121 ( .A1(n15935), .A2(n15934), .B1(n15933), .B2(n15963), .ZN(
        n15936) );
  INV_X1 U19122 ( .A(n15936), .ZN(n15937) );
  OAI211_X1 U19123 ( .C1(n20007), .C2(n15939), .A(n15938), .B(n15937), .ZN(
        P1_U2982) );
  NAND2_X1 U19124 ( .A1(n15941), .A2(n15940), .ZN(n15942) );
  AOI22_X1 U19125 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n9645), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15947) );
  AOI22_X1 U19126 ( .A1(n15945), .A2(n15960), .B1(n15950), .B2(n15944), .ZN(
        n15946) );
  OAI211_X1 U19127 ( .C1(n15993), .C2(n20007), .A(n15947), .B(n15946), .ZN(
        P1_U2984) );
  AOI22_X1 U19128 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16031), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n15953) );
  AOI22_X1 U19129 ( .A1(n15951), .A2(n15960), .B1(n15950), .B2(n15949), .ZN(
        n15952) );
  OAI211_X1 U19130 ( .C1(n20007), .C2(n15954), .A(n15953), .B(n15952), .ZN(
        P1_U2989) );
  AOI22_X1 U19131 ( .A1(n15948), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16031), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15962) );
  NAND2_X1 U19132 ( .A1(n15957), .A2(n15956), .ZN(n15958) );
  XNOR2_X1 U19133 ( .A(n15955), .B(n15958), .ZN(n16034) );
  AOI22_X1 U19134 ( .A1(n20100), .A2(n15960), .B1(n16034), .B2(n15959), .ZN(
        n15961) );
  OAI211_X1 U19135 ( .C1(n15963), .C2(n20034), .A(n15962), .B(n15961), .ZN(
        P1_U2992) );
  OAI222_X1 U19136 ( .A1(n15967), .A2(n20173), .B1(n15966), .B2(n15965), .C1(
        n20164), .C2(n15964), .ZN(n15968) );
  INV_X1 U19137 ( .A(n15968), .ZN(n15970) );
  NAND2_X1 U19138 ( .A1(n9645), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15969) );
  OAI211_X1 U19139 ( .C1(n15972), .C2(n15971), .A(n15970), .B(n15969), .ZN(
        P1_U3012) );
  OAI22_X1 U19140 ( .A1(n15974), .A2(n20164), .B1(n20173), .B2(n15973), .ZN(
        n15975) );
  AOI21_X1 U19141 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15976), .A(
        n15975), .ZN(n15980) );
  NAND3_X1 U19142 ( .A1(n15978), .A2(n15991), .A3(n15977), .ZN(n15979) );
  OAI211_X1 U19143 ( .C1(n20770), .C2(n20073), .A(n15980), .B(n15979), .ZN(
        P1_U3013) );
  OAI222_X1 U19144 ( .A1(n15982), .A2(n20173), .B1(n20073), .B2(n20767), .C1(
        n20164), .C2(n15981), .ZN(n15983) );
  INV_X1 U19145 ( .A(n15983), .ZN(n15986) );
  OAI211_X1 U19146 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15991), .B(n15984), .ZN(
        n15985) );
  OAI211_X1 U19147 ( .C1(n15997), .C2(n15987), .A(n15986), .B(n15985), .ZN(
        P1_U3015) );
  OAI22_X1 U19148 ( .A1(n15989), .A2(n20173), .B1(n15988), .B2(n20073), .ZN(
        n15990) );
  AOI21_X1 U19149 ( .B1(n15991), .B2(n15996), .A(n15990), .ZN(n15992) );
  OAI21_X1 U19150 ( .B1(n15993), .B2(n20164), .A(n15992), .ZN(n15994) );
  INV_X1 U19151 ( .A(n15994), .ZN(n15995) );
  OAI21_X1 U19152 ( .B1(n15997), .B2(n15996), .A(n15995), .ZN(P1_U3016) );
  NAND2_X1 U19153 ( .A1(n15999), .A2(n15998), .ZN(n16016) );
  NAND4_X1 U19154 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n16000), .ZN(n16008) );
  AOI21_X1 U19155 ( .B1(n16002), .B2(n16032), .A(n16001), .ZN(n16007) );
  INV_X1 U19156 ( .A(n16003), .ZN(n16005) );
  AOI22_X1 U19157 ( .A1(n16005), .A2(n16033), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16004), .ZN(n16006) );
  OAI211_X1 U19158 ( .C1(n16016), .C2(n16008), .A(n16007), .B(n16006), .ZN(
        P1_U3017) );
  INV_X1 U19159 ( .A(n16009), .ZN(n16010) );
  AOI21_X1 U19160 ( .B1(n16011), .B2(n16032), .A(n16010), .ZN(n16015) );
  AOI22_X1 U19161 ( .A1(n16013), .A2(n16033), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16012), .ZN(n16014) );
  OAI211_X1 U19162 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16016), .A(
        n16015), .B(n16014), .ZN(P1_U3020) );
  INV_X1 U19163 ( .A(n16017), .ZN(n16023) );
  AOI21_X1 U19164 ( .B1(n16032), .B2(n9757), .A(n16018), .ZN(n16022) );
  AOI22_X1 U19165 ( .A1(n16020), .A2(n16033), .B1(n13971), .B2(n16019), .ZN(
        n16021) );
  OAI211_X1 U19166 ( .C1(n16023), .C2(n13971), .A(n16022), .B(n16021), .ZN(
        P1_U3022) );
  INV_X1 U19167 ( .A(n16024), .ZN(n16025) );
  NAND2_X1 U19168 ( .A1(n16026), .A2(n16025), .ZN(n16029) );
  INV_X1 U19169 ( .A(n16027), .ZN(n16028) );
  AOI21_X1 U19170 ( .B1(n16030), .B2(n16029), .A(n16028), .ZN(n20097) );
  AOI22_X1 U19171 ( .A1(n16032), .A2(n20097), .B1(n16031), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16037) );
  AOI22_X1 U19172 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n16035), .B1(
        n16034), .B2(n16033), .ZN(n16036) );
  OAI211_X1 U19173 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16038), .A(
        n16037), .B(n16036), .ZN(P1_U3024) );
  OAI221_X1 U19174 ( .B1(n20738), .B2(n16039), .C1(P1_STATEBS16_REG_SCAN_IN), 
        .C2(P1_STATE2_REG_0__SCAN_IN), .A(P1_STATE2_REG_1__SCAN_IN), .ZN(
        n20729) );
  INV_X1 U19175 ( .A(n20729), .ZN(n16043) );
  NOR2_X1 U19176 ( .A1(n16040), .A2(n16039), .ZN(n20727) );
  AOI21_X1 U19177 ( .B1(n20727), .B2(n16041), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n16042) );
  AOI221_X1 U19178 ( .B1(n20726), .B2(n16044), .C1(n16043), .C2(n16044), .A(
        n16042), .ZN(P1_U3162) );
  OAI21_X1 U19179 ( .B1(n20727), .B2(n13115), .A(n16045), .ZN(P1_U3466) );
  INV_X1 U19180 ( .A(n16046), .ZN(n16048) );
  AOI22_X1 U19181 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19095), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19102), .ZN(n16047) );
  OAI21_X1 U19182 ( .B1(n16048), .B2(n19099), .A(n16047), .ZN(n16049) );
  AOI21_X1 U19183 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19096), .A(n16049), .ZN(
        n16056) );
  NOR2_X1 U19184 ( .A1(n19021), .A2(n16058), .ZN(n16051) );
  XNOR2_X1 U19185 ( .A(n16051), .B(n16050), .ZN(n16054) );
  AOI21_X1 U19186 ( .B1(n16054), .B2(n19089), .A(n16053), .ZN(n16055) );
  OAI211_X1 U19187 ( .C1(n16057), .C2(n19098), .A(n16056), .B(n16055), .ZN(
        P2_U2825) );
  AOI21_X1 U19188 ( .B1(n16060), .B2(n16059), .A(n16058), .ZN(n16068) );
  INV_X1 U19189 ( .A(n16061), .ZN(n16064) );
  AOI22_X1 U19190 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19096), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19102), .ZN(n16062) );
  OAI21_X1 U19191 ( .B1(n10125), .B2(n19093), .A(n16062), .ZN(n16063) );
  AOI21_X1 U19192 ( .B1(n16064), .B2(n19076), .A(n16063), .ZN(n16065) );
  OAI21_X1 U19193 ( .B1(n16066), .B2(n19099), .A(n16065), .ZN(n16067) );
  AOI21_X1 U19194 ( .B1(n19089), .B2(n16068), .A(n16067), .ZN(n16069) );
  OAI21_X1 U19195 ( .B1(n16070), .B2(n19098), .A(n16069), .ZN(P2_U2826) );
  AOI211_X1 U19196 ( .C1(n16073), .C2(n16072), .A(n16071), .B(n19851), .ZN(
        n16080) );
  AOI22_X1 U19197 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19096), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19102), .ZN(n16074) );
  OAI21_X1 U19198 ( .B1(n10124), .B2(n19093), .A(n16074), .ZN(n16075) );
  AOI21_X1 U19199 ( .B1(n16076), .B2(n19076), .A(n16075), .ZN(n16077) );
  OAI21_X1 U19200 ( .B1(n19099), .B2(n16078), .A(n16077), .ZN(n16079) );
  AOI211_X1 U19201 ( .C1(n18973), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        n16082) );
  INV_X1 U19202 ( .A(n16082), .ZN(P2_U2829) );
  OAI22_X1 U19203 ( .A1(n16084), .A2(n19099), .B1(n19093), .B2(n16083), .ZN(
        n16085) );
  INV_X1 U19204 ( .A(n16085), .ZN(n16097) );
  AOI22_X1 U19205 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19096), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19102), .ZN(n16096) );
  INV_X1 U19206 ( .A(n16086), .ZN(n16087) );
  OAI22_X1 U19207 ( .A1(n16088), .A2(n19107), .B1(n16087), .B2(n19098), .ZN(
        n16089) );
  INV_X1 U19208 ( .A(n16089), .ZN(n16095) );
  AOI21_X1 U19209 ( .B1(n16092), .B2(n16091), .A(n16090), .ZN(n16093) );
  NAND2_X1 U19210 ( .A1(n19089), .A2(n16093), .ZN(n16094) );
  NAND4_X1 U19211 ( .A1(n16097), .A2(n16096), .A3(n16095), .A4(n16094), .ZN(
        P2_U2830) );
  AOI22_X1 U19212 ( .A1(n19148), .A2(n16098), .B1(n12661), .B2(n12991), .ZN(
        P2_U2856) );
  INV_X1 U19213 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16101) );
  AOI22_X1 U19214 ( .A1(n16099), .A2(n19127), .B1(n19148), .B2(n16143), .ZN(
        n16100) );
  OAI21_X1 U19215 ( .B1(n19148), .B2(n16101), .A(n16100), .ZN(P2_U2864) );
  AOI21_X1 U19216 ( .B1(n16102), .B2(n15079), .A(n11728), .ZN(n16113) );
  INV_X1 U19217 ( .A(n16148), .ZN(n16103) );
  AOI22_X1 U19218 ( .A1(n16113), .A2(n19127), .B1(n19148), .B2(n16103), .ZN(
        n16104) );
  OAI21_X1 U19219 ( .B1(n19148), .B2(n15772), .A(n16104), .ZN(P2_U2865) );
  NOR2_X1 U19220 ( .A1(n15086), .A2(n16105), .ZN(n16106) );
  OR2_X1 U19221 ( .A1(n15078), .A2(n16106), .ZN(n16121) );
  OAI22_X1 U19222 ( .A1(n16121), .A2(n19145), .B1(n19148), .B2(n10150), .ZN(
        n16107) );
  INV_X1 U19223 ( .A(n16107), .ZN(n16108) );
  OAI21_X1 U19224 ( .B1(n12991), .B2(n18931), .A(n16108), .ZN(P2_U2867) );
  AOI21_X1 U19225 ( .B1(n16109), .B2(n13838), .A(n10237), .ZN(n16129) );
  AOI22_X1 U19226 ( .A1(n16129), .A2(n19127), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n12991), .ZN(n16110) );
  OAI21_X1 U19227 ( .B1(n12991), .B2(n18954), .A(n16110), .ZN(P2_U2869) );
  AOI22_X1 U19228 ( .A1(n16127), .A2(n16111), .B1(n19169), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16116) );
  AOI22_X1 U19229 ( .A1(n19153), .A2(BUF1_REG_22__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16115) );
  AOI22_X1 U19230 ( .A1(n16113), .A2(n19173), .B1(n19150), .B2(n16112), .ZN(
        n16114) );
  NAND3_X1 U19231 ( .A1(n16116), .A2(n16115), .A3(n16114), .ZN(P2_U2897) );
  AOI22_X1 U19232 ( .A1(n16127), .A2(n16117), .B1(n19169), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16125) );
  AOI22_X1 U19233 ( .A1(n19153), .A2(BUF1_REG_20__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16124) );
  INV_X1 U19234 ( .A(n16118), .ZN(n18930) );
  OAI22_X1 U19235 ( .A1(n16121), .A2(n16120), .B1(n16119), .B2(n18930), .ZN(
        n16122) );
  INV_X1 U19236 ( .A(n16122), .ZN(n16123) );
  NAND3_X1 U19237 ( .A1(n16125), .A2(n16124), .A3(n16123), .ZN(P2_U2899) );
  AOI22_X1 U19238 ( .A1(n16127), .A2(n16126), .B1(n19169), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16132) );
  AOI22_X1 U19239 ( .A1(n19153), .A2(BUF1_REG_18__SCAN_IN), .B1(n19152), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16131) );
  INV_X1 U19240 ( .A(n18953), .ZN(n16128) );
  AOI22_X1 U19241 ( .A1(n16129), .A2(n19173), .B1(n19150), .B2(n16128), .ZN(
        n16130) );
  NAND3_X1 U19242 ( .A1(n16132), .A2(n16131), .A3(n16130), .ZN(P2_U2901) );
  AOI22_X1 U19243 ( .A1(n16187), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n12657), .ZN(n16138) );
  OAI22_X1 U19244 ( .A1(n16134), .A2(n19224), .B1(n19223), .B2(n16133), .ZN(
        n16135) );
  AOI21_X1 U19245 ( .B1(n19227), .B2(n16136), .A(n16135), .ZN(n16137) );
  OAI211_X1 U19246 ( .C1(n16236), .C2(n16139), .A(n16138), .B(n16137), .ZN(
        P2_U2990) );
  OAI22_X1 U19247 ( .A1(n19231), .A2(n16140), .B1(n19904), .B2(n19066), .ZN(
        n16141) );
  AOI21_X1 U19248 ( .B1(n19216), .B2(n16142), .A(n16141), .ZN(n16146) );
  AOI22_X1 U19249 ( .A1(n16144), .A2(n16240), .B1(n16239), .B2(n16143), .ZN(
        n16145) );
  OAI211_X1 U19250 ( .C1(n16251), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        P2_U2991) );
  AOI22_X1 U19251 ( .A1(n16187), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n12657), .ZN(n16153) );
  OAI22_X1 U19252 ( .A1(n16149), .A2(n19224), .B1(n19223), .B2(n16148), .ZN(
        n16150) );
  AOI21_X1 U19253 ( .B1(n19227), .B2(n16151), .A(n16150), .ZN(n16152) );
  OAI211_X1 U19254 ( .C1(n16236), .C2(n16154), .A(n16153), .B(n16152), .ZN(
        P2_U2992) );
  AOI22_X1 U19255 ( .A1(n16187), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n12657), .ZN(n16159) );
  OAI222_X1 U19256 ( .A1(n16156), .A2(n16251), .B1(n16155), .B2(n19224), .C1(
        n19223), .C2(n18954), .ZN(n16157) );
  INV_X1 U19257 ( .A(n16157), .ZN(n16158) );
  OAI211_X1 U19258 ( .C1(n16236), .C2(n16160), .A(n16159), .B(n16158), .ZN(
        P2_U2996) );
  NOR2_X1 U19259 ( .A1(n18982), .A2(n16236), .ZN(n16163) );
  INV_X1 U19260 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18978) );
  OAI21_X1 U19261 ( .B1(n19231), .B2(n18978), .A(n16161), .ZN(n16162) );
  AOI211_X1 U19262 ( .C1(n16164), .C2(n16240), .A(n16163), .B(n16162), .ZN(
        n16168) );
  OAI211_X1 U19263 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16166), .A(
        n19227), .B(n16165), .ZN(n16167) );
  OAI211_X1 U19264 ( .C1(n19120), .C2(n19223), .A(n16168), .B(n16167), .ZN(
        P2_U2998) );
  AOI22_X1 U19265 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n12657), .B1(n19216), 
        .B2(n16169), .ZN(n16175) );
  INV_X1 U19266 ( .A(n16170), .ZN(n16172) );
  OAI22_X1 U19267 ( .A1(n16172), .A2(n16251), .B1(n16171), .B2(n19224), .ZN(
        n16173) );
  AOI21_X1 U19268 ( .B1(n16239), .B2(n18990), .A(n16173), .ZN(n16174) );
  OAI211_X1 U19269 ( .C1(n19231), .C2(n16176), .A(n16175), .B(n16174), .ZN(
        P2_U2999) );
  AOI22_X1 U19270 ( .A1(n16187), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n12657), .ZN(n16185) );
  NAND2_X1 U19271 ( .A1(n16178), .A2(n16177), .ZN(n16179) );
  XNOR2_X1 U19272 ( .A(n16180), .B(n16179), .ZN(n16257) );
  OAI21_X1 U19273 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16182), .A(
        n16181), .ZN(n16183) );
  INV_X1 U19274 ( .A(n16183), .ZN(n16255) );
  AOI222_X1 U19275 ( .A1(n16257), .A2(n16240), .B1(n16239), .B2(n16256), .C1(
        n16255), .C2(n19227), .ZN(n16184) );
  OAI211_X1 U19276 ( .C1(n16236), .C2(n16186), .A(n16185), .B(n16184), .ZN(
        P2_U3000) );
  AOI22_X1 U19277 ( .A1(n16187), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n12657), .ZN(n16191) );
  AOI222_X1 U19278 ( .A1(n16189), .A2(n16240), .B1(n16239), .B2(n19126), .C1(
        n16188), .C2(n19227), .ZN(n16190) );
  OAI211_X1 U19279 ( .C1(n16236), .C2(n16192), .A(n16191), .B(n16190), .ZN(
        P2_U3002) );
  AOI22_X1 U19280 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n12657), .B1(n19216), 
        .B2(n19023), .ZN(n16197) );
  OAI22_X1 U19281 ( .A1(n16194), .A2(n16251), .B1(n16193), .B2(n19224), .ZN(
        n16195) );
  AOI21_X1 U19282 ( .B1(n16239), .B2(n19024), .A(n16195), .ZN(n16196) );
  OAI211_X1 U19283 ( .C1(n19231), .C2(n19017), .A(n16197), .B(n16196), .ZN(
        P2_U3003) );
  AOI22_X1 U19284 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n12657), .B1(n19216), 
        .B2(n19033), .ZN(n16212) );
  AOI21_X1 U19285 ( .B1(n16200), .B2(n16199), .A(n16198), .ZN(n16270) );
  NAND2_X1 U19286 ( .A1(n16202), .A2(n16201), .ZN(n16206) );
  NAND2_X1 U19287 ( .A1(n16204), .A2(n16203), .ZN(n16205) );
  XOR2_X1 U19288 ( .A(n16206), .B(n16205), .Z(n16274) );
  NOR2_X1 U19289 ( .A1(n16207), .A2(n9759), .ZN(n16208) );
  OR2_X1 U19290 ( .A1(n16209), .A2(n16208), .ZN(n19038) );
  OAI22_X1 U19291 ( .A1(n16274), .A2(n19224), .B1(n19223), .B2(n19038), .ZN(
        n16210) );
  AOI21_X1 U19292 ( .B1(n19227), .B2(n16270), .A(n16210), .ZN(n16211) );
  OAI211_X1 U19293 ( .C1(n19231), .C2(n16213), .A(n16212), .B(n16211), .ZN(
        P2_U3004) );
  OAI22_X1 U19294 ( .A1(n19231), .A2(n12587), .B1(n16236), .B2(n19047), .ZN(
        n16214) );
  AOI21_X1 U19295 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n12657), .A(n16214), .ZN(
        n16218) );
  AOI22_X1 U19296 ( .A1(n16216), .A2(n16240), .B1(n16239), .B2(n16215), .ZN(
        n16217) );
  OAI211_X1 U19297 ( .C1(n16251), .C2(n16219), .A(n16218), .B(n16217), .ZN(
        P2_U3005) );
  AOI22_X1 U19298 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n15785), .B1(n19216), 
        .B2(n16220), .ZN(n16234) );
  OAI21_X1 U19299 ( .B1(n16223), .B2(n16222), .A(n16221), .ZN(n16278) );
  NAND2_X1 U19300 ( .A1(n15572), .A2(n16224), .ZN(n16229) );
  INV_X1 U19301 ( .A(n16225), .ZN(n16226) );
  NOR2_X1 U19302 ( .A1(n16227), .A2(n16226), .ZN(n16228) );
  XNOR2_X1 U19303 ( .A(n16229), .B(n16228), .ZN(n16280) );
  INV_X1 U19304 ( .A(n19144), .ZN(n16230) );
  AOI22_X1 U19305 ( .A1(n16280), .A2(n16240), .B1(n16239), .B2(n16230), .ZN(
        n16231) );
  OAI21_X1 U19306 ( .B1(n16278), .B2(n16251), .A(n16231), .ZN(n16232) );
  INV_X1 U19307 ( .A(n16232), .ZN(n16233) );
  OAI211_X1 U19308 ( .C1(n19231), .C2(n16235), .A(n16234), .B(n16233), .ZN(
        P2_U3006) );
  INV_X1 U19309 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16237) );
  OAI22_X1 U19310 ( .A1(n19231), .A2(n16237), .B1(n16236), .B2(n19055), .ZN(
        n16238) );
  AOI21_X1 U19311 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n15785), .A(n16238), .ZN(
        n16243) );
  AOI22_X1 U19312 ( .A1(n16241), .A2(n16240), .B1(n16239), .B2(n19059), .ZN(
        n16242) );
  OAI211_X1 U19313 ( .C1(n16251), .C2(n16244), .A(n16243), .B(n16242), .ZN(
        P2_U3007) );
  OAI22_X1 U19314 ( .A1(n19231), .A2(n19068), .B1(n19877), .B2(n19066), .ZN(
        n16248) );
  OAI22_X1 U19315 ( .A1(n16246), .A2(n19224), .B1(n19223), .B2(n16245), .ZN(
        n16247) );
  AOI211_X1 U19316 ( .C1(n19216), .C2(n19074), .A(n16248), .B(n16247), .ZN(
        n16249) );
  OAI21_X1 U19317 ( .B1(n16251), .B2(n16250), .A(n16249), .ZN(P2_U3008) );
  INV_X1 U19318 ( .A(n16252), .ZN(n16253) );
  AOI22_X1 U19319 ( .A1(n16254), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19262), .B2(n16253), .ZN(n16263) );
  AOI222_X1 U19320 ( .A1(n16257), .A2(n19255), .B1(n19248), .B2(n16256), .C1(
        n16255), .C2(n19250), .ZN(n16262) );
  NAND2_X1 U19321 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n15785), .ZN(n16261) );
  OR3_X1 U19322 ( .A1(n16259), .A2(n16258), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16260) );
  NAND4_X1 U19323 ( .A1(n16263), .A2(n16262), .A3(n16261), .A4(n16260), .ZN(
        P2_U3032) );
  INV_X1 U19324 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19886) );
  NOR2_X1 U19325 ( .A1(n19886), .A2(n19066), .ZN(n16268) );
  XNOR2_X1 U19326 ( .A(n16265), .B(n16264), .ZN(n19162) );
  OAI22_X1 U19327 ( .A1(n19162), .A2(n16290), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16266), .ZN(n16267) );
  AOI211_X1 U19328 ( .C1(n16269), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16268), .B(n16267), .ZN(n16272) );
  INV_X1 U19329 ( .A(n19038), .ZN(n19134) );
  AOI22_X1 U19330 ( .A1(n16270), .A2(n19250), .B1(n19248), .B2(n19134), .ZN(
        n16271) );
  OAI211_X1 U19331 ( .C1(n16274), .C2(n16273), .A(n16272), .B(n16271), .ZN(
        P2_U3036) );
  AOI22_X1 U19332 ( .A1(n16276), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19262), .B2(n16275), .ZN(n16286) );
  OAI22_X1 U19333 ( .A1(n16278), .A2(n16292), .B1(n16277), .B2(n19144), .ZN(
        n16279) );
  AOI21_X1 U19334 ( .B1(n19255), .B2(n16280), .A(n16279), .ZN(n16285) );
  NAND2_X1 U19335 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n15785), .ZN(n16284) );
  OAI211_X1 U19336 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16282), .B(n16281), .ZN(n16283) );
  NAND4_X1 U19337 ( .A1(n16286), .A2(n16285), .A3(n16284), .A4(n16283), .ZN(
        P2_U3038) );
  AOI21_X1 U19338 ( .B1(n16288), .B2(n19248), .A(n16287), .ZN(n16289) );
  OAI21_X1 U19339 ( .B1(n16291), .B2(n16290), .A(n16289), .ZN(n16296) );
  NOR3_X1 U19340 ( .A1(n16294), .A2(n16293), .A3(n16292), .ZN(n16295) );
  AOI211_X1 U19341 ( .C1(n16297), .C2(n19255), .A(n16296), .B(n16295), .ZN(
        n16298) );
  OAI221_X1 U19342 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16301), .C1(
        n16300), .C2(n16299), .A(n16298), .ZN(P2_U3043) );
  INV_X1 U19343 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19941) );
  NAND2_X1 U19344 ( .A1(n16302), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16303) );
  OAI21_X1 U19345 ( .B1(n16304), .B2(n19959), .A(n16303), .ZN(n16306) );
  NAND2_X1 U19346 ( .A1(n16304), .A2(n19959), .ZN(n16305) );
  NAND2_X1 U19347 ( .A1(n16306), .A2(n16305), .ZN(n16307) );
  OAI211_X1 U19348 ( .C1(n16314), .C2(n19941), .A(n16337), .B(n16307), .ZN(
        n16316) );
  NAND2_X1 U19349 ( .A1(n16316), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16311) );
  NOR2_X1 U19350 ( .A1(n16337), .A2(n16308), .ZN(n16309) );
  AOI21_X1 U19351 ( .B1(n16310), .B2(n16337), .A(n16309), .ZN(n16339) );
  NAND2_X1 U19352 ( .A1(n16311), .A2(n16339), .ZN(n16315) );
  INV_X1 U19353 ( .A(n16337), .ZN(n16313) );
  NAND2_X1 U19354 ( .A1(n16313), .A2(n11376), .ZN(n16312) );
  OAI21_X1 U19355 ( .B1(n16314), .B2(n16313), .A(n16312), .ZN(n16319) );
  AOI21_X1 U19356 ( .B1(n16315), .B2(n16319), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16318) );
  NOR2_X1 U19357 ( .A1(n16316), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16317) );
  OAI21_X1 U19358 ( .B1(n16318), .B2(n16317), .A(n15862), .ZN(n16342) );
  INV_X1 U19359 ( .A(n16319), .ZN(n16340) );
  INV_X1 U19360 ( .A(n16320), .ZN(n16326) );
  NAND2_X1 U19361 ( .A1(n16327), .A2(n16321), .ZN(n16325) );
  NAND2_X1 U19362 ( .A1(n16323), .A2(n16322), .ZN(n16324) );
  OAI211_X1 U19363 ( .C1(n16327), .C2(n16326), .A(n16325), .B(n16324), .ZN(
        n19972) );
  NOR2_X1 U19364 ( .A1(P2_MORE_REG_SCAN_IN), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(
        n16333) );
  NOR2_X1 U19365 ( .A1(n16328), .A2(n11415), .ZN(n16329) );
  AOI21_X1 U19366 ( .B1(n16331), .B2(n16330), .A(n16329), .ZN(n16332) );
  OAI21_X1 U19367 ( .B1(n16334), .B2(n16333), .A(n16332), .ZN(n16335) );
  NOR2_X1 U19368 ( .A1(n19972), .A2(n16335), .ZN(n16336) );
  OAI21_X1 U19369 ( .B1(n16337), .B2(n12751), .A(n16336), .ZN(n16338) );
  AOI21_X1 U19370 ( .B1(n16340), .B2(n16339), .A(n16338), .ZN(n16341) );
  NAND2_X1 U19371 ( .A1(n16342), .A2(n16341), .ZN(n16351) );
  AOI211_X1 U19372 ( .C1(n16345), .C2(n16351), .A(n16344), .B(n16343), .ZN(
        n16356) );
  OR2_X1 U19373 ( .A1(n19981), .A2(n19980), .ZN(n16346) );
  AOI21_X1 U19374 ( .B1(n16348), .B2(n16347), .A(n16346), .ZN(n16352) );
  AOI22_X1 U19375 ( .A1(n16350), .A2(n16349), .B1(n19985), .B2(n16352), .ZN(
        n16354) );
  OAI21_X1 U19376 ( .B1(n16351), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16353) );
  AND2_X1 U19377 ( .A1(n16353), .A2(n16352), .ZN(n19850) );
  INV_X1 U19378 ( .A(n19850), .ZN(n19848) );
  NAND2_X1 U19379 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19848), .ZN(n16359) );
  OAI21_X1 U19380 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16354), .A(n16359), 
        .ZN(n16355) );
  OAI211_X1 U19381 ( .C1(n19970), .C2(n16357), .A(n16356), .B(n16355), .ZN(
        P2_U3176) );
  AOI21_X1 U19382 ( .B1(n16359), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16358), 
        .ZN(n16360) );
  INV_X1 U19383 ( .A(n16360), .ZN(P2_U3593) );
  OAI22_X1 U19384 ( .A1(n16386), .A2(n17744), .B1(n16377), .B2(n17904), .ZN(
        n16367) );
  OAI21_X1 U19385 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n9772), .A(
        n16361), .ZN(n16567) );
  NOR2_X1 U19386 ( .A1(n17738), .A2(n16567), .ZN(n16366) );
  OAI221_X1 U19387 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16364), .C1(
        n10065), .C2(n16363), .A(n16362), .ZN(n16365) );
  AOI211_X1 U19388 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n16367), .A(
        n16366), .B(n16365), .ZN(n16374) );
  NAND2_X1 U19389 ( .A1(n16369), .A2(n16368), .ZN(n17967) );
  NOR2_X1 U19390 ( .A1(n16370), .A2(n17619), .ZN(n17560) );
  NAND3_X1 U19391 ( .A1(n16372), .A2(n16371), .A3(n17560), .ZN(n16373) );
  OAI211_X1 U19392 ( .C1(n16375), .C2(n17789), .A(n16374), .B(n16373), .ZN(
        P3_U2800) );
  OAI21_X1 U19393 ( .B1(n18519), .B2(n16376), .A(n16378), .ZN(n16384) );
  AOI211_X1 U19394 ( .C1(n16394), .C2(n16412), .A(n16377), .B(n17904), .ZN(
        n16383) );
  AOI21_X1 U19395 ( .B1(n16378), .B2(n16561), .A(n9772), .ZN(n16577) );
  OAI21_X1 U19396 ( .B1(n16379), .B2(n17756), .A(n16577), .ZN(n16381) );
  NAND2_X1 U19397 ( .A1(n16381), .A2(n16380), .ZN(n16382) );
  AOI211_X1 U19398 ( .C1(n16385), .C2(n16384), .A(n16383), .B(n16382), .ZN(
        n16389) );
  NOR2_X1 U19399 ( .A1(n16386), .A2(n17744), .ZN(n16387) );
  OAI21_X1 U19400 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16410), .A(
        n16387), .ZN(n16388) );
  OAI211_X1 U19401 ( .C1(n16390), .C2(n17789), .A(n16389), .B(n16388), .ZN(
        P3_U2801) );
  OAI211_X1 U19402 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18203), .A(
        n16391), .B(n18205), .ZN(n16397) );
  NOR3_X1 U19403 ( .A1(n16394), .A2(n16393), .A3(n16392), .ZN(n16395) );
  AOI211_X1 U19404 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16397), .A(
        n16396), .B(n16395), .ZN(n16401) );
  AOI22_X1 U19405 ( .A1(n16399), .A2(n18134), .B1(n16398), .B2(n18133), .ZN(
        n16400) );
  OAI211_X1 U19406 ( .C1(n16402), .C2(n18223), .A(n16401), .B(n16400), .ZN(
        P3_U2831) );
  NAND4_X1 U19407 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17813), .A3(
        n16403), .A4(n16416), .ZN(n16420) );
  INV_X1 U19408 ( .A(n18023), .ZN(n17962) );
  AOI21_X1 U19409 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18687), .A(
        n18664), .ZN(n18185) );
  AOI22_X1 U19410 ( .A1(n18706), .A2(n16404), .B1(n18093), .B2(n17940), .ZN(
        n18010) );
  OAI21_X1 U19411 ( .B1(n17962), .B2(n18185), .A(n18010), .ZN(n16405) );
  AOI22_X1 U19412 ( .A1(n18707), .A2(n17964), .B1(n16406), .B2(n16405), .ZN(
        n17961) );
  NOR2_X1 U19413 ( .A1(n17961), .A2(n18126), .ZN(n17977) );
  NOR3_X1 U19414 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16408), .A3(
        n16407), .ZN(n17544) );
  OAI211_X1 U19415 ( .C1(n16410), .C2(n18092), .A(n18215), .B(n16409), .ZN(
        n16411) );
  AOI21_X1 U19416 ( .B1(n18706), .B2(n16412), .A(n16411), .ZN(n16417) );
  AOI22_X1 U19417 ( .A1(n17813), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n16416), .B2(n10010), .ZN(n17547) );
  NAND2_X1 U19418 ( .A1(n17548), .A2(n17547), .ZN(n17546) );
  INV_X1 U19419 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18816) );
  NOR2_X1 U19420 ( .A1(n18108), .A2(n18816), .ZN(n17543) );
  OR3_X1 U19421 ( .A1(n16418), .A2(n18111), .A3(n17547), .ZN(n16419) );
  NOR3_X1 U19422 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16422) );
  NOR4_X1 U19423 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16421) );
  INV_X2 U19424 ( .A(n16509), .ZN(U215) );
  NAND4_X1 U19425 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16422), .A3(n16421), .A4(
        U215), .ZN(U213) );
  INV_X1 U19426 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16511) );
  INV_X2 U19427 ( .A(U214), .ZN(n16472) );
  INV_X1 U19428 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16512) );
  OAI222_X1 U19429 ( .A1(U212), .A2(n16511), .B1(n16474), .B2(n20223), .C1(
        U214), .C2(n16512), .ZN(U216) );
  AOI22_X1 U19430 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16460), .ZN(n16424) );
  OAI21_X1 U19431 ( .B1(n16425), .B2(n16474), .A(n16424), .ZN(U217) );
  INV_X1 U19432 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20212) );
  AOI22_X1 U19433 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16460), .ZN(n16426) );
  OAI21_X1 U19434 ( .B1(n20212), .B2(n16474), .A(n16426), .ZN(U218) );
  AOI22_X1 U19435 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16460), .ZN(n16427) );
  OAI21_X1 U19436 ( .B1(n16428), .B2(n16474), .A(n16427), .ZN(U219) );
  INV_X1 U19437 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20204) );
  AOI22_X1 U19438 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16460), .ZN(n16429) );
  OAI21_X1 U19439 ( .B1(n20204), .B2(n16474), .A(n16429), .ZN(U220) );
  AOI22_X1 U19440 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16460), .ZN(n16430) );
  OAI21_X1 U19441 ( .B1(n20198), .B2(n16474), .A(n16430), .ZN(U221) );
  AOI22_X1 U19442 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16460), .ZN(n16431) );
  OAI21_X1 U19443 ( .B1(n20190), .B2(n16474), .A(n16431), .ZN(U222) );
  AOI22_X1 U19444 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16460), .ZN(n16432) );
  OAI21_X1 U19445 ( .B1(n20183), .B2(n16474), .A(n16432), .ZN(U223) );
  AOI22_X1 U19446 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16460), .ZN(n16433) );
  OAI21_X1 U19447 ( .B1(n20219), .B2(n16474), .A(n16433), .ZN(U224) );
  AOI22_X1 U19448 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16460), .ZN(n16434) );
  OAI21_X1 U19449 ( .B1(n16435), .B2(n16474), .A(n16434), .ZN(U225) );
  INV_X1 U19450 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20215) );
  AOI22_X1 U19451 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16460), .ZN(n16436) );
  OAI21_X1 U19452 ( .B1(n20215), .B2(n16474), .A(n16436), .ZN(U226) );
  AOI22_X1 U19453 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16460), .ZN(n16437) );
  OAI21_X1 U19454 ( .B1(n16438), .B2(n16474), .A(n16437), .ZN(U227) );
  INV_X1 U19455 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20208) );
  AOI22_X1 U19456 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16460), .ZN(n16439) );
  OAI21_X1 U19457 ( .B1(n20208), .B2(n16474), .A(n16439), .ZN(U228) );
  INV_X1 U19458 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20200) );
  AOI22_X1 U19459 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16460), .ZN(n16440) );
  OAI21_X1 U19460 ( .B1(n20200), .B2(n16474), .A(n16440), .ZN(U229) );
  INV_X1 U19461 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20195) );
  AOI22_X1 U19462 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16460), .ZN(n16441) );
  OAI21_X1 U19463 ( .B1(n20195), .B2(n16474), .A(n16441), .ZN(U230) );
  INV_X1 U19464 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20186) );
  AOI22_X1 U19465 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16460), .ZN(n16442) );
  OAI21_X1 U19466 ( .B1(n20186), .B2(n16474), .A(n16442), .ZN(U231) );
  INV_X1 U19467 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16444) );
  AOI22_X1 U19468 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16460), .ZN(n16443) );
  OAI21_X1 U19469 ( .B1(n16444), .B2(n16474), .A(n16443), .ZN(U232) );
  AOI22_X1 U19470 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16460), .ZN(n16445) );
  OAI21_X1 U19471 ( .B1(n16446), .B2(n16474), .A(n16445), .ZN(U233) );
  AOI22_X1 U19472 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16460), .ZN(n16447) );
  OAI21_X1 U19473 ( .B1(n16448), .B2(n16474), .A(n16447), .ZN(U234) );
  AOI22_X1 U19474 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16460), .ZN(n16449) );
  OAI21_X1 U19475 ( .B1(n16450), .B2(n16474), .A(n16449), .ZN(U235) );
  AOI22_X1 U19476 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16460), .ZN(n16451) );
  OAI21_X1 U19477 ( .B1(n13220), .B2(n16474), .A(n16451), .ZN(U236) );
  AOI22_X1 U19478 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16460), .ZN(n16452) );
  OAI21_X1 U19479 ( .B1(n16453), .B2(n16474), .A(n16452), .ZN(U237) );
  AOI22_X1 U19480 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16460), .ZN(n16454) );
  OAI21_X1 U19481 ( .B1(n16455), .B2(n16474), .A(n16454), .ZN(U238) );
  AOI22_X1 U19482 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16460), .ZN(n16456) );
  OAI21_X1 U19483 ( .B1(n16457), .B2(n16474), .A(n16456), .ZN(U239) );
  INV_X1 U19484 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16459) );
  AOI22_X1 U19485 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16460), .ZN(n16458) );
  OAI21_X1 U19486 ( .B1(n16459), .B2(n16474), .A(n16458), .ZN(U240) );
  AOI22_X1 U19487 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16460), .ZN(n16461) );
  OAI21_X1 U19488 ( .B1(n16462), .B2(n16474), .A(n16461), .ZN(U241) );
  AOI22_X1 U19489 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16460), .ZN(n16463) );
  OAI21_X1 U19490 ( .B1(n13207), .B2(n16474), .A(n16463), .ZN(U242) );
  AOI22_X1 U19491 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16460), .ZN(n16464) );
  OAI21_X1 U19492 ( .B1(n16465), .B2(n16474), .A(n16464), .ZN(U243) );
  INV_X1 U19493 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16467) );
  AOI22_X1 U19494 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16460), .ZN(n16466) );
  OAI21_X1 U19495 ( .B1(n16467), .B2(n16474), .A(n16466), .ZN(U244) );
  INV_X1 U19496 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U19497 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16460), .ZN(n16468) );
  OAI21_X1 U19498 ( .B1(n16469), .B2(n16474), .A(n16468), .ZN(U245) );
  INV_X1 U19499 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16471) );
  AOI22_X1 U19500 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16460), .ZN(n16470) );
  OAI21_X1 U19501 ( .B1(n16471), .B2(n16474), .A(n16470), .ZN(U246) );
  INV_X1 U19502 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19503 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16472), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16460), .ZN(n16473) );
  OAI21_X1 U19504 ( .B1(n16475), .B2(n16474), .A(n16473), .ZN(U247) );
  OAI22_X1 U19505 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16509), .ZN(n16476) );
  INV_X1 U19506 ( .A(n16476), .ZN(U251) );
  OAI22_X1 U19507 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16509), .ZN(n16477) );
  INV_X1 U19508 ( .A(n16477), .ZN(U252) );
  OAI22_X1 U19509 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16509), .ZN(n16478) );
  INV_X1 U19510 ( .A(n16478), .ZN(U253) );
  OAI22_X1 U19511 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16509), .ZN(n16479) );
  INV_X1 U19512 ( .A(n16479), .ZN(U254) );
  OAI22_X1 U19513 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16509), .ZN(n16480) );
  INV_X1 U19514 ( .A(n16480), .ZN(U255) );
  OAI22_X1 U19515 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16509), .ZN(n16481) );
  INV_X1 U19516 ( .A(n16481), .ZN(U256) );
  OAI22_X1 U19517 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16509), .ZN(n16482) );
  INV_X1 U19518 ( .A(n16482), .ZN(U257) );
  OAI22_X1 U19519 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16509), .ZN(n16483) );
  INV_X1 U19520 ( .A(n16483), .ZN(U258) );
  OAI22_X1 U19521 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16509), .ZN(n16484) );
  INV_X1 U19522 ( .A(n16484), .ZN(U259) );
  OAI22_X1 U19523 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16503), .ZN(n16485) );
  INV_X1 U19524 ( .A(n16485), .ZN(U260) );
  OAI22_X1 U19525 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16503), .ZN(n16486) );
  INV_X1 U19526 ( .A(n16486), .ZN(U261) );
  OAI22_X1 U19527 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16509), .ZN(n16487) );
  INV_X1 U19528 ( .A(n16487), .ZN(U262) );
  OAI22_X1 U19529 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16509), .ZN(n16488) );
  INV_X1 U19530 ( .A(n16488), .ZN(U263) );
  OAI22_X1 U19531 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16509), .ZN(n16489) );
  INV_X1 U19532 ( .A(n16489), .ZN(U264) );
  OAI22_X1 U19533 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16509), .ZN(n16490) );
  INV_X1 U19534 ( .A(n16490), .ZN(U265) );
  OAI22_X1 U19535 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16503), .ZN(n16491) );
  INV_X1 U19536 ( .A(n16491), .ZN(U266) );
  OAI22_X1 U19537 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16503), .ZN(n16492) );
  INV_X1 U19538 ( .A(n16492), .ZN(U267) );
  OAI22_X1 U19539 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16503), .ZN(n16493) );
  INV_X1 U19540 ( .A(n16493), .ZN(U268) );
  OAI22_X1 U19541 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16503), .ZN(n16494) );
  INV_X1 U19542 ( .A(n16494), .ZN(U269) );
  OAI22_X1 U19543 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16503), .ZN(n16495) );
  INV_X1 U19544 ( .A(n16495), .ZN(U270) );
  OAI22_X1 U19545 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16503), .ZN(n16496) );
  INV_X1 U19546 ( .A(n16496), .ZN(U271) );
  OAI22_X1 U19547 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16509), .ZN(n16497) );
  INV_X1 U19548 ( .A(n16497), .ZN(U272) );
  OAI22_X1 U19549 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16509), .ZN(n16498) );
  INV_X1 U19550 ( .A(n16498), .ZN(U273) );
  OAI22_X1 U19551 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16503), .ZN(n16499) );
  INV_X1 U19552 ( .A(n16499), .ZN(U274) );
  OAI22_X1 U19553 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16509), .ZN(n16500) );
  INV_X1 U19554 ( .A(n16500), .ZN(U275) );
  OAI22_X1 U19555 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16509), .ZN(n16501) );
  INV_X1 U19556 ( .A(n16501), .ZN(U276) );
  OAI22_X1 U19557 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16509), .ZN(n16502) );
  INV_X1 U19558 ( .A(n16502), .ZN(U277) );
  OAI22_X1 U19559 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16503), .ZN(n16504) );
  INV_X1 U19560 ( .A(n16504), .ZN(U278) );
  OAI22_X1 U19561 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16509), .ZN(n16505) );
  INV_X1 U19562 ( .A(n16505), .ZN(U279) );
  OAI22_X1 U19563 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16509), .ZN(n16506) );
  INV_X1 U19564 ( .A(n16506), .ZN(U280) );
  OAI22_X1 U19565 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16509), .ZN(n16508) );
  INV_X1 U19566 ( .A(n16508), .ZN(U281) );
  INV_X1 U19567 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U19568 ( .A1(n16509), .A2(n16511), .B1(n17277), .B2(U215), .ZN(U282) );
  INV_X1 U19569 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16510) );
  AOI222_X1 U19570 ( .A1(n16512), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16511), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16510), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16513) );
  INV_X2 U19571 ( .A(n16515), .ZN(n16514) );
  INV_X1 U19572 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18779) );
  INV_X1 U19573 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U19574 ( .A1(n16514), .A2(n18779), .B1(n19887), .B2(n16515), .ZN(
        U347) );
  INV_X1 U19575 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18777) );
  INV_X1 U19576 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U19577 ( .A1(n16514), .A2(n18777), .B1(n19885), .B2(n16515), .ZN(
        U348) );
  INV_X1 U19578 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18774) );
  INV_X1 U19579 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U19580 ( .A1(n16514), .A2(n18774), .B1(n19883), .B2(n16515), .ZN(
        U349) );
  INV_X1 U19581 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18773) );
  INV_X1 U19582 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U19583 ( .A1(n16514), .A2(n18773), .B1(n19881), .B2(n16515), .ZN(
        U350) );
  INV_X1 U19584 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18771) );
  INV_X1 U19585 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19878) );
  AOI22_X1 U19586 ( .A1(n16514), .A2(n18771), .B1(n19878), .B2(n16515), .ZN(
        U351) );
  INV_X1 U19587 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18768) );
  INV_X1 U19588 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19876) );
  AOI22_X1 U19589 ( .A1(n16514), .A2(n18768), .B1(n19876), .B2(n16515), .ZN(
        U352) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18767) );
  INV_X1 U19591 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19875) );
  AOI22_X1 U19592 ( .A1(n16514), .A2(n18767), .B1(n19875), .B2(n16515), .ZN(
        U353) );
  INV_X1 U19593 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18765) );
  AOI22_X1 U19594 ( .A1(n16514), .A2(n18765), .B1(n19874), .B2(n16515), .ZN(
        U354) );
  INV_X1 U19595 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18818) );
  INV_X1 U19596 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19916) );
  AOI22_X1 U19597 ( .A1(n16514), .A2(n18818), .B1(n19916), .B2(n16515), .ZN(
        U356) );
  INV_X1 U19598 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18815) );
  INV_X1 U19599 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19914) );
  AOI22_X1 U19600 ( .A1(n16514), .A2(n18815), .B1(n19914), .B2(n16515), .ZN(
        U357) );
  INV_X1 U19601 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18814) );
  INV_X1 U19602 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19912) );
  AOI22_X1 U19603 ( .A1(n16514), .A2(n18814), .B1(n19912), .B2(n16515), .ZN(
        U358) );
  INV_X1 U19604 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18812) );
  INV_X1 U19605 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19911) );
  AOI22_X1 U19606 ( .A1(n16514), .A2(n18812), .B1(n19911), .B2(n16515), .ZN(
        U359) );
  INV_X1 U19607 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18809) );
  INV_X1 U19608 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19909) );
  AOI22_X1 U19609 ( .A1(n16514), .A2(n18809), .B1(n19909), .B2(n16515), .ZN(
        U360) );
  INV_X1 U19610 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18806) );
  INV_X1 U19611 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U19612 ( .A1(n16514), .A2(n18806), .B1(n19907), .B2(n16515), .ZN(
        U361) );
  INV_X1 U19613 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18804) );
  INV_X1 U19614 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U19615 ( .A1(n16514), .A2(n18804), .B1(n19905), .B2(n16515), .ZN(
        U362) );
  INV_X1 U19616 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18803) );
  INV_X1 U19617 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19903) );
  AOI22_X1 U19618 ( .A1(n16514), .A2(n18803), .B1(n19903), .B2(n16515), .ZN(
        U363) );
  INV_X1 U19619 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18801) );
  INV_X1 U19620 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19902) );
  AOI22_X1 U19621 ( .A1(n16514), .A2(n18801), .B1(n19902), .B2(n16515), .ZN(
        U364) );
  INV_X1 U19622 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18763) );
  INV_X1 U19623 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19873) );
  AOI22_X1 U19624 ( .A1(n16514), .A2(n18763), .B1(n19873), .B2(n16515), .ZN(
        U365) );
  INV_X1 U19625 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18798) );
  INV_X1 U19626 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U19627 ( .A1(n16514), .A2(n18798), .B1(n19901), .B2(n16515), .ZN(
        U366) );
  INV_X1 U19628 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18797) );
  INV_X1 U19629 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19900) );
  AOI22_X1 U19630 ( .A1(n16514), .A2(n18797), .B1(n19900), .B2(n16515), .ZN(
        U367) );
  INV_X1 U19631 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18795) );
  INV_X1 U19632 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19898) );
  AOI22_X1 U19633 ( .A1(n16514), .A2(n18795), .B1(n19898), .B2(n16515), .ZN(
        U368) );
  INV_X1 U19634 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18793) );
  INV_X1 U19635 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U19636 ( .A1(n16514), .A2(n18793), .B1(n19897), .B2(n16515), .ZN(
        U369) );
  INV_X1 U19637 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18791) );
  INV_X1 U19638 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19895) );
  AOI22_X1 U19639 ( .A1(n16514), .A2(n18791), .B1(n19895), .B2(n16515), .ZN(
        U370) );
  INV_X1 U19640 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18789) );
  INV_X1 U19641 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19893) );
  AOI22_X1 U19642 ( .A1(n16514), .A2(n18789), .B1(n19893), .B2(n16515), .ZN(
        U371) );
  INV_X1 U19643 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18786) );
  INV_X1 U19644 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U19645 ( .A1(n16514), .A2(n18786), .B1(n19891), .B2(n16515), .ZN(
        U372) );
  INV_X1 U19646 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18785) );
  INV_X1 U19647 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U19648 ( .A1(n16514), .A2(n18785), .B1(n19890), .B2(n16515), .ZN(
        U373) );
  INV_X1 U19649 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18783) );
  INV_X1 U19650 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19889) );
  AOI22_X1 U19651 ( .A1(n16514), .A2(n18783), .B1(n19889), .B2(n16515), .ZN(
        U374) );
  INV_X1 U19652 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18781) );
  INV_X1 U19653 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19888) );
  AOI22_X1 U19654 ( .A1(n16514), .A2(n18781), .B1(n19888), .B2(n16515), .ZN(
        U375) );
  INV_X1 U19655 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18761) );
  INV_X1 U19656 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19871) );
  AOI22_X1 U19657 ( .A1(n16514), .A2(n18761), .B1(n19871), .B2(n16515), .ZN(
        U376) );
  INV_X1 U19658 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18760) );
  NAND2_X1 U19659 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18760), .ZN(n18748) );
  AOI22_X1 U19660 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18748), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18758), .ZN(n18830) );
  AOI21_X1 U19661 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18830), .ZN(n16516) );
  INV_X1 U19662 ( .A(n16516), .ZN(P3_U2633) );
  INV_X1 U19663 ( .A(n16522), .ZN(n16518) );
  OAI21_X1 U19664 ( .B1(n16518), .B2(n17466), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16519) );
  OAI21_X1 U19665 ( .B1(n18896), .B2(n18735), .A(n16519), .ZN(P3_U2634) );
  AOI21_X1 U19666 ( .B1(n18758), .B2(n18760), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16520) );
  AOI22_X1 U19667 ( .A1(n18893), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16520), 
        .B2(n18894), .ZN(P3_U2635) );
  NOR2_X1 U19668 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18744) );
  OAI21_X1 U19669 ( .B1(n18744), .B2(BS16), .A(n18830), .ZN(n18828) );
  OAI21_X1 U19670 ( .B1(n18830), .B2(n18883), .A(n18828), .ZN(P3_U2636) );
  AND3_X1 U19671 ( .A1(n18711), .A2(n16522), .A3(n16521), .ZN(n18715) );
  NOR2_X1 U19672 ( .A1(n18715), .A2(n18732), .ZN(n18877) );
  OAI21_X1 U19673 ( .B1(n18877), .B2(n18226), .A(n16523), .ZN(P3_U2637) );
  NOR4_X1 U19674 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16527) );
  NOR4_X1 U19675 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16526) );
  NOR4_X1 U19676 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16525) );
  NOR4_X1 U19677 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16524) );
  NAND4_X1 U19678 ( .A1(n16527), .A2(n16526), .A3(n16525), .A4(n16524), .ZN(
        n16533) );
  NOR4_X1 U19679 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16531) );
  AOI211_X1 U19680 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16530) );
  NOR4_X1 U19681 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16529) );
  NOR4_X1 U19682 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16528) );
  NAND4_X1 U19683 ( .A1(n16531), .A2(n16530), .A3(n16529), .A4(n16528), .ZN(
        n16532) );
  NOR2_X1 U19684 ( .A1(n16533), .A2(n16532), .ZN(n18875) );
  INV_X1 U19685 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16535) );
  NOR3_X1 U19686 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16536) );
  OAI21_X1 U19687 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16536), .A(n18875), .ZN(
        n16534) );
  OAI21_X1 U19688 ( .B1(n18875), .B2(n16535), .A(n16534), .ZN(P3_U2638) );
  INV_X1 U19689 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18868) );
  INV_X1 U19690 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18829) );
  AOI21_X1 U19691 ( .B1(n18868), .B2(n18829), .A(n16536), .ZN(n16538) );
  INV_X1 U19692 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16537) );
  INV_X1 U19693 ( .A(n18875), .ZN(n18870) );
  AOI22_X1 U19694 ( .A1(n18875), .A2(n16538), .B1(n16537), .B2(n18870), .ZN(
        P3_U2639) );
  NAND2_X1 U19695 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16544), .ZN(n16540) );
  AOI211_X4 U19696 ( .C1(n18883), .C2(n18885), .A(n16542), .B(n16540), .ZN(
        n16904) );
  NOR3_X1 U19697 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16877) );
  INV_X1 U19698 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17246) );
  NAND2_X1 U19699 ( .A1(n16877), .A2(n17246), .ZN(n16870) );
  NOR2_X1 U19700 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16870), .ZN(n16851) );
  NAND2_X1 U19701 ( .A1(n16851), .A2(n17240), .ZN(n16844) );
  NAND2_X1 U19702 ( .A1(n16825), .A2(n16821), .ZN(n16820) );
  INV_X1 U19703 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17161) );
  NAND2_X1 U19704 ( .A1(n16803), .A2(n17161), .ZN(n16796) );
  INV_X1 U19705 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16774) );
  NAND2_X1 U19706 ( .A1(n16778), .A2(n16774), .ZN(n16773) );
  INV_X1 U19707 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16749) );
  NAND2_X1 U19708 ( .A1(n16756), .A2(n16749), .ZN(n16746) );
  INV_X1 U19709 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16723) );
  NAND2_X1 U19710 ( .A1(n16733), .A2(n16723), .ZN(n16721) );
  NAND2_X1 U19711 ( .A1(n16710), .A2(n17076), .ZN(n16701) );
  NOR2_X1 U19712 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16701), .ZN(n16691) );
  INV_X1 U19713 ( .A(n16691), .ZN(n16673) );
  NAND2_X1 U19714 ( .A1(n16665), .A2(n17011), .ZN(n16660) );
  NOR2_X1 U19715 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16660), .ZN(n16646) );
  NAND2_X1 U19716 ( .A1(n16646), .A2(n16641), .ZN(n16640) );
  NOR2_X1 U19717 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16640), .ZN(n16614) );
  NAND2_X1 U19718 ( .A1(n16614), .A2(n16623), .ZN(n16607) );
  NOR2_X1 U19719 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16607), .ZN(n16606) );
  NAND2_X1 U19720 ( .A1(n16606), .A2(n16912), .ZN(n16599) );
  NOR2_X1 U19721 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16599), .ZN(n16586) );
  INV_X1 U19722 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16955) );
  NAND2_X1 U19723 ( .A1(n16586), .A2(n16955), .ZN(n16566) );
  NOR2_X1 U19724 ( .A1(n16896), .A2(n16566), .ZN(n16571) );
  INV_X1 U19725 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16918) );
  INV_X1 U19726 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18821) );
  INV_X1 U19727 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18813) );
  NOR2_X1 U19728 ( .A1(n18816), .A2(n18813), .ZN(n16584) );
  INV_X1 U19729 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18811) );
  INV_X1 U19730 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18808) );
  AOI211_X1 U19731 ( .C1(n18882), .C2(n18884), .A(n18751), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16543) );
  INV_X1 U19732 ( .A(n16543), .ZN(n18725) );
  INV_X1 U19733 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18805) );
  INV_X1 U19734 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18796) );
  INV_X1 U19735 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18787) );
  INV_X1 U19736 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18782) );
  INV_X1 U19737 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18766) );
  NAND3_X1 U19738 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16852) );
  NOR2_X1 U19739 ( .A1(n18766), .A2(n16852), .ZN(n16839) );
  NAND2_X1 U19740 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16839), .ZN(n16812) );
  NAND3_X1 U19741 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n16767) );
  NOR2_X1 U19742 ( .A1(n16812), .A2(n16767), .ZN(n16780) );
  NAND4_X1 U19743 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16780), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16761) );
  NOR2_X1 U19744 ( .A1(n18782), .A2(n16761), .ZN(n16745) );
  NAND2_X1 U19745 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16745), .ZN(n16734) );
  NOR2_X1 U19746 ( .A1(n18787), .A2(n16734), .ZN(n16679) );
  NAND3_X1 U19747 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16678) );
  INV_X1 U19748 ( .A(n16678), .ZN(n16680) );
  NAND3_X1 U19749 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16679), .A3(n16680), 
        .ZN(n16674) );
  NOR2_X1 U19750 ( .A1(n18796), .A2(n16674), .ZN(n16664) );
  NAND2_X1 U19751 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16664), .ZN(n16645) );
  NAND2_X1 U19752 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16644) );
  NOR3_X1 U19753 ( .A1(n18805), .A2(n16645), .A3(n16644), .ZN(n16625) );
  NAND3_X1 U19754 ( .A1(n16864), .A2(n16625), .A3(P3_REIP_REG_24__SCAN_IN), 
        .ZN(n16617) );
  NOR3_X1 U19755 ( .A1(n18811), .A2(n18808), .A3(n16617), .ZN(n16598) );
  NAND3_X1 U19756 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16584), .A3(n16598), 
        .ZN(n16548) );
  NOR3_X1 U19757 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18821), .A3(n16548), 
        .ZN(n16547) );
  NAND4_X1 U19758 ( .A1(n18727), .A2(n18735), .A3(n18883), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n16879) );
  NAND2_X1 U19759 ( .A1(n18727), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18606) );
  NOR3_X1 U19760 ( .A1(n18735), .A2(n18606), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n16541) );
  AOI211_X4 U19761 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16544), .A(n16543), .B(
        n16542), .ZN(n16905) );
  AOI22_X1 U19762 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16889), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16905), .ZN(n16545) );
  INV_X1 U19763 ( .A(n16545), .ZN(n16546) );
  AOI211_X1 U19764 ( .C1(n16571), .C2(n16918), .A(n16547), .B(n16546), .ZN(
        n16565) );
  NOR2_X1 U19765 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16548), .ZN(n16570) );
  NOR2_X1 U19766 ( .A1(n16899), .A2(n16864), .ZN(n16681) );
  INV_X1 U19767 ( .A(n16681), .ZN(n16903) );
  NAND2_X1 U19768 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16584), .ZN(n16550) );
  NOR2_X1 U19769 ( .A1(n18811), .A2(n18808), .ZN(n16549) );
  INV_X1 U19770 ( .A(n16899), .ZN(n16906) );
  OAI21_X1 U19771 ( .B1(n16892), .B2(n16625), .A(n16906), .ZN(n16639) );
  INV_X1 U19772 ( .A(n16639), .ZN(n16615) );
  OAI221_X1 U19773 ( .B1(n16681), .B2(P3_REIP_REG_24__SCAN_IN), .C1(n16681), 
        .C2(n16549), .A(n16615), .ZN(n16611) );
  AOI21_X1 U19774 ( .B1(n16903), .B2(n16550), .A(n16611), .ZN(n16568) );
  INV_X1 U19775 ( .A(n16568), .ZN(n16580) );
  OAI21_X1 U19776 ( .B1(n16570), .B2(n16580), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16564) );
  INV_X1 U19777 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17598) );
  INV_X1 U19778 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17585) );
  NAND2_X1 U19779 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17582), .ZN(
        n16558) );
  NOR3_X1 U19780 ( .A1(n17598), .A2(n17585), .A3(n16558), .ZN(n16560) );
  INV_X1 U19781 ( .A(n16560), .ZN(n17538) );
  NOR2_X1 U19782 ( .A1(n17567), .A2(n17538), .ZN(n16552) );
  INV_X1 U19783 ( .A(n16562), .ZN(n16551) );
  OAI21_X1 U19784 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16552), .A(
        n16551), .ZN(n17555) );
  INV_X1 U19785 ( .A(n17555), .ZN(n16595) );
  INV_X1 U19786 ( .A(n16558), .ZN(n16559) );
  NAND2_X1 U19787 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16559), .ZN(
        n16553) );
  AOI21_X1 U19788 ( .B1(n17585), .B2(n16553), .A(n16560), .ZN(n17588) );
  INV_X1 U19789 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17893) );
  NOR2_X1 U19790 ( .A1(n17893), .A2(n17609), .ZN(n17581) );
  OAI21_X1 U19791 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17581), .A(
        n16558), .ZN(n16554) );
  INV_X1 U19792 ( .A(n16554), .ZN(n17612) );
  INV_X1 U19793 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17637) );
  NAND2_X1 U19794 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17622), .ZN(
        n16555) );
  XOR2_X1 U19795 ( .A(n17637), .B(n16555), .Z(n17646) );
  NAND2_X1 U19796 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17669), .ZN(
        n17659) );
  INV_X1 U19797 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17713) );
  NAND2_X1 U19798 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n12570), .ZN(
        n17736) );
  OR2_X1 U19799 ( .A1(n16556), .A2(n17736), .ZN(n17696) );
  NOR2_X1 U19800 ( .A1(n17713), .A2(n17696), .ZN(n16725) );
  INV_X1 U19801 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16861) );
  INV_X1 U19802 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17671) );
  INV_X1 U19803 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17661) );
  NOR2_X1 U19804 ( .A1(n17671), .A2(n17661), .ZN(n17663) );
  NAND2_X1 U19805 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9758), .ZN(
        n17620) );
  AOI22_X1 U19806 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17622), .B1(
        n17623), .B2(n17620), .ZN(n17653) );
  NOR2_X1 U19807 ( .A1(n16684), .A2(n17653), .ZN(n16666) );
  NOR2_X1 U19808 ( .A1(n16666), .A2(n16860), .ZN(n16656) );
  NOR2_X1 U19809 ( .A1(n17646), .A2(n16656), .ZN(n16655) );
  NOR2_X1 U19810 ( .A1(n16655), .A2(n16860), .ZN(n16649) );
  INV_X1 U19811 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17625) );
  NAND3_X1 U19812 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17622), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16557) );
  AOI21_X1 U19813 ( .B1(n17625), .B2(n16557), .A(n17581), .ZN(n17628) );
  NOR2_X1 U19814 ( .A1(n16634), .A2(n16860), .ZN(n16629) );
  AOI22_X1 U19815 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16559), .B1(
        n16558), .B2(n17598), .ZN(n17604) );
  OAI22_X1 U19816 ( .A1(n17567), .A2(n16560), .B1(n17538), .B2(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17568) );
  OAI21_X1 U19817 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16562), .A(
        n16561), .ZN(n17541) );
  INV_X1 U19818 ( .A(n17541), .ZN(n16588) );
  NAND4_X1 U19819 ( .A1(n10056), .A2(n18736), .A3(n16575), .A4(n16567), .ZN(
        n16563) );
  NAND3_X1 U19820 ( .A1(n16565), .A2(n16564), .A3(n16563), .ZN(P3_U2640) );
  NAND2_X1 U19821 ( .A1(n16904), .A2(n16566), .ZN(n16573) );
  OAI22_X1 U19822 ( .A1(n16568), .A2(n18821), .B1(n10065), .B2(n16874), .ZN(
        n16569) );
  OAI21_X1 U19823 ( .B1(n16905), .B2(n16571), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16572) );
  NAND2_X1 U19824 ( .A1(n16584), .A2(n16598), .ZN(n16583) );
  AOI22_X1 U19825 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16889), .B1(
        n16905), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16582) );
  INV_X1 U19826 ( .A(n16586), .ZN(n16574) );
  AOI21_X1 U19827 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16574), .A(n16573), .ZN(
        n16579) );
  AOI211_X1 U19828 ( .C1(n16577), .C2(n16576), .A(n16575), .B(n16879), .ZN(
        n16578) );
  AOI211_X1 U19829 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16580), .A(n16579), 
        .B(n16578), .ZN(n16581) );
  OAI211_X1 U19830 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16583), .A(n16582), 
        .B(n16581), .ZN(P3_U2642) );
  AOI21_X1 U19831 ( .B1(n18816), .B2(n18813), .A(n16584), .ZN(n16585) );
  AOI22_X1 U19832 ( .A1(n16905), .A2(P3_EBX_REG_28__SCAN_IN), .B1(n16598), 
        .B2(n16585), .ZN(n16592) );
  AOI211_X1 U19833 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16599), .A(n16586), .B(
        n16896), .ZN(n16590) );
  AOI211_X1 U19834 ( .C1(n16588), .C2(n16587), .A(n9739), .B(n16879), .ZN(
        n16589) );
  AOI211_X1 U19835 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16611), .A(n16590), 
        .B(n16589), .ZN(n16591) );
  OAI211_X1 U19836 ( .C1(n10064), .C2(n16874), .A(n16592), .B(n16591), .ZN(
        P3_U2643) );
  INV_X1 U19837 ( .A(n16611), .ZN(n16602) );
  AOI211_X1 U19838 ( .C1(n16595), .C2(n16594), .A(n16593), .B(n16879), .ZN(
        n16597) );
  INV_X1 U19839 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17535) );
  OAI22_X1 U19840 ( .A1(n17535), .A2(n16874), .B1(n16891), .B2(n16912), .ZN(
        n16596) );
  AOI211_X1 U19841 ( .C1(n16598), .C2(n18813), .A(n16597), .B(n16596), .ZN(
        n16601) );
  OAI211_X1 U19842 ( .C1(n16606), .C2(n16912), .A(n16904), .B(n16599), .ZN(
        n16600) );
  OAI211_X1 U19843 ( .C1(n16602), .C2(n18813), .A(n16601), .B(n16600), .ZN(
        P3_U2644) );
  AOI22_X1 U19844 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16889), .B1(
        n16905), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16613) );
  OAI21_X1 U19845 ( .B1(n18808), .B2(n16617), .A(n18811), .ZN(n16610) );
  INV_X1 U19846 ( .A(n16603), .ZN(n16604) );
  AOI211_X1 U19847 ( .C1(n17568), .C2(n16605), .A(n16604), .B(n16879), .ZN(
        n16609) );
  AOI211_X1 U19848 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16607), .A(n16606), .B(
        n16896), .ZN(n16608) );
  AOI211_X1 U19849 ( .C1(n16611), .C2(n16610), .A(n16609), .B(n16608), .ZN(
        n16612) );
  NAND2_X1 U19850 ( .A1(n16613), .A2(n16612), .ZN(P3_U2645) );
  OR2_X1 U19851 ( .A1(n16896), .A2(n16614), .ZN(n16626) );
  AOI21_X1 U19852 ( .B1(n16904), .B2(n16614), .A(n16905), .ZN(n16622) );
  OAI21_X1 U19853 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16892), .A(n16615), 
        .ZN(n16620) );
  AOI211_X1 U19854 ( .C1(n17588), .C2(n16616), .A(n9742), .B(n16879), .ZN(
        n16619) );
  OAI22_X1 U19855 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16617), .B1(n17585), 
        .B2(n16874), .ZN(n16618) );
  AOI211_X1 U19856 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16620), .A(n16619), 
        .B(n16618), .ZN(n16621) );
  OAI221_X1 U19857 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16626), .C1(n16623), 
        .C2(n16622), .A(n16621), .ZN(P3_U2646) );
  NOR2_X1 U19858 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16892), .ZN(n16624) );
  AOI22_X1 U19859 ( .A1(n16905), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16625), 
        .B2(n16624), .ZN(n16633) );
  AOI21_X1 U19860 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16640), .A(n16626), .ZN(
        n16631) );
  INV_X1 U19861 ( .A(n16627), .ZN(n16628) );
  AOI211_X1 U19862 ( .C1(n17604), .C2(n16629), .A(n16628), .B(n16879), .ZN(
        n16630) );
  AOI211_X1 U19863 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16639), .A(n16631), 
        .B(n16630), .ZN(n16632) );
  OAI211_X1 U19864 ( .C1(n17598), .C2(n16874), .A(n16633), .B(n16632), .ZN(
        P3_U2647) );
  OAI21_X1 U19865 ( .B1(n16644), .B2(n16663), .A(n18805), .ZN(n16638) );
  AOI211_X1 U19866 ( .C1(n17612), .C2(n16635), .A(n16634), .B(n16879), .ZN(
        n16637) );
  OAI22_X1 U19867 ( .A1(n17584), .A2(n16874), .B1(n16891), .B2(n16641), .ZN(
        n16636) );
  AOI211_X1 U19868 ( .C1(n16639), .C2(n16638), .A(n16637), .B(n16636), .ZN(
        n16643) );
  OAI211_X1 U19869 ( .C1(n16646), .C2(n16641), .A(n16904), .B(n16640), .ZN(
        n16642) );
  NAND2_X1 U19870 ( .A1(n16643), .A2(n16642), .ZN(P3_U2648) );
  OAI21_X1 U19871 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(P3_REIP_REG_21__SCAN_IN), 
        .A(n16644), .ZN(n16654) );
  AOI22_X1 U19872 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16889), .B1(
        n16905), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16653) );
  AOI21_X1 U19873 ( .B1(n16645), .B2(n16864), .A(n16899), .ZN(n16671) );
  INV_X1 U19874 ( .A(n16671), .ZN(n16659) );
  AOI211_X1 U19875 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16660), .A(n16646), .B(
        n16896), .ZN(n16651) );
  INV_X1 U19876 ( .A(n16647), .ZN(n16648) );
  AOI211_X1 U19877 ( .C1(n17628), .C2(n16649), .A(n16648), .B(n16879), .ZN(
        n16650) );
  AOI211_X1 U19878 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16659), .A(n16651), 
        .B(n16650), .ZN(n16652) );
  OAI211_X1 U19879 ( .C1(n16663), .C2(n16654), .A(n16653), .B(n16652), .ZN(
        P3_U2649) );
  AOI211_X1 U19880 ( .C1(n17646), .C2(n16656), .A(n16655), .B(n16879), .ZN(
        n16658) );
  OAI22_X1 U19881 ( .A1(n17637), .A2(n16874), .B1(n16891), .B2(n17011), .ZN(
        n16657) );
  AOI211_X1 U19882 ( .C1(n16659), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16658), 
        .B(n16657), .ZN(n16662) );
  OAI211_X1 U19883 ( .C1(n16665), .C2(n17011), .A(n16904), .B(n16660), .ZN(
        n16661) );
  OAI211_X1 U19884 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16663), .A(n16662), 
        .B(n16661), .ZN(P3_U2650) );
  AOI21_X1 U19885 ( .B1(n16864), .B2(n16664), .A(P3_REIP_REG_20__SCAN_IN), 
        .ZN(n16672) );
  AOI22_X1 U19886 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16889), .B1(
        n16905), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16670) );
  AOI211_X1 U19887 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16676), .A(n16665), .B(
        n16896), .ZN(n16668) );
  AOI211_X1 U19888 ( .C1(n17653), .C2(n16684), .A(n16666), .B(n16879), .ZN(
        n16667) );
  NOR2_X1 U19889 ( .A1(n16668), .A2(n16667), .ZN(n16669) );
  OAI211_X1 U19890 ( .C1(n16672), .C2(n16671), .A(n16670), .B(n16669), .ZN(
        P3_U2651) );
  AOI22_X1 U19891 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16889), .B1(
        n16905), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16689) );
  AOI21_X1 U19892 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16673), .A(n16896), .ZN(
        n16677) );
  NOR3_X1 U19893 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16892), .A3(n16674), 
        .ZN(n16675) );
  AOI211_X1 U19894 ( .C1(n16677), .C2(n16676), .A(n18210), .B(n16675), .ZN(
        n16688) );
  NAND2_X1 U19895 ( .A1(n16864), .A2(n16679), .ZN(n16726) );
  NOR3_X1 U19896 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16678), .A3(n16726), 
        .ZN(n16694) );
  NAND2_X1 U19897 ( .A1(n16679), .A2(n16906), .ZN(n16735) );
  NAND2_X1 U19898 ( .A1(n16903), .A2(n16735), .ZN(n16738) );
  OAI21_X1 U19899 ( .B1(n16681), .B2(n16680), .A(n16738), .ZN(n16690) );
  OAI21_X1 U19900 ( .B1(n16694), .B2(n16690), .A(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n16687) );
  NOR2_X1 U19901 ( .A1(n17671), .A2(n17659), .ZN(n16695) );
  OAI21_X1 U19902 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16695), .A(
        n17620), .ZN(n17660) );
  INV_X1 U19903 ( .A(n17660), .ZN(n16685) );
  INV_X1 U19904 ( .A(n16715), .ZN(n16727) );
  OAI21_X1 U19905 ( .B1(n16860), .B2(n16695), .A(n16727), .ZN(n16682) );
  INV_X1 U19906 ( .A(n16682), .ZN(n16683) );
  OAI221_X1 U19907 ( .B1(n16685), .B2(n16684), .C1(n17660), .C2(n16683), .A(
        n18736), .ZN(n16686) );
  NAND4_X1 U19908 ( .A1(n16689), .A2(n16688), .A3(n16687), .A4(n16686), .ZN(
        P3_U2652) );
  INV_X1 U19909 ( .A(n16690), .ZN(n16709) );
  INV_X1 U19910 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18794) );
  AOI211_X1 U19911 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16701), .A(n16691), .B(
        n16896), .ZN(n16693) );
  OAI22_X1 U19912 ( .A1(n17671), .A2(n16874), .B1(n16891), .B2(n17059), .ZN(
        n16692) );
  NOR4_X1 U19913 ( .A1(n18210), .A2(n16694), .A3(n16693), .A4(n16692), .ZN(
        n16700) );
  AOI21_X1 U19914 ( .B1(n17671), .B2(n17659), .A(n16695), .ZN(n17674) );
  INV_X1 U19915 ( .A(n17674), .ZN(n16697) );
  INV_X1 U19916 ( .A(n16698), .ZN(n16696) );
  OAI221_X1 U19917 ( .B1(n16698), .B2(n16697), .C1(n16696), .C2(n17674), .A(
        n18736), .ZN(n16699) );
  OAI211_X1 U19918 ( .C1(n16709), .C2(n18794), .A(n16700), .B(n16699), .ZN(
        P3_U2653) );
  INV_X1 U19919 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18792) );
  INV_X1 U19920 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18790) );
  INV_X1 U19921 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18788) );
  NOR4_X1 U19922 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n18790), .A3(n18788), 
        .A4(n16726), .ZN(n16704) );
  OAI211_X1 U19923 ( .C1(n16710), .C2(n17076), .A(n16904), .B(n16701), .ZN(
        n16702) );
  OAI211_X1 U19924 ( .C1(n16891), .C2(n17076), .A(n18108), .B(n16702), .ZN(
        n16703) );
  AOI211_X1 U19925 ( .C1(n16889), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16704), .B(n16703), .ZN(n16708) );
  NOR2_X1 U19926 ( .A1(n17893), .A2(n17681), .ZN(n16712) );
  OAI21_X1 U19927 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16712), .A(
        n17659), .ZN(n17683) );
  NOR2_X1 U19928 ( .A1(n17893), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16875) );
  INV_X1 U19929 ( .A(n16875), .ZN(n16848) );
  OAI21_X1 U19930 ( .B1(n17681), .B2(n16848), .A(n10056), .ZN(n16706) );
  AOI21_X1 U19931 ( .B1(n17683), .B2(n16706), .A(n16879), .ZN(n16705) );
  OAI21_X1 U19932 ( .B1(n17683), .B2(n16706), .A(n16705), .ZN(n16707) );
  OAI211_X1 U19933 ( .C1(n16709), .C2(n18792), .A(n16708), .B(n16707), .ZN(
        P3_U2654) );
  INV_X1 U19934 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17698) );
  AOI211_X1 U19935 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16721), .A(n16710), .B(
        n16896), .ZN(n16711) );
  AOI211_X1 U19936 ( .C1(n16905), .C2(P3_EBX_REG_16__SCAN_IN), .A(n18210), .B(
        n16711), .ZN(n16720) );
  NOR2_X1 U19937 ( .A1(n18788), .A2(n16726), .ZN(n16718) );
  OAI21_X1 U19938 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16726), .A(n16738), 
        .ZN(n16717) );
  INV_X1 U19939 ( .A(n16725), .ZN(n16713) );
  AOI21_X1 U19940 ( .B1(n17698), .B2(n16713), .A(n16712), .ZN(n17701) );
  INV_X1 U19941 ( .A(n17701), .ZN(n16714) );
  AOI221_X1 U19942 ( .B1(n16715), .B2(n17701), .C1(n16727), .C2(n16714), .A(
        n16879), .ZN(n16716) );
  AOI221_X1 U19943 ( .B1(n16718), .B2(n18790), .C1(n16717), .C2(
        P3_REIP_REG_16__SCAN_IN), .A(n16716), .ZN(n16719) );
  OAI211_X1 U19944 ( .C1(n17698), .C2(n16874), .A(n16720), .B(n16719), .ZN(
        P3_U2655) );
  OAI211_X1 U19945 ( .C1(n16733), .C2(n16723), .A(n16904), .B(n16721), .ZN(
        n16722) );
  OAI211_X1 U19946 ( .C1(n16891), .C2(n16723), .A(n18108), .B(n16722), .ZN(
        n16724) );
  AOI21_X1 U19947 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n16889), .A(
        n16724), .ZN(n16732) );
  AOI21_X1 U19948 ( .B1(n17713), .B2(n17696), .A(n16725), .ZN(n17716) );
  NOR2_X1 U19949 ( .A1(n16860), .A2(n16861), .ZN(n16890) );
  OR2_X1 U19950 ( .A1(n16879), .A2(n16890), .ZN(n16902) );
  AOI21_X1 U19951 ( .B1(n10056), .B2(n17696), .A(n16902), .ZN(n16730) );
  NOR2_X1 U19952 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16726), .ZN(n16729) );
  NOR3_X1 U19953 ( .A1(n17716), .A2(n16727), .A3(n16879), .ZN(n16728) );
  AOI211_X1 U19954 ( .C1(n17716), .C2(n16730), .A(n16729), .B(n16728), .ZN(
        n16731) );
  OAI211_X1 U19955 ( .C1(n18788), .C2(n16738), .A(n16732), .B(n16731), .ZN(
        P3_U2656) );
  NOR2_X1 U19956 ( .A1(n17742), .A2(n17736), .ZN(n16743) );
  OAI21_X1 U19957 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16743), .A(
        n17696), .ZN(n17726) );
  AOI21_X1 U19958 ( .B1(n16743), .B2(n16861), .A(n16860), .ZN(n16753) );
  XOR2_X1 U19959 ( .A(n17726), .B(n16753), .Z(n16742) );
  AOI211_X1 U19960 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16746), .A(n16733), .B(
        n16896), .ZN(n16740) );
  NOR2_X1 U19961 ( .A1(n16892), .A2(n16734), .ZN(n16736) );
  AOI22_X1 U19962 ( .A1(n16905), .A2(P3_EBX_REG_14__SCAN_IN), .B1(n16736), 
        .B2(n16735), .ZN(n16737) );
  OAI211_X1 U19963 ( .C1(n18787), .C2(n16738), .A(n16737), .B(n18108), .ZN(
        n16739) );
  AOI211_X1 U19964 ( .C1(n16889), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16740), .B(n16739), .ZN(n16741) );
  OAI21_X1 U19965 ( .B1(n16879), .B2(n16742), .A(n16741), .ZN(P3_U2657) );
  INV_X1 U19966 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17739) );
  INV_X1 U19967 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17759) );
  NOR2_X1 U19968 ( .A1(n17759), .A2(n17736), .ZN(n16758) );
  INV_X1 U19969 ( .A(n16743), .ZN(n16744) );
  OAI21_X1 U19970 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16758), .A(
        n16744), .ZN(n17737) );
  AOI211_X1 U19971 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n10056), .A(
        n17737), .B(n16902), .ZN(n16752) );
  AOI21_X1 U19972 ( .B1(n16864), .B2(n16761), .A(n16899), .ZN(n16770) );
  NAND2_X1 U19973 ( .A1(n16864), .A2(n18782), .ZN(n16760) );
  INV_X1 U19974 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18784) );
  AOI21_X1 U19975 ( .B1(n16770), .B2(n16760), .A(n18784), .ZN(n16751) );
  NAND3_X1 U19976 ( .A1(n16864), .A2(n16745), .A3(n18784), .ZN(n16748) );
  OAI211_X1 U19977 ( .C1(n16756), .C2(n16749), .A(n16904), .B(n16746), .ZN(
        n16747) );
  OAI211_X1 U19978 ( .C1(n16749), .C2(n16891), .A(n16748), .B(n16747), .ZN(
        n16750) );
  NOR4_X1 U19979 ( .A1(n18210), .A2(n16752), .A3(n16751), .A4(n16750), .ZN(
        n16755) );
  NAND3_X1 U19980 ( .A1(n18736), .A2(n16753), .A3(n17737), .ZN(n16754) );
  OAI211_X1 U19981 ( .C1(n16874), .C2(n17739), .A(n16755), .B(n16754), .ZN(
        P3_U2658) );
  AOI211_X1 U19982 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16773), .A(n16756), .B(
        n16896), .ZN(n16757) );
  AOI21_X1 U19983 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16905), .A(n16757), .ZN(
        n16765) );
  AOI21_X1 U19984 ( .B1(n17759), .B2(n17736), .A(n16758), .ZN(n17757) );
  OAI21_X1 U19985 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17736), .A(
        n10056), .ZN(n16759) );
  XNOR2_X1 U19986 ( .A(n17757), .B(n16759), .ZN(n16763) );
  OAI22_X1 U19987 ( .A1(n17759), .A2(n16874), .B1(n16761), .B2(n16760), .ZN(
        n16762) );
  AOI211_X1 U19988 ( .C1(n18736), .C2(n16763), .A(n18210), .B(n16762), .ZN(
        n16764) );
  OAI211_X1 U19989 ( .C1(n16770), .C2(n18782), .A(n16765), .B(n16764), .ZN(
        P3_U2659) );
  INV_X1 U19990 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16777) );
  INV_X1 U19991 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18778) );
  INV_X1 U19992 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18776) );
  NOR2_X1 U19993 ( .A1(n18778), .A2(n18776), .ZN(n16782) );
  NOR2_X1 U19994 ( .A1(n16892), .A2(n16812), .ZN(n16831) );
  INV_X1 U19995 ( .A(n16831), .ZN(n16766) );
  NOR2_X1 U19996 ( .A1(n16767), .A2(n16766), .ZN(n16795) );
  AOI21_X1 U19997 ( .B1(n16782), .B2(n16795), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16771) );
  INV_X1 U19998 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17780) );
  INV_X1 U19999 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16826) );
  NOR2_X1 U20000 ( .A1(n17893), .A2(n17847), .ZN(n16847) );
  NAND2_X1 U20001 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16847), .ZN(
        n16835) );
  NOR2_X1 U20002 ( .A1(n16826), .A2(n16835), .ZN(n16829) );
  INV_X1 U20003 ( .A(n16829), .ZN(n16814) );
  NOR2_X1 U20004 ( .A1(n17807), .A2(n16814), .ZN(n16800) );
  NAND2_X1 U20005 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16800), .ZN(
        n16790) );
  NOR2_X1 U20006 ( .A1(n17780), .A2(n16790), .ZN(n16783) );
  AOI21_X1 U20007 ( .B1(n16783), .B2(n16861), .A(n16860), .ZN(n16768) );
  OAI21_X1 U20008 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16783), .A(
        n17736), .ZN(n17767) );
  XOR2_X1 U20009 ( .A(n16768), .B(n17767), .Z(n16769) );
  OAI22_X1 U20010 ( .A1(n16771), .A2(n16770), .B1(n16879), .B2(n16769), .ZN(
        n16772) );
  AOI211_X1 U20011 ( .C1(n16905), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18210), .B(
        n16772), .ZN(n16776) );
  OAI211_X1 U20012 ( .C1(n16778), .C2(n16774), .A(n16904), .B(n16773), .ZN(
        n16775) );
  OAI211_X1 U20013 ( .C1(n16874), .C2(n16777), .A(n16776), .B(n16775), .ZN(
        P3_U2660) );
  AOI211_X1 U20014 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16796), .A(n16778), .B(
        n16896), .ZN(n16779) );
  AOI211_X1 U20015 ( .C1(n16905), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18210), .B(
        n16779), .ZN(n16789) );
  OAI21_X1 U20016 ( .B1(n16780), .B2(n16892), .A(n16906), .ZN(n16808) );
  INV_X1 U20017 ( .A(n16795), .ZN(n16781) );
  AOI211_X1 U20018 ( .C1(n18778), .C2(n18776), .A(n16782), .B(n16781), .ZN(
        n16787) );
  AOI21_X1 U20019 ( .B1(n17780), .B2(n16790), .A(n16783), .ZN(n17783) );
  OAI21_X1 U20020 ( .B1(n16790), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n10056), .ZN(n16793) );
  INV_X1 U20021 ( .A(n16793), .ZN(n16785) );
  OAI21_X1 U20022 ( .B1(n17783), .B2(n16785), .A(n18736), .ZN(n16784) );
  AOI21_X1 U20023 ( .B1(n17783), .B2(n16785), .A(n16784), .ZN(n16786) );
  AOI211_X1 U20024 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n16808), .A(n16787), 
        .B(n16786), .ZN(n16788) );
  OAI211_X1 U20025 ( .C1(n17780), .C2(n16874), .A(n16789), .B(n16788), .ZN(
        P3_U2661) );
  AOI22_X1 U20026 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16889), .B1(
        n16905), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n16799) );
  OAI21_X1 U20027 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16800), .A(
        n16790), .ZN(n17795) );
  INV_X1 U20028 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16791) );
  AOI211_X1 U20029 ( .C1(n16791), .C2(n16861), .A(n16860), .B(n17795), .ZN(
        n16792) );
  AOI211_X1 U20030 ( .C1(n16793), .C2(n17795), .A(n16792), .B(n16879), .ZN(
        n16794) );
  AOI221_X1 U20031 ( .B1(n16795), .B2(n18776), .C1(n16808), .C2(
        P3_REIP_REG_9__SCAN_IN), .A(n16794), .ZN(n16798) );
  OAI211_X1 U20032 ( .C1(n16803), .C2(n17161), .A(n16904), .B(n16796), .ZN(
        n16797) );
  NAND4_X1 U20033 ( .A1(n16799), .A2(n16798), .A3(n18108), .A4(n16797), .ZN(
        P3_U2662) );
  INV_X1 U20034 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17821) );
  NOR3_X1 U20035 ( .A1(n17893), .A2(n17820), .A3(n17821), .ZN(n16813) );
  AOI21_X1 U20036 ( .B1(n16813), .B2(n16861), .A(n16860), .ZN(n16802) );
  INV_X1 U20037 ( .A(n16800), .ZN(n16801) );
  OAI21_X1 U20038 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16813), .A(
        n16801), .ZN(n17810) );
  XOR2_X1 U20039 ( .A(n16802), .B(n17810), .Z(n16811) );
  AOI22_X1 U20040 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16889), .B1(
        n16905), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n16810) );
  AOI211_X1 U20041 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16820), .A(n16803), .B(
        n16896), .ZN(n16807) );
  NAND2_X1 U20042 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16819) );
  INV_X1 U20043 ( .A(n16819), .ZN(n16804) );
  NAND3_X1 U20044 ( .A1(n16804), .A2(n18775), .A3(n16831), .ZN(n16805) );
  NAND2_X1 U20045 ( .A1(n18108), .A2(n16805), .ZN(n16806) );
  AOI211_X1 U20046 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n16808), .A(n16807), .B(
        n16806), .ZN(n16809) );
  OAI211_X1 U20047 ( .C1(n16879), .C2(n16811), .A(n16810), .B(n16809), .ZN(
        P3_U2663) );
  INV_X1 U20048 ( .A(n16812), .ZN(n16837) );
  OAI21_X1 U20049 ( .B1(n16837), .B2(n16892), .A(n16906), .ZN(n16843) );
  AOI21_X1 U20050 ( .B1(n17821), .B2(n16814), .A(n16813), .ZN(n17828) );
  AOI21_X1 U20051 ( .B1(n16829), .B2(n16861), .A(n16860), .ZN(n16816) );
  OAI21_X1 U20052 ( .B1(n17828), .B2(n16816), .A(n18736), .ZN(n16815) );
  AOI21_X1 U20053 ( .B1(n17828), .B2(n16816), .A(n16815), .ZN(n16818) );
  OAI22_X1 U20054 ( .A1(n17821), .A2(n16874), .B1(n16891), .B2(n16821), .ZN(
        n16817) );
  AOI211_X1 U20055 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n16843), .A(n16818), .B(
        n16817), .ZN(n16824) );
  OAI211_X1 U20056 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16831), .B(n16819), .ZN(n16823) );
  OAI211_X1 U20057 ( .C1(n16825), .C2(n16821), .A(n16904), .B(n16820), .ZN(
        n16822) );
  NAND4_X1 U20058 ( .A1(n16824), .A2(n18108), .A3(n16823), .A4(n16822), .ZN(
        P3_U2664) );
  AOI21_X1 U20059 ( .B1(n16826), .B2(n16835), .A(n16829), .ZN(n17840) );
  OAI21_X1 U20060 ( .B1(n16826), .B2(n16860), .A(n17840), .ZN(n16834) );
  AOI211_X1 U20061 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16844), .A(n16825), .B(
        n16896), .ZN(n16828) );
  OAI22_X1 U20062 ( .A1(n16826), .A2(n16874), .B1(n16891), .B2(n17231), .ZN(
        n16827) );
  NOR3_X1 U20063 ( .A1(n18210), .A2(n16828), .A3(n16827), .ZN(n16833) );
  INV_X1 U20064 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18770) );
  NAND2_X1 U20065 ( .A1(n10056), .A2(n18736), .ZN(n16888) );
  AOI211_X1 U20066 ( .C1(n16829), .C2(n16861), .A(n17840), .B(n16888), .ZN(
        n16830) );
  AOI221_X1 U20067 ( .B1(n16831), .B2(n18770), .C1(n16843), .C2(
        P3_REIP_REG_6__SCAN_IN), .A(n16830), .ZN(n16832) );
  OAI211_X1 U20068 ( .C1(n16902), .C2(n16834), .A(n16833), .B(n16832), .ZN(
        P3_U2665) );
  OAI21_X1 U20069 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16847), .A(
        n16835), .ZN(n17850) );
  INV_X1 U20070 ( .A(n16847), .ZN(n16836) );
  OAI21_X1 U20071 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16836), .A(
        n10056), .ZN(n16849) );
  XNOR2_X1 U20072 ( .A(n17850), .B(n16849), .ZN(n16841) );
  NOR2_X1 U20073 ( .A1(n16837), .A2(n16892), .ZN(n16838) );
  AOI22_X1 U20074 ( .A1(n16905), .A2(P3_EBX_REG_5__SCAN_IN), .B1(n16839), .B2(
        n16838), .ZN(n16840) );
  OAI211_X1 U20075 ( .C1(n16879), .C2(n16841), .A(n16840), .B(n18108), .ZN(
        n16842) );
  AOI21_X1 U20076 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n16843), .A(n16842), .ZN(
        n16846) );
  OAI211_X1 U20077 ( .C1(n16851), .C2(n17240), .A(n16904), .B(n16844), .ZN(
        n16845) );
  OAI211_X1 U20078 ( .C1(n16874), .C2(n17846), .A(n16846), .B(n16845), .ZN(
        P3_U2666) );
  AOI21_X1 U20079 ( .B1(n16864), .B2(n16852), .A(n16899), .ZN(n16866) );
  NAND2_X1 U20080 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10042), .ZN(
        n16859) );
  AOI21_X1 U20081 ( .B1(n10045), .B2(n16859), .A(n16847), .ZN(n17863) );
  NAND2_X1 U20082 ( .A1(n10042), .A2(n10045), .ZN(n17860) );
  OAI22_X1 U20083 ( .A1(n17863), .A2(n16849), .B1(n16848), .B2(n17860), .ZN(
        n16850) );
  OAI221_X1 U20084 ( .B1(n16850), .B2(n17863), .C1(n16850), .C2(n16860), .A(
        n18736), .ZN(n16858) );
  AOI211_X1 U20085 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16870), .A(n16851), .B(
        n16896), .ZN(n16856) );
  NAND2_X1 U20086 ( .A1(n18237), .A2(n18899), .ZN(n16895) );
  INV_X1 U20087 ( .A(n16895), .ZN(n18901) );
  NOR3_X1 U20088 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16892), .A3(n16852), .ZN(
        n16853) );
  AOI221_X1 U20089 ( .B1(n17147), .B2(n18901), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18901), .A(n16853), .ZN(
        n16854) );
  OAI211_X1 U20090 ( .C1(n10045), .C2(n16874), .A(n16854), .B(n18108), .ZN(
        n16855) );
  AOI211_X1 U20091 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16905), .A(n16856), .B(
        n16855), .ZN(n16857) );
  OAI211_X1 U20092 ( .C1(n16866), .C2(n18766), .A(n16858), .B(n16857), .ZN(
        P3_U2667) );
  NAND2_X1 U20093 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16876) );
  INV_X1 U20094 ( .A(n16876), .ZN(n16862) );
  OAI21_X1 U20095 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16862), .A(
        n16859), .ZN(n17872) );
  AOI21_X1 U20096 ( .B1(n16862), .B2(n16861), .A(n16860), .ZN(n16863) );
  XNOR2_X1 U20097 ( .A(n17872), .B(n16863), .ZN(n16869) );
  NAND3_X1 U20098 ( .A1(n16864), .A2(P3_REIP_REG_1__SCAN_IN), .A3(
        P3_REIP_REG_2__SCAN_IN), .ZN(n16867) );
  INV_X1 U20099 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18764) );
  NOR2_X1 U20100 ( .A1(n18859), .A2(n18852), .ZN(n18676) );
  NAND2_X1 U20101 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18676), .ZN(
        n18671) );
  AOI21_X1 U20102 ( .B1(n18841), .B2(n18671), .A(n17147), .ZN(n18838) );
  AOI22_X1 U20103 ( .A1(n16905), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n18901), .B2(
        n18838), .ZN(n16865) );
  OAI221_X1 U20104 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n16867), .C1(n18764), 
        .C2(n16866), .A(n16865), .ZN(n16868) );
  AOI21_X1 U20105 ( .B1(n16869), .B2(n18736), .A(n16868), .ZN(n16872) );
  OAI211_X1 U20106 ( .C1(n16877), .C2(n17246), .A(n16904), .B(n16870), .ZN(
        n16871) );
  OAI211_X1 U20107 ( .C1(n16874), .C2(n16873), .A(n16872), .B(n16871), .ZN(
        P3_U2668) );
  OAI21_X1 U20108 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16876), .ZN(n17883) );
  OAI22_X1 U20109 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16876), .B1(
        n16875), .B2(n17883), .ZN(n16887) );
  AOI22_X1 U20110 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16889), .B1(
        n16905), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n16886) );
  NAND2_X1 U20111 ( .A1(n17268), .A2(n17262), .ZN(n16878) );
  AOI211_X1 U20112 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16878), .A(n16877), .B(
        n16896), .ZN(n16884) );
  NOR3_X1 U20113 ( .A1(n10056), .A2(n16879), .A3(n17883), .ZN(n16883) );
  INV_X1 U20114 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18762) );
  AOI221_X1 U20115 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_2__SCAN_IN), 
        .C1(n18868), .C2(n18762), .A(n16892), .ZN(n16882) );
  NAND2_X1 U20116 ( .A1(n18852), .A2(n18675), .ZN(n18669) );
  NAND2_X1 U20117 ( .A1(n18671), .A2(n18669), .ZN(n18845) );
  OAI22_X1 U20118 ( .A1(n16906), .A2(n18762), .B1(n18845), .B2(n16895), .ZN(
        n16881) );
  NOR4_X1 U20119 ( .A1(n16884), .A2(n16883), .A3(n16882), .A4(n16881), .ZN(
        n16885) );
  OAI211_X1 U20120 ( .C1(n16888), .C2(n16887), .A(n16886), .B(n16885), .ZN(
        P3_U2669) );
  AOI21_X1 U20121 ( .B1(n18736), .B2(n16890), .A(n16889), .ZN(n16901) );
  OAI22_X1 U20122 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16892), .B1(n16891), 
        .B2(n17262), .ZN(n16898) );
  AOI21_X1 U20123 ( .B1(n17268), .B2(n17262), .A(n17245), .ZN(n16893) );
  INV_X1 U20124 ( .A(n16893), .ZN(n17263) );
  NAND2_X1 U20125 ( .A1(n16894), .A2(n18675), .ZN(n18853) );
  OAI22_X1 U20126 ( .A1(n16896), .A2(n17263), .B1(n18853), .B2(n16895), .ZN(
        n16897) );
  AOI211_X1 U20127 ( .C1(n16899), .C2(P3_REIP_REG_1__SCAN_IN), .A(n16898), .B(
        n16897), .ZN(n16900) );
  OAI221_X1 U20128 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16902), .C1(
        n17893), .C2(n16901), .A(n16900), .ZN(P3_U2670) );
  AOI22_X1 U20129 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16903), .B1(n18901), 
        .B2(n18866), .ZN(n16909) );
  OAI21_X1 U20130 ( .B1(n16905), .B2(n16904), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16908) );
  INV_X1 U20131 ( .A(n18862), .ZN(n18847) );
  NAND3_X1 U20132 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18847), .A3(
        n16906), .ZN(n16907) );
  NAND3_X1 U20133 ( .A1(n16909), .A2(n16908), .A3(n16907), .ZN(P3_U2671) );
  INV_X1 U20134 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16910) );
  NOR2_X1 U20135 ( .A1(n16910), .A2(n17045), .ZN(n17029) );
  NAND4_X1 U20136 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n16911)
         );
  NOR4_X1 U20137 ( .A1(n16955), .A2(n16913), .A3(n16912), .A4(n16911), .ZN(
        n16914) );
  NAND4_X1 U20138 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17029), .A4(n16914), .ZN(n16917) );
  NOR2_X1 U20139 ( .A1(n16918), .A2(n16917), .ZN(n16947) );
  NAND2_X1 U20140 ( .A1(n17260), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16916) );
  NAND2_X1 U20141 ( .A1(n16947), .A2(n18268), .ZN(n16915) );
  OAI22_X1 U20142 ( .A1(n16947), .A2(n16916), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16915), .ZN(P3_U2672) );
  NAND2_X1 U20143 ( .A1(n16918), .A2(n16917), .ZN(n16919) );
  NAND2_X1 U20144 ( .A1(n16919), .A2(n17256), .ZN(n16946) );
  AOI22_X1 U20145 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16920) );
  OAI21_X1 U20146 ( .B1(n16984), .B2(n17116), .A(n16920), .ZN(n16931) );
  AOI22_X1 U20147 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U20148 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16921) );
  OAI21_X1 U20149 ( .B1(n12307), .B2(n16922), .A(n16921), .ZN(n16927) );
  AOI22_X1 U20150 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16924) );
  AOI22_X1 U20151 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16923) );
  OAI211_X1 U20152 ( .C1(n17172), .C2(n16925), .A(n16924), .B(n16923), .ZN(
        n16926) );
  AOI211_X1 U20153 ( .C1(n17195), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n16927), .B(n16926), .ZN(n16928) );
  OAI211_X1 U20154 ( .C1(n9695), .C2(n17123), .A(n16929), .B(n16928), .ZN(
        n16930) );
  AOI211_X1 U20155 ( .C1(n17173), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n16931), .B(n16930), .ZN(n16951) );
  NOR2_X1 U20156 ( .A1(n16951), .A2(n16950), .ZN(n16949) );
  AOI22_X1 U20157 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17192), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n15698), .ZN(n16943) );
  AOI22_X1 U20158 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17186), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16932) );
  OAI21_X1 U20159 ( .B1(n12308), .B2(n16933), .A(n16932), .ZN(n16941) );
  OAI22_X1 U20160 ( .A1(n16934), .A2(n12307), .B1(n17235), .B2(n17181), .ZN(
        n16935) );
  AOI21_X1 U20161 ( .B1(n17030), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n16935), .ZN(n16939) );
  AOI22_X1 U20162 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17165), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n9646), .ZN(n16938) );
  AOI22_X1 U20163 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17194), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17147), .ZN(n16937) );
  AOI22_X1 U20164 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17195), .B1(
        n9659), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16936) );
  NAND4_X1 U20165 ( .A1(n16939), .A2(n16938), .A3(n16937), .A4(n16936), .ZN(
        n16940) );
  AOI211_X1 U20166 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n16941), .B(n16940), .ZN(n16942) );
  OAI211_X1 U20167 ( .C1(n16944), .C2(n17172), .A(n16943), .B(n16942), .ZN(
        n16945) );
  XNOR2_X1 U20168 ( .A(n16949), .B(n16945), .ZN(n17279) );
  OAI22_X1 U20169 ( .A1(n16947), .A2(n16946), .B1(n17279), .B2(n17256), .ZN(
        P3_U2673) );
  INV_X1 U20170 ( .A(n16948), .ZN(n16954) );
  AOI21_X1 U20171 ( .B1(n16951), .B2(n16950), .A(n16949), .ZN(n17283) );
  AOI22_X1 U20172 ( .A1(n17266), .A2(n17283), .B1(n16952), .B2(n16955), .ZN(
        n16953) );
  OAI21_X1 U20173 ( .B1(n16955), .B2(n16954), .A(n16953), .ZN(P3_U2674) );
  INV_X1 U20174 ( .A(n16956), .ZN(n16965) );
  AOI21_X1 U20175 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17256), .A(n16965), .ZN(
        n16960) );
  AOI21_X1 U20176 ( .B1(n16958), .B2(n16962), .A(n16957), .ZN(n17291) );
  INV_X1 U20177 ( .A(n17291), .ZN(n16959) );
  OAI22_X1 U20178 ( .A1(n16961), .A2(n16960), .B1(n16959), .B2(n17256), .ZN(
        P3_U2676) );
  AOI21_X1 U20179 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17256), .A(n16971), .ZN(
        n16964) );
  OAI21_X1 U20180 ( .B1(n16967), .B2(n16963), .A(n16962), .ZN(n17299) );
  OAI22_X1 U20181 ( .A1(n16965), .A2(n16964), .B1(n17299), .B2(n17256), .ZN(
        P3_U2677) );
  INV_X1 U20182 ( .A(n16966), .ZN(n16975) );
  AOI21_X1 U20183 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17256), .A(n16975), .ZN(
        n16970) );
  AOI21_X1 U20184 ( .B1(n16968), .B2(n16972), .A(n16967), .ZN(n17300) );
  INV_X1 U20185 ( .A(n17300), .ZN(n16969) );
  OAI22_X1 U20186 ( .A1(n16971), .A2(n16970), .B1(n16969), .B2(n17256), .ZN(
        P3_U2678) );
  AOI21_X1 U20187 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17260), .A(n16982), .ZN(
        n16974) );
  OAI21_X1 U20188 ( .B1(n16977), .B2(n16973), .A(n16972), .ZN(n17310) );
  OAI22_X1 U20189 ( .A1(n16975), .A2(n16974), .B1(n17310), .B2(n17256), .ZN(
        P3_U2679) );
  INV_X1 U20190 ( .A(n16976), .ZN(n16997) );
  AOI21_X1 U20191 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17260), .A(n16997), .ZN(
        n16981) );
  AOI21_X1 U20192 ( .B1(n16979), .B2(n16978), .A(n16977), .ZN(n17314) );
  INV_X1 U20193 ( .A(n17314), .ZN(n16980) );
  OAI22_X1 U20194 ( .A1(n16982), .A2(n16981), .B1(n16980), .B2(n17260), .ZN(
        P3_U2680) );
  AOI21_X1 U20195 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17260), .A(n16983), .ZN(
        n16996) );
  AOI22_X1 U20196 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20197 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20198 ( .A1(n9659), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16992) );
  INV_X1 U20199 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17237) );
  OAI22_X1 U20200 ( .A1(n16984), .A2(n17114), .B1(n17133), .B2(n17237), .ZN(
        n16990) );
  AOI22_X1 U20201 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20202 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20203 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16986) );
  NAND2_X1 U20204 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n16985) );
  NAND4_X1 U20205 ( .A1(n16988), .A2(n16987), .A3(n16986), .A4(n16985), .ZN(
        n16989) );
  AOI211_X1 U20206 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n16990), .B(n16989), .ZN(n16991) );
  NAND4_X1 U20207 ( .A1(n16994), .A2(n16993), .A3(n16992), .A4(n16991), .ZN(
        n17317) );
  INV_X1 U20208 ( .A(n17317), .ZN(n16995) );
  OAI22_X1 U20209 ( .A1(n16997), .A2(n16996), .B1(n16995), .B2(n17256), .ZN(
        P3_U2681) );
  AOI22_X1 U20210 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16998) );
  OAI21_X1 U20211 ( .B1(n10260), .B2(n16999), .A(n16998), .ZN(n17010) );
  AOI22_X1 U20212 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17169), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20213 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17000) );
  OAI21_X1 U20214 ( .B1(n17133), .B2(n17242), .A(n17000), .ZN(n17005) );
  AOI22_X1 U20215 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20216 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17001) );
  OAI211_X1 U20217 ( .C1(n17172), .C2(n17003), .A(n17002), .B(n17001), .ZN(
        n17004) );
  AOI211_X1 U20218 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17005), .B(n17004), .ZN(n17006) );
  OAI211_X1 U20219 ( .C1(n21028), .C2(n17008), .A(n17007), .B(n17006), .ZN(
        n17009) );
  AOI211_X1 U20220 ( .C1(n17165), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n17010), .B(n17009), .ZN(n17324) );
  INV_X1 U20221 ( .A(n17324), .ZN(n17013) );
  OAI21_X1 U20222 ( .B1(n17011), .B2(n17029), .A(n17256), .ZN(n17012) );
  OAI21_X1 U20223 ( .B1(n17260), .B2(n17013), .A(n17012), .ZN(n17014) );
  OAI21_X1 U20224 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17015), .A(n17014), .ZN(
        P3_U2682) );
  AOI21_X1 U20225 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17260), .A(n17016), .ZN(
        n17028) );
  AOI22_X1 U20226 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17017) );
  OAI21_X1 U20227 ( .B1(n9695), .B2(n17131), .A(n17017), .ZN(n17027) );
  AOI22_X1 U20228 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17024) );
  OAI22_X1 U20229 ( .A1(n17215), .A2(n17130), .B1(n17181), .B2(n17132), .ZN(
        n17022) );
  AOI22_X1 U20230 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17020) );
  AOI22_X1 U20231 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20232 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9659), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17018) );
  NAND3_X1 U20233 ( .A1(n17020), .A2(n17019), .A3(n17018), .ZN(n17021) );
  AOI211_X1 U20234 ( .C1(n17169), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n17022), .B(n17021), .ZN(n17023) );
  OAI211_X1 U20235 ( .C1(n12308), .C2(n17025), .A(n17024), .B(n17023), .ZN(
        n17026) );
  AOI211_X1 U20236 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n17027), .B(n17026), .ZN(n17331) );
  OAI22_X1 U20237 ( .A1(n17029), .A2(n17028), .B1(n17331), .B2(n17260), .ZN(
        P3_U2683) );
  AOI22_X1 U20238 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17031) );
  OAI21_X1 U20239 ( .B1(n10260), .B2(n17032), .A(n17031), .ZN(n17043) );
  INV_X1 U20240 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U20241 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17041) );
  OAI22_X1 U20242 ( .A1(n12308), .A2(n17034), .B1(n17172), .B2(n17033), .ZN(
        n17039) );
  AOI22_X1 U20243 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20244 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17036) );
  AOI22_X1 U20245 ( .A1(n9659), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17035) );
  NAND3_X1 U20246 ( .A1(n17037), .A2(n17036), .A3(n17035), .ZN(n17038) );
  AOI211_X1 U20247 ( .C1(n17169), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n17039), .B(n17038), .ZN(n17040) );
  OAI211_X1 U20248 ( .C1(n17133), .C2(n17251), .A(n17041), .B(n17040), .ZN(
        n17042) );
  AOI211_X1 U20249 ( .C1(n17044), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n17043), .B(n17042), .ZN(n17336) );
  OAI21_X1 U20250 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17057), .A(n17045), .ZN(
        n17046) );
  AOI22_X1 U20251 ( .A1(n17266), .A2(n17336), .B1(n17046), .B2(n17256), .ZN(
        P3_U2684) );
  AOI22_X1 U20252 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20253 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20254 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17047) );
  OAI211_X1 U20255 ( .C1(n17215), .C2(n17167), .A(n17048), .B(n17047), .ZN(
        n17054) );
  AOI22_X1 U20256 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20257 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17051) );
  AOI22_X1 U20258 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17169), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17050) );
  NAND2_X1 U20259 ( .A1(n9659), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n17049) );
  NAND4_X1 U20260 ( .A1(n17052), .A2(n17051), .A3(n17050), .A4(n17049), .ZN(
        n17053) );
  AOI211_X1 U20261 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17054), .B(n17053), .ZN(n17055) );
  OAI211_X1 U20262 ( .C1(n17133), .C2(n17257), .A(n17056), .B(n17055), .ZN(
        n17338) );
  AOI21_X1 U20263 ( .B1(n17059), .B2(n17058), .A(n17057), .ZN(n17060) );
  MUX2_X1 U20264 ( .A(n17338), .B(n17060), .S(n17256), .Z(P3_U2685) );
  AOI22_X1 U20265 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20266 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20267 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17061) );
  OAI211_X1 U20268 ( .C1(n17215), .C2(n17063), .A(n17062), .B(n17061), .ZN(
        n17069) );
  AOI22_X1 U20269 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20270 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20271 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17065) );
  NAND2_X1 U20272 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n17064) );
  NAND4_X1 U20273 ( .A1(n17067), .A2(n17066), .A3(n17065), .A4(n17064), .ZN(
        n17068) );
  AOI211_X1 U20274 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n17069), .B(n17068), .ZN(n17070) );
  OAI211_X1 U20275 ( .C1(n17133), .C2(n17261), .A(n17071), .B(n17070), .ZN(
        n17346) );
  NAND2_X1 U20276 ( .A1(n18268), .A2(n17269), .ZN(n17264) );
  INV_X1 U20277 ( .A(n17264), .ZN(n17265) );
  AOI21_X1 U20278 ( .B1(n17076), .B2(n17073), .A(n17072), .ZN(n17074) );
  AOI22_X1 U20279 ( .A1(n17266), .A2(n17346), .B1(n17265), .B2(n17074), .ZN(
        n17075) );
  OAI21_X1 U20280 ( .B1(n17269), .B2(n17076), .A(n17075), .ZN(P3_U2686) );
  AOI22_X1 U20281 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17077) );
  OAI21_X1 U20282 ( .B1(n10260), .B2(n17078), .A(n17077), .ZN(n17090) );
  AOI22_X1 U20283 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17088) );
  OAI22_X1 U20284 ( .A1(n17080), .A2(n17079), .B1(n10251), .B2(n17226), .ZN(
        n17085) );
  AOI22_X1 U20285 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20286 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20287 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9659), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17081) );
  NAND3_X1 U20288 ( .A1(n17083), .A2(n17082), .A3(n17081), .ZN(n17084) );
  AOI211_X1 U20289 ( .C1(n17086), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n17085), .B(n17084), .ZN(n17087) );
  OAI211_X1 U20290 ( .C1(n17133), .C2(n17214), .A(n17088), .B(n17087), .ZN(
        n17089) );
  AOI211_X1 U20291 ( .C1(n17187), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17090), .B(n17089), .ZN(n17354) );
  NOR2_X1 U20292 ( .A1(n17240), .A2(n17239), .ZN(n17244) );
  NAND3_X1 U20293 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(n17244), .ZN(n17232) );
  NOR2_X1 U20294 ( .A1(n17091), .A2(n17232), .ZN(n17163) );
  NAND2_X1 U20295 ( .A1(n17092), .A2(n17163), .ZN(n17093) );
  NAND2_X1 U20296 ( .A1(n17260), .A2(n17093), .ZN(n17110) );
  INV_X1 U20297 ( .A(n17110), .ZN(n17095) );
  NOR3_X1 U20298 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17365), .A3(n17093), .ZN(
        n17094) );
  AOI21_X1 U20299 ( .B1(n17095), .B2(P3_EBX_REG_16__SCAN_IN), .A(n17094), .ZN(
        n17096) );
  OAI21_X1 U20300 ( .B1(n17354), .B2(n17256), .A(n17096), .ZN(P3_U2687) );
  AOI22_X1 U20301 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17147), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17191), .ZN(n17109) );
  AOI22_X1 U20302 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9646), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17108) );
  OAI22_X1 U20303 ( .A1(n17172), .A2(n17098), .B1(n17133), .B2(n17097), .ZN(
        n17106) );
  AOI22_X1 U20304 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17169), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17103) );
  AOI22_X1 U20305 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17194), .ZN(n17100) );
  AOI22_X1 U20306 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17186), .ZN(n17099) );
  OAI211_X1 U20307 ( .C1(n17215), .C2(n17235), .A(n17100), .B(n17099), .ZN(
        n17101) );
  AOI21_X1 U20308 ( .B1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n9659), .A(
        n17101), .ZN(n17102) );
  OAI211_X1 U20309 ( .C1(n12308), .C2(n17104), .A(n17103), .B(n17102), .ZN(
        n17105) );
  AOI211_X1 U20310 ( .C1(n17187), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n17106), .B(n17105), .ZN(n17107) );
  NAND3_X1 U20311 ( .A1(n17109), .A2(n17108), .A3(n17107), .ZN(n17355) );
  INV_X1 U20312 ( .A(n17355), .ZN(n17112) );
  AND3_X1 U20313 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n17163), .ZN(n17126) );
  AND2_X1 U20314 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17126), .ZN(n17128) );
  NOR2_X1 U20315 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17128), .ZN(n17111) );
  OAI22_X1 U20316 ( .A1(n17112), .A2(n17260), .B1(n17111), .B2(n17110), .ZN(
        P3_U2688) );
  AOI22_X1 U20317 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17113) );
  OAI21_X1 U20318 ( .B1(n10251), .B2(n17114), .A(n17113), .ZN(n17125) );
  AOI22_X1 U20319 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20320 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17115) );
  OAI21_X1 U20321 ( .B1(n12307), .B2(n17116), .A(n17115), .ZN(n17120) );
  AOI22_X1 U20322 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20323 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17117) );
  OAI211_X1 U20324 ( .C1(n17215), .C2(n17237), .A(n17118), .B(n17117), .ZN(
        n17119) );
  AOI211_X1 U20325 ( .C1(n9659), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17120), .B(n17119), .ZN(n17121) );
  OAI211_X1 U20326 ( .C1(n17133), .C2(n17123), .A(n17122), .B(n17121), .ZN(
        n17124) );
  AOI211_X1 U20327 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n17125), .B(n17124), .ZN(n17363) );
  OAI21_X1 U20328 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17126), .A(n17256), .ZN(
        n17127) );
  OAI22_X1 U20329 ( .A1(n17363), .A2(n17256), .B1(n17128), .B2(n17127), .ZN(
        P3_U2689) );
  AOI22_X1 U20330 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17129) );
  OAI21_X1 U20331 ( .B1(n17168), .B2(n17130), .A(n17129), .ZN(n17143) );
  AOI22_X1 U20332 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17140) );
  OAI22_X1 U20333 ( .A1(n17133), .A2(n17132), .B1(n17181), .B2(n17131), .ZN(
        n17138) );
  AOI22_X1 U20334 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20335 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20336 ( .A1(n9659), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17134) );
  NAND3_X1 U20337 ( .A1(n17136), .A2(n17135), .A3(n17134), .ZN(n17137) );
  AOI211_X1 U20338 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17138), .B(n17137), .ZN(n17139) );
  OAI211_X1 U20339 ( .C1(n12307), .C2(n17141), .A(n17140), .B(n17139), .ZN(
        n17142) );
  AOI211_X1 U20340 ( .C1(n17186), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n17143), .B(n17142), .ZN(n17372) );
  NOR2_X1 U20341 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17163), .ZN(n17146) );
  NAND2_X1 U20342 ( .A1(n17260), .A2(n17144), .ZN(n17145) );
  OAI22_X1 U20343 ( .A1(n17372), .A2(n17256), .B1(n17146), .B2(n17145), .ZN(
        P3_U2691) );
  AOI22_X1 U20344 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20345 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20346 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17148) );
  OAI211_X1 U20347 ( .C1(n17215), .C2(n17251), .A(n17149), .B(n17148), .ZN(
        n17157) );
  AOI22_X1 U20348 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20349 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20350 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17153) );
  NAND2_X1 U20351 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n17152) );
  NAND4_X1 U20352 ( .A1(n17155), .A2(n17154), .A3(n17153), .A4(n17152), .ZN(
        n17156) );
  AOI211_X1 U20353 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17157), .B(n17156), .ZN(n17158) );
  OAI211_X1 U20354 ( .C1(n10260), .C2(n17160), .A(n17159), .B(n17158), .ZN(
        n17376) );
  INV_X1 U20355 ( .A(n17376), .ZN(n17164) );
  INV_X1 U20356 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17228) );
  NOR3_X1 U20357 ( .A1(n17161), .A2(n17228), .A3(n17232), .ZN(n17206) );
  AND2_X1 U20358 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17206), .ZN(n17185) );
  OAI21_X1 U20359 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17185), .A(n17256), .ZN(
        n17162) );
  OAI22_X1 U20360 ( .A1(n17164), .A2(n17260), .B1(n17163), .B2(n17162), .ZN(
        P3_U2692) );
  AOI22_X1 U20361 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15698), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17166) );
  OAI21_X1 U20362 ( .B1(n17168), .B2(n17167), .A(n17166), .ZN(n17183) );
  AOI22_X1 U20363 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17169), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17179) );
  INV_X1 U20364 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17171) );
  AOI22_X1 U20365 ( .A1(n9657), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17170) );
  OAI21_X1 U20366 ( .B1(n17172), .B2(n17171), .A(n17170), .ZN(n17177) );
  AOI22_X1 U20367 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20368 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9646), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17174) );
  OAI211_X1 U20369 ( .C1(n17215), .C2(n17257), .A(n17175), .B(n17174), .ZN(
        n17176) );
  AOI211_X1 U20370 ( .C1(n9658), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17177), .B(n17176), .ZN(n17178) );
  OAI211_X1 U20371 ( .C1(n17181), .C2(n17180), .A(n17179), .B(n17178), .ZN(
        n17182) );
  AOI211_X1 U20372 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n17183), .B(n17182), .ZN(n17379) );
  OAI21_X1 U20373 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17206), .A(n17256), .ZN(
        n17184) );
  OAI22_X1 U20374 ( .A1(n17379), .A2(n17260), .B1(n17185), .B2(n17184), .ZN(
        P3_U2693) );
  AOI22_X1 U20375 ( .A1(n17187), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17186), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17188) );
  OAI21_X1 U20376 ( .B1(n17190), .B2(n17189), .A(n17188), .ZN(n17205) );
  AOI22_X1 U20377 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20378 ( .A1(n17169), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9659), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17193) );
  INV_X1 U20379 ( .A(n17193), .ZN(n17200) );
  AOI22_X1 U20380 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U20381 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20382 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17196) );
  NAND3_X1 U20383 ( .A1(n17198), .A2(n17197), .A3(n17196), .ZN(n17199) );
  AOI211_X1 U20384 ( .C1(n17210), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n17200), .B(n17199), .ZN(n17201) );
  OAI211_X1 U20385 ( .C1(n21028), .C2(n17203), .A(n17202), .B(n17201), .ZN(
        n17204) );
  AOI211_X1 U20386 ( .C1(n17030), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n17205), .B(n17204), .ZN(n17386) );
  NOR2_X1 U20387 ( .A1(n17228), .A2(n17232), .ZN(n17208) );
  INV_X1 U20388 ( .A(n17206), .ZN(n17207) );
  OAI21_X1 U20389 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17208), .A(n17207), .ZN(
        n17209) );
  AOI22_X1 U20390 ( .A1(n17266), .A2(n17386), .B1(n17209), .B2(n17256), .ZN(
        P3_U2694) );
  AOI22_X1 U20391 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20392 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20393 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17212) );
  OAI211_X1 U20394 ( .C1(n17215), .C2(n17214), .A(n17213), .B(n17212), .ZN(
        n17223) );
  AOI22_X1 U20395 ( .A1(n15698), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17216), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20396 ( .A1(n9646), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17220) );
  AOI22_X1 U20397 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17219) );
  NAND2_X1 U20398 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n17218) );
  NAND4_X1 U20399 ( .A1(n17221), .A2(n17220), .A3(n17219), .A4(n17218), .ZN(
        n17222) );
  AOI211_X1 U20400 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17223), .B(n17222), .ZN(n17224) );
  OAI211_X1 U20401 ( .C1(n12307), .C2(n17226), .A(n17225), .B(n17224), .ZN(
        n17390) );
  INV_X1 U20402 ( .A(n17232), .ZN(n17227) );
  OAI33_X1 U20403 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17365), .A3(n17232), .B1(
        n17228), .B2(n17266), .B3(n17227), .ZN(n17229) );
  AOI21_X1 U20404 ( .B1(n17266), .B2(n17390), .A(n17229), .ZN(n17230) );
  INV_X1 U20405 ( .A(n17230), .ZN(P3_U2695) );
  NAND2_X1 U20406 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17249), .ZN(n17238) );
  NOR2_X1 U20407 ( .A1(n17231), .A2(n17238), .ZN(n17233) );
  OAI211_X1 U20408 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n17233), .A(n17232), .B(
        n17256), .ZN(n17234) );
  OAI21_X1 U20409 ( .B1(n17260), .B2(n17235), .A(n17234), .ZN(P3_U2696) );
  NAND3_X1 U20410 ( .A1(n17238), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17260), .ZN(
        n17236) );
  OAI221_X1 U20411 ( .B1(n17238), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17260), 
        .C2(n17237), .A(n17236), .ZN(P3_U2697) );
  AOI21_X1 U20412 ( .B1(n17240), .B2(n17239), .A(n17266), .ZN(n17241) );
  INV_X1 U20413 ( .A(n17241), .ZN(n17243) );
  OAI22_X1 U20414 ( .A1(n17244), .A2(n17243), .B1(n17242), .B2(n17256), .ZN(
        P3_U2698) );
  INV_X1 U20415 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17250) );
  NAND2_X1 U20416 ( .A1(n17245), .A2(n17265), .ZN(n17254) );
  NOR3_X1 U20417 ( .A1(n17246), .A2(n17250), .A3(n17254), .ZN(n17253) );
  AOI21_X1 U20418 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17260), .A(n17253), .ZN(
        n17248) );
  OAI22_X1 U20419 ( .A1(n17249), .A2(n17248), .B1(n17247), .B2(n17256), .ZN(
        P3_U2699) );
  NOR2_X1 U20420 ( .A1(n17250), .A2(n17254), .ZN(n17259) );
  AOI21_X1 U20421 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17260), .A(n17259), .ZN(
        n17252) );
  OAI22_X1 U20422 ( .A1(n17253), .A2(n17252), .B1(n17251), .B2(n17256), .ZN(
        P3_U2700) );
  INV_X1 U20423 ( .A(n17254), .ZN(n17255) );
  AOI21_X1 U20424 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17256), .A(n17255), .ZN(
        n17258) );
  OAI22_X1 U20425 ( .A1(n17259), .A2(n17258), .B1(n17257), .B2(n17256), .ZN(
        P3_U2701) );
  OAI222_X1 U20426 ( .A1(n17264), .A2(n17263), .B1(n17262), .B2(n17269), .C1(
        n17261), .C2(n17260), .ZN(P3_U2702) );
  AOI22_X1 U20427 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17266), .B1(
        n17265), .B2(n17268), .ZN(n17267) );
  OAI21_X1 U20428 ( .B1(n17269), .B2(n17268), .A(n17267), .ZN(P3_U2703) );
  INV_X1 U20429 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17492) );
  INV_X1 U20430 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17488) );
  INV_X1 U20431 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17486) );
  INV_X1 U20432 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17484) );
  INV_X1 U20433 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17470) );
  INV_X1 U20434 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17529) );
  NAND3_X1 U20435 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n17272) );
  NAND4_X1 U20436 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17271) );
  INV_X1 U20437 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17527) );
  INV_X1 U20438 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17525) );
  INV_X1 U20439 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17517) );
  INV_X1 U20440 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17515) );
  NOR4_X1 U20441 ( .A1(n17527), .A2(n17525), .A3(n17517), .A4(n17515), .ZN(
        n17273) );
  INV_X1 U20442 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17482) );
  INV_X1 U20443 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17480) );
  INV_X1 U20444 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17478) );
  INV_X1 U20445 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17472) );
  NAND2_X1 U20446 ( .A1(n18268), .A2(n17311), .ZN(n17305) );
  NOR2_X1 U20447 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n9693), .ZN(n17275) );
  NAND2_X1 U20448 ( .A1(n17412), .A2(n9693), .ZN(n17282) );
  OAI21_X1 U20449 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17421), .A(n17282), .ZN(
        n17274) );
  AOI22_X1 U20450 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17275), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17274), .ZN(n17276) );
  OAI21_X1 U20451 ( .B1(n17277), .B2(n17322), .A(n17276), .ZN(P3_U2704) );
  INV_X1 U20452 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17498) );
  NOR2_X2 U20453 ( .A1(n17278), .A2(n17412), .ZN(n17350) );
  INV_X1 U20454 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18260) );
  OAI22_X1 U20455 ( .A1(n17279), .A2(n17414), .B1(n18260), .B2(n17322), .ZN(
        n17280) );
  AOI21_X1 U20456 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17350), .A(n17280), .ZN(
        n17281) );
  OAI221_X1 U20457 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n9693), .C1(n17498), 
        .C2(n17282), .A(n17281), .ZN(P3_U2705) );
  INV_X1 U20458 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19298) );
  AOI22_X1 U20459 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17350), .B1(n17419), .B2(
        n17283), .ZN(n17286) );
  OAI211_X1 U20460 ( .C1(n17284), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17412), .B(
        n9693), .ZN(n17285) );
  OAI211_X1 U20461 ( .C1(n17322), .C2(n19298), .A(n17286), .B(n17285), .ZN(
        P3_U2706) );
  AOI22_X1 U20462 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17349), .ZN(n17289) );
  OAI211_X1 U20463 ( .C1(n17292), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17412), .B(
        n17287), .ZN(n17288) );
  OAI211_X1 U20464 ( .C1(n17290), .C2(n17414), .A(n17289), .B(n17288), .ZN(
        P3_U2707) );
  INV_X1 U20465 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18247) );
  AOI22_X1 U20466 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17350), .B1(n17419), .B2(
        n17291), .ZN(n17295) );
  AOI211_X1 U20467 ( .C1(n17492), .C2(n17296), .A(n17292), .B(n17384), .ZN(
        n17293) );
  INV_X1 U20468 ( .A(n17293), .ZN(n17294) );
  OAI211_X1 U20469 ( .C1(n17322), .C2(n18247), .A(n17295), .B(n17294), .ZN(
        P3_U2708) );
  AOI22_X1 U20470 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17349), .ZN(n17298) );
  OAI211_X1 U20471 ( .C1(n17301), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17412), .B(
        n17296), .ZN(n17297) );
  OAI211_X1 U20472 ( .C1(n17299), .C2(n17414), .A(n17298), .B(n17297), .ZN(
        P3_U2709) );
  INV_X1 U20473 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n19283) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17350), .B1(n17419), .B2(
        n17300), .ZN(n17304) );
  AOI211_X1 U20475 ( .C1(n17488), .C2(n17306), .A(n17301), .B(n17384), .ZN(
        n17302) );
  INV_X1 U20476 ( .A(n17302), .ZN(n17303) );
  OAI211_X1 U20477 ( .C1(n17322), .C2(n19283), .A(n17304), .B(n17303), .ZN(
        P3_U2710) );
  AOI22_X1 U20478 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17349), .ZN(n17309) );
  OAI21_X1 U20479 ( .B1(n17486), .B2(n17384), .A(n17305), .ZN(n17307) );
  NAND2_X1 U20480 ( .A1(n17307), .A2(n17306), .ZN(n17308) );
  OAI211_X1 U20481 ( .C1(n17310), .C2(n17414), .A(n17309), .B(n17308), .ZN(
        P3_U2711) );
  AOI22_X1 U20482 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17349), .ZN(n17316) );
  AOI211_X1 U20483 ( .C1(n17484), .C2(n17312), .A(n17384), .B(n17311), .ZN(
        n17313) );
  AOI21_X1 U20484 ( .B1(n17314), .B2(n17419), .A(n17313), .ZN(n17315) );
  NAND2_X1 U20485 ( .A1(n17316), .A2(n17315), .ZN(P3_U2712) );
  INV_X1 U20486 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17476) );
  INV_X1 U20487 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17474) );
  NAND2_X1 U20488 ( .A1(n18268), .A2(n9698), .ZN(n17343) );
  NAND2_X1 U20489 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17332), .ZN(n17328) );
  OR2_X1 U20490 ( .A1(n17480), .A2(n17328), .ZN(n17321) );
  AOI22_X1 U20491 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17349), .B1(n17419), .B2(
        n17317), .ZN(n17320) );
  NAND2_X1 U20492 ( .A1(n17412), .A2(n17328), .ZN(n17327) );
  OAI21_X1 U20493 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17421), .A(n17327), .ZN(
        n17318) );
  AOI22_X1 U20494 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17350), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17318), .ZN(n17319) );
  OAI211_X1 U20495 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17321), .A(n17320), .B(
        n17319), .ZN(P3_U2713) );
  INV_X1 U20496 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n17323) );
  OAI22_X1 U20497 ( .A1(n17324), .A2(n17414), .B1(n17323), .B2(n17322), .ZN(
        n17325) );
  AOI21_X1 U20498 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17350), .A(n17325), .ZN(
        n17326) );
  OAI221_X1 U20499 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17328), .C1(n17480), 
        .C2(n17327), .A(n17326), .ZN(P3_U2714) );
  AOI22_X1 U20500 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17349), .ZN(n17330) );
  OAI211_X1 U20501 ( .C1(n17332), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17412), .B(
        n17328), .ZN(n17329) );
  OAI211_X1 U20502 ( .C1(n17331), .C2(n17414), .A(n17330), .B(n17329), .ZN(
        P3_U2715) );
  AOI22_X1 U20503 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17349), .ZN(n17335) );
  NOR2_X1 U20504 ( .A1(n17474), .A2(n17345), .ZN(n17342) );
  INV_X1 U20505 ( .A(n17332), .ZN(n17333) );
  OAI211_X1 U20506 ( .C1(n17342), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17412), .B(
        n17333), .ZN(n17334) );
  OAI211_X1 U20507 ( .C1(n17336), .C2(n17414), .A(n17335), .B(n17334), .ZN(
        P3_U2716) );
  AOI21_X1 U20508 ( .B1(P3_EAX_REG_18__SCAN_IN), .B2(n17412), .A(n17337), .ZN(
        n17341) );
  AOI22_X1 U20509 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17349), .B1(n17419), .B2(
        n17338), .ZN(n17340) );
  NAND2_X1 U20510 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17350), .ZN(n17339) );
  OAI211_X1 U20511 ( .C1(n17342), .C2(n17341), .A(n17340), .B(n17339), .ZN(
        P3_U2717) );
  OAI21_X1 U20512 ( .B1(n17384), .B2(n17472), .A(n17343), .ZN(n17344) );
  AOI22_X1 U20513 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n17349), .B1(n17345), .B2(
        n17344), .ZN(n17348) );
  AOI22_X1 U20514 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17350), .B1(n17419), .B2(
        n17346), .ZN(n17347) );
  NAND2_X1 U20515 ( .A1(n17348), .A2(n17347), .ZN(P3_U2718) );
  AOI22_X1 U20516 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17350), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17349), .ZN(n17353) );
  AOI211_X1 U20517 ( .C1(n17470), .C2(n17356), .A(n17384), .B(n9698), .ZN(
        n17351) );
  INV_X1 U20518 ( .A(n17351), .ZN(n17352) );
  OAI211_X1 U20519 ( .C1(n17354), .C2(n17414), .A(n17353), .B(n17352), .ZN(
        P3_U2719) );
  AOI22_X1 U20520 ( .A1(n17419), .A2(n17355), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n17420), .ZN(n17359) );
  OAI211_X1 U20521 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17357), .A(n17412), .B(
        n17356), .ZN(n17358) );
  NAND2_X1 U20522 ( .A1(n17359), .A2(n17358), .ZN(P3_U2720) );
  NOR2_X1 U20523 ( .A1(n17365), .A2(n17360), .ZN(n17367) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17420), .B1(n17367), .B2(
        n17529), .ZN(n17362) );
  NAND3_X1 U20525 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17412), .A3(n17360), 
        .ZN(n17361) );
  OAI211_X1 U20526 ( .C1(n17363), .C2(n17414), .A(n17362), .B(n17361), .ZN(
        P3_U2721) );
  INV_X1 U20527 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17369) );
  NOR2_X1 U20528 ( .A1(n17365), .A2(n9983), .ZN(n17396) );
  NAND2_X1 U20529 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17396), .ZN(n17383) );
  NAND3_X1 U20530 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(n17388), .ZN(n17370) );
  NOR2_X1 U20531 ( .A1(n17525), .A2(n17370), .ZN(n17374) );
  AOI21_X1 U20532 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17412), .A(n17374), .ZN(
        n17368) );
  OAI222_X1 U20533 ( .A1(n17417), .A2(n17369), .B1(n17368), .B2(n17367), .C1(
        n17414), .C2(n17366), .ZN(P3_U2722) );
  OAI21_X1 U20534 ( .B1(n17525), .B2(n17384), .A(n17370), .ZN(n17371) );
  INV_X1 U20535 ( .A(n17371), .ZN(n17373) );
  OAI222_X1 U20536 ( .A1(n17417), .A2(n17375), .B1(n17374), .B2(n17373), .C1(
        n17414), .C2(n17372), .ZN(P3_U2723) );
  NAND2_X1 U20537 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17388), .ZN(n17378) );
  INV_X1 U20538 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17521) );
  NAND2_X1 U20539 ( .A1(n17412), .A2(n17378), .ZN(n17381) );
  AOI22_X1 U20540 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17420), .B1(n17419), .B2(
        n17376), .ZN(n17377) );
  OAI221_X1 U20541 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17378), .C1(n17521), 
        .C2(n17381), .A(n17377), .ZN(P3_U2724) );
  INV_X1 U20542 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17382) );
  NOR2_X1 U20543 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17388), .ZN(n17380) );
  OAI222_X1 U20544 ( .A1(n17417), .A2(n17382), .B1(n17381), .B2(n17380), .C1(
        n17414), .C2(n17379), .ZN(P3_U2725) );
  INV_X1 U20545 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17389) );
  OAI21_X1 U20546 ( .B1(n17517), .B2(n17384), .A(n17383), .ZN(n17385) );
  INV_X1 U20547 ( .A(n17385), .ZN(n17387) );
  OAI222_X1 U20548 ( .A1(n17417), .A2(n17389), .B1(n17388), .B2(n17387), .C1(
        n17414), .C2(n17386), .ZN(P3_U2726) );
  AOI22_X1 U20549 ( .A1(n17419), .A2(n17390), .B1(n17396), .B2(n17515), .ZN(
        n17392) );
  NAND3_X1 U20550 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17412), .A3(n9983), .ZN(
        n17391) );
  OAI211_X1 U20551 ( .C1(n17417), .C2(n17393), .A(n17392), .B(n17391), .ZN(
        P3_U2727) );
  INV_X1 U20552 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18265) );
  INV_X1 U20553 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17511) );
  INV_X1 U20554 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17507) );
  NOR3_X1 U20555 ( .A1(n9986), .A2(n17500), .A3(n17421), .ZN(n17411) );
  NAND2_X1 U20556 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17416), .ZN(n17404) );
  NOR2_X1 U20557 ( .A1(n17507), .A2(n17404), .ZN(n17407) );
  NAND2_X1 U20558 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17407), .ZN(n17397) );
  NOR2_X1 U20559 ( .A1(n17511), .A2(n17397), .ZN(n17400) );
  AOI21_X1 U20560 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17412), .A(n17400), .ZN(
        n17395) );
  OAI222_X1 U20561 ( .A1(n17417), .A2(n18265), .B1(n17396), .B2(n17395), .C1(
        n17414), .C2(n17394), .ZN(P3_U2728) );
  INV_X1 U20562 ( .A(n17397), .ZN(n17403) );
  AOI21_X1 U20563 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17412), .A(n17403), .ZN(
        n17399) );
  OAI222_X1 U20564 ( .A1(n17417), .A2(n18261), .B1(n17400), .B2(n17399), .C1(
        n17414), .C2(n17398), .ZN(P3_U2729) );
  INV_X1 U20565 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18256) );
  AOI21_X1 U20566 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17412), .A(n17407), .ZN(
        n17402) );
  OAI222_X1 U20567 ( .A1(n18256), .A2(n17417), .B1(n17403), .B2(n17402), .C1(
        n17414), .C2(n17401), .ZN(P3_U2730) );
  INV_X1 U20568 ( .A(n17404), .ZN(n17410) );
  AOI21_X1 U20569 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17412), .A(n17410), .ZN(
        n17406) );
  OAI222_X1 U20570 ( .A1(n18252), .A2(n17417), .B1(n17407), .B2(n17406), .C1(
        n17414), .C2(n17405), .ZN(P3_U2731) );
  INV_X1 U20571 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18248) );
  AOI21_X1 U20572 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17412), .A(n17416), .ZN(
        n17409) );
  OAI222_X1 U20573 ( .A1(n18248), .A2(n17417), .B1(n17410), .B2(n17409), .C1(
        n17414), .C2(n17408), .ZN(P3_U2732) );
  INV_X1 U20574 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18243) );
  AOI21_X1 U20575 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17412), .A(n17411), .ZN(
        n17415) );
  OAI222_X1 U20576 ( .A1(n18243), .A2(n17417), .B1(n17416), .B2(n17415), .C1(
        n17414), .C2(n17413), .ZN(P3_U2733) );
  AOI22_X1 U20577 ( .A1(n17420), .A2(BUF2_REG_1__SCAN_IN), .B1(n17419), .B2(
        n17418), .ZN(n17426) );
  NOR2_X1 U20578 ( .A1(n17500), .A2(n17421), .ZN(n17424) );
  NOR2_X1 U20579 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17421), .ZN(n17423) );
  OAI22_X1 U20580 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17424), .B1(n17423), .B2(
        n17422), .ZN(n17425) );
  NAND2_X1 U20581 ( .A1(n17426), .A2(n17425), .ZN(P3_U2734) );
  NOR2_X1 U20582 ( .A1(n18844), .A2(n18742), .ZN(n18881) );
  AND2_X1 U20583 ( .A1(n17443), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20584 ( .A1(n17446), .A2(n17428), .ZN(n17445) );
  AOI22_X1 U20585 ( .A1(n18881), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17462), .ZN(n17429) );
  OAI21_X1 U20586 ( .B1(n17498), .B2(n17445), .A(n17429), .ZN(P3_U2737) );
  INV_X1 U20587 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U20588 ( .A1(n18881), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17430) );
  OAI21_X1 U20589 ( .B1(n17496), .B2(n17445), .A(n17430), .ZN(P3_U2738) );
  INV_X1 U20590 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U20591 ( .A1(n18881), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17431) );
  OAI21_X1 U20592 ( .B1(n17494), .B2(n17445), .A(n17431), .ZN(P3_U2739) );
  AOI22_X1 U20593 ( .A1(n18881), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17432) );
  OAI21_X1 U20594 ( .B1(n17492), .B2(n17445), .A(n17432), .ZN(P3_U2740) );
  INV_X1 U20595 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17490) );
  AOI22_X1 U20596 ( .A1(n18881), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17433) );
  OAI21_X1 U20597 ( .B1(n17490), .B2(n17445), .A(n17433), .ZN(P3_U2741) );
  AOI22_X1 U20598 ( .A1(n18881), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17434) );
  OAI21_X1 U20599 ( .B1(n17488), .B2(n17445), .A(n17434), .ZN(P3_U2742) );
  AOI22_X1 U20600 ( .A1(n18881), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20601 ( .B1(n17486), .B2(n17445), .A(n17435), .ZN(P3_U2743) );
  CLKBUF_X1 U20602 ( .A(n18881), .Z(n17463) );
  AOI22_X1 U20603 ( .A1(n17463), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17436) );
  OAI21_X1 U20604 ( .B1(n17484), .B2(n17445), .A(n17436), .ZN(P3_U2744) );
  AOI22_X1 U20605 ( .A1(n17463), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17437) );
  OAI21_X1 U20606 ( .B1(n17482), .B2(n17445), .A(n17437), .ZN(P3_U2745) );
  AOI22_X1 U20607 ( .A1(n17463), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17438) );
  OAI21_X1 U20608 ( .B1(n17480), .B2(n17445), .A(n17438), .ZN(P3_U2746) );
  AOI22_X1 U20609 ( .A1(n17463), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17439) );
  OAI21_X1 U20610 ( .B1(n17478), .B2(n17445), .A(n17439), .ZN(P3_U2747) );
  AOI22_X1 U20611 ( .A1(n17463), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17440) );
  OAI21_X1 U20612 ( .B1(n17476), .B2(n17445), .A(n17440), .ZN(P3_U2748) );
  AOI22_X1 U20613 ( .A1(n17463), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17441) );
  OAI21_X1 U20614 ( .B1(n17474), .B2(n17445), .A(n17441), .ZN(P3_U2749) );
  AOI22_X1 U20615 ( .A1(n17463), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17442) );
  OAI21_X1 U20616 ( .B1(n17472), .B2(n17445), .A(n17442), .ZN(P3_U2750) );
  AOI22_X1 U20617 ( .A1(n17463), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17443), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17444) );
  OAI21_X1 U20618 ( .B1(n17470), .B2(n17445), .A(n17444), .ZN(P3_U2751) );
  AOI22_X1 U20619 ( .A1(n17463), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20620 ( .B1(n9992), .B2(n17465), .A(n17447), .ZN(P3_U2752) );
  AOI22_X1 U20621 ( .A1(n17463), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17448) );
  OAI21_X1 U20622 ( .B1(n17529), .B2(n17465), .A(n17448), .ZN(P3_U2753) );
  AOI22_X1 U20623 ( .A1(n17463), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20624 ( .B1(n17527), .B2(n17465), .A(n17449), .ZN(P3_U2754) );
  AOI22_X1 U20625 ( .A1(n17463), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17450) );
  OAI21_X1 U20626 ( .B1(n17525), .B2(n17465), .A(n17450), .ZN(P3_U2755) );
  AOI22_X1 U20627 ( .A1(n17463), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17451) );
  OAI21_X1 U20628 ( .B1(n17521), .B2(n17465), .A(n17451), .ZN(P3_U2756) );
  INV_X1 U20629 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U20630 ( .A1(n17463), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U20631 ( .B1(n17519), .B2(n17465), .A(n17452), .ZN(P3_U2757) );
  AOI22_X1 U20632 ( .A1(n17463), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17453) );
  OAI21_X1 U20633 ( .B1(n17517), .B2(n17465), .A(n17453), .ZN(P3_U2758) );
  AOI22_X1 U20634 ( .A1(n17463), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17454) );
  OAI21_X1 U20635 ( .B1(n17515), .B2(n17465), .A(n17454), .ZN(P3_U2759) );
  INV_X1 U20636 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U20637 ( .A1(n17463), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17455) );
  OAI21_X1 U20638 ( .B1(n17513), .B2(n17465), .A(n17455), .ZN(P3_U2760) );
  AOI22_X1 U20639 ( .A1(n17463), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17456) );
  OAI21_X1 U20640 ( .B1(n17511), .B2(n17465), .A(n17456), .ZN(P3_U2761) );
  INV_X1 U20641 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U20642 ( .A1(n17463), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17457) );
  OAI21_X1 U20643 ( .B1(n17509), .B2(n17465), .A(n17457), .ZN(P3_U2762) );
  AOI22_X1 U20644 ( .A1(n17463), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17458) );
  OAI21_X1 U20645 ( .B1(n17507), .B2(n17465), .A(n17458), .ZN(P3_U2763) );
  INV_X1 U20646 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17505) );
  AOI22_X1 U20647 ( .A1(n17463), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20648 ( .B1(n17505), .B2(n17465), .A(n17459), .ZN(P3_U2764) );
  INV_X1 U20649 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17503) );
  AOI22_X1 U20650 ( .A1(n17463), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17460) );
  OAI21_X1 U20651 ( .B1(n17503), .B2(n17465), .A(n17460), .ZN(P3_U2765) );
  AOI22_X1 U20652 ( .A1(n17463), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17461) );
  OAI21_X1 U20653 ( .B1(n9986), .B2(n17465), .A(n17461), .ZN(P3_U2766) );
  AOI22_X1 U20654 ( .A1(n17463), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17462), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17464) );
  OAI21_X1 U20655 ( .B1(n17500), .B2(n17465), .A(n17464), .ZN(P3_U2767) );
  NAND2_X1 U20656 ( .A1(n18884), .A2(n17468), .ZN(n18724) );
  INV_X1 U20657 ( .A(n17466), .ZN(n17467) );
  AOI22_X1 U20658 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17531), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17522), .ZN(n17469) );
  OAI21_X1 U20659 ( .B1(n17470), .B2(n17533), .A(n17469), .ZN(P3_U2768) );
  AOI22_X1 U20660 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17531), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17522), .ZN(n17471) );
  OAI21_X1 U20661 ( .B1(n17472), .B2(n17533), .A(n17471), .ZN(P3_U2769) );
  AOI22_X1 U20662 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17531), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17522), .ZN(n17473) );
  OAI21_X1 U20663 ( .B1(n17474), .B2(n17533), .A(n17473), .ZN(P3_U2770) );
  AOI22_X1 U20664 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17523), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17522), .ZN(n17475) );
  OAI21_X1 U20665 ( .B1(n17476), .B2(n17533), .A(n17475), .ZN(P3_U2771) );
  AOI22_X1 U20666 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17523), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17522), .ZN(n17477) );
  OAI21_X1 U20667 ( .B1(n17478), .B2(n17533), .A(n17477), .ZN(P3_U2772) );
  AOI22_X1 U20668 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17523), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17522), .ZN(n17479) );
  OAI21_X1 U20669 ( .B1(n17480), .B2(n17533), .A(n17479), .ZN(P3_U2773) );
  AOI22_X1 U20670 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17523), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17522), .ZN(n17481) );
  OAI21_X1 U20671 ( .B1(n17482), .B2(n17533), .A(n17481), .ZN(P3_U2774) );
  AOI22_X1 U20672 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17523), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17522), .ZN(n17483) );
  OAI21_X1 U20673 ( .B1(n17484), .B2(n17533), .A(n17483), .ZN(P3_U2775) );
  AOI22_X1 U20674 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17523), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17522), .ZN(n17485) );
  OAI21_X1 U20675 ( .B1(n17486), .B2(n17533), .A(n17485), .ZN(P3_U2776) );
  AOI22_X1 U20676 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17523), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17522), .ZN(n17487) );
  OAI21_X1 U20677 ( .B1(n17488), .B2(n17533), .A(n17487), .ZN(P3_U2777) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17523), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17522), .ZN(n17489) );
  OAI21_X1 U20679 ( .B1(n17490), .B2(n17533), .A(n17489), .ZN(P3_U2778) );
  AOI22_X1 U20680 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17523), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17522), .ZN(n17491) );
  OAI21_X1 U20681 ( .B1(n17492), .B2(n17533), .A(n17491), .ZN(P3_U2779) );
  AOI22_X1 U20682 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17531), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17522), .ZN(n17493) );
  OAI21_X1 U20683 ( .B1(n17494), .B2(n17533), .A(n17493), .ZN(P3_U2780) );
  AOI22_X1 U20684 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17531), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17522), .ZN(n17495) );
  OAI21_X1 U20685 ( .B1(n17496), .B2(n17533), .A(n17495), .ZN(P3_U2781) );
  AOI22_X1 U20686 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17531), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17522), .ZN(n17497) );
  OAI21_X1 U20687 ( .B1(n17498), .B2(n17533), .A(n17497), .ZN(P3_U2782) );
  AOI22_X1 U20688 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17522), .ZN(n17499) );
  OAI21_X1 U20689 ( .B1(n17500), .B2(n17533), .A(n17499), .ZN(P3_U2783) );
  AOI22_X1 U20690 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17522), .ZN(n17501) );
  OAI21_X1 U20691 ( .B1(n9986), .B2(n17533), .A(n17501), .ZN(P3_U2784) );
  AOI22_X1 U20692 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17522), .ZN(n17502) );
  OAI21_X1 U20693 ( .B1(n17503), .B2(n17533), .A(n17502), .ZN(P3_U2785) );
  AOI22_X1 U20694 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17522), .ZN(n17504) );
  OAI21_X1 U20695 ( .B1(n17505), .B2(n17533), .A(n17504), .ZN(P3_U2786) );
  AOI22_X1 U20696 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17530), .ZN(n17506) );
  OAI21_X1 U20697 ( .B1(n17507), .B2(n17533), .A(n17506), .ZN(P3_U2787) );
  AOI22_X1 U20698 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17530), .ZN(n17508) );
  OAI21_X1 U20699 ( .B1(n17509), .B2(n17533), .A(n17508), .ZN(P3_U2788) );
  AOI22_X1 U20700 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17530), .ZN(n17510) );
  OAI21_X1 U20701 ( .B1(n17511), .B2(n17533), .A(n17510), .ZN(P3_U2789) );
  AOI22_X1 U20702 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17530), .ZN(n17512) );
  OAI21_X1 U20703 ( .B1(n17513), .B2(n17533), .A(n17512), .ZN(P3_U2790) );
  AOI22_X1 U20704 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17530), .ZN(n17514) );
  OAI21_X1 U20705 ( .B1(n17515), .B2(n17533), .A(n17514), .ZN(P3_U2791) );
  AOI22_X1 U20706 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17530), .ZN(n17516) );
  OAI21_X1 U20707 ( .B1(n17517), .B2(n17533), .A(n17516), .ZN(P3_U2792) );
  AOI22_X1 U20708 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17523), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17522), .ZN(n17518) );
  OAI21_X1 U20709 ( .B1(n17519), .B2(n17533), .A(n17518), .ZN(P3_U2793) );
  AOI22_X1 U20710 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17530), .ZN(n17520) );
  OAI21_X1 U20711 ( .B1(n17521), .B2(n17533), .A(n17520), .ZN(P3_U2794) );
  AOI22_X1 U20712 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17523), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17522), .ZN(n17524) );
  OAI21_X1 U20713 ( .B1(n17525), .B2(n17533), .A(n17524), .ZN(P3_U2795) );
  AOI22_X1 U20714 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17530), .ZN(n17526) );
  OAI21_X1 U20715 ( .B1(n17527), .B2(n17533), .A(n17526), .ZN(P3_U2796) );
  AOI22_X1 U20716 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17530), .ZN(n17528) );
  OAI21_X1 U20717 ( .B1(n17529), .B2(n17533), .A(n17528), .ZN(P3_U2797) );
  AOI22_X1 U20718 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17531), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17530), .ZN(n17532) );
  OAI21_X1 U20719 ( .B1(n9992), .B2(n17533), .A(n17532), .ZN(P3_U2798) );
  NAND3_X1 U20720 ( .A1(n17534), .A2(n17710), .A3(n10064), .ZN(n17540) );
  AND3_X1 U20721 ( .A1(n17710), .A2(n17535), .A3(n17536), .ZN(n17557) );
  OAI21_X1 U20722 ( .B1(n17536), .B2(n17862), .A(n17900), .ZN(n17537) );
  AOI21_X1 U20723 ( .B1(n17697), .B2(n17538), .A(n17537), .ZN(n17565) );
  OAI21_X1 U20724 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17682), .A(
        n17565), .ZN(n17558) );
  OAI21_X1 U20725 ( .B1(n17557), .B2(n17558), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17539) );
  OAI211_X1 U20726 ( .C1(n17738), .C2(n17541), .A(n17540), .B(n17539), .ZN(
        n17542) );
  AOI211_X1 U20727 ( .C1(n17702), .C2(n17544), .A(n17543), .B(n17542), .ZN(
        n17551) );
  NAND2_X1 U20728 ( .A1(n17744), .A2(n17904), .ZN(n17650) );
  AOI22_X1 U20729 ( .A1(n17815), .A2(n17912), .B1(n17892), .B2(n17545), .ZN(
        n17571) );
  NAND2_X1 U20730 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17571), .ZN(
        n17559) );
  NAND3_X1 U20731 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17650), .A3(
        n17559), .ZN(n17550) );
  OAI211_X1 U20732 ( .C1(n17548), .C2(n17547), .A(n17814), .B(n17546), .ZN(
        n17549) );
  NAND3_X1 U20733 ( .A1(n17551), .A2(n17550), .A3(n17549), .ZN(P3_U2802) );
  NOR2_X1 U20734 ( .A1(n17553), .A2(n17552), .ZN(n17554) );
  XOR2_X1 U20735 ( .A(n17554), .B(n17813), .Z(n17918) );
  OAI22_X1 U20736 ( .A1(n18108), .A2(n18813), .B1(n17738), .B2(n17555), .ZN(
        n17556) );
  AOI211_X1 U20737 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17558), .A(
        n17557), .B(n17556), .ZN(n17562) );
  OAI21_X1 U20738 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17560), .A(
        n17559), .ZN(n17561) );
  OAI211_X1 U20739 ( .C1(n17918), .C2(n17789), .A(n17562), .B(n17561), .ZN(
        P3_U2803) );
  AOI21_X1 U20740 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17564), .A(
        n17563), .ZN(n17925) );
  NOR2_X1 U20741 ( .A1(n18108), .A2(n18811), .ZN(n17923) );
  AOI221_X1 U20742 ( .B1(n18519), .B2(n17567), .C1(n17566), .C2(n17567), .A(
        n17565), .ZN(n17576) );
  INV_X1 U20743 ( .A(n17568), .ZN(n17569) );
  AOI21_X1 U20744 ( .B1(n17738), .B2(n17682), .A(n17569), .ZN(n17575) );
  NOR2_X1 U20745 ( .A1(n17570), .A2(n17619), .ZN(n17573) );
  INV_X1 U20746 ( .A(n17571), .ZN(n17572) );
  MUX2_X1 U20747 ( .A(n17573), .B(n17572), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17574) );
  NOR4_X1 U20748 ( .A1(n17923), .A2(n17576), .A3(n17575), .A4(n17574), .ZN(
        n17577) );
  OAI21_X1 U20749 ( .B1(n17925), .B2(n17789), .A(n17577), .ZN(P3_U2804) );
  INV_X1 U20750 ( .A(n18035), .ZN(n17579) );
  OAI22_X1 U20751 ( .A1(n17580), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n17579), .B2(n17578), .ZN(n17939) );
  NAND2_X1 U20752 ( .A1(n17582), .A2(n17710), .ZN(n17599) );
  AOI221_X1 U20753 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C1(n17598), .C2(n17585), .A(
        n17599), .ZN(n17587) );
  OAI22_X1 U20754 ( .A1(n18519), .A2(n17582), .B1(n18742), .B2(n17581), .ZN(
        n17583) );
  OR2_X1 U20755 ( .A1(n17583), .A2(n17886), .ZN(n17610) );
  AOI21_X1 U20756 ( .B1(n17624), .B2(n17584), .A(n17610), .ZN(n17597) );
  OAI22_X1 U20757 ( .A1(n17597), .A2(n17585), .B1(n18108), .B2(n18808), .ZN(
        n17586) );
  AOI211_X1 U20758 ( .C1(n17588), .C2(n17756), .A(n17587), .B(n17586), .ZN(
        n17594) );
  NAND2_X1 U20759 ( .A1(n17951), .A2(n18034), .ZN(n17945) );
  AOI221_X1 U20760 ( .B1(n17949), .B2(n17927), .C1(n17945), .C2(n17927), .A(
        n17589), .ZN(n17936) );
  AOI21_X1 U20761 ( .B1(n17591), .B2(n10010), .A(n17590), .ZN(n17592) );
  XOR2_X1 U20762 ( .A(n17592), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17935) );
  AOI22_X1 U20763 ( .A1(n17892), .A2(n17936), .B1(n17814), .B2(n17935), .ZN(
        n17593) );
  OAI211_X1 U20764 ( .C1(n17744), .C2(n17939), .A(n17594), .B(n17593), .ZN(
        P3_U2805) );
  AOI21_X1 U20765 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17596), .A(
        n17595), .ZN(n17954) );
  NAND2_X1 U20766 ( .A1(n18210), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17952) );
  OAI221_X1 U20767 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17599), .C1(
        n17598), .C2(n17597), .A(n17952), .ZN(n17603) );
  NOR2_X1 U20768 ( .A1(n17618), .A2(n17619), .ZN(n17601) );
  AOI22_X1 U20769 ( .A1(n17815), .A2(n17941), .B1(n17892), .B2(n17945), .ZN(
        n17617) );
  INV_X1 U20770 ( .A(n17617), .ZN(n17600) );
  MUX2_X1 U20771 ( .A(n17601), .B(n17600), .S(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n17602) );
  AOI211_X1 U20772 ( .C1(n17756), .C2(n17604), .A(n17603), .B(n17602), .ZN(
        n17605) );
  OAI21_X1 U20773 ( .B1(n17954), .B2(n17789), .A(n17605), .ZN(P3_U2806) );
  INV_X1 U20774 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17975) );
  OAI21_X1 U20775 ( .B1(n17677), .B2(n17606), .A(n17630), .ZN(n17607) );
  OAI211_X1 U20776 ( .C1(n17813), .C2(n17975), .A(n17607), .B(n17648), .ZN(
        n17608) );
  XOR2_X1 U20777 ( .A(n17618), .B(n17608), .Z(n17956) );
  INV_X1 U20778 ( .A(n17609), .ZN(n17611) );
  OAI221_X1 U20779 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17611), .C1(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n18548), .A(n17610), .ZN(
        n17614) );
  OAI21_X1 U20780 ( .B1(n17756), .B2(n17624), .A(n17612), .ZN(n17613) );
  OAI211_X1 U20781 ( .C1(n18805), .C2(n18108), .A(n17614), .B(n17613), .ZN(
        n17615) );
  AOI21_X1 U20782 ( .B1(n17814), .B2(n17956), .A(n17615), .ZN(n17616) );
  OAI221_X1 U20783 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17619), 
        .C1(n17618), .C2(n17617), .A(n17616), .ZN(P3_U2807) );
  OAI22_X1 U20784 ( .A1(n18035), .A2(n17744), .B1(n18034), .B2(n17904), .ZN(
        n17703) );
  AOI21_X1 U20785 ( .B1(n17967), .B2(n17650), .A(n17703), .ZN(n17643) );
  NAND2_X1 U20786 ( .A1(n17622), .A2(n17710), .ZN(n17638) );
  AOI221_X1 U20787 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17637), .C2(n17625), .A(
        n17638), .ZN(n17627) );
  NAND2_X1 U20788 ( .A1(n17697), .A2(n17620), .ZN(n17621) );
  OAI211_X1 U20789 ( .C1(n17622), .C2(n17862), .A(n17900), .B(n17621), .ZN(
        n17652) );
  AOI21_X1 U20790 ( .B1(n17624), .B2(n17623), .A(n17652), .ZN(n17636) );
  INV_X1 U20791 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18802) );
  OAI22_X1 U20792 ( .A1(n17636), .A2(n17625), .B1(n18108), .B2(n18802), .ZN(
        n17626) );
  AOI211_X1 U20793 ( .C1(n17628), .C2(n17756), .A(n17627), .B(n17626), .ZN(
        n17635) );
  AOI221_X1 U20794 ( .B1(n17631), .B2(n17630), .C1(n17967), .C2(n17630), .A(
        n17629), .ZN(n17632) );
  XOR2_X1 U20795 ( .A(n17632), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n17960) );
  AOI22_X1 U20796 ( .A1(n17960), .A2(n17814), .B1(n17633), .B2(n17975), .ZN(
        n17634) );
  OAI211_X1 U20797 ( .C1(n17643), .C2(n17975), .A(n17635), .B(n17634), .ZN(
        P3_U2808) );
  NAND2_X1 U20798 ( .A1(n17641), .A2(n17982), .ZN(n17989) );
  NOR2_X1 U20799 ( .A1(n18005), .A2(n18017), .ZN(n17976) );
  NAND2_X1 U20800 ( .A1(n17702), .A2(n17976), .ZN(n17668) );
  NAND2_X1 U20801 ( .A1(n18210), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17987) );
  OAI221_X1 U20802 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17638), .C1(
        n17637), .C2(n17636), .A(n17987), .ZN(n17645) );
  AND3_X1 U20803 ( .A1(n17813), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17639), .ZN(n17657) );
  AOI22_X1 U20804 ( .A1(n17641), .A2(n17657), .B1(n17677), .B2(n17640), .ZN(
        n17642) );
  XOR2_X1 U20805 ( .A(n17642), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n17978) );
  OAI22_X1 U20806 ( .A1(n17643), .A2(n17982), .B1(n17978), .B2(n17789), .ZN(
        n17644) );
  AOI211_X1 U20807 ( .C1(n17756), .C2(n17646), .A(n17645), .B(n17644), .ZN(
        n17647) );
  OAI21_X1 U20808 ( .B1(n17989), .B2(n17668), .A(n17647), .ZN(P3_U2809) );
  INV_X1 U20809 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17968) );
  OAI221_X1 U20810 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17675), 
        .C1(n18001), .C2(n17657), .A(n17648), .ZN(n17649) );
  XOR2_X1 U20811 ( .A(n17968), .B(n17649), .Z(n17993) );
  NAND2_X1 U20812 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17976), .ZN(
        n17990) );
  AOI21_X1 U20813 ( .B1(n17650), .B2(n17990), .A(n17703), .ZN(n17667) );
  NAND2_X1 U20814 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17968), .ZN(
        n17997) );
  OAI22_X1 U20815 ( .A1(n17667), .A2(n17968), .B1(n17668), .B2(n17997), .ZN(
        n17651) );
  AOI21_X1 U20816 ( .B1(n17814), .B2(n17993), .A(n17651), .ZN(n17656) );
  NAND2_X1 U20817 ( .A1(n18210), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17995) );
  OAI221_X1 U20818 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9758), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18548), .A(n17652), .ZN(
        n17655) );
  OAI21_X1 U20819 ( .B1(n17756), .B2(n17624), .A(n17653), .ZN(n17654) );
  NAND4_X1 U20820 ( .A1(n17656), .A2(n17995), .A3(n17655), .A4(n17654), .ZN(
        P3_U2810) );
  AOI21_X1 U20821 ( .B1(n17675), .B2(n17677), .A(n17657), .ZN(n17658) );
  XOR2_X1 U20822 ( .A(n18001), .B(n17658), .Z(n17998) );
  OAI21_X1 U20823 ( .B1(n17669), .B2(n17862), .A(n17900), .ZN(n17691) );
  AOI21_X1 U20824 ( .B1(n17697), .B2(n17659), .A(n17691), .ZN(n17670) );
  OAI22_X1 U20825 ( .A1(n17670), .A2(n17661), .B1(n17738), .B2(n17660), .ZN(
        n17665) );
  OAI211_X1 U20826 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17669), .B(n17710), .ZN(n17662) );
  OAI22_X1 U20827 ( .A1(n17663), .A2(n17662), .B1(n18108), .B2(n18796), .ZN(
        n17664) );
  AOI211_X1 U20828 ( .C1(n17814), .C2(n17998), .A(n17665), .B(n17664), .ZN(
        n17666) );
  OAI221_X1 U20829 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17668), 
        .C1(n18001), .C2(n17667), .A(n17666), .ZN(P3_U2811) );
  AOI21_X1 U20830 ( .B1(n17702), .B2(n18005), .A(n17703), .ZN(n17693) );
  NAND2_X1 U20831 ( .A1(n17669), .A2(n17710), .ZN(n17672) );
  NAND2_X1 U20832 ( .A1(n18210), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18014) );
  OAI221_X1 U20833 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17672), .C1(
        n17671), .C2(n17670), .A(n18014), .ZN(n17673) );
  AOI21_X1 U20834 ( .B1(n17756), .B2(n17674), .A(n17673), .ZN(n17679) );
  AOI21_X1 U20835 ( .B1(n17813), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17675), .ZN(n17676) );
  XOR2_X1 U20836 ( .A(n17677), .B(n17676), .Z(n18013) );
  NOR2_X1 U20837 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18005), .ZN(
        n18012) );
  AOI22_X1 U20838 ( .A1(n17814), .A2(n18013), .B1(n17702), .B2(n18012), .ZN(
        n17678) );
  OAI211_X1 U20839 ( .C1(n17693), .C2(n18017), .A(n17679), .B(n17678), .ZN(
        P3_U2812) );
  OAI21_X1 U20840 ( .B1(n17681), .B2(n18519), .A(n17680), .ZN(n17690) );
  OAI22_X1 U20841 ( .A1(n17884), .A2(n17683), .B1(n18108), .B2(n18792), .ZN(
        n17689) );
  AOI21_X1 U20842 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17685), .A(
        n17684), .ZN(n18022) );
  NOR2_X1 U20843 ( .A1(n18029), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18018) );
  INV_X1 U20844 ( .A(n18018), .ZN(n17686) );
  OAI22_X1 U20845 ( .A1(n18022), .A2(n17789), .B1(n17687), .B2(n17686), .ZN(
        n17688) );
  AOI211_X1 U20846 ( .C1(n17691), .C2(n17690), .A(n17689), .B(n17688), .ZN(
        n17692) );
  OAI21_X1 U20847 ( .B1(n17693), .B2(n18008), .A(n17692), .ZN(P3_U2813) );
  NOR2_X1 U20848 ( .A1(n10010), .A2(n17773), .ZN(n17777) );
  OAI22_X1 U20849 ( .A1(n17813), .A2(n17694), .B1(n17790), .B2(n18011), .ZN(
        n17695) );
  XOR2_X1 U20850 ( .A(n18029), .B(n17695), .Z(n18033) );
  NOR2_X1 U20851 ( .A1(n18108), .A2(n18790), .ZN(n18028) );
  OAI211_X1 U20852 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17711), .B(n17710), .ZN(n17699) );
  OAI21_X1 U20853 ( .B1(n17711), .B2(n17862), .A(n17900), .ZN(n17723) );
  AOI21_X1 U20854 ( .B1(n17697), .B2(n17696), .A(n17723), .ZN(n17712) );
  OAI22_X1 U20855 ( .A1(n10256), .A2(n17699), .B1(n17712), .B2(n17698), .ZN(
        n17700) );
  AOI211_X1 U20856 ( .C1(n17756), .C2(n17701), .A(n18028), .B(n17700), .ZN(
        n17705) );
  AOI22_X1 U20857 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17703), .B1(
        n17702), .B2(n18029), .ZN(n17704) );
  OAI211_X1 U20858 ( .C1(n18033), .C2(n17789), .A(n17705), .B(n17704), .ZN(
        P3_U2814) );
  NOR3_X1 U20859 ( .A1(n18057), .A2(n18077), .A3(n17706), .ZN(n17707) );
  NOR3_X1 U20860 ( .A1(n17813), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17791), .ZN(n17776) );
  NAND2_X1 U20861 ( .A1(n17776), .A2(n18104), .ZN(n17765) );
  AOI22_X1 U20862 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17707), .B1(
        n17750), .B2(n17747), .ZN(n17708) );
  AOI221_X1 U20863 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18081), 
        .C1(n10010), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17708), .ZN(
        n17709) );
  XOR2_X1 U20864 ( .A(n18048), .B(n17709), .Z(n18041) );
  NAND2_X1 U20865 ( .A1(n17711), .A2(n17710), .ZN(n17714) );
  NAND2_X1 U20866 ( .A1(n18210), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18046) );
  OAI221_X1 U20867 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17714), .C1(
        n17713), .C2(n17712), .A(n18046), .ZN(n17715) );
  AOI21_X1 U20868 ( .B1(n17756), .B2(n17716), .A(n17715), .ZN(n17720) );
  NOR2_X1 U20869 ( .A1(n18035), .A2(n17744), .ZN(n17718) );
  NAND2_X1 U20870 ( .A1(n17729), .A2(n18048), .ZN(n18039) );
  NOR2_X1 U20871 ( .A1(n18034), .A2(n17904), .ZN(n17717) );
  INV_X1 U20872 ( .A(n17734), .ZN(n18051) );
  NOR3_X1 U20873 ( .A1(n18090), .A2(n17747), .A3(n18051), .ZN(n17722) );
  NAND2_X1 U20874 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17722), .ZN(
        n17721) );
  NAND2_X1 U20875 ( .A1(n18048), .A2(n17721), .ZN(n18044) );
  AOI22_X1 U20876 ( .A1(n17718), .A2(n18039), .B1(n17717), .B2(n18044), .ZN(
        n17719) );
  OAI211_X1 U20877 ( .C1(n17789), .C2(n18041), .A(n17720), .B(n17719), .ZN(
        P3_U2815) );
  OAI21_X1 U20878 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17722), .A(
        n17721), .ZN(n18065) );
  NOR2_X1 U20879 ( .A1(n18519), .A2(n17753), .ZN(n17769) );
  OAI221_X1 U20880 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17724), .C1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n17769), .A(n17723), .ZN(
        n17725) );
  OAI21_X1 U20881 ( .B1(n17884), .B2(n17726), .A(n17725), .ZN(n17732) );
  NOR2_X1 U20882 ( .A1(n18051), .A2(n17790), .ZN(n17745) );
  NOR2_X1 U20883 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17727) );
  AOI22_X1 U20884 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17745), .B1(
        n17727), .B2(n17750), .ZN(n17728) );
  XOR2_X1 U20885 ( .A(n17728), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18060) );
  OAI21_X1 U20886 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17730), .A(
        n17729), .ZN(n18058) );
  OAI22_X1 U20887 ( .A1(n18060), .A2(n17789), .B1(n17744), .B2(n18058), .ZN(
        n17731) );
  AOI211_X1 U20888 ( .C1(n18210), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17732), 
        .B(n17731), .ZN(n17733) );
  OAI21_X1 U20889 ( .B1(n17904), .B2(n18065), .A(n17733), .ZN(P3_U2816) );
  NAND2_X1 U20890 ( .A1(n17734), .A2(n17747), .ZN(n18076) );
  AOI211_X1 U20891 ( .C1(n17759), .C2(n17739), .A(n17754), .B(n17753), .ZN(
        n17743) );
  NOR2_X1 U20892 ( .A1(n18108), .A2(n18784), .ZN(n17741) );
  OAI21_X1 U20893 ( .B1(n12570), .B2(n17862), .A(n18742), .ZN(n17735) );
  AOI21_X1 U20894 ( .B1(n17736), .B2(n17735), .A(n17886), .ZN(n17760) );
  OAI22_X1 U20895 ( .A1(n17760), .A2(n17739), .B1(n17738), .B2(n17737), .ZN(
        n17740) );
  AOI211_X1 U20896 ( .C1(n17743), .C2(n17742), .A(n17741), .B(n17740), .ZN(
        n17749) );
  NOR2_X1 U20897 ( .A1(n18051), .A2(n18090), .ZN(n18067) );
  NOR2_X1 U20898 ( .A1(n17773), .A2(n18051), .ZN(n18069) );
  OAI22_X1 U20899 ( .A1(n18067), .A2(n17904), .B1(n18069), .B2(n17744), .ZN(
        n17762) );
  AOI21_X1 U20900 ( .B1(n17750), .B2(n18081), .A(n17745), .ZN(n17746) );
  XOR2_X1 U20901 ( .A(n17747), .B(n17746), .Z(n18066) );
  AOI22_X1 U20902 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17762), .B1(
        n17814), .B2(n18066), .ZN(n17748) );
  OAI211_X1 U20903 ( .C1(n17802), .C2(n18076), .A(n17749), .B(n17748), .ZN(
        P3_U2817) );
  INV_X1 U20904 ( .A(n17772), .ZN(n18096) );
  NOR2_X1 U20905 ( .A1(n18096), .A2(n17790), .ZN(n17751) );
  AOI21_X1 U20906 ( .B1(n17751), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17750), .ZN(n17752) );
  XOR2_X1 U20907 ( .A(n17752), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18087) );
  NOR2_X1 U20908 ( .A1(n17802), .A2(n18077), .ZN(n17763) );
  NOR2_X1 U20909 ( .A1(n17754), .A2(n17753), .ZN(n17755) );
  AOI22_X1 U20910 ( .A1(n17757), .A2(n17756), .B1(n17755), .B2(n17759), .ZN(
        n17758) );
  NAND2_X1 U20911 ( .A1(n18210), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18085) );
  OAI211_X1 U20912 ( .C1(n17760), .C2(n17759), .A(n17758), .B(n18085), .ZN(
        n17761) );
  AOI221_X1 U20913 ( .B1(n17763), .B2(n18081), .C1(n17762), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17761), .ZN(n17764) );
  OAI21_X1 U20914 ( .B1(n18087), .B2(n17789), .A(n17764), .ZN(P3_U2818) );
  OR2_X1 U20915 ( .A1(n18096), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18101) );
  OAI21_X1 U20916 ( .B1(n17790), .B2(n18096), .A(n17765), .ZN(n17766) );
  XOR2_X1 U20917 ( .A(n17766), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18088) );
  INV_X1 U20918 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18780) );
  NOR2_X1 U20919 ( .A1(n18108), .A2(n18780), .ZN(n17771) );
  INV_X1 U20920 ( .A(n17838), .ZN(n17895) );
  NOR3_X1 U20921 ( .A1(n18519), .A2(n17820), .A3(n17807), .ZN(n17794) );
  NAND2_X1 U20922 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17794), .ZN(
        n17793) );
  NOR2_X1 U20923 ( .A1(n17780), .A2(n17793), .ZN(n17779) );
  AOI21_X1 U20924 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17895), .A(
        n17779), .ZN(n17768) );
  OAI22_X1 U20925 ( .A1(n17769), .A2(n17768), .B1(n17884), .B2(n17767), .ZN(
        n17770) );
  AOI211_X1 U20926 ( .C1(n17814), .C2(n18088), .A(n17771), .B(n17770), .ZN(
        n17775) );
  NOR2_X1 U20927 ( .A1(n17772), .A2(n17802), .ZN(n17785) );
  AOI22_X1 U20928 ( .A1(n17773), .A2(n17815), .B1(n17892), .B2(n18090), .ZN(
        n17801) );
  INV_X1 U20929 ( .A(n17801), .ZN(n17786) );
  OAI21_X1 U20930 ( .B1(n17785), .B2(n17786), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17774) );
  OAI211_X1 U20931 ( .C1(n17802), .C2(n18101), .A(n17775), .B(n17774), .ZN(
        P3_U2819) );
  AOI21_X1 U20932 ( .B1(n17777), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17776), .ZN(n17778) );
  XOR2_X1 U20933 ( .A(n17778), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n18112) );
  AOI211_X1 U20934 ( .C1(n17793), .C2(n17780), .A(n17838), .B(n17779), .ZN(
        n17782) );
  NOR2_X1 U20935 ( .A1(n18108), .A2(n18778), .ZN(n17781) );
  AOI211_X1 U20936 ( .C1(n17783), .C2(n17894), .A(n17782), .B(n17781), .ZN(
        n17788) );
  NAND2_X1 U20937 ( .A1(n18120), .A2(n18104), .ZN(n17784) );
  AOI22_X1 U20938 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17786), .B1(
        n17785), .B2(n17784), .ZN(n17787) );
  OAI211_X1 U20939 ( .C1(n18112), .C2(n17789), .A(n17788), .B(n17787), .ZN(
        P3_U2820) );
  OAI21_X1 U20940 ( .B1(n17791), .B2(n17813), .A(n17790), .ZN(n17792) );
  XOR2_X1 U20941 ( .A(n17792), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18117) );
  NOR2_X1 U20942 ( .A1(n18108), .A2(n18776), .ZN(n17799) );
  INV_X1 U20943 ( .A(n17793), .ZN(n17797) );
  AOI21_X1 U20944 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17895), .A(
        n17794), .ZN(n17796) );
  OAI22_X1 U20945 ( .A1(n17797), .A2(n17796), .B1(n17884), .B2(n17795), .ZN(
        n17798) );
  AOI211_X1 U20946 ( .C1(n17814), .C2(n18117), .A(n17799), .B(n17798), .ZN(
        n17800) );
  OAI221_X1 U20947 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17802), .C1(
        n18120), .C2(n17801), .A(n17800), .ZN(P3_U2821) );
  OAI21_X1 U20948 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17804), .A(
        n17803), .ZN(n18137) );
  AOI21_X1 U20949 ( .B1(n17820), .B2(n17805), .A(n17886), .ZN(n17806) );
  INV_X1 U20950 ( .A(n17806), .ZN(n17823) );
  NOR2_X1 U20951 ( .A1(n17820), .A2(n17821), .ZN(n17808) );
  OAI211_X1 U20952 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17808), .A(
        n18548), .B(n17807), .ZN(n17809) );
  NAND2_X1 U20953 ( .A1(n18210), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18128) );
  OAI211_X1 U20954 ( .C1(n17884), .C2(n17810), .A(n17809), .B(n18128), .ZN(
        n17811) );
  AOI21_X1 U20955 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17823), .A(
        n17811), .ZN(n17817) );
  AOI22_X1 U20956 ( .A1(n17815), .A2(n17812), .B1(n17814), .B2(n18132), .ZN(
        n17816) );
  OAI211_X1 U20957 ( .C1(n17904), .C2(n18137), .A(n17817), .B(n17816), .ZN(
        P3_U2822) );
  OAI21_X1 U20958 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17819), .A(
        n17818), .ZN(n18145) );
  NOR2_X1 U20959 ( .A1(n18519), .A2(n17820), .ZN(n17822) );
  INV_X1 U20960 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18772) );
  NOR2_X1 U20961 ( .A1(n18108), .A2(n18772), .ZN(n18142) );
  AOI221_X1 U20962 ( .B1(n17823), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17822), .C2(n17821), .A(n18142), .ZN(n17830) );
  AOI21_X1 U20963 ( .B1(n17826), .B2(n17825), .A(n17824), .ZN(n17827) );
  XOR2_X1 U20964 ( .A(n17827), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18143) );
  AOI22_X1 U20965 ( .A1(n17892), .A2(n18143), .B1(n17828), .B2(n17894), .ZN(
        n17829) );
  OAI211_X1 U20966 ( .C1(n17903), .C2(n18145), .A(n17830), .B(n17829), .ZN(
        P3_U2823) );
  OAI21_X1 U20967 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17832), .A(
        n17831), .ZN(n18153) );
  NAND2_X1 U20968 ( .A1(n18548), .A2(n17839), .ZN(n17836) );
  OAI21_X1 U20969 ( .B1(n17835), .B2(n17834), .A(n17833), .ZN(n18147) );
  OAI22_X1 U20970 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17836), .B1(
        n17903), .B2(n18147), .ZN(n17837) );
  AOI21_X1 U20971 ( .B1(n18210), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17837), .ZN(
        n17842) );
  AOI21_X1 U20972 ( .B1(n17839), .B2(n18548), .A(n17838), .ZN(n17853) );
  AOI22_X1 U20973 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17853), .B1(
        n17840), .B2(n17894), .ZN(n17841) );
  OAI211_X1 U20974 ( .C1(n17904), .C2(n18153), .A(n17842), .B(n17841), .ZN(
        P3_U2824) );
  OAI21_X1 U20975 ( .B1(n17845), .B2(n17844), .A(n17843), .ZN(n18156) );
  OAI21_X1 U20976 ( .B1(n17886), .B2(n17847), .A(n17846), .ZN(n17852) );
  OAI21_X1 U20977 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17849), .A(
        n17848), .ZN(n18161) );
  OAI22_X1 U20978 ( .A1(n17884), .A2(n17850), .B1(n17903), .B2(n18161), .ZN(
        n17851) );
  AOI21_X1 U20979 ( .B1(n17853), .B2(n17852), .A(n17851), .ZN(n17854) );
  NAND2_X1 U20980 ( .A1(n18210), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18155) );
  OAI211_X1 U20981 ( .C1(n17904), .C2(n18156), .A(n17854), .B(n18155), .ZN(
        P3_U2825) );
  OAI21_X1 U20982 ( .B1(n17857), .B2(n17856), .A(n17855), .ZN(n18174) );
  OAI21_X1 U20983 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17859), .A(
        n17858), .ZN(n18168) );
  OAI22_X1 U20984 ( .A1(n17904), .A2(n18168), .B1(n18519), .B2(n17860), .ZN(
        n17861) );
  AOI21_X1 U20985 ( .B1(n18210), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17861), .ZN(
        n17865) );
  OAI21_X1 U20986 ( .B1(n10042), .B2(n17862), .A(n17900), .ZN(n17875) );
  AOI22_X1 U20987 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17875), .B1(
        n17863), .B2(n17894), .ZN(n17864) );
  OAI211_X1 U20988 ( .C1(n17903), .C2(n18174), .A(n17865), .B(n17864), .ZN(
        P3_U2826) );
  OAI21_X1 U20989 ( .B1(n17868), .B2(n17867), .A(n17866), .ZN(n18176) );
  NOR2_X1 U20990 ( .A1(n17886), .A2(n17887), .ZN(n17874) );
  OAI21_X1 U20991 ( .B1(n17871), .B2(n17870), .A(n17869), .ZN(n18183) );
  OAI22_X1 U20992 ( .A1(n17884), .A2(n17872), .B1(n17903), .B2(n18183), .ZN(
        n17873) );
  AOI221_X1 U20993 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17875), .C1(
        n17874), .C2(n17875), .A(n17873), .ZN(n17876) );
  NAND2_X1 U20994 ( .A1(n18210), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18181) );
  OAI211_X1 U20995 ( .C1(n17904), .C2(n18176), .A(n17876), .B(n18181), .ZN(
        P3_U2827) );
  OAI21_X1 U20996 ( .B1(n17879), .B2(n17878), .A(n17877), .ZN(n18196) );
  OAI21_X1 U20997 ( .B1(n17882), .B2(n17881), .A(n17880), .ZN(n18186) );
  OAI22_X1 U20998 ( .A1(n17884), .A2(n17883), .B1(n17904), .B2(n18186), .ZN(
        n17885) );
  AOI221_X1 U20999 ( .B1(n18548), .B2(n17887), .C1(n17886), .C2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17885), .ZN(n17888) );
  NAND2_X1 U21000 ( .A1(n18210), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18200) );
  OAI211_X1 U21001 ( .C1(n17903), .C2(n18196), .A(n17888), .B(n18200), .ZN(
        P3_U2828) );
  OAI21_X1 U21002 ( .B1(n17898), .B2(n17890), .A(n17889), .ZN(n18213) );
  NAND2_X1 U21003 ( .A1(n18863), .A2(n17899), .ZN(n17891) );
  XNOR2_X1 U21004 ( .A(n17891), .B(n17890), .ZN(n18208) );
  AOI22_X1 U21005 ( .A1(n17892), .A2(n18208), .B1(n18210), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17897) );
  AOI22_X1 U21006 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17895), .B1(
        n17894), .B2(n17893), .ZN(n17896) );
  OAI211_X1 U21007 ( .C1(n17903), .C2(n18213), .A(n17897), .B(n17896), .ZN(
        P3_U2829) );
  AOI21_X1 U21008 ( .B1(n17899), .B2(n18863), .A(n17898), .ZN(n18224) );
  INV_X1 U21009 ( .A(n18224), .ZN(n18222) );
  NAND3_X1 U21010 ( .A1(n18844), .A2(n18742), .A3(n17900), .ZN(n17901) );
  AOI22_X1 U21011 ( .A1(n18210), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17901), .ZN(n17902) );
  OAI221_X1 U21012 ( .B1(n18224), .B2(n17904), .C1(n18222), .C2(n17903), .A(
        n17902), .ZN(P3_U2830) );
  NOR3_X1 U21013 ( .A1(n17961), .A2(n17967), .A3(n17975), .ZN(n17955) );
  NAND2_X1 U21014 ( .A1(n17905), .A2(n17955), .ZN(n17920) );
  NOR2_X1 U21015 ( .A1(n17921), .A2(n17920), .ZN(n17914) );
  NOR2_X1 U21016 ( .A1(n17906), .A2(n18187), .ZN(n17911) );
  INV_X1 U21017 ( .A(n18165), .ZN(n18191) );
  INV_X1 U21018 ( .A(n17929), .ZN(n17908) );
  NOR2_X1 U21019 ( .A1(n18679), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18193) );
  INV_X1 U21020 ( .A(n18193), .ZN(n18162) );
  OAI21_X1 U21021 ( .B1(n18191), .B2(n17907), .A(n18162), .ZN(n17944) );
  AOI21_X1 U21022 ( .B1(n18165), .B2(n17908), .A(n17944), .ZN(n17932) );
  OAI211_X1 U21023 ( .C1(n18191), .C2(n9777), .A(n17932), .B(n17909), .ZN(
        n17910) );
  INV_X1 U21024 ( .A(n17919), .ZN(n17913) );
  MUX2_X1 U21025 ( .A(n17914), .B(n17913), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17915) );
  AOI22_X1 U21026 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18084), .B1(
        n18215), .B2(n17915), .ZN(n17917) );
  NAND2_X1 U21027 ( .A1(n18210), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17916) );
  OAI211_X1 U21028 ( .C1(n17918), .C2(n18111), .A(n17917), .B(n17916), .ZN(
        P3_U2835) );
  AOI211_X1 U21029 ( .C1(n17921), .C2(n17920), .A(n17919), .B(n18126), .ZN(
        n17922) );
  AOI211_X1 U21030 ( .C1(n18084), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17923), .B(n17922), .ZN(n17924) );
  OAI21_X1 U21031 ( .B1(n17925), .B2(n18111), .A(n17924), .ZN(P3_U2836) );
  NOR2_X1 U21032 ( .A1(n18108), .A2(n18808), .ZN(n17934) );
  OAI21_X1 U21033 ( .B1(n18707), .B2(n17927), .A(n17926), .ZN(n17931) );
  AOI21_X1 U21034 ( .B1(n17929), .B2(n17928), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17930) );
  AOI211_X1 U21035 ( .C1(n17932), .C2(n17931), .A(n17930), .B(n18126), .ZN(
        n17933) );
  AOI211_X1 U21036 ( .C1(n18084), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17934), .B(n17933), .ZN(n17938) );
  AOI22_X1 U21037 ( .A1(n18209), .A2(n17936), .B1(n18133), .B2(n17935), .ZN(
        n17937) );
  OAI211_X1 U21038 ( .C1(n18059), .C2(n17939), .A(n17938), .B(n17937), .ZN(
        P3_U2837) );
  AOI21_X1 U21039 ( .B1(n17941), .B2(n17940), .A(n18084), .ZN(n17942) );
  INV_X1 U21040 ( .A(n17942), .ZN(n17943) );
  AOI211_X1 U21041 ( .C1(n18706), .C2(n17945), .A(n17944), .B(n17943), .ZN(
        n17948) );
  OAI211_X1 U21042 ( .C1(n17946), .C2(n18190), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17948), .ZN(n17947) );
  NAND2_X1 U21043 ( .A1(n18108), .A2(n17947), .ZN(n17958) );
  AOI21_X1 U21044 ( .B1(n18167), .B2(n17948), .A(n17958), .ZN(n17950) );
  OAI222_X1 U21045 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17951), 
        .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17977), .C1(n17950), 
        .C2(n17949), .ZN(n17953) );
  OAI211_X1 U21046 ( .C1(n17954), .C2(n18111), .A(n17953), .B(n17952), .ZN(
        P3_U2838) );
  AOI21_X1 U21047 ( .B1(n17955), .B2(n18205), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17959) );
  AOI22_X1 U21048 ( .A1(n18210), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18133), 
        .B2(n17956), .ZN(n17957) );
  OAI21_X1 U21049 ( .B1(n17959), .B2(n17958), .A(n17957), .ZN(P3_U2839) );
  AOI22_X1 U21050 ( .A1(n18210), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n18133), 
        .B2(n17960), .ZN(n17974) );
  NOR2_X1 U21051 ( .A1(n17961), .A2(n17967), .ZN(n17972) );
  NOR2_X1 U21052 ( .A1(n18863), .A2(n17962), .ZN(n18114) );
  INV_X1 U21053 ( .A(n18114), .ZN(n18050) );
  NOR2_X1 U21054 ( .A1(n18011), .A2(n18050), .ZN(n18024) );
  AOI21_X1 U21055 ( .B1(n17976), .B2(n18024), .A(n18679), .ZN(n17966) );
  OAI21_X1 U21056 ( .B1(n18003), .B2(n17990), .A(n18664), .ZN(n17963) );
  OAI221_X1 U21057 ( .B1(n18190), .B2(n17964), .C1(n18190), .C2(n17976), .A(
        n17963), .ZN(n17965) );
  NOR2_X1 U21058 ( .A1(n17966), .A2(n17965), .ZN(n17980) );
  NAND2_X1 U21059 ( .A1(n18187), .A2(n18092), .ZN(n18095) );
  AOI22_X1 U21060 ( .A1(n18664), .A2(n17968), .B1(n17967), .B2(n18095), .ZN(
        n17984) );
  OAI22_X1 U21061 ( .A1(n18035), .A2(n18092), .B1(n18034), .B2(n18187), .ZN(
        n17979) );
  AOI21_X1 U21062 ( .B1(n18122), .B2(n17969), .A(n17979), .ZN(n17970) );
  NAND4_X1 U21063 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17980), .A3(
        n17984), .A4(n17970), .ZN(n17971) );
  OAI211_X1 U21064 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17972), .A(
        n18215), .B(n17971), .ZN(n17973) );
  OAI211_X1 U21065 ( .C1(n18205), .C2(n17975), .A(n17974), .B(n17973), .ZN(
        P3_U2840) );
  NAND2_X1 U21066 ( .A1(n17977), .A2(n17976), .ZN(n18002) );
  INV_X1 U21067 ( .A(n17978), .ZN(n17986) );
  NAND2_X1 U21068 ( .A1(n18027), .A2(n17980), .ZN(n17991) );
  AOI21_X1 U21069 ( .B1(n17981), .B2(n18204), .A(n17991), .ZN(n17983) );
  AOI211_X1 U21070 ( .C1(n17984), .C2(n17983), .A(n18210), .B(n17982), .ZN(
        n17985) );
  AOI21_X1 U21071 ( .B1(n18133), .B2(n17986), .A(n17985), .ZN(n17988) );
  OAI211_X1 U21072 ( .C1(n17989), .C2(n18002), .A(n17988), .B(n17987), .ZN(
        P3_U2841) );
  NAND3_X1 U21073 ( .A1(n18001), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18204), 
        .ZN(n17992) );
  OAI221_X1 U21074 ( .B1(n17991), .B2(n17990), .C1(n17991), .C2(n18095), .A(
        n18108), .ZN(n18000) );
  NAND2_X1 U21075 ( .A1(n17992), .A2(n18000), .ZN(n17994) );
  AOI22_X1 U21076 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17994), .B1(
        n18133), .B2(n17993), .ZN(n17996) );
  OAI211_X1 U21077 ( .C1(n18002), .C2(n17997), .A(n17996), .B(n17995), .ZN(
        P3_U2842) );
  AOI22_X1 U21078 ( .A1(n18210), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n18133), 
        .B2(n17998), .ZN(n17999) );
  OAI221_X1 U21079 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18002), 
        .C1(n18001), .C2(n18000), .A(n17999), .ZN(P3_U2843) );
  NOR3_X1 U21080 ( .A1(n18193), .A2(n18003), .A3(n18029), .ZN(n18007) );
  AOI222_X1 U21081 ( .A1(n18707), .A2(n18005), .B1(n18707), .B2(n18004), .C1(
        n18005), .C2(n18095), .ZN(n18006) );
  OAI211_X1 U21082 ( .C1(n18191), .C2(n18007), .A(n18027), .B(n18006), .ZN(
        n18019) );
  OAI221_X1 U21083 ( .B1(n18019), .B2(n18165), .C1(n18019), .C2(n18008), .A(
        n18108), .ZN(n18016) );
  NAND2_X1 U21084 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18164) );
  OAI22_X1 U21085 ( .A1(n18188), .A2(n18190), .B1(n18164), .B2(n18185), .ZN(
        n18179) );
  NAND3_X1 U21086 ( .A1(n18009), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18179), .ZN(n18140) );
  NOR2_X1 U21087 ( .A1(n9879), .A2(n18140), .ZN(n18130) );
  NAND2_X1 U21088 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18130), .ZN(
        n18049) );
  NAND2_X1 U21089 ( .A1(n18010), .A2(n18049), .ZN(n18078) );
  NAND2_X1 U21090 ( .A1(n18215), .A2(n18078), .ZN(n18121) );
  NOR2_X1 U21091 ( .A1(n18011), .A2(n18121), .ZN(n18030) );
  AOI22_X1 U21092 ( .A1(n18133), .A2(n18013), .B1(n18012), .B2(n18030), .ZN(
        n18015) );
  OAI211_X1 U21093 ( .C1(n18017), .C2(n18016), .A(n18015), .B(n18014), .ZN(
        P3_U2844) );
  AOI22_X1 U21094 ( .A1(n18210), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18030), 
        .B2(n18018), .ZN(n18021) );
  NAND3_X1 U21095 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18108), .A3(
        n18019), .ZN(n18020) );
  OAI211_X1 U21096 ( .C1(n18022), .C2(n18111), .A(n18021), .B(n18020), .ZN(
        P3_U2845) );
  NOR2_X1 U21097 ( .A1(n18689), .A2(n18023), .ZN(n18103) );
  NOR2_X1 U21098 ( .A1(n18103), .A2(n18687), .ZN(n18113) );
  AOI21_X1 U21099 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18113), .A(
        n18024), .ZN(n18026) );
  NOR2_X1 U21100 ( .A1(n18025), .A2(n18190), .ZN(n18089) );
  AOI211_X1 U21101 ( .C1(n18037), .C2(n18102), .A(n18026), .B(n18089), .ZN(
        n18036) );
  AOI221_X1 U21102 ( .B1(n18167), .B2(n18027), .C1(n18036), .C2(n18027), .A(
        n18210), .ZN(n18031) );
  AOI221_X1 U21103 ( .B1(n18031), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), 
        .C1(n18030), .C2(n18029), .A(n18028), .ZN(n18032) );
  OAI21_X1 U21104 ( .B1(n18033), .B2(n18111), .A(n18032), .ZN(P3_U2846) );
  NOR2_X1 U21105 ( .A1(n18034), .A2(n18223), .ZN(n18045) );
  NOR2_X1 U21106 ( .A1(n18035), .A2(n18092), .ZN(n18040) );
  AOI221_X1 U21107 ( .B1(n18037), .B2(n18048), .C1(n18049), .C2(n18048), .A(
        n18036), .ZN(n18038) );
  AOI21_X1 U21108 ( .B1(n18040), .B2(n18039), .A(n18038), .ZN(n18042) );
  OAI22_X1 U21109 ( .A1(n18042), .A2(n18126), .B1(n18111), .B2(n18041), .ZN(
        n18043) );
  AOI21_X1 U21110 ( .B1(n18045), .B2(n18044), .A(n18043), .ZN(n18047) );
  OAI211_X1 U21111 ( .C1(n18205), .C2(n18048), .A(n18047), .B(n18046), .ZN(
        P3_U2847) );
  NOR2_X1 U21112 ( .A1(n18053), .A2(n18049), .ZN(n18056) );
  INV_X1 U21113 ( .A(n18068), .ZN(n18052) );
  AOI211_X1 U21114 ( .C1(n18122), .C2(n18053), .A(n18103), .B(n18052), .ZN(
        n18054) );
  INV_X1 U21115 ( .A(n18054), .ZN(n18055) );
  MUX2_X1 U21116 ( .A(n18056), .B(n18055), .S(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n18063) );
  OAI22_X1 U21117 ( .A1(n18057), .A2(n18205), .B1(n18108), .B2(n18787), .ZN(
        n18062) );
  OAI22_X1 U21118 ( .A1(n18060), .A2(n18111), .B1(n18059), .B2(n18058), .ZN(
        n18061) );
  AOI211_X1 U21119 ( .C1(n18215), .C2(n18063), .A(n18062), .B(n18061), .ZN(
        n18064) );
  OAI21_X1 U21120 ( .B1(n18223), .B2(n18065), .A(n18064), .ZN(P3_U2848) );
  AOI22_X1 U21121 ( .A1(n18210), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18133), 
        .B2(n18066), .ZN(n18075) );
  INV_X1 U21122 ( .A(n18067), .ZN(n18071) );
  OAI21_X1 U21123 ( .B1(n18103), .B2(n18077), .A(n18102), .ZN(n18097) );
  OAI211_X1 U21124 ( .C1(n18069), .C2(n18092), .A(n18068), .B(n18097), .ZN(
        n18070) );
  AOI21_X1 U21125 ( .B1(n18706), .B2(n18071), .A(n18070), .ZN(n18082) );
  OAI211_X1 U21126 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18072), .A(
        n18215), .B(n18082), .ZN(n18073) );
  NAND3_X1 U21127 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18108), .A3(
        n18073), .ZN(n18074) );
  OAI211_X1 U21128 ( .C1(n18121), .C2(n18076), .A(n18075), .B(n18074), .ZN(
        P3_U2849) );
  INV_X1 U21129 ( .A(n18077), .ZN(n18079) );
  NAND3_X1 U21130 ( .A1(n18079), .A2(n18078), .A3(n18081), .ZN(n18080) );
  OAI21_X1 U21131 ( .B1(n18082), .B2(n18081), .A(n18080), .ZN(n18083) );
  AOI22_X1 U21132 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18084), .B1(
        n18215), .B2(n18083), .ZN(n18086) );
  OAI211_X1 U21133 ( .C1(n18087), .C2(n18111), .A(n18086), .B(n18085), .ZN(
        P3_U2850) );
  AOI22_X1 U21134 ( .A1(n18210), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18133), 
        .B2(n18088), .ZN(n18100) );
  AOI21_X1 U21135 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18114), .A(
        n18679), .ZN(n18094) );
  AOI211_X1 U21136 ( .C1(n18090), .C2(n18706), .A(n18089), .B(n18126), .ZN(
        n18091) );
  OAI21_X1 U21137 ( .B1(n18093), .B2(n18092), .A(n18091), .ZN(n18116) );
  AOI211_X1 U21138 ( .C1(n18096), .C2(n18095), .A(n18094), .B(n18116), .ZN(
        n18106) );
  OAI211_X1 U21139 ( .C1(n18679), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18106), .B(n18097), .ZN(n18098) );
  NAND3_X1 U21140 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18108), .A3(
        n18098), .ZN(n18099) );
  OAI211_X1 U21141 ( .C1(n18121), .C2(n18101), .A(n18100), .B(n18099), .ZN(
        P3_U2851) );
  OAI21_X1 U21142 ( .B1(n18103), .B2(n18120), .A(n18102), .ZN(n18105) );
  AOI21_X1 U21143 ( .B1(n18106), .B2(n18105), .A(n18104), .ZN(n18109) );
  NOR3_X1 U21144 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18120), .A3(
        n18121), .ZN(n18107) );
  AOI221_X1 U21145 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n18210), .C1(n18109), 
        .C2(n18108), .A(n18107), .ZN(n18110) );
  OAI21_X1 U21146 ( .B1(n18112), .B2(n18111), .A(n18110), .ZN(P3_U2852) );
  NOR2_X1 U21147 ( .A1(n18114), .A2(n18113), .ZN(n18115) );
  OAI21_X1 U21148 ( .B1(n18116), .B2(n18115), .A(n18108), .ZN(n18119) );
  AOI22_X1 U21149 ( .A1(n18210), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18133), 
        .B2(n18117), .ZN(n18118) );
  OAI221_X1 U21150 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18121), .C1(
        n18120), .C2(n18119), .A(n18118), .ZN(P3_U2853) );
  NOR2_X1 U21151 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18126), .ZN(
        n18131) );
  INV_X1 U21152 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18148) );
  OAI211_X1 U21153 ( .C1(n18148), .C2(n9879), .A(n18122), .B(n18215), .ZN(
        n18139) );
  OR2_X1 U21154 ( .A1(n18193), .A2(n18123), .ZN(n18124) );
  AOI22_X1 U21155 ( .A1(n18707), .A2(n18125), .B1(n18165), .B2(n18124), .ZN(
        n18127) );
  OAI21_X1 U21156 ( .B1(n18127), .B2(n18126), .A(n18205), .ZN(n18159) );
  INV_X1 U21157 ( .A(n18159), .ZN(n18149) );
  AND2_X1 U21158 ( .A1(n18139), .A2(n18149), .ZN(n18138) );
  OAI21_X1 U21159 ( .B1(n18138), .B2(n9878), .A(n18128), .ZN(n18129) );
  AOI21_X1 U21160 ( .B1(n18131), .B2(n18130), .A(n18129), .ZN(n18136) );
  AOI22_X1 U21161 ( .A1(n17812), .A2(n18134), .B1(n18133), .B2(n18132), .ZN(
        n18135) );
  OAI211_X1 U21162 ( .C1(n18223), .C2(n18137), .A(n18136), .B(n18135), .ZN(
        P3_U2854) );
  AOI221_X1 U21163 ( .B1(n18140), .B2(n9879), .C1(n18139), .C2(n9879), .A(
        n18138), .ZN(n18141) );
  AOI211_X1 U21164 ( .C1(n18143), .C2(n18209), .A(n18142), .B(n18141), .ZN(
        n18144) );
  OAI21_X1 U21165 ( .B1(n18221), .B2(n18145), .A(n18144), .ZN(P3_U2855) );
  NAND3_X1 U21166 ( .A1(n18215), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18179), .ZN(n18169) );
  NOR3_X1 U21167 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18146), .A3(
        n18169), .ZN(n18151) );
  OAI22_X1 U21168 ( .A1(n18149), .A2(n18148), .B1(n18221), .B2(n18147), .ZN(
        n18150) );
  AOI211_X1 U21169 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n18210), .A(n18151), .B(
        n18150), .ZN(n18152) );
  OAI21_X1 U21170 ( .B1(n18223), .B2(n18153), .A(n18152), .ZN(P3_U2856) );
  INV_X1 U21171 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18154) );
  NOR3_X1 U21172 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18154), .A3(
        n18169), .ZN(n18158) );
  OAI21_X1 U21173 ( .B1(n18223), .B2(n18156), .A(n18155), .ZN(n18157) );
  AOI211_X1 U21174 ( .C1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n18159), .A(
        n18158), .B(n18157), .ZN(n18160) );
  OAI21_X1 U21175 ( .B1(n18221), .B2(n18161), .A(n18160), .ZN(P3_U2857) );
  OAI211_X1 U21176 ( .C1(n18190), .C2(n18163), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18162), .ZN(n18166) );
  OAI221_X1 U21177 ( .B1(n18166), .B2(n18165), .C1(n18166), .C2(n18164), .A(
        n18215), .ZN(n18175) );
  OAI21_X1 U21178 ( .B1(n18167), .B2(n18175), .A(n18205), .ZN(n18171) );
  OAI22_X1 U21179 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18169), .B1(
        n18168), .B2(n18223), .ZN(n18170) );
  AOI21_X1 U21180 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18171), .A(
        n18170), .ZN(n18173) );
  NAND2_X1 U21181 ( .A1(n18210), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18172) );
  OAI211_X1 U21182 ( .C1(n18174), .C2(n18221), .A(n18173), .B(n18172), .ZN(
        P3_U2858) );
  INV_X1 U21183 ( .A(n18175), .ZN(n18180) );
  OAI22_X1 U21184 ( .A1(n18177), .A2(n18205), .B1(n18223), .B2(n18176), .ZN(
        n18178) );
  AOI221_X1 U21185 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18180), .C1(
        n18179), .C2(n18180), .A(n18178), .ZN(n18182) );
  OAI211_X1 U21186 ( .C1(n18183), .C2(n18221), .A(n18182), .B(n18181), .ZN(
        P3_U2859) );
  NAND2_X1 U21187 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18201), .ZN(
        n18184) );
  OAI22_X1 U21188 ( .A1(n18187), .A2(n18186), .B1(n18185), .B2(n18184), .ZN(
        n18198) );
  NAND2_X1 U21189 ( .A1(n18707), .A2(n18188), .ZN(n18195) );
  NAND2_X1 U21190 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18189) );
  OAI22_X1 U21191 ( .A1(n18191), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n18190), .B2(n18189), .ZN(n18192) );
  OAI21_X1 U21192 ( .B1(n18193), .B2(n18192), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18194) );
  OAI211_X1 U21193 ( .C1(n18196), .C2(n18713), .A(n18195), .B(n18194), .ZN(
        n18197) );
  OAI21_X1 U21194 ( .B1(n18198), .B2(n18197), .A(n18215), .ZN(n18199) );
  OAI211_X1 U21195 ( .C1(n18205), .C2(n18201), .A(n18200), .B(n18199), .ZN(
        P3_U2860) );
  NOR2_X1 U21196 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18664), .ZN(
        n18202) );
  NOR2_X1 U21197 ( .A1(n18203), .A2(n18202), .ZN(n18206) );
  NAND2_X1 U21198 ( .A1(n18204), .A2(n18215), .ZN(n18216) );
  OAI21_X1 U21199 ( .B1(n18216), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18205), .ZN(n18214) );
  MUX2_X1 U21200 ( .A(n18206), .B(n18214), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n18207) );
  AOI21_X1 U21201 ( .B1(n18209), .B2(n18208), .A(n18207), .ZN(n18212) );
  NAND2_X1 U21202 ( .A1(n18210), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18211) );
  OAI211_X1 U21203 ( .C1(n18213), .C2(n18221), .A(n18212), .B(n18211), .ZN(
        P3_U2861) );
  INV_X1 U21204 ( .A(n18214), .ZN(n18218) );
  NAND2_X1 U21205 ( .A1(n18215), .A2(n18664), .ZN(n18217) );
  AOI22_X1 U21206 ( .A1(n18218), .A2(n18217), .B1(n18863), .B2(n18216), .ZN(
        n18219) );
  AOI21_X1 U21207 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n18210), .A(n18219), .ZN(
        n18220) );
  OAI221_X1 U21208 ( .B1(n18224), .B2(n18223), .C1(n18222), .C2(n18221), .A(
        n18220), .ZN(P3_U2862) );
  AOI211_X1 U21209 ( .C1(n18226), .C2(n18225), .A(n18727), .B(n18844), .ZN(
        n18729) );
  OAI21_X1 U21210 ( .B1(n18729), .B2(n18272), .A(n18231), .ZN(n18227) );
  OAI221_X1 U21211 ( .B1(n18469), .B2(n18879), .C1(n18469), .C2(n18231), .A(
        n18227), .ZN(P3_U2863) );
  NAND2_X1 U21212 ( .A1(n18698), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18494) );
  INV_X1 U21213 ( .A(n18494), .ZN(n18493) );
  NAND2_X1 U21214 ( .A1(n18701), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18403) );
  INV_X1 U21215 ( .A(n18403), .ZN(n18402) );
  NOR2_X1 U21216 ( .A1(n18493), .A2(n18402), .ZN(n18229) );
  OAI22_X1 U21217 ( .A1(n18230), .A2(n18701), .B1(n18229), .B2(n18228), .ZN(
        P3_U2866) );
  NOR2_X1 U21218 ( .A1(n18702), .A2(n18231), .ZN(P3_U2867) );
  INV_X1 U21219 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18232) );
  NOR2_X1 U21220 ( .A1(n18519), .A2(n18232), .ZN(n18608) );
  INV_X1 U21221 ( .A(n18608), .ZN(n18497) );
  NOR2_X1 U21222 ( .A1(n18701), .A2(n18446), .ZN(n18605) );
  NAND2_X1 U21223 ( .A1(n18605), .A2(n18469), .ZN(n18291) );
  NOR2_X1 U21224 ( .A1(n18698), .A2(n18701), .ZN(n18610) );
  INV_X1 U21225 ( .A(n18610), .ZN(n18545) );
  NAND2_X1 U21226 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18693), .ZN(
        n18448) );
  NOR2_X2 U21227 ( .A1(n18545), .A2(n18448), .ZN(n18647) );
  NAND2_X1 U21228 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18548), .ZN(n18614) );
  INV_X1 U21229 ( .A(n18614), .ZN(n18492) );
  INV_X1 U21230 ( .A(n18518), .ZN(n18577) );
  AND2_X1 U21231 ( .A1(n18577), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18607) );
  INV_X1 U21232 ( .A(n18606), .ZN(n18726) );
  NAND2_X1 U21233 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18692) );
  NOR2_X2 U21234 ( .A1(n18692), .A2(n18545), .ZN(n18658) );
  NAND2_X1 U21235 ( .A1(n18693), .A2(n18469), .ZN(n18694) );
  NOR2_X1 U21236 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18315) );
  INV_X1 U21237 ( .A(n18315), .ZN(n18316) );
  NOR2_X2 U21238 ( .A1(n18694), .A2(n18316), .ZN(n18329) );
  NOR2_X1 U21239 ( .A1(n18658), .A2(n18329), .ZN(n18292) );
  NOR2_X1 U21240 ( .A1(n18726), .A2(n18292), .ZN(n18266) );
  AOI22_X1 U21241 ( .A1(n18647), .A2(n18492), .B1(n18607), .B2(n18266), .ZN(
        n18239) );
  INV_X1 U21242 ( .A(n18291), .ZN(n18602) );
  NOR2_X1 U21243 ( .A1(n18602), .A2(n18647), .ZN(n18573) );
  INV_X1 U21244 ( .A(n18573), .ZN(n18234) );
  AOI211_X1 U21245 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18292), .B(n18518), .ZN(
        n18233) );
  AOI21_X1 U21246 ( .B1(n18548), .B2(n18234), .A(n18233), .ZN(n18269) );
  NAND2_X1 U21247 ( .A1(n18236), .A2(n18235), .ZN(n18267) );
  NOR2_X2 U21248 ( .A1(n18237), .A2(n18267), .ZN(n18611) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18269), .B1(
        n18329), .B2(n18611), .ZN(n18238) );
  OAI211_X1 U21250 ( .C1(n18497), .C2(n18291), .A(n18239), .B(n18238), .ZN(
        P3_U2868) );
  INV_X1 U21251 ( .A(n18647), .ZN(n18663) );
  NOR2_X1 U21252 ( .A1(n19283), .A2(n18519), .ZN(n18551) );
  INV_X1 U21253 ( .A(n18551), .ZN(n18620) );
  NAND2_X1 U21254 ( .A1(n18548), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18554) );
  INV_X1 U21255 ( .A(n18554), .ZN(n18616) );
  AND2_X1 U21256 ( .A1(n18577), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18615) );
  AOI22_X1 U21257 ( .A1(n18602), .A2(n18616), .B1(n18266), .B2(n18615), .ZN(
        n18241) );
  NOR2_X2 U21258 ( .A1(n18884), .A2(n18267), .ZN(n18617) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18269), .B1(
        n18329), .B2(n18617), .ZN(n18240) );
  OAI211_X1 U21260 ( .C1(n18663), .C2(n18620), .A(n18241), .B(n18240), .ZN(
        P3_U2869) );
  INV_X1 U21261 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18242) );
  NOR2_X1 U21262 ( .A1(n18242), .A2(n18519), .ZN(n18582) );
  INV_X1 U21263 ( .A(n18582), .ZN(n18626) );
  NAND2_X1 U21264 ( .A1(n18548), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18585) );
  INV_X1 U21265 ( .A(n18585), .ZN(n18622) );
  NOR2_X2 U21266 ( .A1(n18518), .A2(n18243), .ZN(n18621) );
  AOI22_X1 U21267 ( .A1(n18602), .A2(n18622), .B1(n18266), .B2(n18621), .ZN(
        n18246) );
  NOR2_X2 U21268 ( .A1(n18244), .A2(n18267), .ZN(n18623) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18269), .B1(
        n18329), .B2(n18623), .ZN(n18245) );
  OAI211_X1 U21270 ( .C1(n18663), .C2(n18626), .A(n18246), .B(n18245), .ZN(
        P3_U2870) );
  NOR2_X1 U21271 ( .A1(n18247), .A2(n18519), .ZN(n18628) );
  INV_X1 U21272 ( .A(n18628), .ZN(n18589) );
  NAND2_X1 U21273 ( .A1(n18548), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18632) );
  INV_X1 U21274 ( .A(n18632), .ZN(n18586) );
  NOR2_X2 U21275 ( .A1(n18518), .A2(n18248), .ZN(n18627) );
  AOI22_X1 U21276 ( .A1(n18602), .A2(n18586), .B1(n18266), .B2(n18627), .ZN(
        n18251) );
  NOR2_X2 U21277 ( .A1(n18249), .A2(n18267), .ZN(n18629) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18269), .B1(
        n18329), .B2(n18629), .ZN(n18250) );
  OAI211_X1 U21279 ( .C1(n18663), .C2(n18589), .A(n18251), .B(n18250), .ZN(
        P3_U2871) );
  NAND2_X1 U21280 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18548), .ZN(n18533) );
  NAND2_X1 U21281 ( .A1(n18548), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18638) );
  INV_X1 U21282 ( .A(n18638), .ZN(n18530) );
  NOR2_X2 U21283 ( .A1(n18518), .A2(n18252), .ZN(n18633) );
  AOI22_X1 U21284 ( .A1(n18602), .A2(n18530), .B1(n18266), .B2(n18633), .ZN(
        n18255) );
  NOR2_X2 U21285 ( .A1(n18253), .A2(n18267), .ZN(n18635) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18269), .B1(
        n18329), .B2(n18635), .ZN(n18254) );
  OAI211_X1 U21287 ( .C1(n18663), .C2(n18533), .A(n18255), .B(n18254), .ZN(
        P3_U2872) );
  NOR2_X1 U21288 ( .A1(n19298), .A2(n18519), .ZN(n18592) );
  INV_X1 U21289 ( .A(n18592), .ZN(n18644) );
  NAND2_X1 U21290 ( .A1(n18548), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18595) );
  INV_X1 U21291 ( .A(n18595), .ZN(n18640) );
  NOR2_X2 U21292 ( .A1(n18518), .A2(n18256), .ZN(n18639) );
  AOI22_X1 U21293 ( .A1(n18602), .A2(n18640), .B1(n18266), .B2(n18639), .ZN(
        n18259) );
  NOR2_X2 U21294 ( .A1(n18257), .A2(n18267), .ZN(n18641) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18269), .B1(
        n18329), .B2(n18641), .ZN(n18258) );
  OAI211_X1 U21296 ( .C1(n18663), .C2(n18644), .A(n18259), .B(n18258), .ZN(
        P3_U2873) );
  NOR2_X1 U21297 ( .A1(n18260), .A2(n18519), .ZN(n18564) );
  INV_X1 U21298 ( .A(n18564), .ZN(n18652) );
  NAND2_X1 U21299 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18548), .ZN(n18567) );
  INV_X1 U21300 ( .A(n18567), .ZN(n18646) );
  NOR2_X2 U21301 ( .A1(n18261), .A2(n18518), .ZN(n18645) );
  AOI22_X1 U21302 ( .A1(n18602), .A2(n18646), .B1(n18266), .B2(n18645), .ZN(
        n18264) );
  NOR2_X2 U21303 ( .A1(n18262), .A2(n18267), .ZN(n18648) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18269), .B1(
        n18329), .B2(n18648), .ZN(n18263) );
  OAI211_X1 U21305 ( .C1(n18663), .C2(n18652), .A(n18264), .B(n18263), .ZN(
        P3_U2874) );
  NAND2_X1 U21306 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18548), .ZN(n18662) );
  NAND2_X1 U21307 ( .A1(n18548), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18517) );
  INV_X1 U21308 ( .A(n18517), .ZN(n18656) );
  NOR2_X2 U21309 ( .A1(n18265), .A2(n18518), .ZN(n18654) );
  AOI22_X1 U21310 ( .A1(n18647), .A2(n18656), .B1(n18266), .B2(n18654), .ZN(
        n18271) );
  NOR2_X2 U21311 ( .A1(n18268), .A2(n18267), .ZN(n18657) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18269), .B1(
        n18329), .B2(n18657), .ZN(n18270) );
  OAI211_X1 U21313 ( .C1(n18291), .C2(n18662), .A(n18271), .B(n18270), .ZN(
        P3_U2875) );
  INV_X1 U21314 ( .A(n18658), .ZN(n18312) );
  NAND2_X1 U21315 ( .A1(n18693), .A2(n18606), .ZN(n18544) );
  NOR2_X1 U21316 ( .A1(n18316), .A2(n18544), .ZN(n18287) );
  AOI22_X1 U21317 ( .A1(n18602), .A2(n18492), .B1(n18607), .B2(n18287), .ZN(
        n18274) );
  NOR3_X1 U21318 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18272), .A3(
        n18518), .ZN(n18546) );
  AOI22_X1 U21319 ( .A1(n18548), .A2(n18605), .B1(n18315), .B2(n18546), .ZN(
        n18288) );
  NOR2_X2 U21320 ( .A1(n18448), .A2(n18316), .ZN(n18355) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18288), .B1(
        n18611), .B2(n18355), .ZN(n18273) );
  OAI211_X1 U21322 ( .C1(n18497), .C2(n18312), .A(n18274), .B(n18273), .ZN(
        P3_U2876) );
  AOI22_X1 U21323 ( .A1(n18602), .A2(n18551), .B1(n18615), .B2(n18287), .ZN(
        n18276) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18288), .B1(
        n18617), .B2(n18355), .ZN(n18275) );
  OAI211_X1 U21325 ( .C1(n18312), .C2(n18554), .A(n18276), .B(n18275), .ZN(
        P3_U2877) );
  AOI22_X1 U21326 ( .A1(n18658), .A2(n18622), .B1(n18621), .B2(n18287), .ZN(
        n18278) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18288), .B1(
        n18623), .B2(n18355), .ZN(n18277) );
  OAI211_X1 U21328 ( .C1(n18291), .C2(n18626), .A(n18278), .B(n18277), .ZN(
        P3_U2878) );
  AOI22_X1 U21329 ( .A1(n18658), .A2(n18586), .B1(n18627), .B2(n18287), .ZN(
        n18280) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18288), .B1(
        n18629), .B2(n18355), .ZN(n18279) );
  OAI211_X1 U21331 ( .C1(n18291), .C2(n18589), .A(n18280), .B(n18279), .ZN(
        P3_U2879) );
  AOI22_X1 U21332 ( .A1(n18658), .A2(n18530), .B1(n18633), .B2(n18287), .ZN(
        n18282) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18288), .B1(
        n18635), .B2(n18355), .ZN(n18281) );
  OAI211_X1 U21334 ( .C1(n18291), .C2(n18533), .A(n18282), .B(n18281), .ZN(
        P3_U2880) );
  AOI22_X1 U21335 ( .A1(n18602), .A2(n18592), .B1(n18639), .B2(n18287), .ZN(
        n18284) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18288), .B1(
        n18641), .B2(n18355), .ZN(n18283) );
  OAI211_X1 U21337 ( .C1(n18312), .C2(n18595), .A(n18284), .B(n18283), .ZN(
        P3_U2881) );
  AOI22_X1 U21338 ( .A1(n18602), .A2(n18564), .B1(n18645), .B2(n18287), .ZN(
        n18286) );
  AOI22_X1 U21339 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18288), .B1(
        n18648), .B2(n18355), .ZN(n18285) );
  OAI211_X1 U21340 ( .C1(n18312), .C2(n18567), .A(n18286), .B(n18285), .ZN(
        P3_U2882) );
  INV_X1 U21341 ( .A(n18662), .ZN(n18512) );
  AOI22_X1 U21342 ( .A1(n18658), .A2(n18512), .B1(n18654), .B2(n18287), .ZN(
        n18290) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18288), .B1(
        n18657), .B2(n18355), .ZN(n18289) );
  OAI211_X1 U21344 ( .C1(n18291), .C2(n18517), .A(n18290), .B(n18289), .ZN(
        P3_U2883) );
  INV_X1 U21345 ( .A(n18329), .ZN(n18336) );
  NOR2_X1 U21346 ( .A1(n18693), .A2(n18316), .ZN(n18359) );
  NAND2_X1 U21347 ( .A1(n18469), .A2(n18359), .ZN(n18374) );
  NOR2_X1 U21348 ( .A1(n18355), .A2(n18376), .ZN(n18337) );
  NOR2_X1 U21349 ( .A1(n18726), .A2(n18337), .ZN(n18308) );
  AOI22_X1 U21350 ( .A1(n18658), .A2(n18492), .B1(n18607), .B2(n18308), .ZN(
        n18295) );
  OAI21_X1 U21351 ( .B1(n18292), .B2(n18574), .A(n18337), .ZN(n18293) );
  OAI211_X1 U21352 ( .C1(n18376), .C2(n18833), .A(n18577), .B(n18293), .ZN(
        n18309) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18309), .B1(
        n18611), .B2(n18376), .ZN(n18294) );
  OAI211_X1 U21354 ( .C1(n18497), .C2(n18336), .A(n18295), .B(n18294), .ZN(
        P3_U2884) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18309), .B1(
        n18615), .B2(n18308), .ZN(n18297) );
  AOI22_X1 U21356 ( .A1(n18658), .A2(n18551), .B1(n18617), .B2(n18376), .ZN(
        n18296) );
  OAI211_X1 U21357 ( .C1(n18336), .C2(n18554), .A(n18297), .B(n18296), .ZN(
        P3_U2885) );
  AOI22_X1 U21358 ( .A1(n18658), .A2(n18582), .B1(n18621), .B2(n18308), .ZN(
        n18299) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18309), .B1(
        n18623), .B2(n18376), .ZN(n18298) );
  OAI211_X1 U21360 ( .C1(n18336), .C2(n18585), .A(n18299), .B(n18298), .ZN(
        P3_U2886) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18309), .B1(
        n18627), .B2(n18308), .ZN(n18301) );
  AOI22_X1 U21362 ( .A1(n18329), .A2(n18586), .B1(n18629), .B2(n18376), .ZN(
        n18300) );
  OAI211_X1 U21363 ( .C1(n18312), .C2(n18589), .A(n18301), .B(n18300), .ZN(
        P3_U2887) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18309), .B1(
        n18633), .B2(n18308), .ZN(n18303) );
  AOI22_X1 U21365 ( .A1(n18329), .A2(n18530), .B1(n18635), .B2(n18376), .ZN(
        n18302) );
  OAI211_X1 U21366 ( .C1(n18312), .C2(n18533), .A(n18303), .B(n18302), .ZN(
        P3_U2888) );
  AOI22_X1 U21367 ( .A1(n18658), .A2(n18592), .B1(n18639), .B2(n18308), .ZN(
        n18305) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18309), .B1(
        n18641), .B2(n18376), .ZN(n18304) );
  OAI211_X1 U21369 ( .C1(n18336), .C2(n18595), .A(n18305), .B(n18304), .ZN(
        P3_U2889) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18309), .B1(
        n18645), .B2(n18308), .ZN(n18307) );
  AOI22_X1 U21371 ( .A1(n18329), .A2(n18646), .B1(n18648), .B2(n18376), .ZN(
        n18306) );
  OAI211_X1 U21372 ( .C1(n18312), .C2(n18652), .A(n18307), .B(n18306), .ZN(
        P3_U2890) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18309), .B1(
        n18654), .B2(n18308), .ZN(n18311) );
  AOI22_X1 U21374 ( .A1(n18329), .A2(n18512), .B1(n18657), .B2(n18376), .ZN(
        n18310) );
  OAI211_X1 U21375 ( .C1(n18312), .C2(n18517), .A(n18311), .B(n18310), .ZN(
        P3_U2891) );
  INV_X1 U21376 ( .A(n18355), .ZN(n18353) );
  AND2_X1 U21377 ( .A1(n18606), .A2(n18359), .ZN(n18332) );
  AOI22_X1 U21378 ( .A1(n18329), .A2(n18492), .B1(n18607), .B2(n18332), .ZN(
        n18318) );
  NAND2_X1 U21379 ( .A1(n18577), .A2(n18313), .ZN(n18314) );
  OAI21_X1 U21380 ( .B1(n18693), .B2(n18314), .A(n18519), .ZN(n18609) );
  NAND2_X1 U21381 ( .A1(n18315), .A2(n18609), .ZN(n18333) );
  NOR2_X2 U21382 ( .A1(n18692), .A2(n18316), .ZN(n18398) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18333), .B1(
        n18611), .B2(n18398), .ZN(n18317) );
  OAI211_X1 U21384 ( .C1(n18497), .C2(n18353), .A(n18318), .B(n18317), .ZN(
        P3_U2892) );
  AOI22_X1 U21385 ( .A1(n18616), .A2(n18355), .B1(n18615), .B2(n18332), .ZN(
        n18320) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18333), .B1(
        n18617), .B2(n18398), .ZN(n18319) );
  OAI211_X1 U21387 ( .C1(n18336), .C2(n18620), .A(n18320), .B(n18319), .ZN(
        P3_U2893) );
  AOI22_X1 U21388 ( .A1(n18329), .A2(n18582), .B1(n18621), .B2(n18332), .ZN(
        n18322) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18333), .B1(
        n18623), .B2(n18398), .ZN(n18321) );
  OAI211_X1 U21390 ( .C1(n18585), .C2(n18353), .A(n18322), .B(n18321), .ZN(
        P3_U2894) );
  AOI22_X1 U21391 ( .A1(n18586), .A2(n18355), .B1(n18627), .B2(n18332), .ZN(
        n18324) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18333), .B1(
        n18629), .B2(n18398), .ZN(n18323) );
  OAI211_X1 U21393 ( .C1(n18336), .C2(n18589), .A(n18324), .B(n18323), .ZN(
        P3_U2895) );
  INV_X1 U21394 ( .A(n18533), .ZN(n18634) );
  AOI22_X1 U21395 ( .A1(n18329), .A2(n18634), .B1(n18633), .B2(n18332), .ZN(
        n18326) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18333), .B1(
        n18635), .B2(n18398), .ZN(n18325) );
  OAI211_X1 U21397 ( .C1(n18638), .C2(n18353), .A(n18326), .B(n18325), .ZN(
        P3_U2896) );
  AOI22_X1 U21398 ( .A1(n18329), .A2(n18592), .B1(n18639), .B2(n18332), .ZN(
        n18328) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18333), .B1(
        n18641), .B2(n18398), .ZN(n18327) );
  OAI211_X1 U21400 ( .C1(n18595), .C2(n18353), .A(n18328), .B(n18327), .ZN(
        P3_U2897) );
  AOI22_X1 U21401 ( .A1(n18329), .A2(n18564), .B1(n18645), .B2(n18332), .ZN(
        n18331) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18333), .B1(
        n18648), .B2(n18398), .ZN(n18330) );
  OAI211_X1 U21403 ( .C1(n18567), .C2(n18353), .A(n18331), .B(n18330), .ZN(
        P3_U2898) );
  AOI22_X1 U21404 ( .A1(n18512), .A2(n18355), .B1(n18654), .B2(n18332), .ZN(
        n18335) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18333), .B1(
        n18657), .B2(n18398), .ZN(n18334) );
  OAI211_X1 U21406 ( .C1(n18336), .C2(n18517), .A(n18335), .B(n18334), .ZN(
        P3_U2899) );
  NOR2_X2 U21407 ( .A1(n18694), .A2(n18403), .ZN(n18421) );
  NOR2_X1 U21408 ( .A1(n18398), .A2(n18421), .ZN(n18380) );
  NOR2_X1 U21409 ( .A1(n18726), .A2(n18380), .ZN(n18354) );
  AOI22_X1 U21410 ( .A1(n18492), .A2(n18355), .B1(n18607), .B2(n18354), .ZN(
        n18340) );
  OAI22_X1 U21411 ( .A1(n18337), .A2(n18519), .B1(n18380), .B2(n18518), .ZN(
        n18338) );
  OAI21_X1 U21412 ( .B1(n18421), .B2(n18833), .A(n18338), .ZN(n18356) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18356), .B1(
        n18611), .B2(n18421), .ZN(n18339) );
  OAI211_X1 U21414 ( .C1(n18497), .C2(n18374), .A(n18340), .B(n18339), .ZN(
        P3_U2900) );
  AOI22_X1 U21415 ( .A1(n18551), .A2(n18355), .B1(n18615), .B2(n18354), .ZN(
        n18342) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18356), .B1(
        n18617), .B2(n18421), .ZN(n18341) );
  OAI211_X1 U21417 ( .C1(n18554), .C2(n18374), .A(n18342), .B(n18341), .ZN(
        P3_U2901) );
  AOI22_X1 U21418 ( .A1(n18582), .A2(n18355), .B1(n18621), .B2(n18354), .ZN(
        n18344) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18356), .B1(
        n18623), .B2(n18421), .ZN(n18343) );
  OAI211_X1 U21420 ( .C1(n18585), .C2(n18374), .A(n18344), .B(n18343), .ZN(
        P3_U2902) );
  AOI22_X1 U21421 ( .A1(n18586), .A2(n18376), .B1(n18627), .B2(n18354), .ZN(
        n18346) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18356), .B1(
        n18629), .B2(n18421), .ZN(n18345) );
  OAI211_X1 U21423 ( .C1(n18589), .C2(n18353), .A(n18346), .B(n18345), .ZN(
        P3_U2903) );
  AOI22_X1 U21424 ( .A1(n18530), .A2(n18376), .B1(n18633), .B2(n18354), .ZN(
        n18348) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18356), .B1(
        n18635), .B2(n18421), .ZN(n18347) );
  OAI211_X1 U21426 ( .C1(n18533), .C2(n18353), .A(n18348), .B(n18347), .ZN(
        P3_U2904) );
  AOI22_X1 U21427 ( .A1(n18592), .A2(n18355), .B1(n18639), .B2(n18354), .ZN(
        n18350) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18356), .B1(
        n18641), .B2(n18421), .ZN(n18349) );
  OAI211_X1 U21429 ( .C1(n18595), .C2(n18374), .A(n18350), .B(n18349), .ZN(
        P3_U2905) );
  AOI22_X1 U21430 ( .A1(n18646), .A2(n18376), .B1(n18645), .B2(n18354), .ZN(
        n18352) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18356), .B1(
        n18648), .B2(n18421), .ZN(n18351) );
  OAI211_X1 U21432 ( .C1(n18652), .C2(n18353), .A(n18352), .B(n18351), .ZN(
        P3_U2906) );
  AOI22_X1 U21433 ( .A1(n18656), .A2(n18355), .B1(n18654), .B2(n18354), .ZN(
        n18358) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18356), .B1(
        n18657), .B2(n18421), .ZN(n18357) );
  OAI211_X1 U21435 ( .C1(n18662), .C2(n18374), .A(n18358), .B(n18357), .ZN(
        P3_U2907) );
  INV_X1 U21436 ( .A(n18398), .ZN(n18390) );
  NOR2_X1 U21437 ( .A1(n18403), .A2(n18544), .ZN(n18375) );
  AOI22_X1 U21438 ( .A1(n18492), .A2(n18376), .B1(n18607), .B2(n18375), .ZN(
        n18361) );
  AOI22_X1 U21439 ( .A1(n18548), .A2(n18359), .B1(n18402), .B2(n18546), .ZN(
        n18377) );
  NOR2_X2 U21440 ( .A1(n18403), .A2(n18448), .ZN(n18416) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18377), .B1(
        n18611), .B2(n18416), .ZN(n18360) );
  OAI211_X1 U21442 ( .C1(n18497), .C2(n18390), .A(n18361), .B(n18360), .ZN(
        P3_U2908) );
  AOI22_X1 U21443 ( .A1(n18551), .A2(n18376), .B1(n18615), .B2(n18375), .ZN(
        n18363) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18377), .B1(
        n18617), .B2(n18416), .ZN(n18362) );
  OAI211_X1 U21445 ( .C1(n18554), .C2(n18390), .A(n18363), .B(n18362), .ZN(
        P3_U2909) );
  AOI22_X1 U21446 ( .A1(n18621), .A2(n18375), .B1(n18622), .B2(n18398), .ZN(
        n18365) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18377), .B1(
        n18623), .B2(n18416), .ZN(n18364) );
  OAI211_X1 U21448 ( .C1(n18626), .C2(n18374), .A(n18365), .B(n18364), .ZN(
        P3_U2910) );
  AOI22_X1 U21449 ( .A1(n18628), .A2(n18376), .B1(n18627), .B2(n18375), .ZN(
        n18367) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18377), .B1(
        n18629), .B2(n18416), .ZN(n18366) );
  OAI211_X1 U21451 ( .C1(n18632), .C2(n18390), .A(n18367), .B(n18366), .ZN(
        P3_U2911) );
  AOI22_X1 U21452 ( .A1(n18634), .A2(n18376), .B1(n18633), .B2(n18375), .ZN(
        n18369) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18377), .B1(
        n18635), .B2(n18416), .ZN(n18368) );
  OAI211_X1 U21454 ( .C1(n18638), .C2(n18390), .A(n18369), .B(n18368), .ZN(
        P3_U2912) );
  AOI22_X1 U21455 ( .A1(n18592), .A2(n18376), .B1(n18639), .B2(n18375), .ZN(
        n18371) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18377), .B1(
        n18641), .B2(n18416), .ZN(n18370) );
  OAI211_X1 U21457 ( .C1(n18595), .C2(n18390), .A(n18371), .B(n18370), .ZN(
        P3_U2913) );
  AOI22_X1 U21458 ( .A1(n18646), .A2(n18398), .B1(n18645), .B2(n18375), .ZN(
        n18373) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18377), .B1(
        n18648), .B2(n18416), .ZN(n18372) );
  OAI211_X1 U21460 ( .C1(n18652), .C2(n18374), .A(n18373), .B(n18372), .ZN(
        P3_U2914) );
  AOI22_X1 U21461 ( .A1(n18656), .A2(n18376), .B1(n18654), .B2(n18375), .ZN(
        n18379) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18377), .B1(
        n18657), .B2(n18416), .ZN(n18378) );
  OAI211_X1 U21463 ( .C1(n18662), .C2(n18390), .A(n18379), .B(n18378), .ZN(
        P3_U2915) );
  OR3_X1 U21464 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18446), .ZN(n18468) );
  INV_X1 U21465 ( .A(n18468), .ZN(n18459) );
  NOR2_X1 U21466 ( .A1(n18416), .A2(n18459), .ZN(n18425) );
  NOR2_X1 U21467 ( .A1(n18726), .A2(n18425), .ZN(n18397) );
  AOI22_X1 U21468 ( .A1(n18608), .A2(n18421), .B1(n18607), .B2(n18397), .ZN(
        n18383) );
  OAI21_X1 U21469 ( .B1(n18380), .B2(n18574), .A(n18425), .ZN(n18381) );
  OAI211_X1 U21470 ( .C1(n18459), .C2(n18833), .A(n18577), .B(n18381), .ZN(
        n18399) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18399), .B1(
        n18611), .B2(n18459), .ZN(n18382) );
  OAI211_X1 U21472 ( .C1(n18614), .C2(n18390), .A(n18383), .B(n18382), .ZN(
        P3_U2916) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18399), .B1(
        n18615), .B2(n18397), .ZN(n18385) );
  AOI22_X1 U21474 ( .A1(n18617), .A2(n18459), .B1(n18616), .B2(n18421), .ZN(
        n18384) );
  OAI211_X1 U21475 ( .C1(n18620), .C2(n18390), .A(n18385), .B(n18384), .ZN(
        P3_U2917) );
  INV_X1 U21476 ( .A(n18421), .ZN(n18419) );
  AOI22_X1 U21477 ( .A1(n18582), .A2(n18398), .B1(n18621), .B2(n18397), .ZN(
        n18387) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18399), .B1(
        n18623), .B2(n18459), .ZN(n18386) );
  OAI211_X1 U21479 ( .C1(n18585), .C2(n18419), .A(n18387), .B(n18386), .ZN(
        P3_U2918) );
  AOI22_X1 U21480 ( .A1(n18586), .A2(n18421), .B1(n18627), .B2(n18397), .ZN(
        n18389) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18399), .B1(
        n18629), .B2(n18459), .ZN(n18388) );
  OAI211_X1 U21482 ( .C1(n18589), .C2(n18390), .A(n18389), .B(n18388), .ZN(
        P3_U2919) );
  AOI22_X1 U21483 ( .A1(n18634), .A2(n18398), .B1(n18633), .B2(n18397), .ZN(
        n18392) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18399), .B1(
        n18635), .B2(n18459), .ZN(n18391) );
  OAI211_X1 U21485 ( .C1(n18638), .C2(n18419), .A(n18392), .B(n18391), .ZN(
        P3_U2920) );
  AOI22_X1 U21486 ( .A1(n18592), .A2(n18398), .B1(n18639), .B2(n18397), .ZN(
        n18394) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18399), .B1(
        n18641), .B2(n18459), .ZN(n18393) );
  OAI211_X1 U21488 ( .C1(n18595), .C2(n18419), .A(n18394), .B(n18393), .ZN(
        P3_U2921) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18399), .B1(
        n18645), .B2(n18397), .ZN(n18396) );
  AOI22_X1 U21490 ( .A1(n18564), .A2(n18398), .B1(n18648), .B2(n18459), .ZN(
        n18395) );
  OAI211_X1 U21491 ( .C1(n18567), .C2(n18419), .A(n18396), .B(n18395), .ZN(
        P3_U2922) );
  AOI22_X1 U21492 ( .A1(n18656), .A2(n18398), .B1(n18654), .B2(n18397), .ZN(
        n18401) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18399), .B1(
        n18657), .B2(n18459), .ZN(n18400) );
  OAI211_X1 U21494 ( .C1(n18662), .C2(n18419), .A(n18401), .B(n18400), .ZN(
        P3_U2923) );
  AOI22_X1 U21495 ( .A1(n18608), .A2(n18416), .B1(n18607), .B2(n18420), .ZN(
        n18405) );
  NAND2_X1 U21496 ( .A1(n18402), .A2(n18609), .ZN(n18422) );
  NOR2_X2 U21497 ( .A1(n18692), .A2(n18403), .ZN(n18488) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18422), .B1(
        n18611), .B2(n18488), .ZN(n18404) );
  OAI211_X1 U21499 ( .C1(n18614), .C2(n18419), .A(n18405), .B(n18404), .ZN(
        P3_U2924) );
  INV_X1 U21500 ( .A(n18416), .ZN(n18445) );
  AOI22_X1 U21501 ( .A1(n18551), .A2(n18421), .B1(n18615), .B2(n18420), .ZN(
        n18407) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18422), .B1(
        n18617), .B2(n18488), .ZN(n18406) );
  OAI211_X1 U21503 ( .C1(n18554), .C2(n18445), .A(n18407), .B(n18406), .ZN(
        P3_U2925) );
  AOI22_X1 U21504 ( .A1(n18582), .A2(n18421), .B1(n18621), .B2(n18420), .ZN(
        n18409) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18422), .B1(
        n18623), .B2(n18488), .ZN(n18408) );
  OAI211_X1 U21506 ( .C1(n18585), .C2(n18445), .A(n18409), .B(n18408), .ZN(
        P3_U2926) );
  AOI22_X1 U21507 ( .A1(n18586), .A2(n18416), .B1(n18627), .B2(n18420), .ZN(
        n18411) );
  AOI22_X1 U21508 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18422), .B1(
        n18629), .B2(n18488), .ZN(n18410) );
  OAI211_X1 U21509 ( .C1(n18589), .C2(n18419), .A(n18411), .B(n18410), .ZN(
        P3_U2927) );
  AOI22_X1 U21510 ( .A1(n18530), .A2(n18416), .B1(n18633), .B2(n18420), .ZN(
        n18413) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18422), .B1(
        n18635), .B2(n18488), .ZN(n18412) );
  OAI211_X1 U21512 ( .C1(n18533), .C2(n18419), .A(n18413), .B(n18412), .ZN(
        P3_U2928) );
  AOI22_X1 U21513 ( .A1(n18592), .A2(n18421), .B1(n18639), .B2(n18420), .ZN(
        n18415) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18422), .B1(
        n18641), .B2(n18488), .ZN(n18414) );
  OAI211_X1 U21515 ( .C1(n18595), .C2(n18445), .A(n18415), .B(n18414), .ZN(
        P3_U2929) );
  AOI22_X1 U21516 ( .A1(n18646), .A2(n18416), .B1(n18645), .B2(n18420), .ZN(
        n18418) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18422), .B1(
        n18648), .B2(n18488), .ZN(n18417) );
  OAI211_X1 U21518 ( .C1(n18652), .C2(n18419), .A(n18418), .B(n18417), .ZN(
        P3_U2930) );
  AOI22_X1 U21519 ( .A1(n18656), .A2(n18421), .B1(n18654), .B2(n18420), .ZN(
        n18424) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18422), .B1(
        n18657), .B2(n18488), .ZN(n18423) );
  OAI211_X1 U21521 ( .C1(n18662), .C2(n18445), .A(n18424), .B(n18423), .ZN(
        P3_U2931) );
  NOR2_X2 U21522 ( .A1(n18694), .A2(n18494), .ZN(n18506) );
  NOR2_X1 U21523 ( .A1(n18488), .A2(n18506), .ZN(n18470) );
  NOR2_X1 U21524 ( .A1(n18726), .A2(n18470), .ZN(n18441) );
  AOI22_X1 U21525 ( .A1(n18608), .A2(n18459), .B1(n18607), .B2(n18441), .ZN(
        n18428) );
  OAI22_X1 U21526 ( .A1(n18425), .A2(n18519), .B1(n18470), .B2(n18518), .ZN(
        n18426) );
  OAI21_X1 U21527 ( .B1(n18506), .B2(n18833), .A(n18426), .ZN(n18442) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18442), .B1(
        n18611), .B2(n18506), .ZN(n18427) );
  OAI211_X1 U21529 ( .C1(n18614), .C2(n18445), .A(n18428), .B(n18427), .ZN(
        P3_U2932) );
  AOI22_X1 U21530 ( .A1(n18616), .A2(n18459), .B1(n18615), .B2(n18441), .ZN(
        n18430) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18442), .B1(
        n18617), .B2(n18506), .ZN(n18429) );
  OAI211_X1 U21532 ( .C1(n18620), .C2(n18445), .A(n18430), .B(n18429), .ZN(
        P3_U2933) );
  AOI22_X1 U21533 ( .A1(n18621), .A2(n18441), .B1(n18622), .B2(n18459), .ZN(
        n18432) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18442), .B1(
        n18623), .B2(n18506), .ZN(n18431) );
  OAI211_X1 U21535 ( .C1(n18626), .C2(n18445), .A(n18432), .B(n18431), .ZN(
        P3_U2934) );
  AOI22_X1 U21536 ( .A1(n18586), .A2(n18459), .B1(n18627), .B2(n18441), .ZN(
        n18434) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18442), .B1(
        n18629), .B2(n18506), .ZN(n18433) );
  OAI211_X1 U21538 ( .C1(n18589), .C2(n18445), .A(n18434), .B(n18433), .ZN(
        P3_U2935) );
  AOI22_X1 U21539 ( .A1(n18530), .A2(n18459), .B1(n18633), .B2(n18441), .ZN(
        n18436) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18442), .B1(
        n18635), .B2(n18506), .ZN(n18435) );
  OAI211_X1 U21541 ( .C1(n18533), .C2(n18445), .A(n18436), .B(n18435), .ZN(
        P3_U2936) );
  AOI22_X1 U21542 ( .A1(n18639), .A2(n18441), .B1(n18640), .B2(n18459), .ZN(
        n18438) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18442), .B1(
        n18641), .B2(n18506), .ZN(n18437) );
  OAI211_X1 U21544 ( .C1(n18644), .C2(n18445), .A(n18438), .B(n18437), .ZN(
        P3_U2937) );
  AOI22_X1 U21545 ( .A1(n18646), .A2(n18459), .B1(n18645), .B2(n18441), .ZN(
        n18440) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18442), .B1(
        n18648), .B2(n18506), .ZN(n18439) );
  OAI211_X1 U21547 ( .C1(n18652), .C2(n18445), .A(n18440), .B(n18439), .ZN(
        P3_U2938) );
  AOI22_X1 U21548 ( .A1(n18512), .A2(n18459), .B1(n18654), .B2(n18441), .ZN(
        n18444) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18442), .B1(
        n18657), .B2(n18506), .ZN(n18443) );
  OAI211_X1 U21550 ( .C1(n18517), .C2(n18445), .A(n18444), .B(n18443), .ZN(
        P3_U2939) );
  INV_X1 U21551 ( .A(n18488), .ZN(n18486) );
  NOR2_X1 U21552 ( .A1(n18494), .A2(n18544), .ZN(n18464) );
  AOI22_X1 U21553 ( .A1(n18492), .A2(n18459), .B1(n18607), .B2(n18464), .ZN(
        n18450) );
  NOR2_X1 U21554 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18446), .ZN(
        n18447) );
  AOI22_X1 U21555 ( .A1(n18548), .A2(n18447), .B1(n18493), .B2(n18546), .ZN(
        n18465) );
  NOR2_X2 U21556 ( .A1(n18494), .A2(n18448), .ZN(n18540) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18465), .B1(
        n18611), .B2(n18540), .ZN(n18449) );
  OAI211_X1 U21558 ( .C1(n18497), .C2(n18486), .A(n18450), .B(n18449), .ZN(
        P3_U2940) );
  AOI22_X1 U21559 ( .A1(n18551), .A2(n18459), .B1(n18615), .B2(n18464), .ZN(
        n18452) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18465), .B1(
        n18617), .B2(n18540), .ZN(n18451) );
  OAI211_X1 U21561 ( .C1(n18554), .C2(n18486), .A(n18452), .B(n18451), .ZN(
        P3_U2941) );
  AOI22_X1 U21562 ( .A1(n18621), .A2(n18464), .B1(n18622), .B2(n18488), .ZN(
        n18454) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18465), .B1(
        n18623), .B2(n18540), .ZN(n18453) );
  OAI211_X1 U21564 ( .C1(n18626), .C2(n18468), .A(n18454), .B(n18453), .ZN(
        P3_U2942) );
  AOI22_X1 U21565 ( .A1(n18628), .A2(n18459), .B1(n18627), .B2(n18464), .ZN(
        n18456) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18465), .B1(
        n18629), .B2(n18540), .ZN(n18455) );
  OAI211_X1 U21567 ( .C1(n18632), .C2(n18486), .A(n18456), .B(n18455), .ZN(
        P3_U2943) );
  AOI22_X1 U21568 ( .A1(n18634), .A2(n18459), .B1(n18633), .B2(n18464), .ZN(
        n18458) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18465), .B1(
        n18635), .B2(n18540), .ZN(n18457) );
  OAI211_X1 U21570 ( .C1(n18638), .C2(n18486), .A(n18458), .B(n18457), .ZN(
        P3_U2944) );
  AOI22_X1 U21571 ( .A1(n18592), .A2(n18459), .B1(n18639), .B2(n18464), .ZN(
        n18461) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18465), .B1(
        n18641), .B2(n18540), .ZN(n18460) );
  OAI211_X1 U21573 ( .C1(n18595), .C2(n18486), .A(n18461), .B(n18460), .ZN(
        P3_U2945) );
  AOI22_X1 U21574 ( .A1(n18646), .A2(n18488), .B1(n18645), .B2(n18464), .ZN(
        n18463) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18465), .B1(
        n18648), .B2(n18540), .ZN(n18462) );
  OAI211_X1 U21576 ( .C1(n18652), .C2(n18468), .A(n18463), .B(n18462), .ZN(
        P3_U2946) );
  AOI22_X1 U21577 ( .A1(n18512), .A2(n18488), .B1(n18654), .B2(n18464), .ZN(
        n18467) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18465), .B1(
        n18657), .B2(n18540), .ZN(n18466) );
  OAI211_X1 U21579 ( .C1(n18517), .C2(n18468), .A(n18467), .B(n18466), .ZN(
        P3_U2947) );
  NOR2_X1 U21580 ( .A1(n18693), .A2(n18494), .ZN(n18547) );
  NAND2_X1 U21581 ( .A1(n18469), .A2(n18547), .ZN(n18563) );
  NOR2_X1 U21582 ( .A1(n18540), .A2(n18569), .ZN(n18520) );
  OAI21_X1 U21583 ( .B1(n18470), .B2(n18574), .A(n18520), .ZN(n18471) );
  OAI211_X1 U21584 ( .C1(n18569), .C2(n18833), .A(n18577), .B(n18471), .ZN(
        n18489) );
  NOR2_X1 U21585 ( .A1(n18726), .A2(n18520), .ZN(n18487) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18489), .B1(
        n18607), .B2(n18487), .ZN(n18473) );
  AOI22_X1 U21587 ( .A1(n18608), .A2(n18506), .B1(n18611), .B2(n18569), .ZN(
        n18472) );
  OAI211_X1 U21588 ( .C1(n18614), .C2(n18486), .A(n18473), .B(n18472), .ZN(
        P3_U2948) );
  INV_X1 U21589 ( .A(n18506), .ZN(n18516) );
  AOI22_X1 U21590 ( .A1(n18551), .A2(n18488), .B1(n18615), .B2(n18487), .ZN(
        n18475) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18489), .B1(
        n18617), .B2(n18569), .ZN(n18474) );
  OAI211_X1 U21592 ( .C1(n18554), .C2(n18516), .A(n18475), .B(n18474), .ZN(
        P3_U2949) );
  AOI22_X1 U21593 ( .A1(n18582), .A2(n18488), .B1(n18621), .B2(n18487), .ZN(
        n18477) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18489), .B1(
        n18623), .B2(n18569), .ZN(n18476) );
  OAI211_X1 U21595 ( .C1(n18585), .C2(n18516), .A(n18477), .B(n18476), .ZN(
        P3_U2950) );
  AOI22_X1 U21596 ( .A1(n18586), .A2(n18506), .B1(n18627), .B2(n18487), .ZN(
        n18479) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18489), .B1(
        n18629), .B2(n18569), .ZN(n18478) );
  OAI211_X1 U21598 ( .C1(n18589), .C2(n18486), .A(n18479), .B(n18478), .ZN(
        P3_U2951) );
  AOI22_X1 U21599 ( .A1(n18530), .A2(n18506), .B1(n18633), .B2(n18487), .ZN(
        n18481) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18489), .B1(
        n18635), .B2(n18569), .ZN(n18480) );
  OAI211_X1 U21601 ( .C1(n18533), .C2(n18486), .A(n18481), .B(n18480), .ZN(
        P3_U2952) );
  AOI22_X1 U21602 ( .A1(n18592), .A2(n18488), .B1(n18639), .B2(n18487), .ZN(
        n18483) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18489), .B1(
        n18641), .B2(n18569), .ZN(n18482) );
  OAI211_X1 U21604 ( .C1(n18595), .C2(n18516), .A(n18483), .B(n18482), .ZN(
        P3_U2953) );
  AOI22_X1 U21605 ( .A1(n18646), .A2(n18506), .B1(n18645), .B2(n18487), .ZN(
        n18485) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18489), .B1(
        n18648), .B2(n18569), .ZN(n18484) );
  OAI211_X1 U21607 ( .C1(n18652), .C2(n18486), .A(n18485), .B(n18484), .ZN(
        P3_U2954) );
  AOI22_X1 U21608 ( .A1(n18656), .A2(n18488), .B1(n18654), .B2(n18487), .ZN(
        n18491) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18489), .B1(
        n18657), .B2(n18569), .ZN(n18490) );
  OAI211_X1 U21610 ( .C1(n18662), .C2(n18516), .A(n18491), .B(n18490), .ZN(
        P3_U2955) );
  INV_X1 U21611 ( .A(n18540), .ZN(n18536) );
  AND2_X1 U21612 ( .A1(n18606), .A2(n18547), .ZN(n18511) );
  AOI22_X1 U21613 ( .A1(n18492), .A2(n18506), .B1(n18607), .B2(n18511), .ZN(
        n18496) );
  NAND2_X1 U21614 ( .A1(n18493), .A2(n18609), .ZN(n18513) );
  NOR2_X2 U21615 ( .A1(n18692), .A2(n18494), .ZN(n18601) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18513), .B1(
        n18611), .B2(n18601), .ZN(n18495) );
  OAI211_X1 U21617 ( .C1(n18497), .C2(n18536), .A(n18496), .B(n18495), .ZN(
        P3_U2956) );
  AOI22_X1 U21618 ( .A1(n18616), .A2(n18540), .B1(n18615), .B2(n18511), .ZN(
        n18499) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18513), .B1(
        n18617), .B2(n18601), .ZN(n18498) );
  OAI211_X1 U21620 ( .C1(n18620), .C2(n18516), .A(n18499), .B(n18498), .ZN(
        P3_U2957) );
  AOI22_X1 U21621 ( .A1(n18582), .A2(n18506), .B1(n18621), .B2(n18511), .ZN(
        n18501) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18513), .B1(
        n18623), .B2(n18601), .ZN(n18500) );
  OAI211_X1 U21623 ( .C1(n18585), .C2(n18536), .A(n18501), .B(n18500), .ZN(
        P3_U2958) );
  AOI22_X1 U21624 ( .A1(n18586), .A2(n18540), .B1(n18627), .B2(n18511), .ZN(
        n18503) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18513), .B1(
        n18629), .B2(n18601), .ZN(n18502) );
  OAI211_X1 U21626 ( .C1(n18589), .C2(n18516), .A(n18503), .B(n18502), .ZN(
        P3_U2959) );
  AOI22_X1 U21627 ( .A1(n18530), .A2(n18540), .B1(n18633), .B2(n18511), .ZN(
        n18505) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18513), .B1(
        n18635), .B2(n18601), .ZN(n18504) );
  OAI211_X1 U21629 ( .C1(n18533), .C2(n18516), .A(n18505), .B(n18504), .ZN(
        P3_U2960) );
  AOI22_X1 U21630 ( .A1(n18592), .A2(n18506), .B1(n18639), .B2(n18511), .ZN(
        n18508) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18513), .B1(
        n18641), .B2(n18601), .ZN(n18507) );
  OAI211_X1 U21632 ( .C1(n18595), .C2(n18536), .A(n18508), .B(n18507), .ZN(
        P3_U2961) );
  AOI22_X1 U21633 ( .A1(n18646), .A2(n18540), .B1(n18645), .B2(n18511), .ZN(
        n18510) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18513), .B1(
        n18648), .B2(n18601), .ZN(n18509) );
  OAI211_X1 U21635 ( .C1(n18652), .C2(n18516), .A(n18510), .B(n18509), .ZN(
        P3_U2962) );
  AOI22_X1 U21636 ( .A1(n18512), .A2(n18540), .B1(n18654), .B2(n18511), .ZN(
        n18515) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18513), .B1(
        n18657), .B2(n18601), .ZN(n18514) );
  OAI211_X1 U21638 ( .C1(n18517), .C2(n18516), .A(n18515), .B(n18514), .ZN(
        P3_U2963) );
  NOR2_X2 U21639 ( .A1(n18694), .A2(n18545), .ZN(n18655) );
  NOR2_X1 U21640 ( .A1(n18601), .A2(n18655), .ZN(n18575) );
  NOR2_X1 U21641 ( .A1(n18726), .A2(n18575), .ZN(n18539) );
  AOI22_X1 U21642 ( .A1(n18608), .A2(n18569), .B1(n18607), .B2(n18539), .ZN(
        n18523) );
  OAI22_X1 U21643 ( .A1(n18520), .A2(n18519), .B1(n18575), .B2(n18518), .ZN(
        n18521) );
  OAI21_X1 U21644 ( .B1(n18655), .B2(n18833), .A(n18521), .ZN(n18541) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18541), .B1(
        n18611), .B2(n18655), .ZN(n18522) );
  OAI211_X1 U21646 ( .C1(n18614), .C2(n18536), .A(n18523), .B(n18522), .ZN(
        P3_U2964) );
  AOI22_X1 U21647 ( .A1(n18551), .A2(n18540), .B1(n18615), .B2(n18539), .ZN(
        n18525) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18541), .B1(
        n18617), .B2(n18655), .ZN(n18524) );
  OAI211_X1 U21649 ( .C1(n18554), .C2(n18563), .A(n18525), .B(n18524), .ZN(
        P3_U2965) );
  AOI22_X1 U21650 ( .A1(n18621), .A2(n18539), .B1(n18622), .B2(n18569), .ZN(
        n18527) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18541), .B1(
        n18623), .B2(n18655), .ZN(n18526) );
  OAI211_X1 U21652 ( .C1(n18626), .C2(n18536), .A(n18527), .B(n18526), .ZN(
        P3_U2966) );
  AOI22_X1 U21653 ( .A1(n18628), .A2(n18540), .B1(n18627), .B2(n18539), .ZN(
        n18529) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18541), .B1(
        n18629), .B2(n18655), .ZN(n18528) );
  OAI211_X1 U21655 ( .C1(n18632), .C2(n18563), .A(n18529), .B(n18528), .ZN(
        P3_U2967) );
  AOI22_X1 U21656 ( .A1(n18530), .A2(n18569), .B1(n18633), .B2(n18539), .ZN(
        n18532) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18541), .B1(
        n18635), .B2(n18655), .ZN(n18531) );
  OAI211_X1 U21658 ( .C1(n18533), .C2(n18536), .A(n18532), .B(n18531), .ZN(
        P3_U2968) );
  AOI22_X1 U21659 ( .A1(n18639), .A2(n18539), .B1(n18640), .B2(n18569), .ZN(
        n18535) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18541), .B1(
        n18641), .B2(n18655), .ZN(n18534) );
  OAI211_X1 U21661 ( .C1(n18644), .C2(n18536), .A(n18535), .B(n18534), .ZN(
        P3_U2969) );
  AOI22_X1 U21662 ( .A1(n18564), .A2(n18540), .B1(n18645), .B2(n18539), .ZN(
        n18538) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18541), .B1(
        n18648), .B2(n18655), .ZN(n18537) );
  OAI211_X1 U21664 ( .C1(n18567), .C2(n18563), .A(n18538), .B(n18537), .ZN(
        P3_U2970) );
  AOI22_X1 U21665 ( .A1(n18656), .A2(n18540), .B1(n18654), .B2(n18539), .ZN(
        n18543) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18541), .B1(
        n18657), .B2(n18655), .ZN(n18542) );
  OAI211_X1 U21667 ( .C1(n18662), .C2(n18563), .A(n18543), .B(n18542), .ZN(
        P3_U2971) );
  NOR2_X1 U21668 ( .A1(n18545), .A2(n18544), .ZN(n18568) );
  AOI22_X1 U21669 ( .A1(n18608), .A2(n18601), .B1(n18607), .B2(n18568), .ZN(
        n18550) );
  AOI22_X1 U21670 ( .A1(n18548), .A2(n18547), .B1(n18610), .B2(n18546), .ZN(
        n18570) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18570), .B1(
        n18647), .B2(n18611), .ZN(n18549) );
  OAI211_X1 U21672 ( .C1(n18614), .C2(n18563), .A(n18550), .B(n18549), .ZN(
        P3_U2972) );
  INV_X1 U21673 ( .A(n18601), .ZN(n18598) );
  AOI22_X1 U21674 ( .A1(n18551), .A2(n18569), .B1(n18615), .B2(n18568), .ZN(
        n18553) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18570), .B1(
        n18647), .B2(n18617), .ZN(n18552) );
  OAI211_X1 U21676 ( .C1(n18554), .C2(n18598), .A(n18553), .B(n18552), .ZN(
        P3_U2973) );
  AOI22_X1 U21677 ( .A1(n18621), .A2(n18568), .B1(n18622), .B2(n18601), .ZN(
        n18556) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18570), .B1(
        n18647), .B2(n18623), .ZN(n18555) );
  OAI211_X1 U21679 ( .C1(n18626), .C2(n18563), .A(n18556), .B(n18555), .ZN(
        P3_U2974) );
  AOI22_X1 U21680 ( .A1(n18586), .A2(n18601), .B1(n18627), .B2(n18568), .ZN(
        n18558) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18570), .B1(
        n18647), .B2(n18629), .ZN(n18557) );
  OAI211_X1 U21682 ( .C1(n18589), .C2(n18563), .A(n18558), .B(n18557), .ZN(
        P3_U2975) );
  AOI22_X1 U21683 ( .A1(n18634), .A2(n18569), .B1(n18633), .B2(n18568), .ZN(
        n18560) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18570), .B1(
        n18647), .B2(n18635), .ZN(n18559) );
  OAI211_X1 U21685 ( .C1(n18638), .C2(n18598), .A(n18560), .B(n18559), .ZN(
        P3_U2976) );
  AOI22_X1 U21686 ( .A1(n18639), .A2(n18568), .B1(n18640), .B2(n18601), .ZN(
        n18562) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18570), .B1(
        n18647), .B2(n18641), .ZN(n18561) );
  OAI211_X1 U21688 ( .C1(n18644), .C2(n18563), .A(n18562), .B(n18561), .ZN(
        P3_U2977) );
  AOI22_X1 U21689 ( .A1(n18564), .A2(n18569), .B1(n18645), .B2(n18568), .ZN(
        n18566) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18570), .B1(
        n18647), .B2(n18648), .ZN(n18565) );
  OAI211_X1 U21691 ( .C1(n18567), .C2(n18598), .A(n18566), .B(n18565), .ZN(
        P3_U2978) );
  AOI22_X1 U21692 ( .A1(n18656), .A2(n18569), .B1(n18654), .B2(n18568), .ZN(
        n18572) );
  AOI22_X1 U21693 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18570), .B1(
        n18647), .B2(n18657), .ZN(n18571) );
  OAI211_X1 U21694 ( .C1(n18662), .C2(n18598), .A(n18572), .B(n18571), .ZN(
        P3_U2979) );
  NOR2_X1 U21695 ( .A1(n18726), .A2(n18573), .ZN(n18599) );
  AOI22_X1 U21696 ( .A1(n18608), .A2(n18655), .B1(n18607), .B2(n18599), .ZN(
        n18579) );
  OAI21_X1 U21697 ( .B1(n18575), .B2(n18574), .A(n18573), .ZN(n18576) );
  OAI211_X1 U21698 ( .C1(n18602), .C2(n18833), .A(n18577), .B(n18576), .ZN(
        n18600) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18600), .B1(
        n18602), .B2(n18611), .ZN(n18578) );
  OAI211_X1 U21700 ( .C1(n18614), .C2(n18598), .A(n18579), .B(n18578), .ZN(
        P3_U2980) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18600), .B1(
        n18615), .B2(n18599), .ZN(n18581) );
  AOI22_X1 U21702 ( .A1(n18602), .A2(n18617), .B1(n18616), .B2(n18655), .ZN(
        n18580) );
  OAI211_X1 U21703 ( .C1(n18620), .C2(n18598), .A(n18581), .B(n18580), .ZN(
        P3_U2981) );
  INV_X1 U21704 ( .A(n18655), .ZN(n18651) );
  AOI22_X1 U21705 ( .A1(n18582), .A2(n18601), .B1(n18621), .B2(n18599), .ZN(
        n18584) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18600), .B1(
        n18602), .B2(n18623), .ZN(n18583) );
  OAI211_X1 U21707 ( .C1(n18585), .C2(n18651), .A(n18584), .B(n18583), .ZN(
        P3_U2982) );
  AOI22_X1 U21708 ( .A1(n18586), .A2(n18655), .B1(n18627), .B2(n18599), .ZN(
        n18588) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18600), .B1(
        n18602), .B2(n18629), .ZN(n18587) );
  OAI211_X1 U21710 ( .C1(n18589), .C2(n18598), .A(n18588), .B(n18587), .ZN(
        P3_U2983) );
  AOI22_X1 U21711 ( .A1(n18634), .A2(n18601), .B1(n18633), .B2(n18599), .ZN(
        n18591) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18600), .B1(
        n18602), .B2(n18635), .ZN(n18590) );
  OAI211_X1 U21713 ( .C1(n18638), .C2(n18651), .A(n18591), .B(n18590), .ZN(
        P3_U2984) );
  AOI22_X1 U21714 ( .A1(n18592), .A2(n18601), .B1(n18639), .B2(n18599), .ZN(
        n18594) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18600), .B1(
        n18602), .B2(n18641), .ZN(n18593) );
  OAI211_X1 U21716 ( .C1(n18595), .C2(n18651), .A(n18594), .B(n18593), .ZN(
        P3_U2985) );
  AOI22_X1 U21717 ( .A1(n18646), .A2(n18655), .B1(n18645), .B2(n18599), .ZN(
        n18597) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18600), .B1(
        n18602), .B2(n18648), .ZN(n18596) );
  OAI211_X1 U21719 ( .C1(n18652), .C2(n18598), .A(n18597), .B(n18596), .ZN(
        P3_U2986) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18600), .B1(
        n18654), .B2(n18599), .ZN(n18604) );
  AOI22_X1 U21721 ( .A1(n18602), .A2(n18657), .B1(n18656), .B2(n18601), .ZN(
        n18603) );
  OAI211_X1 U21722 ( .C1(n18662), .C2(n18651), .A(n18604), .B(n18603), .ZN(
        P3_U2987) );
  AND2_X1 U21723 ( .A1(n18606), .A2(n18605), .ZN(n18653) );
  AOI22_X1 U21724 ( .A1(n18608), .A2(n18647), .B1(n18607), .B2(n18653), .ZN(
        n18613) );
  NAND2_X1 U21725 ( .A1(n18610), .A2(n18609), .ZN(n18659) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18659), .B1(
        n18658), .B2(n18611), .ZN(n18612) );
  OAI211_X1 U21727 ( .C1(n18614), .C2(n18651), .A(n18613), .B(n18612), .ZN(
        P3_U2988) );
  AOI22_X1 U21728 ( .A1(n18647), .A2(n18616), .B1(n18615), .B2(n18653), .ZN(
        n18619) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18659), .B1(
        n18658), .B2(n18617), .ZN(n18618) );
  OAI211_X1 U21730 ( .C1(n18620), .C2(n18651), .A(n18619), .B(n18618), .ZN(
        P3_U2989) );
  AOI22_X1 U21731 ( .A1(n18647), .A2(n18622), .B1(n18621), .B2(n18653), .ZN(
        n18625) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18659), .B1(
        n18658), .B2(n18623), .ZN(n18624) );
  OAI211_X1 U21733 ( .C1(n18626), .C2(n18651), .A(n18625), .B(n18624), .ZN(
        P3_U2990) );
  AOI22_X1 U21734 ( .A1(n18628), .A2(n18655), .B1(n18627), .B2(n18653), .ZN(
        n18631) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18659), .B1(
        n18658), .B2(n18629), .ZN(n18630) );
  OAI211_X1 U21736 ( .C1(n18663), .C2(n18632), .A(n18631), .B(n18630), .ZN(
        P3_U2991) );
  AOI22_X1 U21737 ( .A1(n18634), .A2(n18655), .B1(n18633), .B2(n18653), .ZN(
        n18637) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18659), .B1(
        n18658), .B2(n18635), .ZN(n18636) );
  OAI211_X1 U21739 ( .C1(n18663), .C2(n18638), .A(n18637), .B(n18636), .ZN(
        P3_U2992) );
  AOI22_X1 U21740 ( .A1(n18647), .A2(n18640), .B1(n18639), .B2(n18653), .ZN(
        n18643) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18659), .B1(
        n18658), .B2(n18641), .ZN(n18642) );
  OAI211_X1 U21742 ( .C1(n18644), .C2(n18651), .A(n18643), .B(n18642), .ZN(
        P3_U2993) );
  AOI22_X1 U21743 ( .A1(n18647), .A2(n18646), .B1(n18645), .B2(n18653), .ZN(
        n18650) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18659), .B1(
        n18658), .B2(n18648), .ZN(n18649) );
  OAI211_X1 U21745 ( .C1(n18652), .C2(n18651), .A(n18650), .B(n18649), .ZN(
        P3_U2994) );
  AOI22_X1 U21746 ( .A1(n18656), .A2(n18655), .B1(n18654), .B2(n18653), .ZN(
        n18661) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18659), .B1(
        n18658), .B2(n18657), .ZN(n18660) );
  OAI211_X1 U21748 ( .C1(n18663), .C2(n18662), .A(n18661), .B(n18660), .ZN(
        P3_U2995) );
  NOR2_X1 U21749 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18664), .ZN(
        n18690) );
  INV_X1 U21750 ( .A(n18690), .ZN(n18665) );
  AOI22_X1 U21751 ( .A1(n18707), .A2(n18669), .B1(n18676), .B2(n18665), .ZN(
        n18836) );
  NOR2_X1 U21752 ( .A1(n18696), .A2(n18836), .ZN(n18673) );
  OAI21_X1 U21753 ( .B1(n18668), .B2(n18667), .A(n18666), .ZN(n18674) );
  OAI21_X1 U21754 ( .B1(n18689), .B2(n18676), .A(n18669), .ZN(n18670) );
  AOI21_X1 U21755 ( .B1(n18671), .B2(n18674), .A(n18670), .ZN(n18834) );
  NAND2_X1 U21756 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18834), .ZN(
        n18672) );
  OAI22_X1 U21757 ( .A1(n18673), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18696), .B2(n18672), .ZN(n18703) );
  AOI21_X1 U21758 ( .B1(n18859), .B2(n18680), .A(n18674), .ZN(n18685) );
  NAND2_X1 U21759 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18675), .ZN(
        n18684) );
  INV_X1 U21760 ( .A(n18676), .ZN(n18677) );
  OAI211_X1 U21761 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18678), .B(n18677), .ZN(
        n18683) );
  NOR2_X1 U21762 ( .A1(n18679), .A2(n18866), .ZN(n18681) );
  OAI211_X1 U21763 ( .C1(n18681), .C2(n18680), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18852), .ZN(n18682) );
  OAI211_X1 U21764 ( .C1(n18685), .C2(n18684), .A(n18683), .B(n18682), .ZN(
        n18686) );
  AOI21_X1 U21765 ( .B1(n18707), .B2(n18845), .A(n18686), .ZN(n18848) );
  INV_X1 U21766 ( .A(n18696), .ZN(n18718) );
  AOI22_X1 U21767 ( .A1(n18696), .A2(n18852), .B1(n18848), .B2(n18718), .ZN(
        n18700) );
  NOR2_X1 U21768 ( .A1(n18688), .A2(n18687), .ZN(n18691) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18689), .B1(
        n18691), .B2(n18866), .ZN(n18861) );
  OAI22_X1 U21770 ( .A1(n18691), .A2(n18853), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18690), .ZN(n18857) );
  AOI222_X1 U21771 ( .A1(n18861), .A2(n18857), .B1(n18861), .B2(n18693), .C1(
        n18857), .C2(n18692), .ZN(n18695) );
  OAI21_X1 U21772 ( .B1(n18696), .B2(n18695), .A(n18694), .ZN(n18697) );
  AOI222_X1 U21773 ( .A1(n18698), .A2(n18700), .B1(n18698), .B2(n18697), .C1(
        n18700), .C2(n18697), .ZN(n18699) );
  AOI211_X1 U21774 ( .C1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n18703), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n18699), .ZN(n18722) );
  INV_X1 U21775 ( .A(n18700), .ZN(n18705) );
  NAND2_X1 U21776 ( .A1(n18702), .A2(n18701), .ZN(n18704) );
  AOI21_X1 U21777 ( .B1(n18705), .B2(n18704), .A(n18703), .ZN(n18721) );
  NOR2_X1 U21778 ( .A1(n18707), .A2(n18706), .ZN(n18709) );
  OAI222_X1 U21779 ( .A1(n18713), .A2(n18712), .B1(n18711), .B2(n18710), .C1(
        n18709), .C2(n18708), .ZN(n18878) );
  AOI221_X1 U21780 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n18715), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n18715), .A(n18714), .ZN(n18716) );
  OAI211_X1 U21781 ( .C1(n18719), .C2(n18718), .A(n18717), .B(n18716), .ZN(
        n18720) );
  NOR4_X1 U21782 ( .A1(n18722), .A2(n18721), .A3(n18878), .A4(n18720), .ZN(
        n18733) );
  AOI22_X1 U21783 ( .A1(n18860), .A2(n18888), .B1(n18751), .B2(n18881), .ZN(
        n18730) );
  OAI211_X1 U21784 ( .C1(n18725), .C2(n18724), .A(n18723), .B(n18733), .ZN(
        n18832) );
  NAND2_X1 U21785 ( .A1(n18726), .A2(n18844), .ZN(n18728) );
  NAND2_X1 U21786 ( .A1(n18751), .A2(n18727), .ZN(n18734) );
  NAND4_X1 U21787 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18832), .A3(n18728), 
        .A4(n18734), .ZN(n18738) );
  OAI22_X1 U21788 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18730), .B1(n18729), 
        .B2(n18738), .ZN(n18731) );
  OAI21_X1 U21789 ( .B1(n18733), .B2(n18732), .A(n18731), .ZN(P3_U2996) );
  NOR3_X1 U21790 ( .A1(n18844), .A2(n18735), .A3(n18734), .ZN(n18740) );
  AOI211_X1 U21791 ( .C1(n18751), .C2(n18881), .A(n18736), .B(n18740), .ZN(
        n18737) );
  OAI21_X1 U21792 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18738), .A(n18737), 
        .ZN(P3_U2997) );
  OAI21_X1 U21793 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18739), .ZN(n18741) );
  AOI21_X1 U21794 ( .B1(n18742), .B2(n18741), .A(n18740), .ZN(P3_U2998) );
  INV_X1 U21795 ( .A(n18830), .ZN(n18743) );
  AND2_X1 U21796 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18743), .ZN(
        P3_U2999) );
  AND2_X1 U21797 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18743), .ZN(
        P3_U3000) );
  AND2_X1 U21798 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18743), .ZN(
        P3_U3001) );
  AND2_X1 U21799 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18743), .ZN(
        P3_U3002) );
  AND2_X1 U21800 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18743), .ZN(
        P3_U3003) );
  AND2_X1 U21801 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18743), .ZN(
        P3_U3004) );
  AND2_X1 U21802 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18743), .ZN(
        P3_U3005) );
  AND2_X1 U21803 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18743), .ZN(
        P3_U3006) );
  AND2_X1 U21804 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18743), .ZN(
        P3_U3007) );
  AND2_X1 U21805 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18743), .ZN(
        P3_U3008) );
  AND2_X1 U21806 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18743), .ZN(
        P3_U3009) );
  AND2_X1 U21807 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18743), .ZN(
        P3_U3010) );
  AND2_X1 U21808 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18743), .ZN(
        P3_U3011) );
  AND2_X1 U21809 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18743), .ZN(
        P3_U3012) );
  AND2_X1 U21810 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18743), .ZN(
        P3_U3013) );
  AND2_X1 U21811 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18743), .ZN(
        P3_U3014) );
  AND2_X1 U21812 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18743), .ZN(
        P3_U3015) );
  AND2_X1 U21813 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18743), .ZN(
        P3_U3016) );
  AND2_X1 U21814 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18743), .ZN(
        P3_U3017) );
  AND2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18743), .ZN(
        P3_U3018) );
  AND2_X1 U21816 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18743), .ZN(
        P3_U3019) );
  AND2_X1 U21817 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18743), .ZN(
        P3_U3020) );
  AND2_X1 U21818 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18743), .ZN(P3_U3021) );
  AND2_X1 U21819 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18743), .ZN(P3_U3022) );
  AND2_X1 U21820 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18743), .ZN(P3_U3023) );
  AND2_X1 U21821 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18743), .ZN(P3_U3024) );
  AND2_X1 U21822 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18743), .ZN(P3_U3025) );
  AND2_X1 U21823 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18743), .ZN(P3_U3026) );
  AND2_X1 U21824 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18743), .ZN(P3_U3027) );
  AND2_X1 U21825 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18743), .ZN(P3_U3028) );
  OAI21_X1 U21826 ( .B1(n18744), .B2(n20976), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18745) );
  AOI22_X1 U21827 ( .A1(n18758), .A2(n18760), .B1(n18894), .B2(n18745), .ZN(
        n18747) );
  INV_X1 U21828 ( .A(NA), .ZN(n20958) );
  OR3_X1 U21829 ( .A1(n20958), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18746) );
  OAI211_X1 U21830 ( .C1(n18885), .C2(n18748), .A(n18747), .B(n18746), .ZN(
        P3_U3029) );
  NOR2_X1 U21831 ( .A1(n18760), .A2(n20976), .ZN(n18756) );
  INV_X1 U21832 ( .A(n18756), .ZN(n18750) );
  INV_X1 U21833 ( .A(n18748), .ZN(n18749) );
  AOI22_X1 U21834 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18750), .B1(HOLD), 
        .B2(n18749), .ZN(n18752) );
  NAND2_X1 U21835 ( .A1(n18751), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18754) );
  OAI211_X1 U21836 ( .C1(n18752), .C2(n18758), .A(n18754), .B(n18882), .ZN(
        P3_U3030) );
  INV_X1 U21837 ( .A(n18754), .ZN(n18753) );
  AOI221_X1 U21838 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18758), .C1(n20958), 
        .C2(n18758), .A(n18753), .ZN(n18759) );
  OAI22_X1 U21839 ( .A1(NA), .A2(n18754), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18755) );
  OAI22_X1 U21840 ( .A1(n18756), .A2(n18755), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18757) );
  OAI22_X1 U21841 ( .A1(n18759), .A2(n18760), .B1(n18758), .B2(n18757), .ZN(
        P3_U3031) );
  OAI222_X1 U21842 ( .A1(n18868), .A2(n18822), .B1(n18761), .B2(n18893), .C1(
        n18762), .C2(n18810), .ZN(P3_U3032) );
  OAI222_X1 U21843 ( .A1(n18810), .A2(n18764), .B1(n18763), .B2(n18893), .C1(
        n18762), .C2(n18822), .ZN(P3_U3033) );
  OAI222_X1 U21844 ( .A1(n18810), .A2(n18766), .B1(n18765), .B2(n18893), .C1(
        n18764), .C2(n18822), .ZN(P3_U3034) );
  INV_X1 U21845 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18769) );
  OAI222_X1 U21846 ( .A1(n18810), .A2(n18769), .B1(n18767), .B2(n18893), .C1(
        n18766), .C2(n18822), .ZN(P3_U3035) );
  OAI222_X1 U21847 ( .A1(n18769), .A2(n18822), .B1(n18768), .B2(n18893), .C1(
        n18770), .C2(n18810), .ZN(P3_U3036) );
  OAI222_X1 U21848 ( .A1(n18810), .A2(n18772), .B1(n18771), .B2(n18893), .C1(
        n18770), .C2(n18822), .ZN(P3_U3037) );
  INV_X1 U21849 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18775) );
  OAI222_X1 U21850 ( .A1(n18810), .A2(n18775), .B1(n18773), .B2(n18893), .C1(
        n18772), .C2(n18822), .ZN(P3_U3038) );
  OAI222_X1 U21851 ( .A1(n18775), .A2(n18822), .B1(n18774), .B2(n18893), .C1(
        n18776), .C2(n18810), .ZN(P3_U3039) );
  OAI222_X1 U21852 ( .A1(n18810), .A2(n18778), .B1(n18777), .B2(n18893), .C1(
        n18776), .C2(n18822), .ZN(P3_U3040) );
  OAI222_X1 U21853 ( .A1(n18810), .A2(n18780), .B1(n18779), .B2(n18893), .C1(
        n18778), .C2(n18822), .ZN(P3_U3041) );
  OAI222_X1 U21854 ( .A1(n18810), .A2(n18782), .B1(n18781), .B2(n18893), .C1(
        n18780), .C2(n18822), .ZN(P3_U3042) );
  OAI222_X1 U21855 ( .A1(n18810), .A2(n18784), .B1(n18783), .B2(n18893), .C1(
        n18782), .C2(n18822), .ZN(P3_U3043) );
  OAI222_X1 U21856 ( .A1(n18810), .A2(n18787), .B1(n18785), .B2(n18893), .C1(
        n18784), .C2(n18822), .ZN(P3_U3044) );
  OAI222_X1 U21857 ( .A1(n18787), .A2(n18822), .B1(n18786), .B2(n18893), .C1(
        n18788), .C2(n18810), .ZN(P3_U3045) );
  OAI222_X1 U21858 ( .A1(n18810), .A2(n18790), .B1(n18789), .B2(n18893), .C1(
        n18788), .C2(n18822), .ZN(P3_U3046) );
  OAI222_X1 U21859 ( .A1(n18810), .A2(n18792), .B1(n18791), .B2(n18893), .C1(
        n18790), .C2(n18822), .ZN(P3_U3047) );
  OAI222_X1 U21860 ( .A1(n18810), .A2(n18794), .B1(n18793), .B2(n18893), .C1(
        n18792), .C2(n18822), .ZN(P3_U3048) );
  OAI222_X1 U21861 ( .A1(n18810), .A2(n18796), .B1(n18795), .B2(n18893), .C1(
        n18794), .C2(n18822), .ZN(P3_U3049) );
  INV_X1 U21862 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18799) );
  OAI222_X1 U21863 ( .A1(n18810), .A2(n18799), .B1(n18797), .B2(n18893), .C1(
        n18796), .C2(n18822), .ZN(P3_U3050) );
  INV_X1 U21864 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18800) );
  OAI222_X1 U21865 ( .A1(n18799), .A2(n18822), .B1(n18798), .B2(n18893), .C1(
        n18800), .C2(n18810), .ZN(P3_U3051) );
  OAI222_X1 U21866 ( .A1(n18810), .A2(n18802), .B1(n18801), .B2(n18893), .C1(
        n18800), .C2(n18822), .ZN(P3_U3052) );
  OAI222_X1 U21867 ( .A1(n18810), .A2(n18805), .B1(n18803), .B2(n18893), .C1(
        n18802), .C2(n18822), .ZN(P3_U3053) );
  INV_X1 U21868 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18807) );
  OAI222_X1 U21869 ( .A1(n18805), .A2(n18822), .B1(n18804), .B2(n18893), .C1(
        n18807), .C2(n18810), .ZN(P3_U3054) );
  OAI222_X1 U21870 ( .A1(n18807), .A2(n18822), .B1(n18806), .B2(n18893), .C1(
        n18808), .C2(n18810), .ZN(P3_U3055) );
  OAI222_X1 U21871 ( .A1(n18810), .A2(n18811), .B1(n18809), .B2(n18893), .C1(
        n18808), .C2(n18822), .ZN(P3_U3056) );
  OAI222_X1 U21872 ( .A1(n18810), .A2(n18813), .B1(n18812), .B2(n18893), .C1(
        n18811), .C2(n18822), .ZN(P3_U3057) );
  OAI222_X1 U21873 ( .A1(n18810), .A2(n18816), .B1(n18814), .B2(n18893), .C1(
        n18813), .C2(n18822), .ZN(P3_U3058) );
  INV_X1 U21874 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18817) );
  OAI222_X1 U21875 ( .A1(n18816), .A2(n18822), .B1(n18815), .B2(n18893), .C1(
        n18817), .C2(n18810), .ZN(P3_U3059) );
  OAI222_X1 U21876 ( .A1(n18810), .A2(n18821), .B1(n18818), .B2(n18893), .C1(
        n18817), .C2(n18822), .ZN(P3_U3060) );
  INV_X1 U21877 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18820) );
  OAI222_X1 U21878 ( .A1(n18822), .A2(n18821), .B1(n18820), .B2(n18893), .C1(
        n18819), .C2(n18810), .ZN(P3_U3061) );
  OAI22_X1 U21879 ( .A1(n18894), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18893), .ZN(n18823) );
  INV_X1 U21880 ( .A(n18823), .ZN(P3_U3274) );
  OAI22_X1 U21881 ( .A1(n18894), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18893), .ZN(n18824) );
  INV_X1 U21882 ( .A(n18824), .ZN(P3_U3275) );
  OAI22_X1 U21883 ( .A1(n18894), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18893), .ZN(n18825) );
  INV_X1 U21884 ( .A(n18825), .ZN(P3_U3276) );
  OAI22_X1 U21885 ( .A1(n18894), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18893), .ZN(n18826) );
  INV_X1 U21886 ( .A(n18826), .ZN(P3_U3277) );
  OAI21_X1 U21887 ( .B1(n18830), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18828), 
        .ZN(n18827) );
  INV_X1 U21888 ( .A(n18827), .ZN(P3_U3280) );
  OAI21_X1 U21889 ( .B1(n18830), .B2(n18829), .A(n18828), .ZN(P3_U3281) );
  OAI221_X1 U21890 ( .B1(n18833), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18833), 
        .C2(n18832), .A(n18831), .ZN(P3_U3282) );
  NOR2_X1 U21891 ( .A1(n18834), .A2(n18847), .ZN(n18835) );
  NOR2_X1 U21892 ( .A1(n18835), .A2(n18867), .ZN(n18840) );
  NOR3_X1 U21893 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18836), .A3(
        n18847), .ZN(n18837) );
  AOI21_X1 U21894 ( .B1(n18838), .B2(n18860), .A(n18837), .ZN(n18839) );
  OAI22_X1 U21895 ( .A1(n18841), .A2(n18840), .B1(n18867), .B2(n18839), .ZN(
        P3_U3285) );
  OAI22_X1 U21896 ( .A1(n18843), .A2(n18842), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18855) );
  INV_X1 U21897 ( .A(n18855), .ZN(n18850) );
  NOR2_X1 U21898 ( .A1(n18844), .A2(n18863), .ZN(n18854) );
  OAI22_X1 U21899 ( .A1(n18848), .A2(n18847), .B1(n18846), .B2(n18845), .ZN(
        n18849) );
  AOI21_X1 U21900 ( .B1(n18850), .B2(n18854), .A(n18849), .ZN(n18851) );
  AOI22_X1 U21901 ( .A1(n18867), .A2(n18852), .B1(n18851), .B2(n18864), .ZN(
        P3_U3288) );
  INV_X1 U21902 ( .A(n18853), .ZN(n18856) );
  AOI222_X1 U21903 ( .A1(n18857), .A2(n18862), .B1(n18860), .B2(n18856), .C1(
        n18855), .C2(n18854), .ZN(n18858) );
  AOI22_X1 U21904 ( .A1(n18867), .A2(n18859), .B1(n18858), .B2(n18864), .ZN(
        P3_U3289) );
  AOI222_X1 U21905 ( .A1(n18863), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18862), 
        .B2(n18861), .C1(n18866), .C2(n18860), .ZN(n18865) );
  AOI22_X1 U21906 ( .A1(n18867), .A2(n18866), .B1(n18865), .B2(n18864), .ZN(
        P3_U3290) );
  AOI21_X1 U21907 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18869) );
  AOI22_X1 U21908 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18869), .B2(n18868), .ZN(n18872) );
  INV_X1 U21909 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18871) );
  AOI22_X1 U21910 ( .A1(n18875), .A2(n18872), .B1(n18871), .B2(n18870), .ZN(
        P3_U3292) );
  INV_X1 U21911 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18874) );
  OAI21_X1 U21912 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18875), .ZN(n18873) );
  OAI21_X1 U21913 ( .B1(n18875), .B2(n18874), .A(n18873), .ZN(P3_U3293) );
  INV_X1 U21914 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18900) );
  OAI22_X1 U21915 ( .A1(n18894), .A2(n18900), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18893), .ZN(n18876) );
  INV_X1 U21916 ( .A(n18876), .ZN(P3_U3294) );
  MUX2_X1 U21917 ( .A(P3_MORE_REG_SCAN_IN), .B(n18878), .S(n18877), .Z(
        P3_U3295) );
  AOI21_X1 U21918 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_0__SCAN_IN), .A(n18879), .ZN(n18880) );
  AOI211_X1 U21919 ( .C1(n18881), .C2(n18885), .A(n18880), .B(n18899), .ZN(
        n18892) );
  AOI21_X1 U21920 ( .B1(n18884), .B2(n18883), .A(n18882), .ZN(n18886) );
  OAI211_X1 U21921 ( .C1(n18887), .C2(n18886), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18885), .ZN(n18889) );
  AOI21_X1 U21922 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18889), .A(n18888), 
        .ZN(n18891) );
  NAND2_X1 U21923 ( .A1(n18892), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18890) );
  OAI21_X1 U21924 ( .B1(n18892), .B2(n18891), .A(n18890), .ZN(P3_U3296) );
  OAI22_X1 U21925 ( .A1(n18894), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18893), .ZN(n18895) );
  INV_X1 U21926 ( .A(n18895), .ZN(P3_U3297) );
  INV_X1 U21927 ( .A(n18896), .ZN(n18897) );
  NOR2_X1 U21928 ( .A1(n18897), .A2(n18899), .ZN(n18903) );
  AOI22_X1 U21929 ( .A1(n18903), .A2(n18900), .B1(n18899), .B2(n18898), .ZN(
        P3_U3298) );
  INV_X1 U21930 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18902) );
  AOI21_X1 U21931 ( .B1(n18903), .B2(n18902), .A(n18901), .ZN(P3_U3299) );
  NAND2_X1 U21932 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19869), .ZN(n19862) );
  NAND2_X1 U21933 ( .A1(n19858), .A2(n18904), .ZN(n19859) );
  OAI21_X1 U21934 ( .B1(n19858), .B2(n19862), .A(n19859), .ZN(n19931) );
  AOI21_X1 U21935 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19931), .ZN(n18905) );
  INV_X1 U21936 ( .A(n18905), .ZN(P2_U2815) );
  INV_X1 U21937 ( .A(n18906), .ZN(n19982) );
  AOI22_X1 U21938 ( .A1(n19982), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19933), 
        .B2(n19849), .ZN(n18907) );
  INV_X1 U21939 ( .A(n18907), .ZN(P2_U2816) );
  AOI21_X1 U21940 ( .B1(n19858), .B2(n19869), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18908) );
  AOI22_X1 U21941 ( .A1(n19880), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18908), 
        .B2(n19998), .ZN(P2_U2817) );
  INV_X1 U21942 ( .A(BS16), .ZN(n20955) );
  AOI21_X1 U21943 ( .B1(n19863), .B2(n20955), .A(n19928), .ZN(n19926) );
  INV_X1 U21944 ( .A(n19926), .ZN(n19929) );
  OAI21_X1 U21945 ( .B1(n19931), .B2(n19989), .A(n19929), .ZN(P2_U2818) );
  NOR4_X1 U21946 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18912) );
  NOR4_X1 U21947 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18911) );
  NOR4_X1 U21948 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18910) );
  NOR4_X1 U21949 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18909) );
  NAND4_X1 U21950 ( .A1(n18912), .A2(n18911), .A3(n18910), .A4(n18909), .ZN(
        n18918) );
  NOR4_X1 U21951 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18916) );
  AOI211_X1 U21952 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18915) );
  NOR4_X1 U21953 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18914) );
  NOR4_X1 U21954 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18913) );
  NAND4_X1 U21955 ( .A1(n18916), .A2(n18915), .A3(n18914), .A4(n18913), .ZN(
        n18917) );
  NOR2_X1 U21956 ( .A1(n18918), .A2(n18917), .ZN(n18929) );
  INV_X1 U21957 ( .A(n18929), .ZN(n18927) );
  NOR2_X1 U21958 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18927), .ZN(n18921) );
  INV_X1 U21959 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18919) );
  AOI22_X1 U21960 ( .A1(n18921), .A2(n18922), .B1(n18927), .B2(n18919), .ZN(
        P2_U2820) );
  INV_X1 U21961 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19930) );
  INV_X1 U21962 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19927) );
  NAND3_X1 U21963 ( .A1(n18922), .A2(n19930), .A3(n19927), .ZN(n18926) );
  INV_X1 U21964 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18920) );
  AOI22_X1 U21965 ( .A1(n18921), .A2(n18926), .B1(n18927), .B2(n18920), .ZN(
        P2_U2821) );
  NAND2_X1 U21966 ( .A1(n18921), .A2(n19930), .ZN(n18925) );
  OAI21_X1 U21967 ( .B1(n19870), .B2(n18922), .A(n18929), .ZN(n18923) );
  OAI21_X1 U21968 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18929), .A(n18923), 
        .ZN(n18924) );
  OAI221_X1 U21969 ( .B1(n18925), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18925), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18924), .ZN(P2_U2822) );
  INV_X1 U21970 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18928) );
  OAI221_X1 U21971 ( .B1(n18929), .B2(n18928), .C1(n18927), .C2(n18926), .A(
        n18925), .ZN(P2_U2823) );
  OAI22_X1 U21972 ( .A1(n18931), .A2(n19107), .B1(n19098), .B2(n18930), .ZN(
        n18932) );
  INV_X1 U21973 ( .A(n18932), .ZN(n18941) );
  AOI211_X1 U21974 ( .C1(n18935), .C2(n18934), .A(n18933), .B(n19851), .ZN(
        n18939) );
  AOI22_X1 U21975 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19096), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19102), .ZN(n18936) );
  OAI21_X1 U21976 ( .B1(n18937), .B2(n19099), .A(n18936), .ZN(n18938) );
  AOI211_X1 U21977 ( .C1(n19095), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n18939), .B(n18938), .ZN(n18940) );
  NAND2_X1 U21978 ( .A1(n18941), .A2(n18940), .ZN(P2_U2835) );
  OAI22_X1 U21979 ( .A1(n18943), .A2(n19107), .B1(n19098), .B2(n18942), .ZN(
        n18944) );
  INV_X1 U21980 ( .A(n18944), .ZN(n18952) );
  AOI211_X1 U21981 ( .C1(n18946), .C2(n9769), .A(n18945), .B(n19851), .ZN(
        n18950) );
  AOI22_X1 U21982 ( .A1(n18947), .A2(n19056), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19095), .ZN(n18948) );
  OAI211_X1 U21983 ( .C1(n19899), .C2(n19067), .A(n18948), .B(n19066), .ZN(
        n18949) );
  AOI211_X1 U21984 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19096), .A(n18950), .B(
        n18949), .ZN(n18951) );
  NAND2_X1 U21985 ( .A1(n18952), .A2(n18951), .ZN(P2_U2836) );
  OAI22_X1 U21986 ( .A1(n18954), .A2(n19107), .B1(n19098), .B2(n18953), .ZN(
        n18955) );
  INV_X1 U21987 ( .A(n18955), .ZN(n18964) );
  AOI211_X1 U21988 ( .C1(n18958), .C2(n18957), .A(n18956), .B(n19851), .ZN(
        n18962) );
  AOI22_X1 U21989 ( .A1(n18959), .A2(n19056), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19096), .ZN(n18960) );
  OAI211_X1 U21990 ( .C1(n11972), .C2(n19067), .A(n18960), .B(n19066), .ZN(
        n18961) );
  AOI211_X1 U21991 ( .C1(n19095), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n18962), .B(n18961), .ZN(n18963) );
  NAND2_X1 U21992 ( .A1(n18964), .A2(n18963), .ZN(P2_U2837) );
  NOR2_X1 U21993 ( .A1(n19021), .A2(n18965), .ZN(n18967) );
  XOR2_X1 U21994 ( .A(n18967), .B(n18966), .Z(n18977) );
  OAI21_X1 U21995 ( .B1(n19896), .B2(n19067), .A(n19066), .ZN(n18971) );
  OAI22_X1 U21996 ( .A1(n18969), .A2(n19099), .B1(n19093), .B2(n18968), .ZN(
        n18970) );
  AOI211_X1 U21997 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19096), .A(n18971), .B(
        n18970), .ZN(n18976) );
  AOI22_X1 U21998 ( .A1(n18974), .A2(n19076), .B1(n18973), .B2(n18972), .ZN(
        n18975) );
  OAI211_X1 U21999 ( .C1(n19851), .C2(n18977), .A(n18976), .B(n18975), .ZN(
        P2_U2838) );
  OAI22_X1 U22000 ( .A1(n18979), .A2(n19099), .B1(n18978), .B2(n19093), .ZN(
        n18980) );
  AOI211_X1 U22001 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19102), .A(n12657), 
        .B(n18980), .ZN(n18987) );
  NAND2_X1 U22002 ( .A1(n9634), .A2(n18994), .ZN(n18981) );
  XOR2_X1 U22003 ( .A(n18982), .B(n18981), .Z(n18985) );
  OAI22_X1 U22004 ( .A1(n19120), .A2(n19107), .B1(n19098), .B2(n18983), .ZN(
        n18984) );
  AOI21_X1 U22005 ( .B1(n19089), .B2(n18985), .A(n18984), .ZN(n18986) );
  OAI211_X1 U22006 ( .C1(n19082), .C2(n14163), .A(n18987), .B(n18986), .ZN(
        P2_U2839) );
  AOI22_X1 U22007 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19095), .B1(
        P2_EBX_REG_15__SCAN_IN), .B2(n19096), .ZN(n18988) );
  OAI211_X1 U22008 ( .C1(n19067), .C2(n19892), .A(n18988), .B(n19066), .ZN(
        n18989) );
  AOI21_X1 U22009 ( .B1(n18990), .B2(n19076), .A(n18989), .ZN(n18991) );
  OAI21_X1 U22010 ( .B1(n18992), .B2(n19099), .A(n18991), .ZN(n18993) );
  AOI21_X1 U22011 ( .B1(n19009), .B2(n16169), .A(n18993), .ZN(n18999) );
  OAI211_X1 U22012 ( .C1(n18997), .C2(n18996), .A(n18995), .B(n18994), .ZN(
        n18998) );
  OAI211_X1 U22013 ( .C1(n19098), .C2(n19000), .A(n18999), .B(n18998), .ZN(
        P2_U2840) );
  INV_X1 U22014 ( .A(n19001), .ZN(n19004) );
  AOI22_X1 U22015 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n19096), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19095), .ZN(n19002) );
  OAI211_X1 U22016 ( .C1(n19067), .C2(n15297), .A(n19002), .B(n19066), .ZN(
        n19003) );
  AOI21_X1 U22017 ( .B1(n19004), .B2(n19076), .A(n19003), .ZN(n19005) );
  OAI21_X1 U22018 ( .B1(n19006), .B2(n19099), .A(n19005), .ZN(n19007) );
  AOI21_X1 U22019 ( .B1(n19009), .B2(n19008), .A(n19007), .ZN(n19015) );
  INV_X1 U22020 ( .A(n19010), .ZN(n19011) );
  OAI211_X1 U22021 ( .C1(n19013), .C2(n19012), .A(n19089), .B(n19011), .ZN(
        n19014) );
  OAI211_X1 U22022 ( .C1(n19098), .C2(n19016), .A(n19015), .B(n19014), .ZN(
        P2_U2842) );
  OAI22_X1 U22023 ( .A1(n19018), .A2(n19099), .B1(n19093), .B2(n19017), .ZN(
        n19019) );
  AOI211_X1 U22024 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19102), .A(n12657), 
        .B(n19019), .ZN(n19030) );
  NOR2_X1 U22025 ( .A1(n19021), .A2(n19020), .ZN(n19022) );
  XOR2_X1 U22026 ( .A(n19023), .B(n19022), .Z(n19028) );
  INV_X1 U22027 ( .A(n19024), .ZN(n19026) );
  OAI22_X1 U22028 ( .A1(n19026), .A2(n19107), .B1(n19098), .B2(n19025), .ZN(
        n19027) );
  AOI21_X1 U22029 ( .B1(n19028), .B2(n19089), .A(n19027), .ZN(n19029) );
  OAI211_X1 U22030 ( .C1(n19082), .C2(n19031), .A(n19030), .B(n19029), .ZN(
        P2_U2844) );
  NAND2_X1 U22031 ( .A1(n9634), .A2(n19032), .ZN(n19034) );
  XOR2_X1 U22032 ( .A(n19034), .B(n19033), .Z(n19042) );
  INV_X1 U22033 ( .A(n19035), .ZN(n19036) );
  AOI22_X1 U22034 ( .A1(n19036), .A2(n19056), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19096), .ZN(n19037) );
  OAI211_X1 U22035 ( .C1(n19886), .C2(n19067), .A(n19037), .B(n19066), .ZN(
        n19040) );
  OAI22_X1 U22036 ( .A1(n19162), .A2(n19098), .B1(n19107), .B2(n19038), .ZN(
        n19039) );
  AOI211_X1 U22037 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19095), .A(
        n19040), .B(n19039), .ZN(n19041) );
  OAI21_X1 U22038 ( .B1(n19042), .B2(n19851), .A(n19041), .ZN(P2_U2845) );
  OAI22_X1 U22039 ( .A1(n19043), .A2(n19099), .B1(n19082), .B2(n12644), .ZN(
        n19044) );
  AOI211_X1 U22040 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19102), .A(n12657), .B(
        n19044), .ZN(n19052) );
  NOR2_X1 U22041 ( .A1(n19021), .A2(n19045), .ZN(n19046) );
  XNOR2_X1 U22042 ( .A(n19047), .B(n19046), .ZN(n19050) );
  OAI22_X1 U22043 ( .A1(n19165), .A2(n19098), .B1(n19107), .B2(n19048), .ZN(
        n19049) );
  AOI21_X1 U22044 ( .B1(n19050), .B2(n19089), .A(n19049), .ZN(n19051) );
  OAI211_X1 U22045 ( .C1(n12587), .C2(n19093), .A(n19052), .B(n19051), .ZN(
        P2_U2846) );
  NOR2_X1 U22046 ( .A1(n19021), .A2(n19053), .ZN(n19054) );
  XOR2_X1 U22047 ( .A(n19055), .B(n19054), .Z(n19065) );
  AOI22_X1 U22048 ( .A1(n19057), .A2(n19056), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19096), .ZN(n19058) );
  OAI211_X1 U22049 ( .C1(n19879), .C2(n19067), .A(n19058), .B(n19066), .ZN(
        n19063) );
  INV_X1 U22050 ( .A(n19059), .ZN(n19061) );
  OAI22_X1 U22051 ( .A1(n19061), .A2(n19107), .B1(n19098), .B2(n19060), .ZN(
        n19062) );
  AOI211_X1 U22052 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19095), .A(
        n19063), .B(n19062), .ZN(n19064) );
  OAI21_X1 U22053 ( .B1(n19851), .B2(n19065), .A(n19064), .ZN(P2_U2848) );
  OAI21_X1 U22054 ( .B1(n19877), .B2(n19067), .A(n19066), .ZN(n19071) );
  OAI22_X1 U22055 ( .A1(n19069), .A2(n19099), .B1(n19093), .B2(n19068), .ZN(
        n19070) );
  AOI211_X1 U22056 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19096), .A(n19071), .B(
        n19070), .ZN(n19079) );
  NAND2_X1 U22057 ( .A1(n9634), .A2(n19072), .ZN(n19073) );
  XNOR2_X1 U22058 ( .A(n19074), .B(n19073), .ZN(n19077) );
  AOI22_X1 U22059 ( .A1(n19077), .A2(n19089), .B1(n19076), .B2(n19075), .ZN(
        n19078) );
  OAI211_X1 U22060 ( .C1(n19098), .C2(n19080), .A(n19079), .B(n19078), .ZN(
        P2_U2849) );
  OAI22_X1 U22061 ( .A1(n19082), .A2(n12642), .B1(n19081), .B2(n19099), .ZN(
        n19083) );
  AOI211_X1 U22062 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19102), .A(n12657), .B(
        n19083), .ZN(n19092) );
  NOR2_X1 U22063 ( .A1(n19021), .A2(n19084), .ZN(n19085) );
  XNOR2_X1 U22064 ( .A(n19086), .B(n19085), .ZN(n19090) );
  OAI22_X1 U22065 ( .A1(n19087), .A2(n19107), .B1(n19178), .B2(n19098), .ZN(
        n19088) );
  AOI21_X1 U22066 ( .B1(n19090), .B2(n19089), .A(n19088), .ZN(n19091) );
  OAI211_X1 U22067 ( .C1(n19094), .C2(n19093), .A(n19092), .B(n19091), .ZN(
        P2_U2850) );
  AOI22_X1 U22068 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19096), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19095), .ZN(n19117) );
  OAI22_X1 U22069 ( .A1(n19100), .A2(n19099), .B1(n19098), .B2(n19097), .ZN(
        n19101) );
  AOI211_X1 U22070 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19102), .A(n12657), .B(
        n19101), .ZN(n19116) );
  OR2_X1 U22071 ( .A1(n19104), .A2(n19103), .ZN(n19106) );
  NAND2_X1 U22072 ( .A1(n19106), .A2(n19105), .ZN(n19232) );
  OAI22_X1 U22073 ( .A1(n19172), .A2(n19108), .B1(n19107), .B2(n19232), .ZN(
        n19109) );
  INV_X1 U22074 ( .A(n19109), .ZN(n19115) );
  AND2_X1 U22075 ( .A1(n9634), .A2(n19110), .ZN(n19113) );
  AOI21_X1 U22076 ( .B1(n19215), .B2(n19113), .A(n19851), .ZN(n19112) );
  OAI21_X1 U22077 ( .B1(n19215), .B2(n19113), .A(n19112), .ZN(n19114) );
  NAND4_X1 U22078 ( .A1(n19117), .A2(n19116), .A3(n19115), .A4(n19114), .ZN(
        P2_U2851) );
  AOI22_X1 U22079 ( .A1(n19118), .A2(n19127), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n12991), .ZN(n19119) );
  OAI21_X1 U22080 ( .B1(n12991), .B2(n19120), .A(n19119), .ZN(P2_U2871) );
  XNOR2_X1 U22081 ( .A(n13477), .B(n19121), .ZN(n19122) );
  AOI22_X1 U22082 ( .A1(n19122), .A2(n19127), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n12991), .ZN(n19123) );
  OAI21_X1 U22083 ( .B1(n19124), .B2(n12991), .A(n19123), .ZN(P2_U2873) );
  XNOR2_X1 U22084 ( .A(n13469), .B(n19125), .ZN(n19128) );
  AOI22_X1 U22085 ( .A1(n19128), .A2(n19127), .B1(n19148), .B2(n19126), .ZN(
        n19129) );
  OAI21_X1 U22086 ( .B1(n19148), .B2(n19130), .A(n19129), .ZN(P2_U2875) );
  INV_X1 U22087 ( .A(n13467), .ZN(n19131) );
  NOR2_X1 U22088 ( .A1(n19131), .A2(n19145), .ZN(n19136) );
  OAI21_X1 U22089 ( .B1(n13256), .B2(n19133), .A(n19132), .ZN(n19135) );
  AOI22_X1 U22090 ( .A1(n19136), .A2(n19135), .B1(n19148), .B2(n19134), .ZN(
        n19137) );
  OAI21_X1 U22091 ( .B1(n19148), .B2(n19138), .A(n19137), .ZN(P2_U2877) );
  INV_X1 U22092 ( .A(n19139), .ZN(n19141) );
  AOI21_X1 U22093 ( .B1(n19141), .B2(n19140), .A(n19145), .ZN(n19142) );
  AOI22_X1 U22094 ( .A1(n19142), .A2(n13256), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n12991), .ZN(n19143) );
  OAI21_X1 U22095 ( .B1(n19144), .B2(n12991), .A(n19143), .ZN(P2_U2879) );
  OAI22_X1 U22096 ( .A1(n19172), .A2(n19145), .B1(n12991), .B2(n19232), .ZN(
        n19146) );
  INV_X1 U22097 ( .A(n19146), .ZN(n19147) );
  OAI21_X1 U22098 ( .B1(n19148), .B2(n12640), .A(n19147), .ZN(P2_U2883) );
  INV_X1 U22099 ( .A(n19149), .ZN(n19151) );
  AOI22_X1 U22100 ( .A1(n19152), .A2(BUF2_REG_31__SCAN_IN), .B1(n19151), .B2(
        n19150), .ZN(n19155) );
  AOI22_X1 U22101 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19169), .B1(n19153), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19154) );
  NAND2_X1 U22102 ( .A1(n19155), .A2(n19154), .ZN(P2_U2888) );
  INV_X1 U22103 ( .A(n19156), .ZN(n19159) );
  AOI22_X1 U22104 ( .A1(n19171), .A2(n19157), .B1(n19169), .B2(
        P2_EAX_REG_12__SCAN_IN), .ZN(n19158) );
  OAI21_X1 U22105 ( .B1(n19179), .B2(n19159), .A(n19158), .ZN(P2_U2907) );
  AOI22_X1 U22106 ( .A1(n19171), .A2(n19160), .B1(n19169), .B2(
        P2_EAX_REG_10__SCAN_IN), .ZN(n19161) );
  OAI21_X1 U22107 ( .B1(n19179), .B2(n19162), .A(n19161), .ZN(P2_U2909) );
  AOI22_X1 U22108 ( .A1(n19171), .A2(n19163), .B1(n19169), .B2(
        P2_EAX_REG_9__SCAN_IN), .ZN(n19164) );
  OAI21_X1 U22109 ( .B1(n19179), .B2(n19165), .A(n19164), .ZN(P2_U2910) );
  AOI22_X1 U22110 ( .A1(n19171), .A2(n19166), .B1(n19169), .B2(
        P2_EAX_REG_8__SCAN_IN), .ZN(n19167) );
  OAI21_X1 U22111 ( .B1(n19179), .B2(n19168), .A(n19167), .ZN(P2_U2911) );
  AOI22_X1 U22112 ( .A1(n19171), .A2(n19170), .B1(n19169), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n19177) );
  INV_X1 U22113 ( .A(n19172), .ZN(n19174) );
  NAND3_X1 U22114 ( .A1(n19175), .A2(n19174), .A3(n19173), .ZN(n19176) );
  OAI211_X1 U22115 ( .C1(n19179), .C2(n19178), .A(n19177), .B(n19176), .ZN(
        P2_U2914) );
  AND2_X1 U22116 ( .A1(n19198), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22117 ( .A1(n19212), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19181) );
  OAI21_X1 U22118 ( .B1(n12732), .B2(n19214), .A(n19181), .ZN(P2_U2936) );
  AOI22_X1 U22119 ( .A1(n19212), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19182) );
  OAI21_X1 U22120 ( .B1(n19183), .B2(n19214), .A(n19182), .ZN(P2_U2937) );
  AOI22_X1 U22121 ( .A1(n19212), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19184) );
  OAI21_X1 U22122 ( .B1(n19185), .B2(n19214), .A(n19184), .ZN(P2_U2938) );
  AOI22_X1 U22123 ( .A1(n19212), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19186) );
  OAI21_X1 U22124 ( .B1(n19187), .B2(n19214), .A(n19186), .ZN(P2_U2939) );
  AOI22_X1 U22125 ( .A1(n19212), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19198), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19188) );
  OAI21_X1 U22126 ( .B1(n19189), .B2(n19214), .A(n19188), .ZN(P2_U2940) );
  AOI22_X1 U22127 ( .A1(n19212), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19198), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19190) );
  OAI21_X1 U22128 ( .B1(n19191), .B2(n19214), .A(n19190), .ZN(P2_U2941) );
  AOI22_X1 U22129 ( .A1(n19212), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19198), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19192) );
  OAI21_X1 U22130 ( .B1(n19193), .B2(n19214), .A(n19192), .ZN(P2_U2942) );
  AOI22_X1 U22131 ( .A1(n19212), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19198), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U22132 ( .B1(n19195), .B2(n19214), .A(n19194), .ZN(P2_U2943) );
  AOI22_X1 U22133 ( .A1(n19212), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19198), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19196) );
  OAI21_X1 U22134 ( .B1(n19197), .B2(n19214), .A(n19196), .ZN(P2_U2944) );
  AOI22_X1 U22135 ( .A1(n19212), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19198), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19199) );
  OAI21_X1 U22136 ( .B1(n19200), .B2(n19214), .A(n19199), .ZN(P2_U2945) );
  INV_X1 U22137 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19202) );
  AOI22_X1 U22138 ( .A1(n19212), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19201) );
  OAI21_X1 U22139 ( .B1(n19202), .B2(n19214), .A(n19201), .ZN(P2_U2946) );
  INV_X1 U22140 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19204) );
  AOI22_X1 U22141 ( .A1(n19212), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19203) );
  OAI21_X1 U22142 ( .B1(n19204), .B2(n19214), .A(n19203), .ZN(P2_U2947) );
  INV_X1 U22143 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19206) );
  AOI22_X1 U22144 ( .A1(n19212), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19205) );
  OAI21_X1 U22145 ( .B1(n19206), .B2(n19214), .A(n19205), .ZN(P2_U2948) );
  INV_X1 U22146 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19208) );
  AOI22_X1 U22147 ( .A1(n19212), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22148 ( .B1(n19208), .B2(n19214), .A(n19207), .ZN(P2_U2949) );
  AOI22_X1 U22149 ( .A1(n19212), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U22150 ( .B1(n19210), .B2(n19214), .A(n19209), .ZN(P2_U2950) );
  AOI22_X1 U22151 ( .A1(n19212), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U22152 ( .B1(n12100), .B2(n19214), .A(n19213), .ZN(P2_U2951) );
  AOI22_X1 U22153 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n15785), .B1(n19216), 
        .B2(n19215), .ZN(n19229) );
  INV_X1 U22154 ( .A(n19217), .ZN(n19218) );
  NOR2_X1 U22155 ( .A1(n19219), .A2(n19218), .ZN(n19220) );
  XNOR2_X1 U22156 ( .A(n19220), .B(n19234), .ZN(n19239) );
  XOR2_X1 U22157 ( .A(n19221), .B(n19222), .Z(n19238) );
  INV_X1 U22158 ( .A(n19238), .ZN(n19225) );
  OAI22_X1 U22159 ( .A1(n19225), .A2(n19224), .B1(n19223), .B2(n19232), .ZN(
        n19226) );
  AOI21_X1 U22160 ( .B1(n19227), .B2(n19239), .A(n19226), .ZN(n19228) );
  OAI211_X1 U22161 ( .C1(n19231), .C2(n19230), .A(n19229), .B(n19228), .ZN(
        P2_U3010) );
  INV_X1 U22162 ( .A(n19232), .ZN(n19233) );
  AOI22_X1 U22163 ( .A1(n19235), .A2(n19234), .B1(n19233), .B2(n19248), .ZN(
        n19243) );
  AOI22_X1 U22164 ( .A1(n19237), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19262), .B2(n19236), .ZN(n19242) );
  AOI22_X1 U22165 ( .A1(n19239), .A2(n19250), .B1(n19255), .B2(n19238), .ZN(
        n19241) );
  NAND2_X1 U22166 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n12657), .ZN(n19240) );
  NAND4_X1 U22167 ( .A1(n19243), .A2(n19242), .A3(n19241), .A4(n19240), .ZN(
        P2_U3042) );
  AOI221_X1 U22168 ( .B1(n19253), .B2(n19246), .C1(n19245), .C2(n19252), .A(
        n19244), .ZN(n19266) );
  AOI21_X1 U22169 ( .B1(n19248), .B2(n12843), .A(n19247), .ZN(n19260) );
  AOI21_X1 U22170 ( .B1(n19251), .B2(n19250), .A(n19249), .ZN(n19259) );
  NAND3_X1 U22171 ( .A1(n19253), .A2(n19252), .A3(n19265), .ZN(n19258) );
  NAND3_X1 U22172 ( .A1(n19256), .A2(n19255), .A3(n19254), .ZN(n19257) );
  NAND4_X1 U22173 ( .A1(n19260), .A2(n19259), .A3(n19258), .A4(n19257), .ZN(
        n19261) );
  AOI21_X1 U22174 ( .B1(n19263), .B2(n19262), .A(n19261), .ZN(n19264) );
  OAI21_X1 U22175 ( .B1(n19266), .B2(n19265), .A(n19264), .ZN(P2_U3044) );
  AOI22_X1 U22176 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19313), .ZN(n19716) );
  NOR2_X1 U22177 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19379) );
  NAND2_X1 U22178 ( .A1(n19959), .A2(n19379), .ZN(n19319) );
  NOR2_X1 U22179 ( .A1(n19319), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19311) );
  INV_X1 U22180 ( .A(n19311), .ZN(n19270) );
  AND2_X1 U22181 ( .A1(n19786), .A2(n19270), .ZN(n19273) );
  INV_X1 U22182 ( .A(n19938), .ZN(n19789) );
  INV_X1 U22183 ( .A(n13658), .ZN(n19271) );
  OAI21_X1 U22184 ( .B1(n19271), .B2(n19311), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19272) );
  OAI21_X1 U22185 ( .B1(n19273), .B2(n19789), .A(n19272), .ZN(n19312) );
  NOR2_X2 U22186 ( .A1(n19274), .A2(n19708), .ZN(n19792) );
  NOR2_X2 U22187 ( .A1(n11415), .A2(n19309), .ZN(n19791) );
  AOI22_X1 U22188 ( .A1(n19312), .A2(n19792), .B1(n19791), .B2(n19311), .ZN(
        n19280) );
  INV_X1 U22189 ( .A(n19786), .ZN(n19276) );
  AOI221_X1 U22190 ( .B1(n19841), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19337), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19276), .ZN(n19277) );
  AOI211_X1 U22191 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n13658), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19277), .ZN(n19278) );
  AOI22_X1 U22192 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19313), .ZN(n19749) );
  AOI22_X1 U22193 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19315), .B1(
        n19337), .B2(n19794), .ZN(n19279) );
  OAI211_X1 U22194 ( .C1(n19716), .C2(n19829), .A(n19280), .B(n19279), .ZN(
        P2_U3048) );
  AOI22_X2 U22195 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19313), .ZN(n19803) );
  NOR2_X2 U22196 ( .A1(n19281), .A2(n19708), .ZN(n19799) );
  NOR2_X2 U22197 ( .A1(n19282), .A2(n19309), .ZN(n19798) );
  AOI22_X1 U22198 ( .A1(n19312), .A2(n19799), .B1(n19798), .B2(n19311), .ZN(
        n19285) );
  INV_X1 U22199 ( .A(n19314), .ZN(n19299) );
  INV_X1 U22200 ( .A(n19313), .ZN(n19297) );
  OAI22_X2 U22201 ( .A1(n20190), .A2(n19299), .B1(n19283), .B2(n19297), .ZN(
        n19800) );
  AOI22_X1 U22202 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19315), .B1(
        n19841), .B2(n19800), .ZN(n19284) );
  OAI211_X1 U22203 ( .C1(n19803), .C2(n19345), .A(n19285), .B(n19284), .ZN(
        P2_U3049) );
  AOI22_X1 U22204 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19313), .ZN(n19688) );
  NOR2_X2 U22205 ( .A1(n19286), .A2(n19708), .ZN(n19805) );
  NOR2_X2 U22206 ( .A1(n19287), .A2(n19309), .ZN(n19804) );
  AOI22_X1 U22207 ( .A1(n19312), .A2(n19805), .B1(n19804), .B2(n19311), .ZN(
        n19289) );
  AOI22_X1 U22208 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19313), .ZN(n19754) );
  INV_X1 U22209 ( .A(n19754), .ZN(n19807) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19315), .B1(
        n19841), .B2(n19807), .ZN(n19288) );
  OAI211_X1 U22211 ( .C1(n19688), .C2(n19345), .A(n19289), .B(n19288), .ZN(
        P2_U3050) );
  NOR2_X2 U22212 ( .A1(n19290), .A2(n19708), .ZN(n19812) );
  INV_X1 U22213 ( .A(n19309), .ZN(n19301) );
  AOI22_X1 U22214 ( .A1(n19312), .A2(n19812), .B1(n19811), .B2(n19311), .ZN(
        n19293) );
  AOI22_X1 U22215 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19313), .ZN(n19724) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19315), .B1(
        n19841), .B2(n19813), .ZN(n19292) );
  OAI211_X1 U22217 ( .C1(n19816), .C2(n19345), .A(n19293), .B(n19292), .ZN(
        P2_U3051) );
  AOI22_X1 U22218 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19313), .ZN(n19760) );
  NOR2_X2 U22219 ( .A1(n19294), .A2(n19708), .ZN(n19818) );
  NOR2_X2 U22220 ( .A1(n11430), .A2(n19309), .ZN(n19817) );
  AOI22_X1 U22221 ( .A1(n19312), .A2(n19818), .B1(n19817), .B2(n19311), .ZN(
        n19296) );
  AOI22_X1 U22222 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19313), .ZN(n19822) );
  AOI22_X1 U22223 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19315), .B1(
        n19337), .B2(n19757), .ZN(n19295) );
  OAI211_X1 U22224 ( .C1(n19760), .C2(n19829), .A(n19296), .B(n19295), .ZN(
        P2_U3052) );
  OAI22_X1 U22225 ( .A1(n20212), .A2(n19299), .B1(n19298), .B2(n19297), .ZN(
        n19825) );
  NOR2_X2 U22226 ( .A1(n19300), .A2(n19708), .ZN(n19824) );
  AOI22_X1 U22227 ( .A1(n19312), .A2(n19824), .B1(n19823), .B2(n19311), .ZN(
        n19303) );
  AOI22_X1 U22228 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19313), .ZN(n19830) );
  AOI22_X1 U22229 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19315), .B1(
        n19337), .B2(n19761), .ZN(n19302) );
  OAI211_X1 U22230 ( .C1(n19764), .C2(n19829), .A(n19303), .B(n19302), .ZN(
        P2_U3053) );
  AOI22_X1 U22231 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19313), .ZN(n19732) );
  NOR2_X2 U22232 ( .A1(n19304), .A2(n19708), .ZN(n19832) );
  AOI22_X1 U22233 ( .A1(n19312), .A2(n19832), .B1(n19831), .B2(n19311), .ZN(
        n19307) );
  AOI22_X1 U22234 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19313), .ZN(n19768) );
  AOI22_X1 U22235 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19315), .B1(
        n19841), .B2(n19834), .ZN(n19306) );
  OAI211_X1 U22236 ( .C1(n19732), .C2(n19345), .A(n19307), .B(n19306), .ZN(
        P2_U3054) );
  AOI22_X1 U22237 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19313), .ZN(n19776) );
  NOR2_X2 U22238 ( .A1(n19308), .A2(n19708), .ZN(n19838) );
  NOR2_X2 U22239 ( .A1(n19310), .A2(n19309), .ZN(n19837) );
  AOI22_X1 U22240 ( .A1(n19312), .A2(n19838), .B1(n19837), .B2(n19311), .ZN(
        n19317) );
  AOI22_X1 U22241 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19314), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19313), .ZN(n19605) );
  AOI22_X1 U22242 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19315), .B1(
        n19841), .B2(n19842), .ZN(n19316) );
  OAI211_X1 U22243 ( .C1(n19776), .C2(n19345), .A(n19317), .B(n19316), .ZN(
        P2_U3055) );
  INV_X1 U22244 ( .A(n19379), .ZN(n19376) );
  NOR2_X1 U22245 ( .A1(n19570), .A2(n19376), .ZN(n19340) );
  NOR3_X1 U22246 ( .A1(n19318), .A2(n19340), .A3(n19980), .ZN(n19321) );
  INV_X1 U22247 ( .A(n19319), .ZN(n19324) );
  AOI21_X1 U22248 ( .B1(n19324), .B2(n19979), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19320) );
  NOR2_X1 U22249 ( .A1(n19321), .A2(n19320), .ZN(n19341) );
  AOI22_X1 U22250 ( .A1(n19341), .A2(n19792), .B1(n19791), .B2(n19340), .ZN(
        n19326) );
  INV_X1 U22251 ( .A(n19340), .ZN(n19322) );
  AOI211_X1 U22252 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19322), .A(n19708), 
        .B(n19321), .ZN(n19323) );
  OAI221_X1 U22253 ( .B1(n19324), .B2(n19567), .C1(n19324), .C2(n19500), .A(
        n19323), .ZN(n19342) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19342), .B1(
        n19367), .B2(n19794), .ZN(n19325) );
  OAI211_X1 U22255 ( .C1(n19716), .C2(n19345), .A(n19326), .B(n19325), .ZN(
        P2_U3056) );
  AOI22_X1 U22256 ( .A1(n19341), .A2(n19799), .B1(n19798), .B2(n19340), .ZN(
        n19328) );
  AOI22_X1 U22257 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19342), .B1(
        n19337), .B2(n19800), .ZN(n19327) );
  OAI211_X1 U22258 ( .C1(n19803), .C2(n19375), .A(n19328), .B(n19327), .ZN(
        P2_U3057) );
  AOI22_X1 U22259 ( .A1(n19341), .A2(n19805), .B1(n19804), .B2(n19340), .ZN(
        n19330) );
  AOI22_X1 U22260 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19342), .B1(
        n19367), .B2(n19806), .ZN(n19329) );
  OAI211_X1 U22261 ( .C1(n19754), .C2(n19345), .A(n19330), .B(n19329), .ZN(
        P2_U3058) );
  AOI22_X1 U22262 ( .A1(n19341), .A2(n19812), .B1(n19811), .B2(n19340), .ZN(
        n19332) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19342), .B1(
        n19337), .B2(n19813), .ZN(n19331) );
  OAI211_X1 U22264 ( .C1(n19816), .C2(n19375), .A(n19332), .B(n19331), .ZN(
        P2_U3059) );
  AOI22_X1 U22265 ( .A1(n19341), .A2(n19818), .B1(n19817), .B2(n19340), .ZN(
        n19334) );
  AOI22_X1 U22266 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19342), .B1(
        n19367), .B2(n19757), .ZN(n19333) );
  OAI211_X1 U22267 ( .C1(n19760), .C2(n19345), .A(n19334), .B(n19333), .ZN(
        P2_U3060) );
  AOI22_X1 U22268 ( .A1(n19341), .A2(n19824), .B1(n19823), .B2(n19340), .ZN(
        n19336) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19342), .B1(
        n19367), .B2(n19761), .ZN(n19335) );
  OAI211_X1 U22270 ( .C1(n19764), .C2(n19345), .A(n19336), .B(n19335), .ZN(
        P2_U3061) );
  AOI22_X1 U22271 ( .A1(n19341), .A2(n19832), .B1(n19831), .B2(n19340), .ZN(
        n19339) );
  AOI22_X1 U22272 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19342), .B1(
        n19337), .B2(n19834), .ZN(n19338) );
  OAI211_X1 U22273 ( .C1(n19732), .C2(n19375), .A(n19339), .B(n19338), .ZN(
        P2_U3062) );
  AOI22_X1 U22274 ( .A1(n19341), .A2(n19838), .B1(n19837), .B2(n19340), .ZN(
        n19344) );
  INV_X1 U22275 ( .A(n19776), .ZN(n19840) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19342), .B1(
        n19367), .B2(n19840), .ZN(n19343) );
  OAI211_X1 U22277 ( .C1(n19605), .C2(n19345), .A(n19344), .B(n19343), .ZN(
        P2_U3063) );
  NOR3_X2 U22278 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19959), .A3(
        n19376), .ZN(n19370) );
  OAI21_X1 U22279 ( .B1(n19346), .B2(n19370), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19347) );
  OR2_X1 U22280 ( .A1(n19376), .A2(n19608), .ZN(n19348) );
  NAND2_X1 U22281 ( .A1(n19347), .A2(n19348), .ZN(n19371) );
  AOI22_X1 U22282 ( .A1(n19371), .A2(n19792), .B1(n19791), .B2(n19370), .ZN(
        n19356) );
  OAI21_X1 U22283 ( .B1(n19395), .B2(n19367), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19349) );
  NAND2_X1 U22284 ( .A1(n19349), .A2(n19348), .ZN(n19353) );
  INV_X1 U22285 ( .A(n19370), .ZN(n19350) );
  OAI21_X1 U22286 ( .B1(n19351), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19350), 
        .ZN(n19352) );
  MUX2_X1 U22287 ( .A(n19353), .B(n19352), .S(n19789), .Z(n19354) );
  NAND2_X1 U22288 ( .A1(n19354), .A2(n19781), .ZN(n19372) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19372), .B1(
        n19395), .B2(n19794), .ZN(n19355) );
  OAI211_X1 U22290 ( .C1(n19716), .C2(n19375), .A(n19356), .B(n19355), .ZN(
        P2_U3064) );
  AOI22_X1 U22291 ( .A1(n19371), .A2(n19799), .B1(n19798), .B2(n19370), .ZN(
        n19358) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19372), .B1(
        n19367), .B2(n19800), .ZN(n19357) );
  OAI211_X1 U22293 ( .C1(n19803), .C2(n19405), .A(n19358), .B(n19357), .ZN(
        P2_U3065) );
  AOI22_X1 U22294 ( .A1(n19371), .A2(n19805), .B1(n19804), .B2(n19370), .ZN(
        n19360) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19372), .B1(
        n19395), .B2(n19806), .ZN(n19359) );
  OAI211_X1 U22296 ( .C1(n19754), .C2(n19375), .A(n19360), .B(n19359), .ZN(
        P2_U3066) );
  AOI22_X1 U22297 ( .A1(n19371), .A2(n19812), .B1(n19811), .B2(n19370), .ZN(
        n19362) );
  INV_X1 U22298 ( .A(n19816), .ZN(n19721) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19372), .B1(
        n19395), .B2(n19721), .ZN(n19361) );
  OAI211_X1 U22300 ( .C1(n19724), .C2(n19375), .A(n19362), .B(n19361), .ZN(
        P2_U3067) );
  AOI22_X1 U22301 ( .A1(n19371), .A2(n19818), .B1(n19817), .B2(n19370), .ZN(
        n19364) );
  INV_X1 U22302 ( .A(n19760), .ZN(n19819) );
  AOI22_X1 U22303 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19372), .B1(
        n19367), .B2(n19819), .ZN(n19363) );
  OAI211_X1 U22304 ( .C1(n19822), .C2(n19405), .A(n19364), .B(n19363), .ZN(
        P2_U3068) );
  AOI22_X1 U22305 ( .A1(n19371), .A2(n19824), .B1(n19823), .B2(n19370), .ZN(
        n19366) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19372), .B1(
        n19367), .B2(n19825), .ZN(n19365) );
  OAI211_X1 U22307 ( .C1(n19830), .C2(n19405), .A(n19366), .B(n19365), .ZN(
        P2_U3069) );
  AOI22_X1 U22308 ( .A1(n19371), .A2(n19832), .B1(n19831), .B2(n19370), .ZN(
        n19369) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19372), .B1(
        n19367), .B2(n19834), .ZN(n19368) );
  OAI211_X1 U22310 ( .C1(n19732), .C2(n19405), .A(n19369), .B(n19368), .ZN(
        P2_U3070) );
  AOI22_X1 U22311 ( .A1(n19371), .A2(n19838), .B1(n19837), .B2(n19370), .ZN(
        n19374) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19372), .B1(
        n19395), .B2(n19840), .ZN(n19373) );
  OAI211_X1 U22313 ( .C1(n19605), .C2(n19375), .A(n19374), .B(n19373), .ZN(
        P2_U3071) );
  NOR2_X1 U22314 ( .A1(n19376), .A2(n19636), .ZN(n19400) );
  AOI22_X1 U22315 ( .A1(n19794), .A2(n19430), .B1(n19400), .B2(n19791), .ZN(
        n19386) );
  INV_X1 U22316 ( .A(n19500), .ZN(n19439) );
  OAI21_X1 U22317 ( .B1(n19439), .B2(n19634), .A(n19938), .ZN(n19384) );
  AOI21_X1 U22318 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19379), .A(
        n19384), .ZN(n19377) );
  AOI211_X1 U22319 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19380), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19377), .ZN(n19378) );
  OAI21_X1 U22320 ( .B1(n19378), .B2(n19400), .A(n19781), .ZN(n19402) );
  NAND2_X1 U22321 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19379), .ZN(
        n19383) );
  INV_X1 U22322 ( .A(n19380), .ZN(n19381) );
  OAI21_X1 U22323 ( .B1(n19381), .B2(n19400), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19382) );
  OAI21_X1 U22324 ( .B1(n19384), .B2(n19383), .A(n19382), .ZN(n19401) );
  AOI22_X1 U22325 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19402), .B1(
        n19792), .B2(n19401), .ZN(n19385) );
  OAI211_X1 U22326 ( .C1(n19716), .C2(n19405), .A(n19386), .B(n19385), .ZN(
        P2_U3072) );
  AOI22_X1 U22327 ( .A1(n19800), .A2(n19395), .B1(n19400), .B2(n19798), .ZN(
        n19388) );
  AOI22_X1 U22328 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19402), .B1(
        n19799), .B2(n19401), .ZN(n19387) );
  OAI211_X1 U22329 ( .C1(n19803), .C2(n19438), .A(n19388), .B(n19387), .ZN(
        P2_U3073) );
  AOI22_X1 U22330 ( .A1(n19806), .A2(n19430), .B1(n19400), .B2(n19804), .ZN(
        n19390) );
  AOI22_X1 U22331 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19402), .B1(
        n19805), .B2(n19401), .ZN(n19389) );
  OAI211_X1 U22332 ( .C1(n19754), .C2(n19405), .A(n19390), .B(n19389), .ZN(
        P2_U3074) );
  AOI22_X1 U22333 ( .A1(n19721), .A2(n19430), .B1(n19400), .B2(n19811), .ZN(
        n19392) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19402), .B1(
        n19812), .B2(n19401), .ZN(n19391) );
  OAI211_X1 U22335 ( .C1(n19724), .C2(n19405), .A(n19392), .B(n19391), .ZN(
        P2_U3075) );
  AOI22_X1 U22336 ( .A1(n19819), .A2(n19395), .B1(n19400), .B2(n19817), .ZN(
        n19394) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19402), .B1(
        n19818), .B2(n19401), .ZN(n19393) );
  OAI211_X1 U22338 ( .C1(n19822), .C2(n19438), .A(n19394), .B(n19393), .ZN(
        P2_U3076) );
  AOI22_X1 U22339 ( .A1(n19825), .A2(n19395), .B1(n19400), .B2(n19823), .ZN(
        n19397) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19402), .B1(
        n19824), .B2(n19401), .ZN(n19396) );
  OAI211_X1 U22341 ( .C1(n19830), .C2(n19438), .A(n19397), .B(n19396), .ZN(
        P2_U3077) );
  INV_X1 U22342 ( .A(n19732), .ZN(n19833) );
  AOI22_X1 U22343 ( .A1(n19833), .A2(n19430), .B1(n19400), .B2(n19831), .ZN(
        n19399) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19402), .B1(
        n19832), .B2(n19401), .ZN(n19398) );
  OAI211_X1 U22345 ( .C1(n19768), .C2(n19405), .A(n19399), .B(n19398), .ZN(
        P2_U3078) );
  AOI22_X1 U22346 ( .A1(n19840), .A2(n19430), .B1(n19400), .B2(n19837), .ZN(
        n19404) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19402), .B1(
        n19838), .B2(n19401), .ZN(n19403) );
  OAI211_X1 U22348 ( .C1(n19605), .C2(n19405), .A(n19404), .B(n19403), .ZN(
        P2_U3079) );
  INV_X1 U22349 ( .A(n19406), .ZN(n19408) );
  NOR2_X1 U22350 ( .A1(n19408), .A2(n19407), .ZN(n19680) );
  NAND2_X1 U22351 ( .A1(n19680), .A2(n19941), .ZN(n19415) );
  INV_X1 U22352 ( .A(n19411), .ZN(n19409) );
  NOR3_X1 U22353 ( .A1(n19950), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19443) );
  INV_X1 U22354 ( .A(n19443), .ZN(n19446) );
  NOR2_X1 U22355 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19446), .ZN(
        n19433) );
  OAI21_X1 U22356 ( .B1(n19409), .B2(n19433), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19410) );
  OAI21_X1 U22357 ( .B1(n19415), .B2(n19789), .A(n19410), .ZN(n19434) );
  AOI22_X1 U22358 ( .A1(n19434), .A2(n19792), .B1(n19791), .B2(n19433), .ZN(
        n19419) );
  AOI21_X1 U22359 ( .B1(n19411), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19417) );
  INV_X1 U22360 ( .A(n19468), .ZN(n19413) );
  OAI21_X1 U22361 ( .B1(n19430), .B2(n19460), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19414) );
  AOI21_X1 U22362 ( .B1(n19415), .B2(n19414), .A(n19708), .ZN(n19416) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19435), .B1(
        n19460), .B2(n19794), .ZN(n19418) );
  OAI211_X1 U22364 ( .C1(n19716), .C2(n19438), .A(n19419), .B(n19418), .ZN(
        P2_U3080) );
  AOI22_X1 U22365 ( .A1(n19434), .A2(n19799), .B1(n19798), .B2(n19433), .ZN(
        n19421) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19435), .B1(
        n19430), .B2(n19800), .ZN(n19420) );
  OAI211_X1 U22367 ( .C1(n19803), .C2(n19467), .A(n19421), .B(n19420), .ZN(
        P2_U3081) );
  AOI22_X1 U22368 ( .A1(n19434), .A2(n19805), .B1(n19804), .B2(n19433), .ZN(
        n19423) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19435), .B1(
        n19460), .B2(n19806), .ZN(n19422) );
  OAI211_X1 U22370 ( .C1(n19754), .C2(n19438), .A(n19423), .B(n19422), .ZN(
        P2_U3082) );
  AOI22_X1 U22371 ( .A1(n19434), .A2(n19812), .B1(n19811), .B2(n19433), .ZN(
        n19425) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19435), .B1(
        n19430), .B2(n19813), .ZN(n19424) );
  OAI211_X1 U22373 ( .C1(n19816), .C2(n19467), .A(n19425), .B(n19424), .ZN(
        P2_U3083) );
  AOI22_X1 U22374 ( .A1(n19434), .A2(n19818), .B1(n19817), .B2(n19433), .ZN(
        n19427) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19435), .B1(
        n19460), .B2(n19757), .ZN(n19426) );
  OAI211_X1 U22376 ( .C1(n19760), .C2(n19438), .A(n19427), .B(n19426), .ZN(
        P2_U3084) );
  AOI22_X1 U22377 ( .A1(n19434), .A2(n19824), .B1(n19823), .B2(n19433), .ZN(
        n19429) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19435), .B1(
        n19430), .B2(n19825), .ZN(n19428) );
  OAI211_X1 U22379 ( .C1(n19830), .C2(n19467), .A(n19429), .B(n19428), .ZN(
        P2_U3085) );
  AOI22_X1 U22380 ( .A1(n19434), .A2(n19832), .B1(n19831), .B2(n19433), .ZN(
        n19432) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19435), .B1(
        n19430), .B2(n19834), .ZN(n19431) );
  OAI211_X1 U22382 ( .C1(n19732), .C2(n19467), .A(n19432), .B(n19431), .ZN(
        P2_U3086) );
  AOI22_X1 U22383 ( .A1(n19434), .A2(n19838), .B1(n19837), .B2(n19433), .ZN(
        n19437) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19435), .B1(
        n19460), .B2(n19840), .ZN(n19436) );
  OAI211_X1 U22385 ( .C1(n19605), .C2(n19438), .A(n19437), .B(n19436), .ZN(
        P2_U3087) );
  INV_X1 U22386 ( .A(n19716), .ZN(n19793) );
  NAND2_X1 U22387 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19443), .ZN(
        n19475) );
  INV_X1 U22388 ( .A(n19475), .ZN(n19470) );
  AOI22_X1 U22389 ( .A1(n19793), .A2(n19460), .B1(n19470), .B2(n19791), .ZN(
        n19449) );
  OAI21_X1 U22390 ( .B1(n19439), .B2(n19706), .A(n19938), .ZN(n19447) );
  INV_X1 U22391 ( .A(n19440), .ZN(n19444) );
  OAI21_X1 U22392 ( .B1(n19444), .B2(n19980), .A(n19979), .ZN(n19441) );
  AOI21_X1 U22393 ( .B1(n19441), .B2(n19475), .A(n19708), .ZN(n19442) );
  OAI21_X1 U22394 ( .B1(n19447), .B2(n19443), .A(n19442), .ZN(n19464) );
  OAI21_X1 U22395 ( .B1(n19444), .B2(n19470), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19445) );
  OAI21_X1 U22396 ( .B1(n19447), .B2(n19446), .A(n19445), .ZN(n19463) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19464), .B1(
        n19792), .B2(n19463), .ZN(n19448) );
  OAI211_X1 U22398 ( .C1(n19749), .C2(n19499), .A(n19449), .B(n19448), .ZN(
        P2_U3088) );
  AOI22_X1 U22399 ( .A1(n19800), .A2(n19460), .B1(n19798), .B2(n19470), .ZN(
        n19451) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19464), .B1(
        n19799), .B2(n19463), .ZN(n19450) );
  OAI211_X1 U22401 ( .C1(n19803), .C2(n19499), .A(n19451), .B(n19450), .ZN(
        P2_U3089) );
  AOI22_X1 U22402 ( .A1(n19806), .A2(n19486), .B1(n19470), .B2(n19804), .ZN(
        n19453) );
  AOI22_X1 U22403 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19464), .B1(
        n19805), .B2(n19463), .ZN(n19452) );
  OAI211_X1 U22404 ( .C1(n19754), .C2(n19467), .A(n19453), .B(n19452), .ZN(
        P2_U3090) );
  AOI22_X1 U22405 ( .A1(n19460), .A2(n19813), .B1(n19470), .B2(n19811), .ZN(
        n19455) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19464), .B1(
        n19812), .B2(n19463), .ZN(n19454) );
  OAI211_X1 U22407 ( .C1(n19816), .C2(n19499), .A(n19455), .B(n19454), .ZN(
        P2_U3091) );
  AOI22_X1 U22408 ( .A1(n19757), .A2(n19486), .B1(n19470), .B2(n19817), .ZN(
        n19457) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19464), .B1(
        n19818), .B2(n19463), .ZN(n19456) );
  OAI211_X1 U22410 ( .C1(n19760), .C2(n19467), .A(n19457), .B(n19456), .ZN(
        P2_U3092) );
  AOI22_X1 U22411 ( .A1(n19761), .A2(n19486), .B1(n19823), .B2(n19470), .ZN(
        n19459) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19464), .B1(
        n19824), .B2(n19463), .ZN(n19458) );
  OAI211_X1 U22413 ( .C1(n19764), .C2(n19467), .A(n19459), .B(n19458), .ZN(
        P2_U3093) );
  AOI22_X1 U22414 ( .A1(n19460), .A2(n19834), .B1(n19470), .B2(n19831), .ZN(
        n19462) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19464), .B1(
        n19832), .B2(n19463), .ZN(n19461) );
  OAI211_X1 U22416 ( .C1(n19732), .C2(n19499), .A(n19462), .B(n19461), .ZN(
        P2_U3094) );
  AOI22_X1 U22417 ( .A1(n19840), .A2(n19486), .B1(n19470), .B2(n19837), .ZN(
        n19466) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19464), .B1(
        n19838), .B2(n19463), .ZN(n19465) );
  OAI211_X1 U22419 ( .C1(n19605), .C2(n19467), .A(n19466), .B(n19465), .ZN(
        P2_U3095) );
  NAND2_X1 U22420 ( .A1(n19777), .A2(n19468), .ZN(n19489) );
  NOR2_X1 U22421 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19779), .ZN(
        n19501) );
  NAND2_X1 U22422 ( .A1(n19966), .A2(n19501), .ZN(n19473) );
  NAND3_X1 U22423 ( .A1(n19469), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19473), 
        .ZN(n19476) );
  INV_X1 U22424 ( .A(n19473), .ZN(n19494) );
  NOR2_X1 U22425 ( .A1(n19470), .A2(n19494), .ZN(n19471) );
  OAI21_X1 U22426 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19471), .A(n19980), 
        .ZN(n19472) );
  AND2_X1 U22427 ( .A1(n19476), .A2(n19472), .ZN(n19495) );
  AOI22_X1 U22428 ( .A1(n19495), .A2(n19792), .B1(n19791), .B2(n19494), .ZN(
        n19479) );
  OAI21_X1 U22429 ( .B1(n19486), .B2(n19532), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19474) );
  OAI221_X1 U22430 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19475), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19474), .A(n19473), .ZN(n19477) );
  NAND3_X1 U22431 ( .A1(n19477), .A2(n19781), .A3(n19476), .ZN(n19496) );
  AOI22_X1 U22432 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19496), .B1(
        n19486), .B2(n19793), .ZN(n19478) );
  OAI211_X1 U22433 ( .C1(n19749), .C2(n19489), .A(n19479), .B(n19478), .ZN(
        P2_U3096) );
  AOI22_X1 U22434 ( .A1(n19495), .A2(n19799), .B1(n19798), .B2(n19494), .ZN(
        n19481) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19496), .B1(
        n19486), .B2(n19800), .ZN(n19480) );
  OAI211_X1 U22436 ( .C1(n19803), .C2(n19489), .A(n19481), .B(n19480), .ZN(
        P2_U3097) );
  AOI22_X1 U22437 ( .A1(n19495), .A2(n19805), .B1(n19804), .B2(n19494), .ZN(
        n19483) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19496), .B1(
        n19532), .B2(n19806), .ZN(n19482) );
  OAI211_X1 U22439 ( .C1(n19754), .C2(n19499), .A(n19483), .B(n19482), .ZN(
        P2_U3098) );
  AOI22_X1 U22440 ( .A1(n19495), .A2(n19812), .B1(n19811), .B2(n19494), .ZN(
        n19485) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19496), .B1(
        n19486), .B2(n19813), .ZN(n19484) );
  OAI211_X1 U22442 ( .C1(n19816), .C2(n19489), .A(n19485), .B(n19484), .ZN(
        P2_U3099) );
  AOI22_X1 U22443 ( .A1(n19495), .A2(n19818), .B1(n19817), .B2(n19494), .ZN(
        n19488) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19496), .B1(
        n19486), .B2(n19819), .ZN(n19487) );
  OAI211_X1 U22445 ( .C1(n19822), .C2(n19489), .A(n19488), .B(n19487), .ZN(
        P2_U3100) );
  AOI22_X1 U22446 ( .A1(n19495), .A2(n19824), .B1(n19823), .B2(n19494), .ZN(
        n19491) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19496), .B1(
        n19532), .B2(n19761), .ZN(n19490) );
  OAI211_X1 U22448 ( .C1(n19764), .C2(n19499), .A(n19491), .B(n19490), .ZN(
        P2_U3101) );
  AOI22_X1 U22449 ( .A1(n19495), .A2(n19832), .B1(n19831), .B2(n19494), .ZN(
        n19493) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19496), .B1(
        n19532), .B2(n19833), .ZN(n19492) );
  OAI211_X1 U22451 ( .C1(n19768), .C2(n19499), .A(n19493), .B(n19492), .ZN(
        P2_U3102) );
  AOI22_X1 U22452 ( .A1(n19495), .A2(n19838), .B1(n19837), .B2(n19494), .ZN(
        n19498) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19496), .B1(
        n19532), .B2(n19840), .ZN(n19497) );
  OAI211_X1 U22454 ( .C1(n19605), .C2(n19499), .A(n19498), .B(n19497), .ZN(
        P2_U3103) );
  AND2_X1 U22455 ( .A1(n19500), .A2(n19777), .ZN(n19937) );
  INV_X1 U22456 ( .A(n19937), .ZN(n19502) );
  INV_X1 U22457 ( .A(n19501), .ZN(n19508) );
  NAND2_X1 U22458 ( .A1(n19502), .A2(n19508), .ZN(n19507) );
  NOR2_X1 U22459 ( .A1(n19966), .A2(n19508), .ZN(n19542) );
  INV_X1 U22460 ( .A(n19542), .ZN(n19539) );
  AND2_X1 U22461 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19539), .ZN(n19503) );
  NAND2_X1 U22462 ( .A1(n19504), .A2(n19503), .ZN(n19510) );
  OAI211_X1 U22463 ( .C1(n19542), .C2(n19979), .A(n19510), .B(n19781), .ZN(
        n19505) );
  INV_X1 U22464 ( .A(n19505), .ZN(n19506) );
  INV_X1 U22465 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19515) );
  OAI21_X1 U22466 ( .B1(n19508), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19980), 
        .ZN(n19509) );
  AND2_X1 U22467 ( .A1(n19510), .A2(n19509), .ZN(n19531) );
  AOI22_X1 U22468 ( .A1(n19531), .A2(n19792), .B1(n19791), .B2(n19542), .ZN(
        n19514) );
  AOI22_X1 U22469 ( .A1(n19561), .A2(n19794), .B1(n19532), .B2(n19793), .ZN(
        n19513) );
  OAI211_X1 U22470 ( .C1(n19526), .C2(n19515), .A(n19514), .B(n19513), .ZN(
        P2_U3104) );
  AOI22_X1 U22471 ( .A1(n19531), .A2(n19799), .B1(n19798), .B2(n19542), .ZN(
        n19517) );
  INV_X1 U22472 ( .A(n19526), .ZN(n19533) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19800), .ZN(n19516) );
  OAI211_X1 U22474 ( .C1(n19803), .C2(n19557), .A(n19517), .B(n19516), .ZN(
        P2_U3105) );
  AOI22_X1 U22475 ( .A1(n19531), .A2(n19805), .B1(n19804), .B2(n19542), .ZN(
        n19519) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19807), .ZN(n19518) );
  OAI211_X1 U22477 ( .C1(n19688), .C2(n19557), .A(n19519), .B(n19518), .ZN(
        P2_U3106) );
  AOI22_X1 U22478 ( .A1(n19531), .A2(n19812), .B1(n19811), .B2(n19542), .ZN(
        n19521) );
  AOI22_X1 U22479 ( .A1(n19561), .A2(n19721), .B1(n19532), .B2(n19813), .ZN(
        n19520) );
  OAI211_X1 U22480 ( .C1(n19526), .C2(n19522), .A(n19521), .B(n19520), .ZN(
        P2_U3107) );
  INV_X1 U22481 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n19525) );
  AOI22_X1 U22482 ( .A1(n19531), .A2(n19818), .B1(n19817), .B2(n19542), .ZN(
        n19524) );
  AOI22_X1 U22483 ( .A1(n19561), .A2(n19757), .B1(n19532), .B2(n19819), .ZN(
        n19523) );
  OAI211_X1 U22484 ( .C1(n19526), .C2(n19525), .A(n19524), .B(n19523), .ZN(
        P2_U3108) );
  AOI22_X1 U22485 ( .A1(n19531), .A2(n19824), .B1(n19823), .B2(n19542), .ZN(
        n19528) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19825), .ZN(n19527) );
  OAI211_X1 U22487 ( .C1(n19830), .C2(n19557), .A(n19528), .B(n19527), .ZN(
        P2_U3109) );
  AOI22_X1 U22488 ( .A1(n19531), .A2(n19832), .B1(n19831), .B2(n19542), .ZN(
        n19530) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19834), .ZN(n19529) );
  OAI211_X1 U22490 ( .C1(n19732), .C2(n19557), .A(n19530), .B(n19529), .ZN(
        P2_U3110) );
  AOI22_X1 U22491 ( .A1(n19531), .A2(n19838), .B1(n19837), .B2(n19542), .ZN(
        n19535) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19842), .ZN(n19534) );
  OAI211_X1 U22493 ( .C1(n19776), .C2(n19557), .A(n19535), .B(n19534), .ZN(
        P2_U3111) );
  INV_X1 U22494 ( .A(n19604), .ZN(n19591) );
  NAND2_X1 U22495 ( .A1(n19950), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19641) );
  OR2_X1 U22496 ( .A1(n19641), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19578) );
  NOR2_X1 U22497 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19578), .ZN(
        n19560) );
  AOI22_X1 U22498 ( .A1(n19794), .A2(n19591), .B1(n19560), .B2(n19791), .ZN(
        n19546) );
  NAND2_X1 U22499 ( .A1(n19557), .A2(n19604), .ZN(n19537) );
  AOI21_X1 U22500 ( .B1(n19537), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19789), 
        .ZN(n19541) );
  AOI21_X1 U22501 ( .B1(n13649), .B2(n19979), .A(n19938), .ZN(n19538) );
  AOI21_X1 U22502 ( .B1(n19541), .B2(n19539), .A(n19538), .ZN(n19540) );
  OAI21_X1 U22503 ( .B1(n19560), .B2(n19540), .A(n19781), .ZN(n19563) );
  OAI21_X1 U22504 ( .B1(n19560), .B2(n19542), .A(n19541), .ZN(n19544) );
  OAI21_X1 U22505 ( .B1(n13649), .B2(n19560), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19543) );
  NAND2_X1 U22506 ( .A1(n19544), .A2(n19543), .ZN(n19562) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19563), .B1(
        n19792), .B2(n19562), .ZN(n19545) );
  OAI211_X1 U22508 ( .C1(n19716), .C2(n19557), .A(n19546), .B(n19545), .ZN(
        P2_U3112) );
  AOI22_X1 U22509 ( .A1(n19800), .A2(n19561), .B1(n19798), .B2(n19560), .ZN(
        n19548) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19563), .B1(
        n19562), .B2(n19799), .ZN(n19547) );
  OAI211_X1 U22511 ( .C1(n19803), .C2(n19604), .A(n19548), .B(n19547), .ZN(
        P2_U3113) );
  AOI22_X1 U22512 ( .A1(n19807), .A2(n19561), .B1(n19560), .B2(n19804), .ZN(
        n19550) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19563), .B1(
        n19562), .B2(n19805), .ZN(n19549) );
  OAI211_X1 U22514 ( .C1(n19688), .C2(n19604), .A(n19550), .B(n19549), .ZN(
        P2_U3114) );
  AOI22_X1 U22515 ( .A1(n19813), .A2(n19561), .B1(n19560), .B2(n19811), .ZN(
        n19552) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19563), .B1(
        n19562), .B2(n19812), .ZN(n19551) );
  OAI211_X1 U22517 ( .C1(n19816), .C2(n19604), .A(n19552), .B(n19551), .ZN(
        P2_U3115) );
  AOI22_X1 U22518 ( .A1(n19757), .A2(n19591), .B1(n19560), .B2(n19817), .ZN(
        n19554) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19563), .B1(
        n19562), .B2(n19818), .ZN(n19553) );
  OAI211_X1 U22520 ( .C1(n19760), .C2(n19557), .A(n19554), .B(n19553), .ZN(
        P2_U3116) );
  AOI22_X1 U22521 ( .A1(n19761), .A2(n19591), .B1(n19823), .B2(n19560), .ZN(
        n19556) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19563), .B1(
        n19562), .B2(n19824), .ZN(n19555) );
  OAI211_X1 U22523 ( .C1(n19764), .C2(n19557), .A(n19556), .B(n19555), .ZN(
        P2_U3117) );
  AOI22_X1 U22524 ( .A1(n19834), .A2(n19561), .B1(n19560), .B2(n19831), .ZN(
        n19559) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19563), .B1(
        n19562), .B2(n19832), .ZN(n19558) );
  OAI211_X1 U22526 ( .C1(n19732), .C2(n19604), .A(n19559), .B(n19558), .ZN(
        P2_U3118) );
  AOI22_X1 U22527 ( .A1(n19842), .A2(n19561), .B1(n19560), .B2(n19837), .ZN(
        n19565) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19563), .B1(
        n19562), .B2(n19838), .ZN(n19564) );
  OAI211_X1 U22529 ( .C1(n19776), .C2(n19604), .A(n19565), .B(n19564), .ZN(
        P2_U3119) );
  NOR2_X1 U22530 ( .A1(n19566), .A2(n19989), .ZN(n19778) );
  NAND2_X1 U22531 ( .A1(n19778), .A2(n19567), .ZN(n19568) );
  NAND2_X1 U22532 ( .A1(n19568), .A2(n19938), .ZN(n19579) );
  INV_X1 U22533 ( .A(n19578), .ZN(n19569) );
  OR2_X1 U22534 ( .A1(n19579), .A2(n19569), .ZN(n19575) );
  NOR2_X1 U22535 ( .A1(n19570), .A2(n19641), .ZN(n19609) );
  INV_X1 U22536 ( .A(n19609), .ZN(n19571) );
  OAI211_X1 U22537 ( .C1(n19572), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19571), 
        .B(n19789), .ZN(n19573) );
  AND2_X1 U22538 ( .A1(n19573), .A2(n19781), .ZN(n19574) );
  INV_X1 U22539 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19583) );
  AOI22_X1 U22540 ( .A1(n19793), .A2(n19591), .B1(n19609), .B2(n19791), .ZN(
        n19582) );
  OAI21_X1 U22541 ( .B1(n19576), .B2(n19609), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19577) );
  OAI21_X1 U22542 ( .B1(n19579), .B2(n19578), .A(n19577), .ZN(n19600) );
  AOI22_X1 U22543 ( .A1(n19792), .A2(n19600), .B1(n19630), .B2(n19794), .ZN(
        n19581) );
  OAI211_X1 U22544 ( .C1(n19588), .C2(n19583), .A(n19582), .B(n19581), .ZN(
        P2_U3120) );
  INV_X1 U22545 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n19587) );
  AOI22_X1 U22546 ( .A1(n19800), .A2(n19591), .B1(n19798), .B2(n19609), .ZN(
        n19586) );
  INV_X1 U22547 ( .A(n19803), .ZN(n19584) );
  AOI22_X1 U22548 ( .A1(n19799), .A2(n19600), .B1(n19630), .B2(n19584), .ZN(
        n19585) );
  OAI211_X1 U22549 ( .C1(n19588), .C2(n19587), .A(n19586), .B(n19585), .ZN(
        P2_U3121) );
  AOI22_X1 U22550 ( .A1(n19807), .A2(n19591), .B1(n19609), .B2(n19804), .ZN(
        n19590) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19601), .B1(
        n19805), .B2(n19600), .ZN(n19589) );
  OAI211_X1 U22552 ( .C1(n19688), .C2(n19625), .A(n19590), .B(n19589), .ZN(
        P2_U3122) );
  AOI22_X1 U22553 ( .A1(n19813), .A2(n19591), .B1(n19609), .B2(n19811), .ZN(
        n19593) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19601), .B1(
        n19812), .B2(n19600), .ZN(n19592) );
  OAI211_X1 U22555 ( .C1(n19816), .C2(n19625), .A(n19593), .B(n19592), .ZN(
        P2_U3123) );
  AOI22_X1 U22556 ( .A1(n19630), .A2(n19757), .B1(n19609), .B2(n19817), .ZN(
        n19595) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19601), .B1(
        n19818), .B2(n19600), .ZN(n19594) );
  OAI211_X1 U22558 ( .C1(n19760), .C2(n19604), .A(n19595), .B(n19594), .ZN(
        P2_U3124) );
  AOI22_X1 U22559 ( .A1(n19630), .A2(n19761), .B1(n19823), .B2(n19609), .ZN(
        n19597) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19601), .B1(
        n19824), .B2(n19600), .ZN(n19596) );
  OAI211_X1 U22561 ( .C1(n19764), .C2(n19604), .A(n19597), .B(n19596), .ZN(
        P2_U3125) );
  AOI22_X1 U22562 ( .A1(n19630), .A2(n19833), .B1(n19609), .B2(n19831), .ZN(
        n19599) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19601), .B1(
        n19832), .B2(n19600), .ZN(n19598) );
  OAI211_X1 U22564 ( .C1(n19768), .C2(n19604), .A(n19599), .B(n19598), .ZN(
        P2_U3126) );
  AOI22_X1 U22565 ( .A1(n19630), .A2(n19840), .B1(n19609), .B2(n19837), .ZN(
        n19603) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19601), .B1(
        n19838), .B2(n19600), .ZN(n19602) );
  OAI211_X1 U22567 ( .C1(n19605), .C2(n19604), .A(n19603), .B(n19602), .ZN(
        P2_U3127) );
  NOR3_X2 U22568 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19959), .A3(
        n19641), .ZN(n19628) );
  OAI21_X1 U22569 ( .B1(n19606), .B2(n19628), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19607) );
  OAI21_X1 U22570 ( .B1(n19641), .B2(n19608), .A(n19607), .ZN(n19629) );
  AOI22_X1 U22571 ( .A1(n19629), .A2(n19792), .B1(n19791), .B2(n19628), .ZN(
        n19614) );
  AOI221_X1 U22572 ( .B1(n19630), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19666), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19609), .ZN(n19610) );
  AOI211_X1 U22573 ( .C1(n19611), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19610), .ZN(n19612) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19631), .B1(
        n19666), .B2(n19794), .ZN(n19613) );
  OAI211_X1 U22575 ( .C1(n19716), .C2(n19625), .A(n19614), .B(n19613), .ZN(
        P2_U3128) );
  AOI22_X1 U22576 ( .A1(n19629), .A2(n19799), .B1(n19798), .B2(n19628), .ZN(
        n19616) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n19800), .ZN(n19615) );
  OAI211_X1 U22578 ( .C1(n19803), .C2(n19663), .A(n19616), .B(n19615), .ZN(
        P2_U3129) );
  AOI22_X1 U22579 ( .A1(n19629), .A2(n19805), .B1(n19804), .B2(n19628), .ZN(
        n19618) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n19807), .ZN(n19617) );
  OAI211_X1 U22581 ( .C1(n19688), .C2(n19663), .A(n19618), .B(n19617), .ZN(
        P2_U3130) );
  AOI22_X1 U22582 ( .A1(n19629), .A2(n19812), .B1(n19811), .B2(n19628), .ZN(
        n19620) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n19813), .ZN(n19619) );
  OAI211_X1 U22584 ( .C1(n19816), .C2(n19663), .A(n19620), .B(n19619), .ZN(
        P2_U3131) );
  AOI22_X1 U22585 ( .A1(n19629), .A2(n19818), .B1(n19817), .B2(n19628), .ZN(
        n19622) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19631), .B1(
        n19666), .B2(n19757), .ZN(n19621) );
  OAI211_X1 U22587 ( .C1(n19760), .C2(n19625), .A(n19622), .B(n19621), .ZN(
        P2_U3132) );
  AOI22_X1 U22588 ( .A1(n19629), .A2(n19824), .B1(n19823), .B2(n19628), .ZN(
        n19624) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19631), .B1(
        n19666), .B2(n19761), .ZN(n19623) );
  OAI211_X1 U22590 ( .C1(n19764), .C2(n19625), .A(n19624), .B(n19623), .ZN(
        P2_U3133) );
  AOI22_X1 U22591 ( .A1(n19629), .A2(n19832), .B1(n19831), .B2(n19628), .ZN(
        n19627) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n19834), .ZN(n19626) );
  OAI211_X1 U22593 ( .C1(n19732), .C2(n19663), .A(n19627), .B(n19626), .ZN(
        P2_U3134) );
  AOI22_X1 U22594 ( .A1(n19629), .A2(n19838), .B1(n19837), .B2(n19628), .ZN(
        n19633) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n19842), .ZN(n19632) );
  OAI211_X1 U22596 ( .C1(n19776), .C2(n19663), .A(n19633), .B(n19632), .ZN(
        P2_U3135) );
  INV_X1 U22597 ( .A(n19699), .ZN(n19675) );
  INV_X1 U22598 ( .A(n19636), .ZN(n19638) );
  INV_X1 U22599 ( .A(n19641), .ZN(n19637) );
  NAND2_X1 U22600 ( .A1(n19638), .A2(n19637), .ZN(n19644) );
  AND2_X1 U22601 ( .A1(n19644), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19639) );
  NAND2_X1 U22602 ( .A1(n19640), .A2(n19639), .ZN(n19645) );
  NOR2_X1 U22603 ( .A1(n19959), .A2(n19641), .ZN(n19648) );
  INV_X1 U22604 ( .A(n19648), .ZN(n19642) );
  OAI21_X1 U22605 ( .B1(n19642), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19980), 
        .ZN(n19643) );
  INV_X1 U22606 ( .A(n19644), .ZN(n19664) );
  AOI22_X1 U22607 ( .A1(n19665), .A2(n19792), .B1(n19791), .B2(n19664), .ZN(
        n19650) );
  OAI211_X1 U22608 ( .C1(n19664), .C2(n19979), .A(n19645), .B(n19781), .ZN(
        n19646) );
  INV_X1 U22609 ( .A(n19646), .ZN(n19647) );
  OAI221_X1 U22610 ( .B1(n19648), .B2(n19932), .C1(n19648), .C2(n19778), .A(
        n19647), .ZN(n19667) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19793), .ZN(n19649) );
  OAI211_X1 U22612 ( .C1(n19749), .C2(n19675), .A(n19650), .B(n19649), .ZN(
        P2_U3136) );
  AOI22_X1 U22613 ( .A1(n19665), .A2(n19799), .B1(n19798), .B2(n19664), .ZN(
        n19652) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19800), .ZN(n19651) );
  OAI211_X1 U22615 ( .C1(n19803), .C2(n19675), .A(n19652), .B(n19651), .ZN(
        P2_U3137) );
  AOI22_X1 U22616 ( .A1(n19665), .A2(n19805), .B1(n19804), .B2(n19664), .ZN(
        n19654) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19667), .B1(
        n19699), .B2(n19806), .ZN(n19653) );
  OAI211_X1 U22618 ( .C1(n19754), .C2(n19663), .A(n19654), .B(n19653), .ZN(
        P2_U3138) );
  AOI22_X1 U22619 ( .A1(n19665), .A2(n19812), .B1(n19811), .B2(n19664), .ZN(
        n19656) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19667), .B1(
        n19699), .B2(n19721), .ZN(n19655) );
  OAI211_X1 U22621 ( .C1(n19724), .C2(n19663), .A(n19656), .B(n19655), .ZN(
        P2_U3139) );
  AOI22_X1 U22622 ( .A1(n19665), .A2(n19818), .B1(n19817), .B2(n19664), .ZN(
        n19658) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19667), .B1(
        n19699), .B2(n19757), .ZN(n19657) );
  OAI211_X1 U22624 ( .C1(n19760), .C2(n19663), .A(n19658), .B(n19657), .ZN(
        P2_U3140) );
  AOI22_X1 U22625 ( .A1(n19665), .A2(n19824), .B1(n19823), .B2(n19664), .ZN(
        n19660) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19667), .B1(
        n19699), .B2(n19761), .ZN(n19659) );
  OAI211_X1 U22627 ( .C1(n19764), .C2(n19663), .A(n19660), .B(n19659), .ZN(
        P2_U3141) );
  AOI22_X1 U22628 ( .A1(n19665), .A2(n19832), .B1(n19831), .B2(n19664), .ZN(
        n19662) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19667), .B1(
        n19699), .B2(n19833), .ZN(n19661) );
  OAI211_X1 U22630 ( .C1(n19768), .C2(n19663), .A(n19662), .B(n19661), .ZN(
        P2_U3142) );
  AOI22_X1 U22631 ( .A1(n19665), .A2(n19838), .B1(n19837), .B2(n19664), .ZN(
        n19669) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19842), .ZN(n19668) );
  OAI211_X1 U22633 ( .C1(n19776), .C2(n19675), .A(n19669), .B(n19668), .ZN(
        P2_U3143) );
  INV_X1 U22634 ( .A(n19738), .ZN(n19670) );
  INV_X1 U22635 ( .A(n19680), .ZN(n19673) );
  NAND3_X1 U22636 ( .A1(n19959), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19703) );
  INV_X1 U22637 ( .A(n19703), .ZN(n19711) );
  NAND2_X1 U22638 ( .A1(n19966), .A2(n19711), .ZN(n19676) );
  INV_X1 U22639 ( .A(n19676), .ZN(n19697) );
  OAI21_X1 U22640 ( .B1(n19671), .B2(n19697), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19672) );
  OAI21_X1 U22641 ( .B1(n19674), .B2(n19673), .A(n19672), .ZN(n19698) );
  AOI22_X1 U22642 ( .A1(n19698), .A2(n19792), .B1(n19791), .B2(n19697), .ZN(
        n19683) );
  AOI21_X1 U22643 ( .B1(n19729), .B2(n19675), .A(n19989), .ZN(n19681) );
  OAI211_X1 U22644 ( .C1(n19677), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19676), 
        .B(n19789), .ZN(n19678) );
  AND2_X1 U22645 ( .A1(n19678), .A2(n19781), .ZN(n19679) );
  OAI211_X1 U22646 ( .C1(n19681), .C2(n19680), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19679), .ZN(n19700) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19700), .B1(
        n19699), .B2(n19793), .ZN(n19682) );
  OAI211_X1 U22648 ( .C1(n19749), .C2(n19729), .A(n19683), .B(n19682), .ZN(
        P2_U3144) );
  AOI22_X1 U22649 ( .A1(n19698), .A2(n19799), .B1(n19798), .B2(n19697), .ZN(
        n19685) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19700), .B1(
        n19699), .B2(n19800), .ZN(n19684) );
  OAI211_X1 U22651 ( .C1(n19803), .C2(n19729), .A(n19685), .B(n19684), .ZN(
        P2_U3145) );
  AOI22_X1 U22652 ( .A1(n19698), .A2(n19805), .B1(n19804), .B2(n19697), .ZN(
        n19687) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19700), .B1(
        n19699), .B2(n19807), .ZN(n19686) );
  OAI211_X1 U22654 ( .C1(n19688), .C2(n19729), .A(n19687), .B(n19686), .ZN(
        P2_U3146) );
  AOI22_X1 U22655 ( .A1(n19698), .A2(n19812), .B1(n19811), .B2(n19697), .ZN(
        n19690) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19700), .B1(
        n19699), .B2(n19813), .ZN(n19689) );
  OAI211_X1 U22657 ( .C1(n19816), .C2(n19729), .A(n19690), .B(n19689), .ZN(
        P2_U3147) );
  AOI22_X1 U22658 ( .A1(n19698), .A2(n19818), .B1(n19817), .B2(n19697), .ZN(
        n19692) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19700), .B1(
        n19699), .B2(n19819), .ZN(n19691) );
  OAI211_X1 U22660 ( .C1(n19822), .C2(n19729), .A(n19692), .B(n19691), .ZN(
        P2_U3148) );
  AOI22_X1 U22661 ( .A1(n19698), .A2(n19824), .B1(n19823), .B2(n19697), .ZN(
        n19694) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19700), .B1(
        n19699), .B2(n19825), .ZN(n19693) );
  OAI211_X1 U22663 ( .C1(n19830), .C2(n19729), .A(n19694), .B(n19693), .ZN(
        P2_U3149) );
  AOI22_X1 U22664 ( .A1(n19698), .A2(n19832), .B1(n19831), .B2(n19697), .ZN(
        n19696) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19700), .B1(
        n19699), .B2(n19834), .ZN(n19695) );
  OAI211_X1 U22666 ( .C1(n19732), .C2(n19729), .A(n19696), .B(n19695), .ZN(
        P2_U3150) );
  AOI22_X1 U22667 ( .A1(n19698), .A2(n19838), .B1(n19837), .B2(n19697), .ZN(
        n19702) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19700), .B1(
        n19699), .B2(n19842), .ZN(n19701) );
  OAI211_X1 U22669 ( .C1(n19776), .C2(n19729), .A(n19702), .B(n19701), .ZN(
        P2_U3151) );
  NOR2_X1 U22670 ( .A1(n19966), .A2(n19703), .ZN(n19740) );
  NOR3_X1 U22671 ( .A1(n19704), .A2(n19740), .A3(n19980), .ZN(n19707) );
  AOI21_X1 U22672 ( .B1(n19979), .B2(n19711), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19705) );
  NOR2_X1 U22673 ( .A1(n19707), .A2(n19705), .ZN(n19733) );
  AOI22_X1 U22674 ( .A1(n19733), .A2(n19792), .B1(n19791), .B2(n19740), .ZN(
        n19715) );
  INV_X1 U22675 ( .A(n19706), .ZN(n19712) );
  INV_X1 U22676 ( .A(n19740), .ZN(n19709) );
  AOI211_X1 U22677 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19709), .A(n19708), 
        .B(n19707), .ZN(n19710) );
  OAI221_X1 U22678 ( .B1(n19711), .B2(n19712), .C1(n19711), .C2(n19778), .A(
        n19710), .ZN(n19735) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19735), .B1(
        n19770), .B2(n19794), .ZN(n19714) );
  OAI211_X1 U22680 ( .C1(n19716), .C2(n19729), .A(n19715), .B(n19714), .ZN(
        P2_U3152) );
  INV_X1 U22681 ( .A(n19770), .ZN(n19767) );
  AOI22_X1 U22682 ( .A1(n19733), .A2(n19799), .B1(n19798), .B2(n19740), .ZN(
        n19718) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19800), .ZN(n19717) );
  OAI211_X1 U22684 ( .C1(n19803), .C2(n19767), .A(n19718), .B(n19717), .ZN(
        P2_U3153) );
  AOI22_X1 U22685 ( .A1(n19733), .A2(n19805), .B1(n19804), .B2(n19740), .ZN(
        n19720) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19735), .B1(
        n19770), .B2(n19806), .ZN(n19719) );
  OAI211_X1 U22687 ( .C1(n19754), .C2(n19729), .A(n19720), .B(n19719), .ZN(
        P2_U3154) );
  AOI22_X1 U22688 ( .A1(n19733), .A2(n19812), .B1(n19811), .B2(n19740), .ZN(
        n19723) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19735), .B1(
        n19770), .B2(n19721), .ZN(n19722) );
  OAI211_X1 U22690 ( .C1(n19724), .C2(n19729), .A(n19723), .B(n19722), .ZN(
        P2_U3155) );
  AOI22_X1 U22691 ( .A1(n19733), .A2(n19818), .B1(n19817), .B2(n19740), .ZN(
        n19726) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19735), .B1(
        n19770), .B2(n19757), .ZN(n19725) );
  OAI211_X1 U22693 ( .C1(n19760), .C2(n19729), .A(n19726), .B(n19725), .ZN(
        P2_U3156) );
  AOI22_X1 U22694 ( .A1(n19733), .A2(n19824), .B1(n19823), .B2(n19740), .ZN(
        n19728) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19735), .B1(
        n19770), .B2(n19761), .ZN(n19727) );
  OAI211_X1 U22696 ( .C1(n19764), .C2(n19729), .A(n19728), .B(n19727), .ZN(
        P2_U3157) );
  AOI22_X1 U22697 ( .A1(n19733), .A2(n19832), .B1(n19831), .B2(n19740), .ZN(
        n19731) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19834), .ZN(n19730) );
  OAI211_X1 U22699 ( .C1(n19732), .C2(n19767), .A(n19731), .B(n19730), .ZN(
        P2_U3158) );
  AOI22_X1 U22700 ( .A1(n19733), .A2(n19838), .B1(n19837), .B2(n19740), .ZN(
        n19737) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19842), .ZN(n19736) );
  OAI211_X1 U22702 ( .C1(n19776), .C2(n19767), .A(n19737), .B(n19736), .ZN(
        P2_U3159) );
  INV_X1 U22703 ( .A(n19843), .ZN(n19775) );
  NOR3_X2 U22704 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19941), .A3(
        n19779), .ZN(n19769) );
  AOI22_X1 U22705 ( .A1(n19793), .A2(n19770), .B1(n19769), .B2(n19791), .ZN(
        n19748) );
  OAI21_X1 U22706 ( .B1(n19843), .B2(n19770), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19739) );
  NAND2_X1 U22707 ( .A1(n19739), .A2(n19938), .ZN(n19746) );
  NOR2_X1 U22708 ( .A1(n19769), .A2(n19740), .ZN(n19745) );
  INV_X1 U22709 ( .A(n19745), .ZN(n19742) );
  OAI211_X1 U22710 ( .C1(n19746), .C2(n19742), .A(n19781), .B(n19741), .ZN(
        n19772) );
  OAI21_X1 U22711 ( .B1(n19743), .B2(n19769), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19744) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19772), .B1(
        n19792), .B2(n19771), .ZN(n19747) );
  OAI211_X1 U22713 ( .C1(n19749), .C2(n19775), .A(n19748), .B(n19747), .ZN(
        P2_U3160) );
  AOI22_X1 U22714 ( .A1(n19800), .A2(n19770), .B1(n19798), .B2(n19769), .ZN(
        n19751) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19772), .B1(
        n19799), .B2(n19771), .ZN(n19750) );
  OAI211_X1 U22716 ( .C1(n19803), .C2(n19775), .A(n19751), .B(n19750), .ZN(
        P2_U3161) );
  AOI22_X1 U22717 ( .A1(n19806), .A2(n19843), .B1(n19769), .B2(n19804), .ZN(
        n19753) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19772), .B1(
        n19805), .B2(n19771), .ZN(n19752) );
  OAI211_X1 U22719 ( .C1(n19754), .C2(n19767), .A(n19753), .B(n19752), .ZN(
        P2_U3162) );
  AOI22_X1 U22720 ( .A1(n19813), .A2(n19770), .B1(n19769), .B2(n19811), .ZN(
        n19756) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19772), .B1(
        n19812), .B2(n19771), .ZN(n19755) );
  OAI211_X1 U22722 ( .C1(n19816), .C2(n19775), .A(n19756), .B(n19755), .ZN(
        P2_U3163) );
  AOI22_X1 U22723 ( .A1(n19757), .A2(n19843), .B1(n19769), .B2(n19817), .ZN(
        n19759) );
  AOI22_X1 U22724 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19772), .B1(
        n19818), .B2(n19771), .ZN(n19758) );
  OAI211_X1 U22725 ( .C1(n19760), .C2(n19767), .A(n19759), .B(n19758), .ZN(
        P2_U3164) );
  AOI22_X1 U22726 ( .A1(n19761), .A2(n19843), .B1(n19823), .B2(n19769), .ZN(
        n19763) );
  AOI22_X1 U22727 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19772), .B1(
        n19824), .B2(n19771), .ZN(n19762) );
  OAI211_X1 U22728 ( .C1(n19764), .C2(n19767), .A(n19763), .B(n19762), .ZN(
        P2_U3165) );
  AOI22_X1 U22729 ( .A1(n19833), .A2(n19843), .B1(n19769), .B2(n19831), .ZN(
        n19766) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19772), .B1(
        n19832), .B2(n19771), .ZN(n19765) );
  OAI211_X1 U22731 ( .C1(n19768), .C2(n19767), .A(n19766), .B(n19765), .ZN(
        P2_U3166) );
  AOI22_X1 U22732 ( .A1(n19842), .A2(n19770), .B1(n19769), .B2(n19837), .ZN(
        n19774) );
  AOI22_X1 U22733 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19772), .B1(
        n19838), .B2(n19771), .ZN(n19773) );
  OAI211_X1 U22734 ( .C1(n19776), .C2(n19775), .A(n19774), .B(n19773), .ZN(
        P2_U3167) );
  NAND2_X1 U22735 ( .A1(n19778), .A2(n19777), .ZN(n19780) );
  OR2_X1 U22736 ( .A1(n19941), .A2(n19779), .ZN(n19790) );
  NAND2_X1 U22737 ( .A1(n19780), .A2(n19790), .ZN(n19784) );
  OAI211_X1 U22738 ( .C1(n19785), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19786), 
        .B(n19789), .ZN(n19782) );
  AND2_X1 U22739 ( .A1(n19782), .A2(n19781), .ZN(n19783) );
  AND2_X1 U22740 ( .A1(n19784), .A2(n19783), .ZN(n19847) );
  INV_X1 U22741 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n19797) );
  INV_X1 U22742 ( .A(n19785), .ZN(n19787) );
  OAI21_X1 U22743 ( .B1(n19787), .B2(n19276), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19788) );
  OAI21_X1 U22744 ( .B1(n19790), .B2(n19789), .A(n19788), .ZN(n19839) );
  AOI22_X1 U22745 ( .A1(n19839), .A2(n19792), .B1(n19276), .B2(n19791), .ZN(
        n19796) );
  AOI22_X1 U22746 ( .A1(n19841), .A2(n19794), .B1(n19843), .B2(n19793), .ZN(
        n19795) );
  OAI211_X1 U22747 ( .C1(n19847), .C2(n19797), .A(n19796), .B(n19795), .ZN(
        P2_U3168) );
  AOI22_X1 U22748 ( .A1(n19839), .A2(n19799), .B1(n19276), .B2(n19798), .ZN(
        n19802) );
  INV_X1 U22749 ( .A(n19847), .ZN(n19826) );
  AOI22_X1 U22750 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19826), .B1(
        n19843), .B2(n19800), .ZN(n19801) );
  OAI211_X1 U22751 ( .C1(n19803), .C2(n19829), .A(n19802), .B(n19801), .ZN(
        P2_U3169) );
  INV_X1 U22752 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n19810) );
  AOI22_X1 U22753 ( .A1(n19839), .A2(n19805), .B1(n19276), .B2(n19804), .ZN(
        n19809) );
  AOI22_X1 U22754 ( .A1(n19843), .A2(n19807), .B1(n19841), .B2(n19806), .ZN(
        n19808) );
  OAI211_X1 U22755 ( .C1(n19847), .C2(n19810), .A(n19809), .B(n19808), .ZN(
        P2_U3170) );
  AOI22_X1 U22756 ( .A1(n19839), .A2(n19812), .B1(n19276), .B2(n19811), .ZN(
        n19815) );
  AOI22_X1 U22757 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19826), .B1(
        n19843), .B2(n19813), .ZN(n19814) );
  OAI211_X1 U22758 ( .C1(n19816), .C2(n19829), .A(n19815), .B(n19814), .ZN(
        P2_U3171) );
  AOI22_X1 U22759 ( .A1(n19839), .A2(n19818), .B1(n19276), .B2(n19817), .ZN(
        n19821) );
  AOI22_X1 U22760 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19826), .B1(
        n19843), .B2(n19819), .ZN(n19820) );
  OAI211_X1 U22761 ( .C1(n19822), .C2(n19829), .A(n19821), .B(n19820), .ZN(
        P2_U3172) );
  AOI22_X1 U22762 ( .A1(n19839), .A2(n19824), .B1(n19276), .B2(n19823), .ZN(
        n19828) );
  AOI22_X1 U22763 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19826), .B1(
        n19843), .B2(n19825), .ZN(n19827) );
  OAI211_X1 U22764 ( .C1(n19830), .C2(n19829), .A(n19828), .B(n19827), .ZN(
        P2_U3173) );
  AOI22_X1 U22765 ( .A1(n19839), .A2(n19832), .B1(n19276), .B2(n19831), .ZN(
        n19836) );
  AOI22_X1 U22766 ( .A1(n19843), .A2(n19834), .B1(n19841), .B2(n19833), .ZN(
        n19835) );
  OAI211_X1 U22767 ( .C1(n19847), .C2(n13869), .A(n19836), .B(n19835), .ZN(
        P2_U3174) );
  INV_X1 U22768 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19846) );
  AOI22_X1 U22769 ( .A1(n19839), .A2(n19838), .B1(n19276), .B2(n19837), .ZN(
        n19845) );
  AOI22_X1 U22770 ( .A1(n19843), .A2(n19842), .B1(n19841), .B2(n19840), .ZN(
        n19844) );
  OAI211_X1 U22771 ( .C1(n19847), .C2(n19846), .A(n19845), .B(n19844), .ZN(
        P2_U3175) );
  OAI221_X1 U22772 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19979), .C1(
        P2_STATE2_REG_2__SCAN_IN), .C2(n19990), .A(n19848), .ZN(n19853) );
  OAI211_X1 U22773 ( .C1(n19850), .C2(n19849), .A(n19985), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19852) );
  OAI211_X1 U22774 ( .C1(n19854), .C2(n19853), .A(n19852), .B(n19851), .ZN(
        P2_U3177) );
  AND2_X1 U22775 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19928), .ZN(
        P2_U3179) );
  AND2_X1 U22776 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19928), .ZN(
        P2_U3180) );
  AND2_X1 U22777 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19928), .ZN(
        P2_U3181) );
  AND2_X1 U22778 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19928), .ZN(
        P2_U3182) );
  AND2_X1 U22779 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19928), .ZN(
        P2_U3183) );
  AND2_X1 U22780 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19928), .ZN(
        P2_U3184) );
  AND2_X1 U22781 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19928), .ZN(
        P2_U3185) );
  AND2_X1 U22782 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19928), .ZN(
        P2_U3186) );
  AND2_X1 U22783 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19928), .ZN(
        P2_U3187) );
  AND2_X1 U22784 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19928), .ZN(
        P2_U3188) );
  AND2_X1 U22785 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19928), .ZN(
        P2_U3189) );
  AND2_X1 U22786 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19928), .ZN(
        P2_U3190) );
  AND2_X1 U22787 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19928), .ZN(
        P2_U3191) );
  AND2_X1 U22788 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19928), .ZN(
        P2_U3192) );
  AND2_X1 U22789 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19928), .ZN(
        P2_U3193) );
  AND2_X1 U22790 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19928), .ZN(
        P2_U3194) );
  AND2_X1 U22791 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19928), .ZN(
        P2_U3195) );
  AND2_X1 U22792 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19928), .ZN(
        P2_U3196) );
  AND2_X1 U22793 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19928), .ZN(
        P2_U3197) );
  AND2_X1 U22794 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19928), .ZN(
        P2_U3198) );
  AND2_X1 U22795 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19928), .ZN(
        P2_U3199) );
  AND2_X1 U22796 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19928), .ZN(
        P2_U3200) );
  AND2_X1 U22797 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19928), .ZN(P2_U3201) );
  AND2_X1 U22798 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19928), .ZN(P2_U3202) );
  AND2_X1 U22799 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19928), .ZN(P2_U3203) );
  AND2_X1 U22800 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19928), .ZN(P2_U3204) );
  AND2_X1 U22801 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19928), .ZN(P2_U3205) );
  AND2_X1 U22802 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19928), .ZN(P2_U3206) );
  AND2_X1 U22803 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19928), .ZN(P2_U3207) );
  AND2_X1 U22804 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19928), .ZN(P2_U3208) );
  OAI21_X1 U22805 ( .B1(n20958), .B2(n19859), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19868) );
  INV_X1 U22806 ( .A(n19868), .ZN(n19857) );
  NAND2_X1 U22807 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19985), .ZN(n19866) );
  AND3_X1 U22808 ( .A1(n19866), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .A3(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19856) );
  INV_X1 U22809 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19996) );
  OAI211_X1 U22810 ( .C1(HOLD), .C2(n19996), .A(n19998), .B(n19863), .ZN(
        n19855) );
  OAI21_X1 U22811 ( .B1(n19857), .B2(n19856), .A(n19855), .ZN(P2_U3209) );
  AND2_X1 U22812 ( .A1(n19987), .A2(n19866), .ZN(n19861) );
  NOR2_X1 U22813 ( .A1(HOLD), .A2(n19858), .ZN(n19867) );
  OAI211_X1 U22814 ( .C1(n19867), .C2(n19869), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19859), .ZN(n19860) );
  OAI211_X1 U22815 ( .C1(n19862), .C2(n20976), .A(n19861), .B(n19860), .ZN(
        P2_U3210) );
  OAI22_X1 U22816 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19863), .B1(NA), 
        .B2(n19866), .ZN(n19864) );
  OAI211_X1 U22817 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19864), .ZN(n19865) );
  OAI221_X1 U22818 ( .B1(n19868), .B2(n19867), .C1(n19868), .C2(n19866), .A(
        n19865), .ZN(P2_U3211) );
  OAI222_X1 U22819 ( .A1(n19922), .A2(n19872), .B1(n19871), .B2(n19880), .C1(
        n19870), .C2(n19917), .ZN(P2_U3212) );
  OAI222_X1 U22820 ( .A1(n19922), .A2(n13432), .B1(n19873), .B2(n19880), .C1(
        n19872), .C2(n19917), .ZN(P2_U3213) );
  OAI222_X1 U22821 ( .A1(n19922), .A2(n12097), .B1(n19874), .B2(n19919), .C1(
        n13432), .C2(n19917), .ZN(P2_U3214) );
  OAI222_X1 U22822 ( .A1(n19922), .A2(n13692), .B1(n19875), .B2(n19880), .C1(
        n12097), .C2(n19917), .ZN(P2_U3215) );
  OAI222_X1 U22823 ( .A1(n19922), .A2(n19877), .B1(n19876), .B2(n19919), .C1(
        n13692), .C2(n19917), .ZN(P2_U3216) );
  OAI222_X1 U22824 ( .A1(n19922), .A2(n19879), .B1(n19878), .B2(n19880), .C1(
        n19877), .C2(n19917), .ZN(P2_U3217) );
  INV_X1 U22825 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19882) );
  OAI222_X1 U22826 ( .A1(n19922), .A2(n19882), .B1(n19881), .B2(n19880), .C1(
        n19879), .C2(n19917), .ZN(P2_U3218) );
  INV_X1 U22827 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19884) );
  OAI222_X1 U22828 ( .A1(n19922), .A2(n19884), .B1(n19883), .B2(n19880), .C1(
        n19882), .C2(n19917), .ZN(P2_U3219) );
  OAI222_X1 U22829 ( .A1(n19922), .A2(n19886), .B1(n19885), .B2(n19880), .C1(
        n19884), .C2(n19917), .ZN(P2_U3220) );
  OAI222_X1 U22830 ( .A1(n19922), .A2(n12219), .B1(n19887), .B2(n19880), .C1(
        n19886), .C2(n19917), .ZN(P2_U3221) );
  OAI222_X1 U22831 ( .A1(n19922), .A2(n12223), .B1(n19888), .B2(n19880), .C1(
        n12219), .C2(n19917), .ZN(P2_U3222) );
  OAI222_X1 U22832 ( .A1(n19922), .A2(n15297), .B1(n19889), .B2(n19880), .C1(
        n12223), .C2(n19917), .ZN(P2_U3223) );
  OAI222_X1 U22833 ( .A1(n19922), .A2(n13936), .B1(n19890), .B2(n19880), .C1(
        n15297), .C2(n19917), .ZN(P2_U3224) );
  OAI222_X1 U22834 ( .A1(n19922), .A2(n19892), .B1(n19891), .B2(n19880), .C1(
        n13936), .C2(n19917), .ZN(P2_U3225) );
  INV_X1 U22835 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19894) );
  OAI222_X1 U22836 ( .A1(n19922), .A2(n19894), .B1(n19893), .B2(n19880), .C1(
        n19892), .C2(n19917), .ZN(P2_U3226) );
  OAI222_X1 U22837 ( .A1(n19922), .A2(n19896), .B1(n19895), .B2(n19880), .C1(
        n19894), .C2(n19917), .ZN(P2_U3227) );
  OAI222_X1 U22838 ( .A1(n19922), .A2(n11972), .B1(n19897), .B2(n19880), .C1(
        n19896), .C2(n19917), .ZN(P2_U3228) );
  OAI222_X1 U22839 ( .A1(n19922), .A2(n19899), .B1(n19898), .B2(n19880), .C1(
        n11972), .C2(n19917), .ZN(P2_U3229) );
  OAI222_X1 U22840 ( .A1(n19922), .A2(n12240), .B1(n19900), .B2(n19919), .C1(
        n19899), .C2(n19917), .ZN(P2_U3230) );
  OAI222_X1 U22841 ( .A1(n19922), .A2(n11985), .B1(n19901), .B2(n19919), .C1(
        n12240), .C2(n19917), .ZN(P2_U3231) );
  OAI222_X1 U22842 ( .A1(n19922), .A2(n12243), .B1(n19902), .B2(n19919), .C1(
        n11985), .C2(n19917), .ZN(P2_U3232) );
  OAI222_X1 U22843 ( .A1(n19922), .A2(n19904), .B1(n19903), .B2(n19919), .C1(
        n12243), .C2(n19917), .ZN(P2_U3233) );
  INV_X1 U22844 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19906) );
  OAI222_X1 U22845 ( .A1(n19922), .A2(n19906), .B1(n19905), .B2(n19919), .C1(
        n19904), .C2(n19917), .ZN(P2_U3234) );
  OAI222_X1 U22846 ( .A1(n19922), .A2(n19908), .B1(n19907), .B2(n19919), .C1(
        n19906), .C2(n19917), .ZN(P2_U3235) );
  OAI222_X1 U22847 ( .A1(n19922), .A2(n19910), .B1(n19909), .B2(n19919), .C1(
        n19908), .C2(n19917), .ZN(P2_U3236) );
  OAI222_X1 U22848 ( .A1(n19922), .A2(n19913), .B1(n19911), .B2(n19919), .C1(
        n19910), .C2(n19917), .ZN(P2_U3237) );
  OAI222_X1 U22849 ( .A1(n19917), .A2(n19913), .B1(n19912), .B2(n19919), .C1(
        n15199), .C2(n19922), .ZN(P2_U3238) );
  OAI222_X1 U22850 ( .A1(n19922), .A2(n19915), .B1(n19914), .B2(n19919), .C1(
        n15199), .C2(n19917), .ZN(P2_U3239) );
  OAI222_X1 U22851 ( .A1(n19922), .A2(n19918), .B1(n19916), .B2(n19919), .C1(
        n19915), .C2(n19917), .ZN(P2_U3240) );
  INV_X1 U22852 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19920) );
  OAI222_X1 U22853 ( .A1(n19922), .A2(n19921), .B1(n19920), .B2(n19919), .C1(
        n19918), .C2(n19917), .ZN(P2_U3241) );
  OAI22_X1 U22854 ( .A1(n19998), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19880), .ZN(n19923) );
  INV_X1 U22855 ( .A(n19923), .ZN(P2_U3585) );
  MUX2_X1 U22856 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19998), .Z(P2_U3586) );
  OAI22_X1 U22857 ( .A1(n19998), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19880), .ZN(n19924) );
  INV_X1 U22858 ( .A(n19924), .ZN(P2_U3587) );
  OAI22_X1 U22859 ( .A1(n19998), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19880), .ZN(n19925) );
  INV_X1 U22860 ( .A(n19925), .ZN(P2_U3588) );
  AOI21_X1 U22861 ( .B1(n19928), .B2(n19927), .A(n19926), .ZN(P2_U3591) );
  OAI21_X1 U22862 ( .B1(n19931), .B2(n19930), .A(n19929), .ZN(P2_U3592) );
  AND2_X1 U22863 ( .A1(n19938), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19955) );
  NAND2_X1 U22864 ( .A1(n19932), .A2(n19955), .ZN(n19944) );
  NAND2_X1 U22865 ( .A1(n19953), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19934) );
  AOI21_X1 U22866 ( .B1(n19934), .B2(n19938), .A(n19933), .ZN(n19942) );
  NAND2_X1 U22867 ( .A1(n19944), .A2(n19942), .ZN(n19936) );
  AOI222_X1 U22868 ( .A1(n19939), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19938), 
        .B2(n19937), .C1(n19936), .C2(n19935), .ZN(n19940) );
  AOI22_X1 U22869 ( .A1(n19967), .A2(n19941), .B1(n19940), .B2(n19964), .ZN(
        P2_U3602) );
  INV_X1 U22870 ( .A(n19942), .ZN(n19947) );
  NOR2_X1 U22871 ( .A1(n19943), .A2(n19979), .ZN(n19946) );
  INV_X1 U22872 ( .A(n19944), .ZN(n19945) );
  AOI211_X1 U22873 ( .C1(n19948), .C2(n19947), .A(n19946), .B(n19945), .ZN(
        n19949) );
  AOI22_X1 U22874 ( .A1(n19967), .A2(n19950), .B1(n19949), .B2(n19964), .ZN(
        P2_U3603) );
  INV_X1 U22875 ( .A(n19951), .ZN(n19960) );
  NOR2_X1 U22876 ( .A1(n19960), .A2(n19952), .ZN(n19954) );
  MUX2_X1 U22877 ( .A(n19955), .B(n19954), .S(n19953), .Z(n19956) );
  AOI21_X1 U22878 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19957), .A(n19956), 
        .ZN(n19958) );
  AOI22_X1 U22879 ( .A1(n19967), .A2(n19959), .B1(n19958), .B2(n19964), .ZN(
        P2_U3604) );
  OAI22_X1 U22880 ( .A1(n19961), .A2(n19960), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19979), .ZN(n19962) );
  AOI21_X1 U22881 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19963), .A(n19962), 
        .ZN(n19965) );
  AOI22_X1 U22882 ( .A1(n19967), .A2(n19966), .B1(n19965), .B2(n19964), .ZN(
        P2_U3605) );
  INV_X1 U22883 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19968) );
  AOI22_X1 U22884 ( .A1(n19919), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19968), 
        .B2(n19998), .ZN(P2_U3608) );
  INV_X1 U22885 ( .A(n19969), .ZN(n19978) );
  AND2_X1 U22886 ( .A1(n19971), .A2(n19970), .ZN(n19973) );
  AOI211_X1 U22887 ( .C1(n19975), .C2(n19974), .A(n19973), .B(n19972), .ZN(
        n19977) );
  NAND2_X1 U22888 ( .A1(n19978), .A2(P2_MORE_REG_SCAN_IN), .ZN(n19976) );
  OAI21_X1 U22889 ( .B1(n19978), .B2(n19977), .A(n19976), .ZN(P2_U3609) );
  OAI21_X1 U22890 ( .B1(n19981), .B2(n19980), .A(n19979), .ZN(n19983) );
  OAI211_X1 U22891 ( .C1(n19985), .C2(n19984), .A(n19983), .B(n19982), .ZN(
        n19997) );
  OAI21_X1 U22892 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n19986), .ZN(n19994) );
  AOI21_X1 U22893 ( .B1(n19989), .B2(n19988), .A(n19987), .ZN(n19991) );
  OAI211_X1 U22894 ( .C1(n19992), .C2(n19991), .A(P2_STATE2_REG_2__SCAN_IN), 
        .B(n19990), .ZN(n19993) );
  NAND3_X1 U22895 ( .A1(n19997), .A2(n19994), .A3(n19993), .ZN(n19995) );
  OAI21_X1 U22896 ( .B1(n19997), .B2(n19996), .A(n19995), .ZN(P2_U3610) );
  OAI22_X1 U22897 ( .A1(n19998), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19880), .ZN(n19999) );
  INV_X1 U22898 ( .A(n19999), .ZN(P2_U3611) );
  AOI21_X1 U22899 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20745), .A(n20739), 
        .ZN(n20741) );
  INV_X1 U22900 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20977) );
  NAND2_X1 U22901 ( .A1(n20739), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20832) );
  INV_X1 U22902 ( .A(n20832), .ZN(n20831) );
  AOI21_X1 U22903 ( .B1(n20741), .B2(n20977), .A(n20831), .ZN(P1_U2802) );
  INV_X1 U22904 ( .A(n20000), .ZN(n20002) );
  OAI21_X1 U22905 ( .B1(n20002), .B2(n20001), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20003) );
  OAI21_X1 U22906 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20004), .A(n20003), 
        .ZN(P1_U2803) );
  INV_X1 U22907 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20946) );
  NOR2_X1 U22908 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20006) );
  NOR2_X1 U22909 ( .A1(n20831), .A2(n20006), .ZN(n20005) );
  AOI22_X1 U22910 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n20831), .B1(n20946), 
        .B2(n20005), .ZN(P1_U2804) );
  NOR2_X1 U22911 ( .A1(n20831), .A2(n20741), .ZN(n20794) );
  OAI21_X1 U22912 ( .B1(BS16), .B2(n20006), .A(n20794), .ZN(n20792) );
  OAI21_X1 U22913 ( .B1(n20794), .B2(n20974), .A(n20792), .ZN(P1_U2805) );
  OAI21_X1 U22914 ( .B1(n20008), .B2(n20968), .A(n20007), .ZN(P1_U2806) );
  NOR4_X1 U22915 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20012) );
  NOR4_X1 U22916 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20011) );
  NOR4_X1 U22917 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20010) );
  NOR4_X1 U22918 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20009) );
  NAND4_X1 U22919 ( .A1(n20012), .A2(n20011), .A3(n20010), .A4(n20009), .ZN(
        n20018) );
  NOR4_X1 U22920 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20016) );
  AOI211_X1 U22921 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20015) );
  NOR4_X1 U22922 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20014) );
  NOR4_X1 U22923 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20013) );
  NAND4_X1 U22924 ( .A1(n20016), .A2(n20015), .A3(n20014), .A4(n20013), .ZN(
        n20017) );
  NOR2_X1 U22925 ( .A1(n20018), .A2(n20017), .ZN(n20827) );
  INV_X1 U22926 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20020) );
  NOR3_X1 U22927 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20021) );
  OAI21_X1 U22928 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20021), .A(n20827), .ZN(
        n20019) );
  OAI21_X1 U22929 ( .B1(n20827), .B2(n20020), .A(n20019), .ZN(P1_U2807) );
  INV_X1 U22930 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20793) );
  AOI21_X1 U22931 ( .B1(n20824), .B2(n20793), .A(n20021), .ZN(n20022) );
  INV_X1 U22932 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20926) );
  INV_X1 U22933 ( .A(n20827), .ZN(n20829) );
  AOI22_X1 U22934 ( .A1(n20827), .A2(n20022), .B1(n20926), .B2(n20829), .ZN(
        P1_U2808) );
  AOI22_X1 U22935 ( .A1(n20049), .A2(n20023), .B1(n20077), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n20033) );
  INV_X1 U22936 ( .A(n20042), .ZN(n20081) );
  NOR2_X1 U22937 ( .A1(n20081), .A2(n20078), .ZN(n20066) );
  NAND2_X1 U22938 ( .A1(n20066), .A2(n20756), .ZN(n20025) );
  OAI22_X1 U22939 ( .A1(n20084), .A2(n20026), .B1(n20025), .B2(n20024), .ZN(
        n20027) );
  AOI211_X1 U22940 ( .C1(n20051), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n9645), .B(n20027), .ZN(n20032) );
  INV_X1 U22941 ( .A(n20028), .ZN(n20030) );
  AOI22_X1 U22942 ( .A1(n20030), .A2(n20055), .B1(P1_REIP_REG_8__SCAN_IN), 
        .B2(n20029), .ZN(n20031) );
  NAND3_X1 U22943 ( .A1(n20033), .A2(n20032), .A3(n20031), .ZN(P1_U2832) );
  INV_X1 U22944 ( .A(n20034), .ZN(n20035) );
  AOI22_X1 U22945 ( .A1(n20049), .A2(n20035), .B1(n20053), .B2(n20097), .ZN(
        n20046) );
  INV_X1 U22946 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20072) );
  NOR2_X1 U22947 ( .A1(n20754), .A2(n20072), .ZN(n20043) );
  INV_X1 U22948 ( .A(n20043), .ZN(n20036) );
  NOR2_X1 U22949 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20036), .ZN(n20040) );
  OAI22_X1 U22950 ( .A1(n20038), .A2(n20102), .B1(n20037), .B2(n20075), .ZN(
        n20039) );
  AOI21_X1 U22951 ( .B1(n20040), .B2(n20066), .A(n20039), .ZN(n20045) );
  AOI21_X1 U22952 ( .B1(n20042), .B2(n20078), .A(n20041), .ZN(n20096) );
  OAI21_X1 U22953 ( .B1(n20081), .B2(n20043), .A(n20096), .ZN(n20054) );
  AOI22_X1 U22954 ( .A1(n20100), .A2(n20055), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20054), .ZN(n20044) );
  NAND4_X1 U22955 ( .A1(n20046), .A2(n20045), .A3(n20044), .A4(n20073), .ZN(
        P1_U2833) );
  INV_X1 U22956 ( .A(n20047), .ZN(n20048) );
  AOI22_X1 U22957 ( .A1(n20049), .A2(n20048), .B1(n20077), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n20060) );
  NOR2_X1 U22958 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20072), .ZN(n20050) );
  AOI22_X1 U22959 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20051), .B1(
        n20066), .B2(n20050), .ZN(n20059) );
  AOI21_X1 U22960 ( .B1(n20053), .B2(n20052), .A(n9645), .ZN(n20058) );
  AOI22_X1 U22961 ( .A1(n20056), .A2(n20055), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20054), .ZN(n20057) );
  NAND4_X1 U22962 ( .A1(n20060), .A2(n20059), .A3(n20058), .A4(n20057), .ZN(
        P1_U2834) );
  INV_X1 U22963 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20062) );
  NAND2_X1 U22964 ( .A1(n20077), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n20061) );
  OAI211_X1 U22965 ( .C1(n20062), .C2(n20075), .A(n20061), .B(n20073), .ZN(
        n20065) );
  NOR2_X1 U22966 ( .A1(n20084), .A2(n20063), .ZN(n20064) );
  AOI211_X1 U22967 ( .C1(n20066), .C2(n20072), .A(n20065), .B(n20064), .ZN(
        n20067) );
  OAI21_X1 U22968 ( .B1(n20087), .B2(n20068), .A(n20067), .ZN(n20069) );
  AOI21_X1 U22969 ( .B1(n20070), .B2(n20092), .A(n20069), .ZN(n20071) );
  OAI21_X1 U22970 ( .B1(n20096), .B2(n20072), .A(n20071), .ZN(P1_U2835) );
  OAI21_X1 U22971 ( .B1(n20075), .B2(n20074), .A(n20073), .ZN(n20076) );
  AOI21_X1 U22972 ( .B1(n20077), .B2(P1_EBX_REG_4__SCAN_IN), .A(n20076), .ZN(
        n20083) );
  NAND3_X1 U22973 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20080) );
  INV_X1 U22974 ( .A(n20078), .ZN(n20079) );
  OR3_X1 U22975 ( .A1(n20081), .A2(n20080), .A3(n20079), .ZN(n20082) );
  OAI211_X1 U22976 ( .C1(n20085), .C2(n20084), .A(n20083), .B(n20082), .ZN(
        n20089) );
  NOR2_X1 U22977 ( .A1(n20087), .A2(n20086), .ZN(n20088) );
  AOI211_X1 U22978 ( .C1(n20091), .C2(n20090), .A(n20089), .B(n20088), .ZN(
        n20095) );
  NAND2_X1 U22979 ( .A1(n20093), .A2(n20092), .ZN(n20094) );
  OAI211_X1 U22980 ( .C1(n20096), .C2(n20748), .A(n20095), .B(n20094), .ZN(
        P1_U2836) );
  AOI22_X1 U22981 ( .A1(n20100), .A2(n20099), .B1(n20098), .B2(n20097), .ZN(
        n20101) );
  OAI21_X1 U22982 ( .B1(n20103), .B2(n20102), .A(n20101), .ZN(P1_U2865) );
  AOI22_X1 U22983 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20105) );
  OAI21_X1 U22984 ( .B1(n13040), .B2(n20132), .A(n20105), .ZN(P1_U2921) );
  AOI22_X1 U22985 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20106) );
  OAI21_X1 U22986 ( .B1(n14599), .B2(n20132), .A(n20106), .ZN(P1_U2922) );
  AOI22_X1 U22987 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20107) );
  OAI21_X1 U22988 ( .B1(n14601), .B2(n20132), .A(n20107), .ZN(P1_U2923) );
  AOI22_X1 U22989 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20108) );
  OAI21_X1 U22990 ( .B1(n14604), .B2(n20132), .A(n20108), .ZN(P1_U2924) );
  AOI22_X1 U22991 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20109) );
  OAI21_X1 U22992 ( .B1(n20110), .B2(n20132), .A(n20109), .ZN(P1_U2925) );
  INV_X1 U22993 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20112) );
  AOI22_X1 U22994 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20111) );
  OAI21_X1 U22995 ( .B1(n20112), .B2(n20132), .A(n20111), .ZN(P1_U2926) );
  AOI22_X1 U22996 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20120), .B1(n20129), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20113) );
  OAI21_X1 U22997 ( .B1(n13836), .B2(n20132), .A(n20113), .ZN(P1_U2927) );
  INV_X1 U22998 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20115) );
  AOI22_X1 U22999 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20120), .B1(n20129), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20114) );
  OAI21_X1 U23000 ( .B1(n20115), .B2(n20132), .A(n20114), .ZN(P1_U2928) );
  AOI22_X1 U23001 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20120), .B1(n20129), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20116) );
  OAI21_X1 U23002 ( .B1(n20117), .B2(n20132), .A(n20116), .ZN(P1_U2929) );
  AOI22_X1 U23003 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20120), .B1(n20129), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20118) );
  OAI21_X1 U23004 ( .B1(n10645), .B2(n20132), .A(n20118), .ZN(P1_U2930) );
  AOI22_X1 U23005 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20120), .B1(n20129), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20119) );
  OAI21_X1 U23006 ( .B1(n10634), .B2(n20132), .A(n20119), .ZN(P1_U2931) );
  INV_X1 U23007 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U23008 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20120), .B1(n20129), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20121) );
  OAI21_X1 U23009 ( .B1(n20122), .B2(n20132), .A(n20121), .ZN(P1_U2932) );
  AOI22_X1 U23010 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20123) );
  OAI21_X1 U23011 ( .B1(n20124), .B2(n20132), .A(n20123), .ZN(P1_U2933) );
  AOI22_X1 U23012 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20125) );
  OAI21_X1 U23013 ( .B1(n20126), .B2(n20132), .A(n20125), .ZN(P1_U2934) );
  AOI22_X1 U23014 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20127) );
  OAI21_X1 U23015 ( .B1(n20128), .B2(n20132), .A(n20127), .ZN(P1_U2935) );
  AOI22_X1 U23016 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20130), .B1(n20129), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20131) );
  OAI21_X1 U23017 ( .B1(n20133), .B2(n20132), .A(n20131), .ZN(P1_U2936) );
  AOI22_X1 U23018 ( .A1(n20161), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n9650), .ZN(n20135) );
  NAND2_X1 U23019 ( .A1(n20149), .A2(n20134), .ZN(n20151) );
  NAND2_X1 U23020 ( .A1(n20135), .A2(n20151), .ZN(P1_U2945) );
  AOI22_X1 U23021 ( .A1(n20161), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n9650), .ZN(n20138) );
  INV_X1 U23022 ( .A(n20136), .ZN(n20137) );
  NAND2_X1 U23023 ( .A1(n20149), .A2(n20137), .ZN(n20153) );
  NAND2_X1 U23024 ( .A1(n20138), .A2(n20153), .ZN(P1_U2946) );
  AOI22_X1 U23025 ( .A1(n20161), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n9650), .ZN(n20140) );
  NAND2_X1 U23026 ( .A1(n20149), .A2(n20139), .ZN(n20155) );
  NAND2_X1 U23027 ( .A1(n20140), .A2(n20155), .ZN(P1_U2947) );
  AOI22_X1 U23028 ( .A1(n20161), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n9650), .ZN(n20143) );
  INV_X1 U23029 ( .A(n20141), .ZN(n20142) );
  NAND2_X1 U23030 ( .A1(n20149), .A2(n20142), .ZN(n20157) );
  NAND2_X1 U23031 ( .A1(n20143), .A2(n20157), .ZN(P1_U2949) );
  AOI22_X1 U23032 ( .A1(n20161), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n9650), .ZN(n20146) );
  INV_X1 U23033 ( .A(n20144), .ZN(n20145) );
  NAND2_X1 U23034 ( .A1(n20149), .A2(n20145), .ZN(n20159) );
  NAND2_X1 U23035 ( .A1(n20146), .A2(n20159), .ZN(P1_U2950) );
  AOI22_X1 U23036 ( .A1(n20161), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n9650), .ZN(n20150) );
  INV_X1 U23037 ( .A(n20147), .ZN(n20148) );
  NAND2_X1 U23038 ( .A1(n20149), .A2(n20148), .ZN(n20162) );
  NAND2_X1 U23039 ( .A1(n20150), .A2(n20162), .ZN(P1_U2951) );
  AOI22_X1 U23040 ( .A1(n20161), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n9650), .ZN(n20152) );
  NAND2_X1 U23041 ( .A1(n20152), .A2(n20151), .ZN(P1_U2960) );
  AOI22_X1 U23042 ( .A1(n20161), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n9650), .ZN(n20154) );
  NAND2_X1 U23043 ( .A1(n20154), .A2(n20153), .ZN(P1_U2961) );
  AOI22_X1 U23044 ( .A1(n20161), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n9650), .ZN(n20156) );
  NAND2_X1 U23045 ( .A1(n20156), .A2(n20155), .ZN(P1_U2962) );
  AOI22_X1 U23046 ( .A1(n20161), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n9650), .ZN(n20158) );
  NAND2_X1 U23047 ( .A1(n20158), .A2(n20157), .ZN(P1_U2964) );
  AOI22_X1 U23048 ( .A1(n20161), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n9650), .ZN(n20160) );
  NAND2_X1 U23049 ( .A1(n20160), .A2(n20159), .ZN(P1_U2965) );
  AOI22_X1 U23050 ( .A1(n20161), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n9650), .ZN(n20163) );
  NAND2_X1 U23051 ( .A1(n20163), .A2(n20162), .ZN(P1_U2966) );
  NOR2_X1 U23052 ( .A1(n20165), .A2(n20164), .ZN(n20177) );
  NOR3_X1 U23053 ( .A1(n20168), .A2(n20167), .A3(n20166), .ZN(n20176) );
  INV_X1 U23054 ( .A(n20169), .ZN(n20175) );
  INV_X1 U23055 ( .A(n20170), .ZN(n20171) );
  OAI21_X1 U23056 ( .B1(n20173), .B2(n20172), .A(n20171), .ZN(n20174) );
  NOR4_X1 U23057 ( .A1(n20177), .A2(n20176), .A3(n20175), .A4(n20174), .ZN(
        n20178) );
  OAI221_X1 U23058 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20181), .C1(
        n20180), .C2(n20179), .A(n20178), .ZN(P1_U3029) );
  NOR2_X1 U23059 ( .A1(n20182), .A2(n20823), .ZN(P1_U3032) );
  INV_X1 U23060 ( .A(DATAI_24_), .ZN(n20939) );
  OAI22_X2 U23061 ( .A1(n20939), .A2(n20221), .B1(n20183), .B2(n20222), .ZN(
        n20673) );
  NOR2_X2 U23062 ( .A1(n20225), .A2(n20184), .ZN(n20666) );
  AOI22_X1 U23063 ( .A1(n20710), .A2(n20673), .B1(n20226), .B2(n20666), .ZN(
        n20188) );
  INV_X1 U23064 ( .A(DATAI_16_), .ZN(n20930) );
  OAI22_X1 U23065 ( .A1(n20186), .A2(n20222), .B1(n20930), .B2(n20221), .ZN(
        n20595) );
  AOI22_X1 U23066 ( .A1(n20665), .A2(n20229), .B1(n20257), .B2(n20595), .ZN(
        n20187) );
  OAI211_X1 U23067 ( .C1(n20227), .C2(n20189), .A(n20188), .B(n20187), .ZN(
        P1_U3033) );
  INV_X1 U23068 ( .A(DATAI_25_), .ZN(n20191) );
  OAI22_X2 U23069 ( .A1(n20191), .A2(n20221), .B1(n20190), .B2(n20222), .ZN(
        n20635) );
  NOR2_X2 U23070 ( .A1(n20225), .A2(n20192), .ZN(n20678) );
  AOI22_X1 U23071 ( .A1(n20710), .A2(n20635), .B1(n20226), .B2(n20678), .ZN(
        n20197) );
  INV_X1 U23072 ( .A(DATAI_17_), .ZN(n20194) );
  AOI22_X1 U23073 ( .A1(n20677), .A2(n20229), .B1(n20257), .B2(n20679), .ZN(
        n20196) );
  OAI211_X1 U23074 ( .C1(n20227), .C2(n10323), .A(n20197), .B(n20196), .ZN(
        P1_U3034) );
  INV_X1 U23075 ( .A(DATAI_26_), .ZN(n20957) );
  OAI22_X2 U23076 ( .A1(n20198), .A2(n20222), .B1(n20957), .B2(n20221), .ZN(
        n20685) );
  NOR2_X2 U23077 ( .A1(n20225), .A2(n10359), .ZN(n20684) );
  AOI22_X1 U23078 ( .A1(n20710), .A2(n20685), .B1(n20226), .B2(n20684), .ZN(
        n20202) );
  INV_X1 U23079 ( .A(DATAI_18_), .ZN(n20947) );
  OAI22_X1 U23080 ( .A1(n20200), .A2(n20222), .B1(n20947), .B2(n20221), .ZN(
        n20601) );
  AOI22_X1 U23081 ( .A1(n20683), .A2(n20229), .B1(n20257), .B2(n20601), .ZN(
        n20201) );
  OAI211_X1 U23082 ( .C1(n20227), .C2(n20203), .A(n20202), .B(n20201), .ZN(
        P1_U3035) );
  INV_X1 U23083 ( .A(DATAI_27_), .ZN(n20888) );
  OAI22_X2 U23084 ( .A1(n20204), .A2(n20222), .B1(n20888), .B2(n20221), .ZN(
        n20691) );
  NOR2_X2 U23085 ( .A1(n20225), .A2(n20205), .ZN(n20690) );
  AOI22_X1 U23086 ( .A1(n20710), .A2(n20691), .B1(n20226), .B2(n20690), .ZN(
        n20210) );
  INV_X1 U23087 ( .A(DATAI_19_), .ZN(n20207) );
  OAI22_X1 U23088 ( .A1(n20208), .A2(n20222), .B1(n20207), .B2(n20221), .ZN(
        n20605) );
  AOI22_X1 U23089 ( .A1(n20689), .A2(n20229), .B1(n20257), .B2(n20605), .ZN(
        n20209) );
  OAI211_X1 U23090 ( .C1(n20227), .C2(n20211), .A(n20210), .B(n20209), .ZN(
        P1_U3036) );
  OAI22_X2 U23091 ( .A1(n20212), .A2(n20222), .B1(n14534), .B2(n20221), .ZN(
        n20647) );
  NOR2_X2 U23092 ( .A1(n20225), .A2(n20213), .ZN(n20701) );
  AOI22_X1 U23093 ( .A1(n20710), .A2(n20647), .B1(n20226), .B2(n20701), .ZN(
        n20217) );
  AOI22_X1 U23094 ( .A1(n20702), .A2(n20229), .B1(n20257), .B2(n20703), .ZN(
        n20216) );
  OAI211_X1 U23095 ( .C1(n20227), .C2(n20218), .A(n20217), .B(n20216), .ZN(
        P1_U3038) );
  INV_X1 U23096 ( .A(DATAI_23_), .ZN(n20220) );
  OAI22_X1 U23097 ( .A1(n20220), .A2(n20221), .B1(n20219), .B2(n20222), .ZN(
        n20617) );
  INV_X1 U23098 ( .A(n20617), .ZN(n20725) );
  INV_X1 U23099 ( .A(DATAI_31_), .ZN(n20973) );
  OAI22_X2 U23100 ( .A1(n20223), .A2(n20222), .B1(n20973), .B2(n20221), .ZN(
        n20719) );
  NOR2_X2 U23101 ( .A1(n20225), .A2(n20224), .ZN(n20716) );
  AOI22_X1 U23102 ( .A1(n20710), .A2(n20719), .B1(n20226), .B2(n20716), .ZN(
        n20232) );
  INV_X1 U23103 ( .A(n20227), .ZN(n20230) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20230), .B1(
        n20718), .B2(n20229), .ZN(n20231) );
  OAI211_X1 U23105 ( .C1(n20725), .C2(n20233), .A(n20232), .B(n20231), .ZN(
        P1_U3040) );
  INV_X1 U23106 ( .A(n20595), .ZN(n20676) );
  OR2_X1 U23107 ( .A1(n9656), .A2(n20261), .ZN(n20594) );
  NOR2_X1 U23108 ( .A1(n20588), .A2(n20236), .ZN(n20255) );
  INV_X1 U23109 ( .A(n20293), .ZN(n20235) );
  INV_X1 U23110 ( .A(n20234), .ZN(n20590) );
  AOI21_X1 U23111 ( .B1(n20235), .B2(n20590), .A(n20255), .ZN(n20237) );
  OAI22_X1 U23112 ( .A1(n20237), .A2(n20664), .B1(n20236), .B2(n20728), .ZN(
        n20256) );
  AOI22_X1 U23113 ( .A1(n20666), .A2(n20255), .B1(n20256), .B2(n20665), .ZN(
        n20241) );
  OAI21_X1 U23114 ( .B1(n20302), .B2(n20974), .A(n20237), .ZN(n20238) );
  OAI221_X1 U23115 ( .B1(n20671), .B2(n20239), .C1(n20664), .C2(n20238), .A(
        n20670), .ZN(n20258) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20673), .ZN(n20240) );
  OAI211_X1 U23117 ( .C1(n20676), .C2(n20262), .A(n20241), .B(n20240), .ZN(
        P1_U3041) );
  INV_X1 U23118 ( .A(n20679), .ZN(n20638) );
  AOI22_X1 U23119 ( .A1(n20678), .A2(n20255), .B1(n20256), .B2(n20677), .ZN(
        n20243) );
  AOI22_X1 U23120 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20635), .ZN(n20242) );
  OAI211_X1 U23121 ( .C1(n20638), .C2(n20262), .A(n20243), .B(n20242), .ZN(
        P1_U3042) );
  INV_X1 U23122 ( .A(n20601), .ZN(n20688) );
  AOI22_X1 U23123 ( .A1(n20684), .A2(n20255), .B1(n20256), .B2(n20683), .ZN(
        n20245) );
  AOI22_X1 U23124 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20685), .ZN(n20244) );
  OAI211_X1 U23125 ( .C1(n20688), .C2(n20262), .A(n20245), .B(n20244), .ZN(
        P1_U3043) );
  INV_X1 U23126 ( .A(n20605), .ZN(n20694) );
  AOI22_X1 U23127 ( .A1(n20690), .A2(n20255), .B1(n20256), .B2(n20689), .ZN(
        n20247) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20691), .ZN(n20246) );
  OAI211_X1 U23129 ( .C1(n20694), .C2(n20262), .A(n20247), .B(n20246), .ZN(
        P1_U3044) );
  AOI22_X1 U23130 ( .A1(n20696), .A2(n20255), .B1(n20695), .B2(n20256), .ZN(
        n20250) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20643), .ZN(n20249) );
  OAI211_X1 U23132 ( .C1(n20646), .C2(n20262), .A(n20250), .B(n20249), .ZN(
        P1_U3045) );
  INV_X1 U23133 ( .A(n20703), .ZN(n20650) );
  AOI22_X1 U23134 ( .A1(n20702), .A2(n20256), .B1(n20701), .B2(n20255), .ZN(
        n20252) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20647), .ZN(n20251) );
  OAI211_X1 U23136 ( .C1(n20650), .C2(n20262), .A(n20252), .B(n20251), .ZN(
        P1_U3046) );
  AOI22_X1 U23137 ( .A1(n20708), .A2(n20256), .B1(n20707), .B2(n20255), .ZN(
        n20254) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20651), .ZN(n20253) );
  OAI211_X1 U23139 ( .C1(n9779), .C2(n20262), .A(n20254), .B(n20253), .ZN(
        P1_U3047) );
  AOI22_X1 U23140 ( .A1(n20718), .A2(n20256), .B1(n20716), .B2(n20255), .ZN(
        n20260) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20719), .ZN(n20259) );
  OAI211_X1 U23142 ( .C1(n20725), .C2(n20262), .A(n20260), .B(n20259), .ZN(
        P1_U3048) );
  NOR3_X1 U23143 ( .A1(n20318), .A2(n20285), .A3(n20664), .ZN(n20263) );
  INV_X1 U23144 ( .A(n20484), .ZN(n20815) );
  NOR2_X1 U23145 ( .A1(n20263), .A2(n20815), .ZN(n20269) );
  INV_X1 U23146 ( .A(n20269), .ZN(n20264) );
  NOR2_X1 U23147 ( .A1(n20293), .A2(n9637), .ZN(n20268) );
  INV_X1 U23148 ( .A(n20665), .ZN(n20561) );
  NOR3_X1 U23149 ( .A1(n20489), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20297) );
  NAND2_X1 U23150 ( .A1(n20588), .A2(n20297), .ZN(n20266) );
  INV_X1 U23151 ( .A(n20266), .ZN(n20284) );
  AOI22_X1 U23152 ( .A1(n20285), .A2(n20673), .B1(n20666), .B2(n20284), .ZN(
        n20271) );
  NOR2_X1 U23153 ( .A1(n10245), .A2(n20728), .ZN(n20379) );
  AOI211_X1 U23154 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20266), .A(n20379), 
        .B(n20265), .ZN(n20267) );
  AOI22_X1 U23155 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20286), .B1(
        n20318), .B2(n20595), .ZN(n20270) );
  OAI211_X1 U23156 ( .C1(n20289), .C2(n20561), .A(n20271), .B(n20270), .ZN(
        P1_U3049) );
  INV_X1 U23157 ( .A(n20677), .ZN(n20564) );
  AOI22_X1 U23158 ( .A1(n20318), .A2(n20679), .B1(n20678), .B2(n20284), .ZN(
        n20273) );
  AOI22_X1 U23159 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n20635), .ZN(n20272) );
  OAI211_X1 U23160 ( .C1(n20289), .C2(n20564), .A(n20273), .B(n20272), .ZN(
        P1_U3050) );
  INV_X1 U23161 ( .A(n20683), .ZN(n20567) );
  AOI22_X1 U23162 ( .A1(n20285), .A2(n20685), .B1(n20684), .B2(n20284), .ZN(
        n20275) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20286), .B1(
        n20318), .B2(n20601), .ZN(n20274) );
  OAI211_X1 U23164 ( .C1(n20289), .C2(n20567), .A(n20275), .B(n20274), .ZN(
        P1_U3051) );
  INV_X1 U23165 ( .A(n20689), .ZN(n20570) );
  AOI22_X1 U23166 ( .A1(n20285), .A2(n20691), .B1(n20690), .B2(n20284), .ZN(
        n20277) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20286), .B1(
        n20318), .B2(n20605), .ZN(n20276) );
  OAI211_X1 U23168 ( .C1(n20289), .C2(n20570), .A(n20277), .B(n20276), .ZN(
        P1_U3052) );
  INV_X1 U23169 ( .A(n20695), .ZN(n20573) );
  AOI22_X1 U23170 ( .A1(n20318), .A2(n20697), .B1(n20696), .B2(n20284), .ZN(
        n20279) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n20643), .ZN(n20278) );
  OAI211_X1 U23172 ( .C1(n20289), .C2(n20573), .A(n20279), .B(n20278), .ZN(
        P1_U3053) );
  INV_X1 U23173 ( .A(n20702), .ZN(n20576) );
  AOI22_X1 U23174 ( .A1(n20318), .A2(n20703), .B1(n20701), .B2(n20284), .ZN(
        n20281) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n20647), .ZN(n20280) );
  OAI211_X1 U23176 ( .C1(n20289), .C2(n20576), .A(n20281), .B(n20280), .ZN(
        P1_U3054) );
  INV_X1 U23177 ( .A(n20708), .ZN(n20579) );
  AOI22_X1 U23178 ( .A1(n20285), .A2(n20651), .B1(n20707), .B2(n20284), .ZN(
        n20283) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20286), .B1(
        n20318), .B2(n9780), .ZN(n20282) );
  OAI211_X1 U23180 ( .C1(n20289), .C2(n20579), .A(n20283), .B(n20282), .ZN(
        P1_U3055) );
  INV_X1 U23181 ( .A(n20718), .ZN(n20586) );
  AOI22_X1 U23182 ( .A1(n20285), .A2(n20719), .B1(n20716), .B2(n20284), .ZN(
        n20288) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20286), .B1(
        n20318), .B2(n20617), .ZN(n20287) );
  OAI211_X1 U23184 ( .C1(n20289), .C2(n20586), .A(n20288), .B(n20287), .ZN(
        P1_U3056) );
  INV_X1 U23185 ( .A(n20302), .ZN(n20290) );
  AOI21_X1 U23186 ( .B1(n20290), .B2(n20523), .A(n20664), .ZN(n20299) );
  AND2_X1 U23187 ( .A1(n20291), .A2(n9664), .ZN(n20661) );
  INV_X1 U23188 ( .A(n20661), .ZN(n20292) );
  OR2_X1 U23189 ( .A1(n20293), .A2(n20292), .ZN(n20295) );
  NOR2_X1 U23190 ( .A1(n20520), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20317) );
  INV_X1 U23191 ( .A(n20317), .ZN(n20294) );
  AND2_X1 U23192 ( .A1(n20295), .A2(n20294), .ZN(n20300) );
  INV_X1 U23193 ( .A(n20300), .ZN(n20296) );
  AOI22_X1 U23194 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20297), .B1(n20299), 
        .B2(n20296), .ZN(n20322) );
  AOI22_X1 U23195 ( .A1(n20318), .A2(n20673), .B1(n20666), .B2(n20317), .ZN(
        n20304) );
  OAI21_X1 U23196 ( .B1(n20671), .B2(n20297), .A(n20670), .ZN(n20298) );
  AOI21_X1 U23197 ( .B1(n20300), .B2(n20299), .A(n20298), .ZN(n20301) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20319), .B1(
        n20348), .B2(n20595), .ZN(n20303) );
  OAI211_X1 U23199 ( .C1(n20322), .C2(n20561), .A(n20304), .B(n20303), .ZN(
        P1_U3057) );
  AOI22_X1 U23200 ( .A1(n20318), .A2(n20635), .B1(n20678), .B2(n20317), .ZN(
        n20306) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20319), .B1(
        n20348), .B2(n20679), .ZN(n20305) );
  OAI211_X1 U23202 ( .C1(n20322), .C2(n20564), .A(n20306), .B(n20305), .ZN(
        P1_U3058) );
  AOI22_X1 U23203 ( .A1(n20348), .A2(n20601), .B1(n20684), .B2(n20317), .ZN(
        n20308) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20685), .ZN(n20307) );
  OAI211_X1 U23205 ( .C1(n20322), .C2(n20567), .A(n20308), .B(n20307), .ZN(
        P1_U3059) );
  AOI22_X1 U23206 ( .A1(n20348), .A2(n20605), .B1(n20690), .B2(n20317), .ZN(
        n20310) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20691), .ZN(n20309) );
  OAI211_X1 U23208 ( .C1(n20322), .C2(n20570), .A(n20310), .B(n20309), .ZN(
        P1_U3060) );
  AOI22_X1 U23209 ( .A1(n20348), .A2(n20697), .B1(n20696), .B2(n20317), .ZN(
        n20312) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20643), .ZN(n20311) );
  OAI211_X1 U23211 ( .C1(n20322), .C2(n20573), .A(n20312), .B(n20311), .ZN(
        P1_U3061) );
  AOI22_X1 U23212 ( .A1(n20348), .A2(n20703), .B1(n20701), .B2(n20317), .ZN(
        n20314) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20647), .ZN(n20313) );
  OAI211_X1 U23214 ( .C1(n20322), .C2(n20576), .A(n20314), .B(n20313), .ZN(
        P1_U3062) );
  AOI22_X1 U23215 ( .A1(n20318), .A2(n20651), .B1(n20707), .B2(n20317), .ZN(
        n20316) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20319), .B1(
        n20348), .B2(n9780), .ZN(n20315) );
  OAI211_X1 U23217 ( .C1(n20322), .C2(n20579), .A(n20316), .B(n20315), .ZN(
        P1_U3063) );
  AOI22_X1 U23218 ( .A1(n20348), .A2(n20617), .B1(n20716), .B2(n20317), .ZN(
        n20321) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20719), .ZN(n20320) );
  OAI211_X1 U23220 ( .C1(n20322), .C2(n20586), .A(n20321), .B(n20320), .ZN(
        P1_U3064) );
  INV_X1 U23221 ( .A(n20408), .ZN(n20324) );
  NOR3_X1 U23222 ( .A1(n11119), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20355) );
  INV_X1 U23223 ( .A(n20355), .ZN(n20352) );
  NOR2_X1 U23224 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20352), .ZN(
        n20346) );
  NOR2_X1 U23225 ( .A1(n13095), .A2(n20325), .ZN(n20405) );
  NAND2_X1 U23226 ( .A1(n20405), .A2(n9637), .ZN(n20328) );
  INV_X1 U23227 ( .A(n20552), .ZN(n20626) );
  OAI22_X1 U23228 ( .A1(n20328), .A2(n20664), .B1(n20626), .B2(n20326), .ZN(
        n20347) );
  AOI22_X1 U23229 ( .A1(n20666), .A2(n20346), .B1(n20665), .B2(n20347), .ZN(
        n20333) );
  INV_X1 U23230 ( .A(n20375), .ZN(n20327) );
  OAI21_X1 U23231 ( .B1(n20348), .B2(n20327), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20329) );
  AOI21_X1 U23232 ( .B1(n20329), .B2(n20328), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20331) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20673), .ZN(n20332) );
  OAI211_X1 U23234 ( .C1(n20676), .C2(n20375), .A(n20333), .B(n20332), .ZN(
        P1_U3065) );
  AOI22_X1 U23235 ( .A1(n20678), .A2(n20346), .B1(n20677), .B2(n20347), .ZN(
        n20335) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20635), .ZN(n20334) );
  OAI211_X1 U23237 ( .C1(n20638), .C2(n20375), .A(n20335), .B(n20334), .ZN(
        P1_U3066) );
  AOI22_X1 U23238 ( .A1(n20684), .A2(n20346), .B1(n20683), .B2(n20347), .ZN(
        n20337) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20685), .ZN(n20336) );
  OAI211_X1 U23240 ( .C1(n20688), .C2(n20375), .A(n20337), .B(n20336), .ZN(
        P1_U3067) );
  AOI22_X1 U23241 ( .A1(n20690), .A2(n20346), .B1(n20689), .B2(n20347), .ZN(
        n20339) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20691), .ZN(n20338) );
  OAI211_X1 U23243 ( .C1(n20694), .C2(n20375), .A(n20339), .B(n20338), .ZN(
        P1_U3068) );
  AOI22_X1 U23244 ( .A1(n20696), .A2(n20346), .B1(n20695), .B2(n20347), .ZN(
        n20341) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20643), .ZN(n20340) );
  OAI211_X1 U23246 ( .C1(n20646), .C2(n20375), .A(n20341), .B(n20340), .ZN(
        P1_U3069) );
  AOI22_X1 U23247 ( .A1(n20702), .A2(n20347), .B1(n20701), .B2(n20346), .ZN(
        n20343) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20647), .ZN(n20342) );
  OAI211_X1 U23249 ( .C1(n20650), .C2(n20375), .A(n20343), .B(n20342), .ZN(
        P1_U3070) );
  AOI22_X1 U23250 ( .A1(n20708), .A2(n20347), .B1(n20707), .B2(n20346), .ZN(
        n20345) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20651), .ZN(n20344) );
  OAI211_X1 U23252 ( .C1(n9779), .C2(n20375), .A(n20345), .B(n20344), .ZN(
        P1_U3071) );
  AOI22_X1 U23253 ( .A1(n20718), .A2(n20347), .B1(n20716), .B2(n20346), .ZN(
        n20351) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20719), .ZN(n20350) );
  OAI211_X1 U23255 ( .C1(n20725), .C2(n20375), .A(n20351), .B(n20350), .ZN(
        P1_U3072) );
  INV_X1 U23256 ( .A(n20673), .ZN(n20598) );
  NOR2_X1 U23257 ( .A1(n20588), .A2(n20352), .ZN(n20370) );
  AOI21_X1 U23258 ( .B1(n20405), .B2(n20590), .A(n20370), .ZN(n20353) );
  OAI22_X1 U23259 ( .A1(n20353), .A2(n20664), .B1(n20352), .B2(n20728), .ZN(
        n20371) );
  AOI22_X1 U23260 ( .A1(n20666), .A2(n20370), .B1(n20665), .B2(n20371), .ZN(
        n20357) );
  OAI21_X1 U23261 ( .B1(n20408), .B2(n20974), .A(n20353), .ZN(n20354) );
  OAI221_X1 U23262 ( .B1(n20671), .B2(n20355), .C1(n20664), .C2(n20354), .A(
        n20670), .ZN(n20372) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20372), .B1(
        n20399), .B2(n20595), .ZN(n20356) );
  OAI211_X1 U23264 ( .C1(n20598), .C2(n20375), .A(n20357), .B(n20356), .ZN(
        P1_U3073) );
  INV_X1 U23265 ( .A(n20635), .ZN(n20682) );
  AOI22_X1 U23266 ( .A1(n20678), .A2(n20370), .B1(n20677), .B2(n20371), .ZN(
        n20359) );
  AOI22_X1 U23267 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20372), .B1(
        n20399), .B2(n20679), .ZN(n20358) );
  OAI211_X1 U23268 ( .C1(n20682), .C2(n20375), .A(n20359), .B(n20358), .ZN(
        P1_U3074) );
  INV_X1 U23269 ( .A(n20685), .ZN(n20604) );
  AOI22_X1 U23270 ( .A1(n20684), .A2(n20370), .B1(n20683), .B2(n20371), .ZN(
        n20361) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20372), .B1(
        n20399), .B2(n20601), .ZN(n20360) );
  OAI211_X1 U23272 ( .C1(n20604), .C2(n20375), .A(n20361), .B(n20360), .ZN(
        P1_U3075) );
  INV_X1 U23273 ( .A(n20691), .ZN(n20608) );
  AOI22_X1 U23274 ( .A1(n20690), .A2(n20370), .B1(n20689), .B2(n20371), .ZN(
        n20363) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20372), .B1(
        n20399), .B2(n20605), .ZN(n20362) );
  OAI211_X1 U23276 ( .C1(n20608), .C2(n20375), .A(n20363), .B(n20362), .ZN(
        P1_U3076) );
  INV_X1 U23277 ( .A(n20643), .ZN(n20700) );
  AOI22_X1 U23278 ( .A1(n20696), .A2(n20370), .B1(n20695), .B2(n20371), .ZN(
        n20365) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20372), .B1(
        n20399), .B2(n20697), .ZN(n20364) );
  OAI211_X1 U23280 ( .C1(n20700), .C2(n20375), .A(n20365), .B(n20364), .ZN(
        P1_U3077) );
  INV_X1 U23281 ( .A(n20647), .ZN(n20706) );
  AOI22_X1 U23282 ( .A1(n20702), .A2(n20371), .B1(n20701), .B2(n20370), .ZN(
        n20367) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20372), .B1(
        n20399), .B2(n20703), .ZN(n20366) );
  OAI211_X1 U23284 ( .C1(n20706), .C2(n20375), .A(n20367), .B(n20366), .ZN(
        P1_U3078) );
  AOI22_X1 U23285 ( .A1(n20708), .A2(n20371), .B1(n20707), .B2(n20370), .ZN(
        n20369) );
  AOI22_X1 U23286 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20372), .B1(
        n20399), .B2(n9780), .ZN(n20368) );
  OAI211_X1 U23287 ( .C1(n20714), .C2(n20375), .A(n20369), .B(n20368), .ZN(
        P1_U3079) );
  INV_X1 U23288 ( .A(n20719), .ZN(n20622) );
  AOI22_X1 U23289 ( .A1(n20718), .A2(n20371), .B1(n20716), .B2(n20370), .ZN(
        n20374) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20372), .B1(
        n20399), .B2(n20617), .ZN(n20373) );
  OAI211_X1 U23291 ( .C1(n20622), .C2(n20375), .A(n20374), .B(n20373), .ZN(
        P1_U3080) );
  NAND3_X1 U23292 ( .A1(n20383), .A2(n20376), .A3(n20671), .ZN(n20377) );
  NAND2_X1 U23293 ( .A1(n20377), .A2(n20484), .ZN(n20381) );
  AND2_X1 U23294 ( .A1(n20405), .A2(n20625), .ZN(n20378) );
  NOR2_X1 U23295 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20409), .ZN(
        n20398) );
  AOI22_X1 U23296 ( .A1(n20399), .A2(n20673), .B1(n20666), .B2(n20398), .ZN(
        n20385) );
  INV_X1 U23297 ( .A(n20378), .ZN(n20380) );
  AOI21_X1 U23298 ( .B1(n20381), .B2(n20380), .A(n20379), .ZN(n20382) );
  OAI211_X1 U23299 ( .C1(n20398), .C2(n13115), .A(n20631), .B(n20382), .ZN(
        n20400) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20400), .B1(
        n20426), .B2(n20595), .ZN(n20384) );
  OAI211_X1 U23301 ( .C1(n20403), .C2(n20561), .A(n20385), .B(n20384), .ZN(
        P1_U3081) );
  AOI22_X1 U23302 ( .A1(n20399), .A2(n20635), .B1(n20678), .B2(n20398), .ZN(
        n20387) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20400), .B1(
        n20426), .B2(n20679), .ZN(n20386) );
  OAI211_X1 U23304 ( .C1(n20403), .C2(n20564), .A(n20387), .B(n20386), .ZN(
        P1_U3082) );
  AOI22_X1 U23305 ( .A1(n20399), .A2(n20685), .B1(n20684), .B2(n20398), .ZN(
        n20389) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20400), .B1(
        n20426), .B2(n20601), .ZN(n20388) );
  OAI211_X1 U23307 ( .C1(n20403), .C2(n20567), .A(n20389), .B(n20388), .ZN(
        P1_U3083) );
  AOI22_X1 U23308 ( .A1(n20399), .A2(n20691), .B1(n20690), .B2(n20398), .ZN(
        n20391) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20400), .B1(
        n20426), .B2(n20605), .ZN(n20390) );
  OAI211_X1 U23310 ( .C1(n20403), .C2(n20570), .A(n20391), .B(n20390), .ZN(
        P1_U3084) );
  AOI22_X1 U23311 ( .A1(n20399), .A2(n20643), .B1(n20696), .B2(n20398), .ZN(
        n20393) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20400), .B1(
        n20426), .B2(n20697), .ZN(n20392) );
  OAI211_X1 U23313 ( .C1(n20403), .C2(n20573), .A(n20393), .B(n20392), .ZN(
        P1_U3085) );
  AOI22_X1 U23314 ( .A1(n20399), .A2(n20647), .B1(n20701), .B2(n20398), .ZN(
        n20395) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20400), .B1(
        n20426), .B2(n20703), .ZN(n20394) );
  OAI211_X1 U23316 ( .C1(n20403), .C2(n20576), .A(n20395), .B(n20394), .ZN(
        P1_U3086) );
  AOI22_X1 U23317 ( .A1(n20399), .A2(n20651), .B1(n20707), .B2(n20398), .ZN(
        n20397) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20400), .B1(
        n20426), .B2(n9780), .ZN(n20396) );
  OAI211_X1 U23319 ( .C1(n20403), .C2(n20579), .A(n20397), .B(n20396), .ZN(
        P1_U3087) );
  AOI22_X1 U23320 ( .A1(n20399), .A2(n20719), .B1(n20716), .B2(n20398), .ZN(
        n20402) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20400), .B1(
        n20426), .B2(n20617), .ZN(n20401) );
  OAI211_X1 U23322 ( .C1(n20403), .C2(n20586), .A(n20402), .B(n20401), .ZN(
        P1_U3088) );
  INV_X1 U23323 ( .A(n20404), .ZN(n20424) );
  AOI21_X1 U23324 ( .B1(n20405), .B2(n20661), .A(n20424), .ZN(n20406) );
  OAI22_X1 U23325 ( .A1(n20406), .A2(n20664), .B1(n20409), .B2(n20728), .ZN(
        n20425) );
  AOI22_X1 U23326 ( .A1(n20666), .A2(n20424), .B1(n20665), .B2(n20425), .ZN(
        n20411) );
  INV_X1 U23327 ( .A(n9656), .ZN(n20407) );
  NOR3_X1 U23328 ( .A1(n20408), .A2(n20407), .A3(n20820), .ZN(n20811) );
  OAI21_X1 U23329 ( .B1(n20811), .B2(n10499), .A(n20670), .ZN(n20427) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20673), .ZN(n20410) );
  OAI211_X1 U23331 ( .C1(n20676), .C2(n20434), .A(n20411), .B(n20410), .ZN(
        P1_U3089) );
  AOI22_X1 U23332 ( .A1(n20678), .A2(n20424), .B1(n20677), .B2(n20425), .ZN(
        n20413) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20635), .ZN(n20412) );
  OAI211_X1 U23334 ( .C1(n20638), .C2(n20434), .A(n20413), .B(n20412), .ZN(
        P1_U3090) );
  AOI22_X1 U23335 ( .A1(n20684), .A2(n20424), .B1(n20683), .B2(n20425), .ZN(
        n20415) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20685), .ZN(n20414) );
  OAI211_X1 U23337 ( .C1(n20688), .C2(n20434), .A(n20415), .B(n20414), .ZN(
        P1_U3091) );
  AOI22_X1 U23338 ( .A1(n20690), .A2(n20424), .B1(n20689), .B2(n20425), .ZN(
        n20417) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20691), .ZN(n20416) );
  OAI211_X1 U23340 ( .C1(n20694), .C2(n20434), .A(n20417), .B(n20416), .ZN(
        P1_U3092) );
  AOI22_X1 U23341 ( .A1(n20696), .A2(n20424), .B1(n20695), .B2(n20425), .ZN(
        n20419) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20643), .ZN(n20418) );
  OAI211_X1 U23343 ( .C1(n20646), .C2(n20434), .A(n20419), .B(n20418), .ZN(
        P1_U3093) );
  AOI22_X1 U23344 ( .A1(n20702), .A2(n20425), .B1(n20701), .B2(n20424), .ZN(
        n20421) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20647), .ZN(n20420) );
  OAI211_X1 U23346 ( .C1(n20650), .C2(n20434), .A(n20421), .B(n20420), .ZN(
        P1_U3094) );
  AOI22_X1 U23347 ( .A1(n20708), .A2(n20425), .B1(n20707), .B2(n20424), .ZN(
        n20423) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20651), .ZN(n20422) );
  OAI211_X1 U23349 ( .C1(n9779), .C2(n20434), .A(n20423), .B(n20422), .ZN(
        P1_U3095) );
  AOI22_X1 U23350 ( .A1(n20718), .A2(n20425), .B1(n20716), .B2(n20424), .ZN(
        n20429) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20719), .ZN(n20428) );
  OAI211_X1 U23352 ( .C1(n20725), .C2(n20434), .A(n20429), .B(n20428), .ZN(
        P1_U3096) );
  NOR3_X1 U23353 ( .A1(n20519), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20462) );
  INV_X1 U23354 ( .A(n20462), .ZN(n20459) );
  NOR2_X1 U23355 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20459), .ZN(
        n20453) );
  AND2_X1 U23356 ( .A1(n20813), .A2(n13095), .ZN(n20521) );
  AOI21_X1 U23357 ( .B1(n20521), .B2(n9637), .A(n20453), .ZN(n20436) );
  INV_X1 U23358 ( .A(n20431), .ZN(n20432) );
  NAND2_X1 U23359 ( .A1(n20432), .A2(n20486), .ZN(n20554) );
  OAI22_X1 U23360 ( .A1(n20436), .A2(n20664), .B1(n20554), .B2(n20433), .ZN(
        n20454) );
  AOI22_X1 U23361 ( .A1(n20666), .A2(n20453), .B1(n20665), .B2(n20454), .ZN(
        n20440) );
  INV_X1 U23362 ( .A(n20482), .ZN(n20435) );
  OAI21_X1 U23363 ( .B1(n20435), .B2(n20455), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20437) );
  NAND2_X1 U23364 ( .A1(n20437), .A2(n20436), .ZN(n20438) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20673), .ZN(n20439) );
  OAI211_X1 U23366 ( .C1(n20676), .C2(n20482), .A(n20440), .B(n20439), .ZN(
        P1_U3097) );
  AOI22_X1 U23367 ( .A1(n20678), .A2(n20453), .B1(n20677), .B2(n20454), .ZN(
        n20442) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20635), .ZN(n20441) );
  OAI211_X1 U23369 ( .C1(n20638), .C2(n20482), .A(n20442), .B(n20441), .ZN(
        P1_U3098) );
  AOI22_X1 U23370 ( .A1(n20684), .A2(n20453), .B1(n20683), .B2(n20454), .ZN(
        n20444) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20685), .ZN(n20443) );
  OAI211_X1 U23372 ( .C1(n20688), .C2(n20482), .A(n20444), .B(n20443), .ZN(
        P1_U3099) );
  AOI22_X1 U23373 ( .A1(n20690), .A2(n20453), .B1(n20689), .B2(n20454), .ZN(
        n20446) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20691), .ZN(n20445) );
  OAI211_X1 U23375 ( .C1(n20694), .C2(n20482), .A(n20446), .B(n20445), .ZN(
        P1_U3100) );
  AOI22_X1 U23376 ( .A1(n20696), .A2(n20453), .B1(n20695), .B2(n20454), .ZN(
        n20448) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20643), .ZN(n20447) );
  OAI211_X1 U23378 ( .C1(n20646), .C2(n20482), .A(n20448), .B(n20447), .ZN(
        P1_U3101) );
  AOI22_X1 U23379 ( .A1(n20702), .A2(n20454), .B1(n20701), .B2(n20453), .ZN(
        n20450) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20647), .ZN(n20449) );
  OAI211_X1 U23381 ( .C1(n20650), .C2(n20482), .A(n20450), .B(n20449), .ZN(
        P1_U3102) );
  AOI22_X1 U23382 ( .A1(n20708), .A2(n20454), .B1(n20707), .B2(n20453), .ZN(
        n20452) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20651), .ZN(n20451) );
  OAI211_X1 U23384 ( .C1(n9779), .C2(n20482), .A(n20452), .B(n20451), .ZN(
        P1_U3103) );
  AOI22_X1 U23385 ( .A1(n20718), .A2(n20454), .B1(n20716), .B2(n20453), .ZN(
        n20458) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20719), .ZN(n20457) );
  OAI211_X1 U23387 ( .C1(n20725), .C2(n20482), .A(n20458), .B(n20457), .ZN(
        P1_U3104) );
  NOR2_X1 U23388 ( .A1(n20588), .A2(n20459), .ZN(n20477) );
  AOI21_X1 U23389 ( .B1(n20521), .B2(n20590), .A(n20477), .ZN(n20460) );
  OAI22_X1 U23390 ( .A1(n20460), .A2(n20664), .B1(n20459), .B2(n20728), .ZN(
        n20478) );
  AOI22_X1 U23391 ( .A1(n20666), .A2(n20477), .B1(n20665), .B2(n20478), .ZN(
        n20464) );
  OAI21_X1 U23392 ( .B1(n20819), .B2(n20974), .A(n20460), .ZN(n20461) );
  OAI221_X1 U23393 ( .B1(n20671), .B2(n20462), .C1(n20664), .C2(n20461), .A(
        n20670), .ZN(n20479) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20479), .B1(
        n20511), .B2(n20595), .ZN(n20463) );
  OAI211_X1 U23395 ( .C1(n20598), .C2(n20482), .A(n20464), .B(n20463), .ZN(
        P1_U3105) );
  AOI22_X1 U23396 ( .A1(n20678), .A2(n20477), .B1(n20677), .B2(n20478), .ZN(
        n20466) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20479), .B1(
        n20511), .B2(n20679), .ZN(n20465) );
  OAI211_X1 U23398 ( .C1(n20682), .C2(n20482), .A(n20466), .B(n20465), .ZN(
        P1_U3106) );
  AOI22_X1 U23399 ( .A1(n20684), .A2(n20477), .B1(n20683), .B2(n20478), .ZN(
        n20468) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20479), .B1(
        n20511), .B2(n20601), .ZN(n20467) );
  OAI211_X1 U23401 ( .C1(n20604), .C2(n20482), .A(n20468), .B(n20467), .ZN(
        P1_U3107) );
  AOI22_X1 U23402 ( .A1(n20690), .A2(n20477), .B1(n20689), .B2(n20478), .ZN(
        n20470) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20479), .B1(
        n20511), .B2(n20605), .ZN(n20469) );
  OAI211_X1 U23404 ( .C1(n20608), .C2(n20482), .A(n20470), .B(n20469), .ZN(
        P1_U3108) );
  AOI22_X1 U23405 ( .A1(n20696), .A2(n20477), .B1(n20695), .B2(n20478), .ZN(
        n20472) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20479), .B1(
        n20511), .B2(n20697), .ZN(n20471) );
  OAI211_X1 U23407 ( .C1(n20700), .C2(n20482), .A(n20472), .B(n20471), .ZN(
        P1_U3109) );
  AOI22_X1 U23408 ( .A1(n20702), .A2(n20478), .B1(n20701), .B2(n20477), .ZN(
        n20474) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20479), .B1(
        n20511), .B2(n20703), .ZN(n20473) );
  OAI211_X1 U23410 ( .C1(n20706), .C2(n20482), .A(n20474), .B(n20473), .ZN(
        P1_U3110) );
  AOI22_X1 U23411 ( .A1(n20708), .A2(n20478), .B1(n20707), .B2(n20477), .ZN(
        n20476) );
  AOI22_X1 U23412 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20479), .B1(
        n20511), .B2(n9780), .ZN(n20475) );
  OAI211_X1 U23413 ( .C1(n20714), .C2(n20482), .A(n20476), .B(n20475), .ZN(
        P1_U3111) );
  AOI22_X1 U23414 ( .A1(n20718), .A2(n20478), .B1(n20716), .B2(n20477), .ZN(
        n20481) );
  AOI22_X1 U23415 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20479), .B1(
        n20511), .B2(n20617), .ZN(n20480) );
  OAI211_X1 U23416 ( .C1(n20622), .C2(n20482), .A(n20481), .B(n20480), .ZN(
        P1_U3112) );
  INV_X1 U23417 ( .A(n20511), .ZN(n20483) );
  NAND2_X1 U23418 ( .A1(n20483), .A2(n20671), .ZN(n20485) );
  OAI21_X1 U23419 ( .B1(n20485), .B2(n20544), .A(n20484), .ZN(n20494) );
  AND2_X1 U23420 ( .A1(n20521), .A2(n20625), .ZN(n20490) );
  OR2_X1 U23421 ( .A1(n20486), .A2(n20519), .ZN(n20627) );
  INV_X1 U23422 ( .A(n20627), .ZN(n20487) );
  NOR3_X1 U23423 ( .A1(n20519), .A2(n20489), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20527) );
  INV_X1 U23424 ( .A(n20527), .ZN(n20522) );
  NOR2_X1 U23425 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20522), .ZN(
        n20510) );
  AOI22_X1 U23426 ( .A1(n20511), .A2(n20673), .B1(n20666), .B2(n20510), .ZN(
        n20497) );
  INV_X1 U23427 ( .A(n20490), .ZN(n20493) );
  NAND2_X1 U23428 ( .A1(n20627), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20630) );
  OAI211_X1 U23429 ( .C1(n13115), .C2(n20510), .A(n20630), .B(n20491), .ZN(
        n20492) );
  AOI21_X1 U23430 ( .B1(n20494), .B2(n20493), .A(n20492), .ZN(n20495) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20512), .B1(
        n20544), .B2(n20595), .ZN(n20496) );
  OAI211_X1 U23432 ( .C1(n20515), .C2(n20561), .A(n20497), .B(n20496), .ZN(
        P1_U3113) );
  AOI22_X1 U23433 ( .A1(n20544), .A2(n20679), .B1(n20678), .B2(n20510), .ZN(
        n20499) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20635), .ZN(n20498) );
  OAI211_X1 U23435 ( .C1(n20515), .C2(n20564), .A(n20499), .B(n20498), .ZN(
        P1_U3114) );
  AOI22_X1 U23436 ( .A1(n20511), .A2(n20685), .B1(n20684), .B2(n20510), .ZN(
        n20501) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20512), .B1(
        n20544), .B2(n20601), .ZN(n20500) );
  OAI211_X1 U23438 ( .C1(n20515), .C2(n20567), .A(n20501), .B(n20500), .ZN(
        P1_U3115) );
  AOI22_X1 U23439 ( .A1(n20544), .A2(n20605), .B1(n20690), .B2(n20510), .ZN(
        n20503) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20691), .ZN(n20502) );
  OAI211_X1 U23441 ( .C1(n20515), .C2(n20570), .A(n20503), .B(n20502), .ZN(
        P1_U3116) );
  AOI22_X1 U23442 ( .A1(n20544), .A2(n20697), .B1(n20696), .B2(n20510), .ZN(
        n20505) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20643), .ZN(n20504) );
  OAI211_X1 U23444 ( .C1(n20515), .C2(n20573), .A(n20505), .B(n20504), .ZN(
        P1_U3117) );
  AOI22_X1 U23445 ( .A1(n20544), .A2(n20703), .B1(n20701), .B2(n20510), .ZN(
        n20507) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20647), .ZN(n20506) );
  OAI211_X1 U23447 ( .C1(n20515), .C2(n20576), .A(n20507), .B(n20506), .ZN(
        P1_U3118) );
  AOI22_X1 U23448 ( .A1(n20544), .A2(n9780), .B1(n20707), .B2(n20510), .ZN(
        n20509) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20512), .B1(
        n20511), .B2(n20651), .ZN(n20508) );
  OAI211_X1 U23450 ( .C1(n20515), .C2(n20579), .A(n20509), .B(n20508), .ZN(
        P1_U3119) );
  AOI22_X1 U23451 ( .A1(n20511), .A2(n20719), .B1(n20716), .B2(n20510), .ZN(
        n20514) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20512), .B1(
        n20544), .B2(n20617), .ZN(n20513) );
  OAI211_X1 U23453 ( .C1(n20515), .C2(n20586), .A(n20514), .B(n20513), .ZN(
        P1_U3120) );
  INV_X1 U23454 ( .A(n20516), .ZN(n20517) );
  NOR2_X1 U23455 ( .A1(n20520), .A2(n20519), .ZN(n20542) );
  AOI21_X1 U23456 ( .B1(n20521), .B2(n20661), .A(n20542), .ZN(n20524) );
  OAI22_X1 U23457 ( .A1(n20524), .A2(n20664), .B1(n20522), .B2(n20728), .ZN(
        n20543) );
  AOI22_X1 U23458 ( .A1(n20666), .A2(n20542), .B1(n20665), .B2(n20543), .ZN(
        n20529) );
  INV_X1 U23459 ( .A(n20523), .ZN(n20525) );
  OAI21_X1 U23460 ( .B1(n20819), .B2(n20525), .A(n20524), .ZN(n20526) );
  OAI221_X1 U23461 ( .B1(n20671), .B2(n20527), .C1(n20664), .C2(n20526), .A(
        n20670), .ZN(n20545) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20673), .ZN(n20528) );
  OAI211_X1 U23463 ( .C1(n20676), .C2(n20558), .A(n20529), .B(n20528), .ZN(
        P1_U3121) );
  AOI22_X1 U23464 ( .A1(n20678), .A2(n20542), .B1(n20677), .B2(n20543), .ZN(
        n20531) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20635), .ZN(n20530) );
  OAI211_X1 U23466 ( .C1(n20638), .C2(n20558), .A(n20531), .B(n20530), .ZN(
        P1_U3122) );
  AOI22_X1 U23467 ( .A1(n20684), .A2(n20542), .B1(n20683), .B2(n20543), .ZN(
        n20533) );
  AOI22_X1 U23468 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20685), .ZN(n20532) );
  OAI211_X1 U23469 ( .C1(n20688), .C2(n20558), .A(n20533), .B(n20532), .ZN(
        P1_U3123) );
  AOI22_X1 U23470 ( .A1(n20690), .A2(n20542), .B1(n20689), .B2(n20543), .ZN(
        n20535) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20691), .ZN(n20534) );
  OAI211_X1 U23472 ( .C1(n20694), .C2(n20558), .A(n20535), .B(n20534), .ZN(
        P1_U3124) );
  AOI22_X1 U23473 ( .A1(n20696), .A2(n20542), .B1(n20695), .B2(n20543), .ZN(
        n20537) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20643), .ZN(n20536) );
  OAI211_X1 U23475 ( .C1(n20646), .C2(n20558), .A(n20537), .B(n20536), .ZN(
        P1_U3125) );
  AOI22_X1 U23476 ( .A1(n20702), .A2(n20543), .B1(n20701), .B2(n20542), .ZN(
        n20539) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20647), .ZN(n20538) );
  OAI211_X1 U23478 ( .C1(n20650), .C2(n20558), .A(n20539), .B(n20538), .ZN(
        P1_U3126) );
  AOI22_X1 U23479 ( .A1(n20708), .A2(n20543), .B1(n20707), .B2(n20542), .ZN(
        n20541) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20651), .ZN(n20540) );
  OAI211_X1 U23481 ( .C1(n9779), .C2(n20558), .A(n20541), .B(n20540), .ZN(
        P1_U3127) );
  AOI22_X1 U23482 ( .A1(n20718), .A2(n20543), .B1(n20716), .B2(n20542), .ZN(
        n20547) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20719), .ZN(n20546) );
  OAI211_X1 U23484 ( .C1(n20725), .C2(n20558), .A(n20547), .B(n20546), .ZN(
        P1_U3128) );
  NAND2_X1 U23485 ( .A1(n20558), .A2(n20621), .ZN(n20549) );
  AOI21_X1 U23486 ( .B1(n20549), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20664), 
        .ZN(n20556) );
  OR2_X1 U23487 ( .A1(n13095), .A2(n20550), .ZN(n20589) );
  OR2_X1 U23488 ( .A1(n20589), .A2(n20625), .ZN(n20555) );
  INV_X1 U23489 ( .A(n20555), .ZN(n20553) );
  INV_X1 U23490 ( .A(n20554), .ZN(n20551) );
  NOR3_X1 U23491 ( .A1(n11119), .A2(n20519), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20593) );
  INV_X1 U23492 ( .A(n20593), .ZN(n20591) );
  NOR2_X1 U23493 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20591), .ZN(
        n20580) );
  AOI22_X1 U23494 ( .A1(n20581), .A2(n20595), .B1(n20666), .B2(n20580), .ZN(
        n20560) );
  AOI22_X1 U23495 ( .A1(n20556), .A2(n20555), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20554), .ZN(n20557) );
  OAI211_X1 U23496 ( .C1(n20580), .C2(n13115), .A(n20631), .B(n20557), .ZN(
        n20583) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20673), .ZN(n20559) );
  OAI211_X1 U23498 ( .C1(n20587), .C2(n20561), .A(n20560), .B(n20559), .ZN(
        P1_U3129) );
  AOI22_X1 U23499 ( .A1(n20581), .A2(n20679), .B1(n20678), .B2(n20580), .ZN(
        n20563) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20635), .ZN(n20562) );
  OAI211_X1 U23501 ( .C1(n20587), .C2(n20564), .A(n20563), .B(n20562), .ZN(
        P1_U3130) );
  AOI22_X1 U23502 ( .A1(n20581), .A2(n20601), .B1(n20684), .B2(n20580), .ZN(
        n20566) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20685), .ZN(n20565) );
  OAI211_X1 U23504 ( .C1(n20587), .C2(n20567), .A(n20566), .B(n20565), .ZN(
        P1_U3131) );
  AOI22_X1 U23505 ( .A1(n20581), .A2(n20605), .B1(n20690), .B2(n20580), .ZN(
        n20569) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20691), .ZN(n20568) );
  OAI211_X1 U23507 ( .C1(n20587), .C2(n20570), .A(n20569), .B(n20568), .ZN(
        P1_U3132) );
  AOI22_X1 U23508 ( .A1(n20581), .A2(n20697), .B1(n20696), .B2(n20580), .ZN(
        n20572) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20643), .ZN(n20571) );
  OAI211_X1 U23510 ( .C1(n20587), .C2(n20573), .A(n20572), .B(n20571), .ZN(
        P1_U3133) );
  AOI22_X1 U23511 ( .A1(n20581), .A2(n20703), .B1(n20701), .B2(n20580), .ZN(
        n20575) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20647), .ZN(n20574) );
  OAI211_X1 U23513 ( .C1(n20587), .C2(n20576), .A(n20575), .B(n20574), .ZN(
        P1_U3134) );
  AOI22_X1 U23514 ( .A1(n20581), .A2(n9780), .B1(n20707), .B2(n20580), .ZN(
        n20578) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20651), .ZN(n20577) );
  OAI211_X1 U23516 ( .C1(n20587), .C2(n20579), .A(n20578), .B(n20577), .ZN(
        P1_U3135) );
  AOI22_X1 U23517 ( .A1(n20581), .A2(n20617), .B1(n20716), .B2(n20580), .ZN(
        n20585) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20719), .ZN(n20584) );
  OAI211_X1 U23519 ( .C1(n20587), .C2(n20586), .A(n20585), .B(n20584), .ZN(
        P1_U3136) );
  NOR2_X1 U23520 ( .A1(n20588), .A2(n20591), .ZN(n20615) );
  AOI21_X1 U23521 ( .B1(n20662), .B2(n20590), .A(n20615), .ZN(n20592) );
  OAI22_X1 U23522 ( .A1(n20592), .A2(n20664), .B1(n20591), .B2(n20728), .ZN(
        n20616) );
  AOI22_X1 U23523 ( .A1(n20666), .A2(n20615), .B1(n20665), .B2(n20616), .ZN(
        n20597) );
  NOR3_X1 U23524 ( .A1(n20624), .A2(n9656), .A3(n20820), .ZN(n20810) );
  OAI21_X1 U23525 ( .B1(n20810), .B2(n20593), .A(n20670), .ZN(n20618) );
  NOR2_X2 U23526 ( .A1(n20624), .A2(n20594), .ZN(n20656) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20618), .B1(
        n20656), .B2(n20595), .ZN(n20596) );
  OAI211_X1 U23528 ( .C1(n20598), .C2(n20621), .A(n20597), .B(n20596), .ZN(
        P1_U3137) );
  AOI22_X1 U23529 ( .A1(n20678), .A2(n20615), .B1(n20677), .B2(n20616), .ZN(
        n20600) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20618), .B1(
        n20656), .B2(n20679), .ZN(n20599) );
  OAI211_X1 U23531 ( .C1(n20682), .C2(n20621), .A(n20600), .B(n20599), .ZN(
        P1_U3138) );
  AOI22_X1 U23532 ( .A1(n20684), .A2(n20615), .B1(n20683), .B2(n20616), .ZN(
        n20603) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20618), .B1(
        n20656), .B2(n20601), .ZN(n20602) );
  OAI211_X1 U23534 ( .C1(n20604), .C2(n20621), .A(n20603), .B(n20602), .ZN(
        P1_U3139) );
  AOI22_X1 U23535 ( .A1(n20690), .A2(n20615), .B1(n20689), .B2(n20616), .ZN(
        n20607) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20618), .B1(
        n20656), .B2(n20605), .ZN(n20606) );
  OAI211_X1 U23537 ( .C1(n20608), .C2(n20621), .A(n20607), .B(n20606), .ZN(
        P1_U3140) );
  AOI22_X1 U23538 ( .A1(n20696), .A2(n20615), .B1(n20695), .B2(n20616), .ZN(
        n20610) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20618), .B1(
        n20656), .B2(n20697), .ZN(n20609) );
  OAI211_X1 U23540 ( .C1(n20700), .C2(n20621), .A(n20610), .B(n20609), .ZN(
        P1_U3141) );
  AOI22_X1 U23541 ( .A1(n20702), .A2(n20616), .B1(n20701), .B2(n20615), .ZN(
        n20612) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20618), .B1(
        n20656), .B2(n20703), .ZN(n20611) );
  OAI211_X1 U23543 ( .C1(n20706), .C2(n20621), .A(n20612), .B(n20611), .ZN(
        P1_U3142) );
  AOI22_X1 U23544 ( .A1(n20708), .A2(n20616), .B1(n20707), .B2(n20615), .ZN(
        n20614) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20618), .B1(
        n20656), .B2(n9780), .ZN(n20613) );
  OAI211_X1 U23546 ( .C1(n20714), .C2(n20621), .A(n20614), .B(n20613), .ZN(
        P1_U3143) );
  AOI22_X1 U23547 ( .A1(n20718), .A2(n20616), .B1(n20716), .B2(n20615), .ZN(
        n20620) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20618), .B1(
        n20656), .B2(n20617), .ZN(n20619) );
  OAI211_X1 U23549 ( .C1(n20622), .C2(n20621), .A(n20620), .B(n20619), .ZN(
        P1_U3144) );
  INV_X1 U23550 ( .A(n20672), .ZN(n20663) );
  NOR2_X1 U23551 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20663), .ZN(
        n20654) );
  NAND2_X1 U23552 ( .A1(n20662), .A2(n20625), .ZN(n20628) );
  OAI22_X1 U23553 ( .A1(n20628), .A2(n20664), .B1(n20627), .B2(n20626), .ZN(
        n20655) );
  AOI22_X1 U23554 ( .A1(n20666), .A2(n20654), .B1(n20665), .B2(n20655), .ZN(
        n20634) );
  OAI21_X1 U23555 ( .B1(n20720), .B2(n20656), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20629) );
  AOI21_X1 U23556 ( .B1(n20629), .B2(n20628), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20632) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20673), .ZN(n20633) );
  OAI211_X1 U23558 ( .C1(n20676), .C2(n20713), .A(n20634), .B(n20633), .ZN(
        P1_U3145) );
  AOI22_X1 U23559 ( .A1(n20678), .A2(n20654), .B1(n20677), .B2(n20655), .ZN(
        n20637) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20635), .ZN(n20636) );
  OAI211_X1 U23561 ( .C1(n20638), .C2(n20713), .A(n20637), .B(n20636), .ZN(
        P1_U3146) );
  AOI22_X1 U23562 ( .A1(n20684), .A2(n20654), .B1(n20683), .B2(n20655), .ZN(
        n20640) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20685), .ZN(n20639) );
  OAI211_X1 U23564 ( .C1(n20688), .C2(n20713), .A(n20640), .B(n20639), .ZN(
        P1_U3147) );
  AOI22_X1 U23565 ( .A1(n20690), .A2(n20654), .B1(n20689), .B2(n20655), .ZN(
        n20642) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20691), .ZN(n20641) );
  OAI211_X1 U23567 ( .C1(n20694), .C2(n20713), .A(n20642), .B(n20641), .ZN(
        P1_U3148) );
  AOI22_X1 U23568 ( .A1(n20696), .A2(n20654), .B1(n20695), .B2(n20655), .ZN(
        n20645) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20643), .ZN(n20644) );
  OAI211_X1 U23570 ( .C1(n20646), .C2(n20713), .A(n20645), .B(n20644), .ZN(
        P1_U3149) );
  AOI22_X1 U23571 ( .A1(n20702), .A2(n20655), .B1(n20701), .B2(n20654), .ZN(
        n20649) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20647), .ZN(n20648) );
  OAI211_X1 U23573 ( .C1(n20650), .C2(n20713), .A(n20649), .B(n20648), .ZN(
        P1_U3150) );
  AOI22_X1 U23574 ( .A1(n20708), .A2(n20655), .B1(n20707), .B2(n20654), .ZN(
        n20653) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20651), .ZN(n20652) );
  OAI211_X1 U23576 ( .C1(n9779), .C2(n20713), .A(n20653), .B(n20652), .ZN(
        P1_U3151) );
  AOI22_X1 U23577 ( .A1(n20718), .A2(n20655), .B1(n20716), .B2(n20654), .ZN(
        n20659) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20719), .ZN(n20658) );
  OAI211_X1 U23579 ( .C1(n20725), .C2(n20713), .A(n20659), .B(n20658), .ZN(
        P1_U3152) );
  INV_X1 U23580 ( .A(n20660), .ZN(n20715) );
  AOI21_X1 U23581 ( .B1(n20662), .B2(n20661), .A(n20715), .ZN(n20667) );
  OAI22_X1 U23582 ( .A1(n20667), .A2(n20664), .B1(n20728), .B2(n20663), .ZN(
        n20717) );
  AOI22_X1 U23583 ( .A1(n20666), .A2(n20715), .B1(n20665), .B2(n20717), .ZN(
        n20675) );
  OAI21_X1 U23584 ( .B1(n20811), .B2(n20668), .A(n20667), .ZN(n20669) );
  OAI211_X1 U23585 ( .C1(n20672), .C2(n20671), .A(n20670), .B(n20669), .ZN(
        n20721) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20721), .B1(
        n20720), .B2(n20673), .ZN(n20674) );
  OAI211_X1 U23587 ( .C1(n20676), .C2(n20724), .A(n20675), .B(n20674), .ZN(
        P1_U3153) );
  AOI22_X1 U23588 ( .A1(n20678), .A2(n20715), .B1(n20677), .B2(n20717), .ZN(
        n20681) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20721), .B1(
        n20710), .B2(n20679), .ZN(n20680) );
  OAI211_X1 U23590 ( .C1(n20682), .C2(n20713), .A(n20681), .B(n20680), .ZN(
        P1_U3154) );
  AOI22_X1 U23591 ( .A1(n20684), .A2(n20715), .B1(n20683), .B2(n20717), .ZN(
        n20687) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20721), .B1(
        n20720), .B2(n20685), .ZN(n20686) );
  OAI211_X1 U23593 ( .C1(n20688), .C2(n20724), .A(n20687), .B(n20686), .ZN(
        P1_U3155) );
  AOI22_X1 U23594 ( .A1(n20690), .A2(n20715), .B1(n20689), .B2(n20717), .ZN(
        n20693) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20721), .B1(
        n20720), .B2(n20691), .ZN(n20692) );
  OAI211_X1 U23596 ( .C1(n20694), .C2(n20724), .A(n20693), .B(n20692), .ZN(
        P1_U3156) );
  AOI22_X1 U23597 ( .A1(n20696), .A2(n20715), .B1(n20695), .B2(n20717), .ZN(
        n20699) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20721), .B1(
        n20710), .B2(n20697), .ZN(n20698) );
  OAI211_X1 U23599 ( .C1(n20700), .C2(n20713), .A(n20699), .B(n20698), .ZN(
        P1_U3157) );
  AOI22_X1 U23600 ( .A1(n20702), .A2(n20717), .B1(n20701), .B2(n20715), .ZN(
        n20705) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20721), .B1(
        n20710), .B2(n20703), .ZN(n20704) );
  OAI211_X1 U23602 ( .C1(n20706), .C2(n20713), .A(n20705), .B(n20704), .ZN(
        P1_U3158) );
  AOI22_X1 U23603 ( .A1(n20708), .A2(n20717), .B1(n20707), .B2(n20715), .ZN(
        n20712) );
  AOI22_X1 U23604 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20721), .B1(
        n20710), .B2(n9780), .ZN(n20711) );
  OAI211_X1 U23605 ( .C1(n20714), .C2(n20713), .A(n20712), .B(n20711), .ZN(
        P1_U3159) );
  AOI22_X1 U23606 ( .A1(n20718), .A2(n20717), .B1(n20716), .B2(n20715), .ZN(
        n20723) );
  AOI22_X1 U23607 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20721), .B1(
        n20720), .B2(n20719), .ZN(n20722) );
  OAI211_X1 U23608 ( .C1(n20725), .C2(n20724), .A(n20723), .B(n20722), .ZN(
        P1_U3160) );
  AOI22_X1 U23609 ( .A1(n20729), .A2(n20728), .B1(n20727), .B2(n20726), .ZN(
        P1_U3163) );
  AND2_X1 U23610 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20730), .ZN(
        P1_U3164) );
  AND2_X1 U23611 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20730), .ZN(
        P1_U3165) );
  AND2_X1 U23612 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20730), .ZN(
        P1_U3166) );
  AND2_X1 U23613 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20730), .ZN(
        P1_U3167) );
  AND2_X1 U23614 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20730), .ZN(
        P1_U3168) );
  AND2_X1 U23615 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20730), .ZN(
        P1_U3169) );
  AND2_X1 U23616 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20730), .ZN(
        P1_U3170) );
  AND2_X1 U23617 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20730), .ZN(
        P1_U3171) );
  AND2_X1 U23618 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20730), .ZN(
        P1_U3172) );
  AND2_X1 U23619 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20730), .ZN(
        P1_U3173) );
  AND2_X1 U23620 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20730), .ZN(
        P1_U3174) );
  AND2_X1 U23621 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20730), .ZN(
        P1_U3175) );
  AND2_X1 U23622 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20730), .ZN(
        P1_U3176) );
  AND2_X1 U23623 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20730), .ZN(
        P1_U3177) );
  AND2_X1 U23624 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20730), .ZN(
        P1_U3178) );
  AND2_X1 U23625 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20730), .ZN(
        P1_U3179) );
  AND2_X1 U23626 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20730), .ZN(
        P1_U3180) );
  AND2_X1 U23627 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20730), .ZN(
        P1_U3181) );
  AND2_X1 U23628 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20730), .ZN(
        P1_U3182) );
  AND2_X1 U23629 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20730), .ZN(
        P1_U3183) );
  AND2_X1 U23630 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20730), .ZN(
        P1_U3184) );
  AND2_X1 U23631 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20730), .ZN(
        P1_U3185) );
  AND2_X1 U23632 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20730), .ZN(P1_U3186) );
  AND2_X1 U23633 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20730), .ZN(P1_U3187) );
  AND2_X1 U23634 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20730), .ZN(P1_U3188) );
  AND2_X1 U23635 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20730), .ZN(P1_U3189) );
  AND2_X1 U23636 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20730), .ZN(P1_U3190) );
  AND2_X1 U23637 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20730), .ZN(P1_U3191) );
  AND2_X1 U23638 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20730), .ZN(P1_U3192) );
  AND2_X1 U23639 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20730), .ZN(P1_U3193) );
  NAND2_X1 U23640 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20731), .ZN(n20735) );
  NOR2_X1 U23641 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20732) );
  OAI22_X1 U23642 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20958), .B1(n20732), 
        .B2(n20976), .ZN(n20733) );
  OAI21_X1 U23643 ( .B1(n20953), .B2(n20733), .A(n20832), .ZN(n20734) );
  OAI221_X1 U23644 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(P1_STATE_REG_0__SCAN_IN), .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20735), .A(n20734), .ZN(P1_U3194) );
  INV_X1 U23645 ( .A(n20735), .ZN(n20736) );
  AOI221_X1 U23646 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20739), .C1(n20958), 
        .C2(n20739), .A(n20736), .ZN(n20744) );
  NOR2_X1 U23647 ( .A1(NA), .A2(n20739), .ZN(n20737) );
  AOI21_X1 U23648 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20737), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n20743) );
  NOR3_X1 U23649 ( .A1(NA), .A2(n20739), .A3(n20738), .ZN(n20740) );
  OAI22_X1 U23650 ( .A1(n20741), .A2(n20740), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20953), .ZN(n20742) );
  OAI22_X1 U23651 ( .A1(n20744), .A2(n20743), .B1(n20976), .B2(n20742), .ZN(
        P1_U3196) );
  NOR2_X1 U23652 ( .A1(n20832), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20782) );
  INV_X1 U23653 ( .A(n20782), .ZN(n20769) );
  INV_X1 U23654 ( .A(n20769), .ZN(n20784) );
  INV_X1 U23655 ( .A(n20831), .ZN(n20785) );
  OR2_X1 U23656 ( .A1(n20745), .A2(n20832), .ZN(n20766) );
  AOI222_X1 U23657 ( .A1(n20784), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n9653), .ZN(n20746) );
  INV_X1 U23658 ( .A(n20746), .ZN(P1_U3197) );
  AOI222_X1 U23659 ( .A1(n9653), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20784), .ZN(n20747) );
  INV_X1 U23660 ( .A(n20747), .ZN(P1_U3198) );
  OAI222_X1 U23661 ( .A1(n20766), .A2(n20750), .B1(n20749), .B2(n20831), .C1(
        n20748), .C2(n20769), .ZN(P1_U3199) );
  AOI222_X1 U23662 ( .A1(n20784), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n9653), .ZN(n20751) );
  INV_X1 U23663 ( .A(n20751), .ZN(P1_U3200) );
  AOI222_X1 U23664 ( .A1(n9653), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20784), .ZN(n20752) );
  INV_X1 U23665 ( .A(n20752), .ZN(P1_U3201) );
  AOI22_X1 U23666 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20832), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20782), .ZN(n20753) );
  OAI21_X1 U23667 ( .B1(n20754), .B2(n20766), .A(n20753), .ZN(P1_U3202) );
  AOI22_X1 U23668 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20832), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n9653), .ZN(n20755) );
  OAI21_X1 U23669 ( .B1(n20756), .B2(n20769), .A(n20755), .ZN(P1_U3203) );
  AOI222_X1 U23670 ( .A1(n9653), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20784), .ZN(n20757) );
  INV_X1 U23671 ( .A(n20757), .ZN(P1_U3204) );
  AOI222_X1 U23672 ( .A1(n9653), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20782), .ZN(n20758) );
  INV_X1 U23673 ( .A(n20758), .ZN(P1_U3205) );
  AOI222_X1 U23674 ( .A1(n9653), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20784), .ZN(n20759) );
  INV_X1 U23675 ( .A(n20759), .ZN(P1_U3206) );
  AOI222_X1 U23676 ( .A1(n9653), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20784), .ZN(n20760) );
  INV_X1 U23677 ( .A(n20760), .ZN(P1_U3207) );
  AOI222_X1 U23678 ( .A1(n20782), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n9653), .ZN(n20761) );
  INV_X1 U23679 ( .A(n20761), .ZN(P1_U3208) );
  AOI222_X1 U23680 ( .A1(n9653), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20784), .ZN(n20762) );
  INV_X1 U23681 ( .A(n20762), .ZN(P1_U3209) );
  AOI222_X1 U23682 ( .A1(n20782), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n9653), .ZN(n20763) );
  INV_X1 U23683 ( .A(n20763), .ZN(P1_U3210) );
  AOI222_X1 U23684 ( .A1(n9653), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20784), .ZN(n20764) );
  INV_X1 U23685 ( .A(n20764), .ZN(P1_U3211) );
  AOI22_X1 U23686 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20832), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20782), .ZN(n20765) );
  OAI21_X1 U23687 ( .B1(n20767), .B2(n20766), .A(n20765), .ZN(P1_U3212) );
  AOI22_X1 U23688 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20832), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n9653), .ZN(n20768) );
  OAI21_X1 U23689 ( .B1(n20770), .B2(n20769), .A(n20768), .ZN(P1_U3213) );
  AOI222_X1 U23690 ( .A1(n20782), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n9653), .ZN(n20771) );
  INV_X1 U23691 ( .A(n20771), .ZN(P1_U3214) );
  AOI222_X1 U23692 ( .A1(n9653), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20784), .ZN(n20772) );
  INV_X1 U23693 ( .A(n20772), .ZN(P1_U3215) );
  AOI222_X1 U23694 ( .A1(n20782), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n9653), .ZN(n20773) );
  INV_X1 U23695 ( .A(n20773), .ZN(P1_U3216) );
  AOI222_X1 U23696 ( .A1(n9653), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20784), .ZN(n20774) );
  INV_X1 U23697 ( .A(n20774), .ZN(P1_U3217) );
  AOI222_X1 U23698 ( .A1(n9653), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20784), .ZN(n20775) );
  INV_X1 U23699 ( .A(n20775), .ZN(P1_U3218) );
  AOI222_X1 U23700 ( .A1(n20782), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n9653), .ZN(n20776) );
  INV_X1 U23701 ( .A(n20776), .ZN(P1_U3219) );
  AOI222_X1 U23702 ( .A1(n20784), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n9653), .ZN(n20777) );
  INV_X1 U23703 ( .A(n20777), .ZN(P1_U3220) );
  AOI222_X1 U23704 ( .A1(n9653), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20784), .ZN(n20778) );
  INV_X1 U23705 ( .A(n20778), .ZN(P1_U3221) );
  AOI222_X1 U23706 ( .A1(n9653), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20784), .ZN(n20779) );
  INV_X1 U23707 ( .A(n20779), .ZN(P1_U3222) );
  AOI222_X1 U23708 ( .A1(n9653), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20784), .ZN(n20780) );
  INV_X1 U23709 ( .A(n20780), .ZN(P1_U3223) );
  AOI222_X1 U23710 ( .A1(n20784), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n9653), .ZN(n20781) );
  INV_X1 U23711 ( .A(n20781), .ZN(P1_U3224) );
  AOI222_X1 U23712 ( .A1(n9653), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20782), .ZN(n20783) );
  INV_X1 U23713 ( .A(n20783), .ZN(P1_U3225) );
  AOI222_X1 U23714 ( .A1(n9653), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20785), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20784), .ZN(n20786) );
  INV_X1 U23715 ( .A(n20786), .ZN(P1_U3226) );
  OAI22_X1 U23716 ( .A1(n20832), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20831), .ZN(n20787) );
  INV_X1 U23717 ( .A(n20787), .ZN(P1_U3458) );
  OAI22_X1 U23718 ( .A1(n20832), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20831), .ZN(n20788) );
  INV_X1 U23719 ( .A(n20788), .ZN(P1_U3459) );
  OAI22_X1 U23720 ( .A1(n20832), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20831), .ZN(n20789) );
  INV_X1 U23721 ( .A(n20789), .ZN(P1_U3460) );
  OAI22_X1 U23722 ( .A1(n20832), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20831), .ZN(n20790) );
  INV_X1 U23723 ( .A(n20790), .ZN(P1_U3461) );
  OAI21_X1 U23724 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20794), .A(n20792), 
        .ZN(n20791) );
  INV_X1 U23725 ( .A(n20791), .ZN(P1_U3464) );
  OAI21_X1 U23726 ( .B1(n20794), .B2(n20793), .A(n20792), .ZN(P1_U3465) );
  INV_X1 U23727 ( .A(n20795), .ZN(n20797) );
  OAI22_X1 U23728 ( .A1(n20797), .A2(n20809), .B1(n20796), .B2(n20801), .ZN(
        n20798) );
  MUX2_X1 U23729 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20798), .S(
        n20804), .Z(P1_U3469) );
  INV_X1 U23730 ( .A(n20799), .ZN(n20800) );
  AOI21_X1 U23731 ( .B1(n20800), .B2(n13115), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n20802) );
  OAI22_X1 U23732 ( .A1(n20803), .A2(n20802), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20801), .ZN(n20805) );
  AOI22_X1 U23733 ( .A1(n20806), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20805), .B2(n20804), .ZN(n20807) );
  OAI21_X1 U23734 ( .B1(n20809), .B2(n20808), .A(n20807), .ZN(P1_U3474) );
  NOR2_X1 U23735 ( .A1(n20811), .A2(n20810), .ZN(n20818) );
  INV_X1 U23736 ( .A(n20812), .ZN(n20816) );
  AOI22_X1 U23737 ( .A1(n20816), .A2(n20815), .B1(n20814), .B2(n20813), .ZN(
        n20817) );
  OAI211_X1 U23738 ( .C1(n20820), .C2(n20819), .A(n20818), .B(n20817), .ZN(
        n20821) );
  NAND2_X1 U23739 ( .A1(n20823), .A2(n20821), .ZN(n20822) );
  OAI21_X1 U23740 ( .B1(n20823), .B2(n20519), .A(n20822), .ZN(P1_U3475) );
  AOI21_X1 U23741 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20825) );
  AOI22_X1 U23742 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20825), .B2(n20824), .ZN(n20826) );
  INV_X1 U23743 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20929) );
  AOI22_X1 U23744 ( .A1(n20827), .A2(n20826), .B1(n20929), .B2(n20829), .ZN(
        P1_U3481) );
  INV_X1 U23745 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20830) );
  NOR2_X1 U23746 ( .A1(n20829), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20828) );
  AOI22_X1 U23747 ( .A1(n20830), .A2(n20829), .B1(n13075), .B2(n20828), .ZN(
        P1_U3482) );
  AOI22_X1 U23748 ( .A1(n20831), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20923), 
        .B2(n20832), .ZN(P1_U3483) );
  OAI22_X1 U23749 ( .A1(n20832), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20831), .ZN(n20833) );
  INV_X1 U23750 ( .A(n20833), .ZN(P1_U3486) );
  AOI22_X1 U23751 ( .A1(DATAI_23_), .A2(keyinput_f9), .B1(DATAI_31_), .B2(
        keyinput_f1), .ZN(n20834) );
  OAI221_X1 U23752 ( .B1(DATAI_23_), .B2(keyinput_f9), .C1(DATAI_31_), .C2(
        keyinput_f1), .A(n20834), .ZN(n20841) );
  AOI22_X1 U23753 ( .A1(keyinput_f49), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .ZN(n20835) );
  OAI221_X1 U23754 ( .B1(keyinput_f49), .B2(P1_BYTEENABLE_REG_1__SCAN_IN), 
        .C1(P1_REIP_REG_31__SCAN_IN), .C2(keyinput_f52), .A(n20835), .ZN(
        n20840) );
  AOI22_X1 U23755 ( .A1(DATAI_19_), .A2(keyinput_f13), .B1(DATAI_4_), .B2(
        keyinput_f28), .ZN(n20836) );
  OAI221_X1 U23756 ( .B1(DATAI_19_), .B2(keyinput_f13), .C1(DATAI_4_), .C2(
        keyinput_f28), .A(n20836), .ZN(n20839) );
  AOI22_X1 U23757 ( .A1(keyinput_f41), .A2(P1_M_IO_N_REG_SCAN_IN), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_f54), .ZN(n20837) );
  OAI221_X1 U23758 ( .B1(keyinput_f41), .B2(P1_M_IO_N_REG_SCAN_IN), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_f54), .A(n20837), .ZN(n20838)
         );
  NOR4_X1 U23759 ( .A1(n20841), .A2(n20840), .A3(n20839), .A4(n20838), .ZN(
        n20868) );
  XOR2_X1 U23760 ( .A(READY1), .B(keyinput_f36), .Z(n20848) );
  AOI22_X1 U23761 ( .A1(keyinput_f34), .A2(NA), .B1(DATAI_22_), .B2(
        keyinput_f10), .ZN(n20842) );
  OAI221_X1 U23762 ( .B1(keyinput_f34), .B2(NA), .C1(DATAI_22_), .C2(
        keyinput_f10), .A(n20842), .ZN(n20847) );
  AOI22_X1 U23763 ( .A1(DATAI_17_), .A2(keyinput_f15), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_f55), .ZN(n20843) );
  OAI221_X1 U23764 ( .B1(DATAI_17_), .B2(keyinput_f15), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput_f55), .A(n20843), .ZN(n20846)
         );
  AOI22_X1 U23765 ( .A1(DATAI_1_), .A2(keyinput_f31), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .ZN(n20844) );
  OAI221_X1 U23766 ( .B1(DATAI_1_), .B2(keyinput_f31), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_f53), .A(n20844), .ZN(n20845)
         );
  NOR4_X1 U23767 ( .A1(n20848), .A2(n20847), .A3(n20846), .A4(n20845), .ZN(
        n20867) );
  AOI22_X1 U23768 ( .A1(keyinput_f47), .A2(P1_W_R_N_REG_SCAN_IN), .B1(
        DATAI_10_), .B2(keyinput_f22), .ZN(n20849) );
  OAI221_X1 U23769 ( .B1(keyinput_f47), .B2(P1_W_R_N_REG_SCAN_IN), .C1(
        DATAI_10_), .C2(keyinput_f22), .A(n20849), .ZN(n20856) );
  AOI22_X1 U23770 ( .A1(keyinput_f51), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        DATAI_24_), .B2(keyinput_f8), .ZN(n20850) );
  OAI221_X1 U23771 ( .B1(keyinput_f51), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), 
        .C1(DATAI_24_), .C2(keyinput_f8), .A(n20850), .ZN(n20855) );
  AOI22_X1 U23772 ( .A1(DATAI_21_), .A2(keyinput_f11), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_f59), .ZN(n20851) );
  OAI221_X1 U23773 ( .B1(DATAI_21_), .B2(keyinput_f11), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_f59), .A(n20851), .ZN(n20854)
         );
  AOI22_X1 U23774 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_f45), .B1(DATAI_8_), 
        .B2(keyinput_f24), .ZN(n20852) );
  OAI221_X1 U23775 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_f45), .C1(DATAI_8_), .C2(keyinput_f24), .A(n20852), .ZN(n20853) );
  NOR4_X1 U23776 ( .A1(n20856), .A2(n20855), .A3(n20854), .A4(n20853), .ZN(
        n20866) );
  AOI22_X1 U23777 ( .A1(keyinput_f48), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        DATAI_25_), .B2(keyinput_f7), .ZN(n20857) );
  OAI221_X1 U23778 ( .B1(keyinput_f48), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), 
        .C1(DATAI_25_), .C2(keyinput_f7), .A(n20857), .ZN(n20864) );
  AOI22_X1 U23779 ( .A1(keyinput_f50), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        DATAI_6_), .B2(keyinput_f26), .ZN(n20858) );
  OAI221_X1 U23780 ( .B1(keyinput_f50), .B2(P1_BYTEENABLE_REG_2__SCAN_IN), 
        .C1(DATAI_6_), .C2(keyinput_f26), .A(n20858), .ZN(n20863) );
  AOI22_X1 U23781 ( .A1(DATAI_28_), .A2(keyinput_f4), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_f60), .ZN(n20859) );
  OAI221_X1 U23782 ( .B1(DATAI_28_), .B2(keyinput_f4), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_f60), .A(n20859), .ZN(n20862)
         );
  AOI22_X1 U23783 ( .A1(DATAI_12_), .A2(keyinput_f20), .B1(DATAI_29_), .B2(
        keyinput_f3), .ZN(n20860) );
  OAI221_X1 U23784 ( .B1(DATAI_12_), .B2(keyinput_f20), .C1(DATAI_29_), .C2(
        keyinput_f3), .A(n20860), .ZN(n20861) );
  NOR4_X1 U23785 ( .A1(n20864), .A2(n20863), .A3(n20862), .A4(n20861), .ZN(
        n20865) );
  NAND4_X1 U23786 ( .A1(n20868), .A2(n20867), .A3(n20866), .A4(n20865), .ZN(
        n20920) );
  INV_X1 U23787 ( .A(DATAI_3_), .ZN(n20871) );
  INV_X1 U23788 ( .A(DATAI_0_), .ZN(n20870) );
  AOI22_X1 U23789 ( .A1(n20871), .A2(keyinput_f29), .B1(keyinput_f32), .B2(
        n20870), .ZN(n20869) );
  OAI221_X1 U23790 ( .B1(n20871), .B2(keyinput_f29), .C1(n20870), .C2(
        keyinput_f32), .A(n20869), .ZN(n20880) );
  AOI22_X1 U23791 ( .A1(n20873), .A2(keyinput_f23), .B1(keyinput_f14), .B2(
        n20947), .ZN(n20872) );
  OAI221_X1 U23792 ( .B1(n20873), .B2(keyinput_f23), .C1(n20947), .C2(
        keyinput_f14), .A(n20872), .ZN(n20879) );
  INV_X1 U23793 ( .A(DATAI_2_), .ZN(n20875) );
  AOI22_X1 U23794 ( .A1(n20875), .A2(keyinput_f30), .B1(keyinput_f33), .B2(
        n20976), .ZN(n20874) );
  OAI221_X1 U23795 ( .B1(n20875), .B2(keyinput_f30), .C1(n20976), .C2(
        keyinput_f33), .A(n20874), .ZN(n20878) );
  INV_X1 U23796 ( .A(READY2), .ZN(n20967) );
  AOI22_X1 U23797 ( .A1(n20967), .A2(keyinput_f37), .B1(keyinput_f39), .B2(
        n20977), .ZN(n20876) );
  OAI221_X1 U23798 ( .B1(n20967), .B2(keyinput_f37), .C1(n20977), .C2(
        keyinput_f39), .A(n20876), .ZN(n20877) );
  NOR4_X1 U23799 ( .A1(n20880), .A2(n20879), .A3(n20878), .A4(n20877), .ZN(
        n20918) );
  AOI22_X1 U23800 ( .A1(n20927), .A2(keyinput_f18), .B1(n20882), .B2(
        keyinput_f58), .ZN(n20881) );
  OAI221_X1 U23801 ( .B1(n20927), .B2(keyinput_f18), .C1(n20882), .C2(
        keyinput_f58), .A(n20881), .ZN(n20892) );
  AOI22_X1 U23802 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_f46), .B1(n20884), 
        .B2(keyinput_f63), .ZN(n20883) );
  OAI221_X1 U23803 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .C1(n20884), 
        .C2(keyinput_f63), .A(n20883), .ZN(n20891) );
  AOI22_X1 U23804 ( .A1(n20886), .A2(keyinput_f12), .B1(n20970), .B2(
        keyinput_f19), .ZN(n20885) );
  OAI221_X1 U23805 ( .B1(n20886), .B2(keyinput_f12), .C1(n20970), .C2(
        keyinput_f19), .A(n20885), .ZN(n20890) );
  AOI22_X1 U23806 ( .A1(n20888), .A2(keyinput_f5), .B1(n20943), .B2(
        keyinput_f56), .ZN(n20887) );
  OAI221_X1 U23807 ( .B1(n20888), .B2(keyinput_f5), .C1(n20943), .C2(
        keyinput_f56), .A(n20887), .ZN(n20889) );
  NOR4_X1 U23808 ( .A1(n20892), .A2(n20891), .A3(n20890), .A4(n20889), .ZN(
        n20917) );
  INV_X1 U23809 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n20961) );
  INV_X1 U23810 ( .A(keyinput_f35), .ZN(n20894) );
  AOI22_X1 U23811 ( .A1(n20961), .A2(keyinput_f38), .B1(BS16), .B2(n20894), 
        .ZN(n20893) );
  OAI221_X1 U23812 ( .B1(n20961), .B2(keyinput_f38), .C1(n20894), .C2(BS16), 
        .A(n20893), .ZN(n20903) );
  AOI22_X1 U23813 ( .A1(n20974), .A2(keyinput_f44), .B1(keyinput_f2), .B2(
        n20933), .ZN(n20895) );
  OAI221_X1 U23814 ( .B1(n20974), .B2(keyinput_f44), .C1(n20933), .C2(
        keyinput_f2), .A(n20895), .ZN(n20902) );
  INV_X1 U23815 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20897) );
  AOI22_X1 U23816 ( .A1(n20897), .A2(keyinput_f0), .B1(keyinput_f42), .B2(
        n20946), .ZN(n20896) );
  OAI221_X1 U23817 ( .B1(n20897), .B2(keyinput_f0), .C1(n20946), .C2(
        keyinput_f42), .A(n20896), .ZN(n20901) );
  AOI22_X1 U23818 ( .A1(n20957), .A2(keyinput_f6), .B1(n20899), .B2(
        keyinput_f62), .ZN(n20898) );
  OAI221_X1 U23819 ( .B1(n20957), .B2(keyinput_f6), .C1(n20899), .C2(
        keyinput_f62), .A(n20898), .ZN(n20900) );
  NOR4_X1 U23820 ( .A1(n20903), .A2(n20902), .A3(n20901), .A4(n20900), .ZN(
        n20916) );
  INV_X1 U23821 ( .A(DATAI_15_), .ZN(n20906) );
  AOI22_X1 U23822 ( .A1(n20906), .A2(keyinput_f17), .B1(n20905), .B2(
        keyinput_f57), .ZN(n20904) );
  OAI221_X1 U23823 ( .B1(n20906), .B2(keyinput_f17), .C1(n20905), .C2(
        keyinput_f57), .A(n20904), .ZN(n20914) );
  AOI22_X1 U23824 ( .A1(n13208), .A2(keyinput_f27), .B1(keyinput_f16), .B2(
        n20930), .ZN(n20907) );
  OAI221_X1 U23825 ( .B1(n13208), .B2(keyinput_f27), .C1(n20930), .C2(
        keyinput_f16), .A(n20907), .ZN(n20913) );
  INV_X1 U23826 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n20909) );
  AOI22_X1 U23827 ( .A1(n13215), .A2(keyinput_f25), .B1(keyinput_f40), .B2(
        n20909), .ZN(n20908) );
  OAI221_X1 U23828 ( .B1(n13215), .B2(keyinput_f25), .C1(n20909), .C2(
        keyinput_f40), .A(n20908), .ZN(n20912) );
  INV_X1 U23829 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20932) );
  AOI22_X1 U23830 ( .A1(n20932), .A2(keyinput_f61), .B1(keyinput_f43), .B2(
        n20953), .ZN(n20910) );
  OAI221_X1 U23831 ( .B1(n20932), .B2(keyinput_f61), .C1(n20953), .C2(
        keyinput_f43), .A(n20910), .ZN(n20911) );
  NOR4_X1 U23832 ( .A1(n20914), .A2(n20913), .A3(n20912), .A4(n20911), .ZN(
        n20915) );
  NAND4_X1 U23833 ( .A1(n20918), .A2(n20917), .A3(n20916), .A4(n20915), .ZN(
        n20919) );
  OAI22_X1 U23834 ( .A1(keyinput_f21), .A2(n13221), .B1(n20920), .B2(n20919), 
        .ZN(n20921) );
  AOI21_X1 U23835 ( .B1(keyinput_f21), .B2(n13221), .A(n20921), .ZN(n21025) );
  AOI22_X1 U23836 ( .A1(n20924), .A2(keyinput_g54), .B1(keyinput_g47), .B2(
        n20923), .ZN(n20922) );
  OAI221_X1 U23837 ( .B1(n20924), .B2(keyinput_g54), .C1(n20923), .C2(
        keyinput_g47), .A(n20922), .ZN(n20937) );
  AOI22_X1 U23838 ( .A1(n20927), .A2(keyinput_g18), .B1(keyinput_g51), .B2(
        n20926), .ZN(n20925) );
  OAI221_X1 U23839 ( .B1(n20927), .B2(keyinput_g18), .C1(n20926), .C2(
        keyinput_g51), .A(n20925), .ZN(n20936) );
  AOI22_X1 U23840 ( .A1(n20930), .A2(keyinput_g16), .B1(keyinput_g50), .B2(
        n20929), .ZN(n20928) );
  OAI221_X1 U23841 ( .B1(n20930), .B2(keyinput_g16), .C1(n20929), .C2(
        keyinput_g50), .A(n20928), .ZN(n20935) );
  AOI22_X1 U23842 ( .A1(n20933), .A2(keyinput_g2), .B1(n20932), .B2(
        keyinput_g61), .ZN(n20931) );
  OAI221_X1 U23843 ( .B1(n20933), .B2(keyinput_g2), .C1(n20932), .C2(
        keyinput_g61), .A(n20931), .ZN(n20934) );
  NOR4_X1 U23844 ( .A1(n20937), .A2(n20936), .A3(n20935), .A4(n20934), .ZN(
        n20985) );
  INV_X1 U23845 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20940) );
  AOI22_X1 U23846 ( .A1(n20940), .A2(keyinput_g53), .B1(keyinput_g8), .B2(
        n20939), .ZN(n20938) );
  OAI221_X1 U23847 ( .B1(n20940), .B2(keyinput_g53), .C1(n20939), .C2(
        keyinput_g8), .A(n20938), .ZN(n20951) );
  AOI22_X1 U23848 ( .A1(DATAI_28_), .A2(keyinput_g4), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .ZN(n20941) );
  OAI221_X1 U23849 ( .B1(DATAI_28_), .B2(keyinput_g4), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_g59), .A(n20941), .ZN(n20950)
         );
  AOI22_X1 U23850 ( .A1(n20944), .A2(keyinput_g45), .B1(n20943), .B2(
        keyinput_g56), .ZN(n20942) );
  OAI221_X1 U23851 ( .B1(n20944), .B2(keyinput_g45), .C1(n20943), .C2(
        keyinput_g56), .A(n20942), .ZN(n20949) );
  AOI22_X1 U23852 ( .A1(n20947), .A2(keyinput_g14), .B1(keyinput_g42), .B2(
        n20946), .ZN(n20945) );
  OAI221_X1 U23853 ( .B1(n20947), .B2(keyinput_g14), .C1(n20946), .C2(
        keyinput_g42), .A(n20945), .ZN(n20948) );
  NOR4_X1 U23854 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n20984) );
  AOI22_X1 U23855 ( .A1(n14567), .A2(keyinput_g11), .B1(keyinput_g43), .B2(
        n20953), .ZN(n20952) );
  OAI221_X1 U23856 ( .B1(n14567), .B2(keyinput_g11), .C1(n20953), .C2(
        keyinput_g43), .A(n20952), .ZN(n20965) );
  AOI22_X1 U23857 ( .A1(n13208), .A2(keyinput_g27), .B1(keyinput_g35), .B2(
        n20955), .ZN(n20954) );
  OAI221_X1 U23858 ( .B1(n13208), .B2(keyinput_g27), .C1(n20955), .C2(
        keyinput_g35), .A(n20954), .ZN(n20964) );
  AOI22_X1 U23859 ( .A1(n20958), .A2(keyinput_g34), .B1(n20957), .B2(
        keyinput_g6), .ZN(n20956) );
  OAI221_X1 U23860 ( .B1(n20958), .B2(keyinput_g34), .C1(n20957), .C2(
        keyinput_g6), .A(n20956), .ZN(n20963) );
  AOI22_X1 U23861 ( .A1(n20961), .A2(keyinput_g38), .B1(n20960), .B2(
        keyinput_g60), .ZN(n20959) );
  OAI221_X1 U23862 ( .B1(n20961), .B2(keyinput_g38), .C1(n20960), .C2(
        keyinput_g60), .A(n20959), .ZN(n20962) );
  NOR4_X1 U23863 ( .A1(n20965), .A2(n20964), .A3(n20963), .A4(n20962), .ZN(
        n20983) );
  AOI22_X1 U23864 ( .A1(n20968), .A2(keyinput_g46), .B1(n20967), .B2(
        keyinput_g37), .ZN(n20966) );
  OAI221_X1 U23865 ( .B1(n20968), .B2(keyinput_g46), .C1(n20967), .C2(
        keyinput_g37), .A(n20966), .ZN(n20981) );
  INV_X1 U23866 ( .A(DATAI_1_), .ZN(n20971) );
  AOI22_X1 U23867 ( .A1(n20971), .A2(keyinput_g31), .B1(n20970), .B2(
        keyinput_g19), .ZN(n20969) );
  OAI221_X1 U23868 ( .B1(n20971), .B2(keyinput_g31), .C1(n20970), .C2(
        keyinput_g19), .A(n20969), .ZN(n20980) );
  AOI22_X1 U23869 ( .A1(n20974), .A2(keyinput_g44), .B1(keyinput_g1), .B2(
        n20973), .ZN(n20972) );
  OAI221_X1 U23870 ( .B1(n20974), .B2(keyinput_g44), .C1(n20973), .C2(
        keyinput_g1), .A(n20972), .ZN(n20979) );
  AOI22_X1 U23871 ( .A1(n20977), .A2(keyinput_g39), .B1(keyinput_g33), .B2(
        n20976), .ZN(n20975) );
  OAI221_X1 U23872 ( .B1(n20977), .B2(keyinput_g39), .C1(n20976), .C2(
        keyinput_g33), .A(n20975), .ZN(n20978) );
  NOR4_X1 U23873 ( .A1(n20981), .A2(n20980), .A3(n20979), .A4(n20978), .ZN(
        n20982) );
  NAND4_X1 U23874 ( .A1(n20985), .A2(n20984), .A3(n20983), .A4(n20982), .ZN(
        n21023) );
  AOI22_X1 U23875 ( .A1(DATAI_23_), .A2(keyinput_g9), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .ZN(n20986) );
  OAI221_X1 U23876 ( .B1(DATAI_23_), .B2(keyinput_g9), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_g62), .A(n20986), .ZN(n20993)
         );
  AOI22_X1 U23877 ( .A1(DATAI_17_), .A2(keyinput_g15), .B1(DATAI_27_), .B2(
        keyinput_g5), .ZN(n20987) );
  OAI221_X1 U23878 ( .B1(DATAI_17_), .B2(keyinput_g15), .C1(DATAI_27_), .C2(
        keyinput_g5), .A(n20987), .ZN(n20992) );
  AOI22_X1 U23879 ( .A1(DATAI_22_), .A2(keyinput_g10), .B1(DATAI_8_), .B2(
        keyinput_g24), .ZN(n20988) );
  OAI221_X1 U23880 ( .B1(DATAI_22_), .B2(keyinput_g10), .C1(DATAI_8_), .C2(
        keyinput_g24), .A(n20988), .ZN(n20991) );
  AOI22_X1 U23881 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_g40), .B1(
        DATAI_12_), .B2(keyinput_g20), .ZN(n20989) );
  OAI221_X1 U23882 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_g40), .C1(
        DATAI_12_), .C2(keyinput_g20), .A(n20989), .ZN(n20990) );
  NOR4_X1 U23883 ( .A1(n20993), .A2(n20992), .A3(n20991), .A4(n20990), .ZN(
        n21021) );
  XOR2_X1 U23884 ( .A(n13215), .B(keyinput_g25), .Z(n21001) );
  AOI22_X1 U23885 ( .A1(DATAI_19_), .A2(keyinput_g13), .B1(n20995), .B2(
        keyinput_g22), .ZN(n20994) );
  OAI221_X1 U23886 ( .B1(DATAI_19_), .B2(keyinput_g13), .C1(n20995), .C2(
        keyinput_g22), .A(n20994), .ZN(n21000) );
  AOI22_X1 U23887 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g48), .B1(
        DATAI_20_), .B2(keyinput_g12), .ZN(n20996) );
  OAI221_X1 U23888 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g48), 
        .C1(DATAI_20_), .C2(keyinput_g12), .A(n20996), .ZN(n20999) );
  AOI22_X1 U23889 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        DATAI_0_), .B2(keyinput_g32), .ZN(n20997) );
  OAI221_X1 U23890 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        DATAI_0_), .C2(keyinput_g32), .A(n20997), .ZN(n20998) );
  NOR4_X1 U23891 ( .A1(n21001), .A2(n21000), .A3(n20999), .A4(n20998), .ZN(
        n21020) );
  AOI22_X1 U23892 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        DATAI_4_), .B2(keyinput_g28), .ZN(n21002) );
  OAI221_X1 U23893 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        DATAI_4_), .C2(keyinput_g28), .A(n21002), .ZN(n21009) );
  AOI22_X1 U23894 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g49), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .ZN(n21003) );
  OAI221_X1 U23895 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g49), 
        .C1(P1_REIP_REG_28__SCAN_IN), .C2(keyinput_g55), .A(n21003), .ZN(
        n21008) );
  AOI22_X1 U23896 ( .A1(DATAI_2_), .A2(keyinput_g30), .B1(DATAI_3_), .B2(
        keyinput_g29), .ZN(n21004) );
  OAI221_X1 U23897 ( .B1(DATAI_2_), .B2(keyinput_g30), .C1(DATAI_3_), .C2(
        keyinput_g29), .A(n21004), .ZN(n21007) );
  AOI22_X1 U23898 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_g57), .B1(
        READY1), .B2(keyinput_g36), .ZN(n21005) );
  OAI221_X1 U23899 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .C1(
        READY1), .C2(keyinput_g36), .A(n21005), .ZN(n21006) );
  NOR4_X1 U23900 ( .A1(n21009), .A2(n21008), .A3(n21007), .A4(n21006), .ZN(
        n21019) );
  AOI22_X1 U23901 ( .A1(DATAI_9_), .A2(keyinput_g23), .B1(DATAI_29_), .B2(
        keyinput_g3), .ZN(n21010) );
  OAI221_X1 U23902 ( .B1(DATAI_9_), .B2(keyinput_g23), .C1(DATAI_29_), .C2(
        keyinput_g3), .A(n21010), .ZN(n21017) );
  AOI22_X1 U23903 ( .A1(DATAI_6_), .A2(keyinput_g26), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .ZN(n21011) );
  OAI221_X1 U23904 ( .B1(DATAI_6_), .B2(keyinput_g26), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_g63), .A(n21011), .ZN(n21016)
         );
  AOI22_X1 U23905 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(DATAI_25_), .B2(
        keyinput_g7), .ZN(n21012) );
  OAI221_X1 U23906 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(DATAI_25_), .C2(
        keyinput_g7), .A(n21012), .ZN(n21015) );
  AOI22_X1 U23907 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_g58), .B1(
        P1_REIP_REG_31__SCAN_IN), .B2(keyinput_g52), .ZN(n21013) );
  OAI221_X1 U23908 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_g58), .C1(
        P1_REIP_REG_31__SCAN_IN), .C2(keyinput_g52), .A(n21013), .ZN(n21014)
         );
  NOR4_X1 U23909 ( .A1(n21017), .A2(n21016), .A3(n21015), .A4(n21014), .ZN(
        n21018) );
  NAND4_X1 U23910 ( .A1(n21021), .A2(n21020), .A3(n21019), .A4(n21018), .ZN(
        n21022) );
  OAI22_X1 U23911 ( .A1(keyinput_g21), .A2(n13221), .B1(n21023), .B2(n21022), 
        .ZN(n21024) );
  AOI211_X1 U23912 ( .C1(keyinput_g21), .C2(n13221), .A(n21025), .B(n21024), 
        .ZN(n21027) );
  AOI22_X1 U23913 ( .A1(n16513), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16515), .ZN(n21026) );
  XNOR2_X1 U23914 ( .A(n21027), .B(n21026), .ZN(U355) );
  CLKBUF_X3 U11167 ( .A(n11064), .Z(n9643) );
  CLKBUF_X3 U11168 ( .A(n11064), .Z(n9644) );
  NAND4_X1 U15189 ( .A1(n18852), .A2(n18859), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15668) );
  INV_X1 U13245 ( .A(n13122), .ZN(n10359) );
  BUF_X1 U11221 ( .A(n11829), .Z(n12036) );
  OAI21_X1 U11305 ( .B1(n13176), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10467), 
        .ZN(n10594) );
  CLKBUF_X1 U11093 ( .A(n10330), .Z(n11056) );
  CLKBUF_X1 U11110 ( .A(n11013), .Z(n10908) );
  CLKBUF_X2 U11114 ( .A(n10330), .Z(n11032) );
  CLKBUF_X1 U11131 ( .A(n10603), .Z(n9664) );
  NAND4_X1 U11138 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n10247), .ZN(
        n13426) );
  OR2_X1 U11156 ( .A1(n13388), .A2(n13389), .ZN(n19380) );
  XOR2_X1 U11162 ( .A(n12553), .B(n12552), .Z(n17859) );
  CLKBUF_X1 U11165 ( .A(n13171), .Z(n14068) );
  NAND2_X1 U11171 ( .A1(n14525), .A2(n10423), .ZN(n10409) );
  CLKBUF_X2 U11203 ( .A(n11172), .Z(n13507) );
  CLKBUF_X1 U11207 ( .A(n13601), .Z(n19111) );
  INV_X4 U11212 ( .A(n14206), .ZN(n15154) );
  OR2_X1 U11215 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12269), .ZN(
        n12307) );
  CLKBUF_X1 U11424 ( .A(n12296), .Z(n17190) );
  CLKBUF_X1 U11451 ( .A(n10258), .Z(n17133) );
  INV_X1 U11721 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18866) );
  OR2_X2 U12417 ( .A1(n12268), .A2(n12267), .ZN(n21028) );
endmodule

