

module b20_C_gen_AntiSAT_k_256_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4511, n4514, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684;

  INV_X1 U5017 ( .A(n8664), .ZN(n8645) );
  NAND3_X1 U5018 ( .A1(n6227), .A2(n6226), .A3(n8910), .ZN(n9047) );
  NAND2_X2 U5019 ( .A1(n5474), .A2(n5473), .ZN(n10194) );
  INV_X1 U5020 ( .A(n6873), .ZN(n5591) );
  INV_X1 U5023 ( .A(n6042), .ZN(n6400) );
  AND2_X2 U5025 ( .A1(n8318), .A2(n5285), .ZN(n6876) );
  NAND2_X1 U5026 ( .A1(n5885), .A2(n6542), .ZN(n5943) );
  INV_X1 U5028 ( .A(n6218), .ZN(n5926) );
  CLKBUF_X1 U5029 ( .A(n9979), .Z(n4511) );
  NOR2_X1 U5030 ( .A1(n9991), .A2(n7511), .ZN(n9979) );
  NAND2_X1 U5031 ( .A1(n5918), .A2(n5943), .ZN(n5970) );
  INV_X1 U5032 ( .A(n5285), .ZN(n5287) );
  INV_X1 U5033 ( .A(n6678), .ZN(n5590) );
  NAND2_X1 U5034 ( .A1(n6222), .A2(n6225), .ZN(n9044) );
  OR2_X1 U5035 ( .A1(n9623), .A2(n9613), .ZN(n9609) );
  INV_X2 U5037 ( .A(n8281), .ZN(n7421) );
  INV_X1 U5038 ( .A(n6876), .ZN(n5343) );
  BUF_X1 U5039 ( .A(n6965), .Z(n4637) );
  NAND2_X1 U5040 ( .A1(n7999), .A2(n8000), .ZN(n7998) );
  INV_X1 U5041 ( .A(n9352), .ZN(n7594) );
  NAND2_X1 U5042 ( .A1(n6990), .A2(n9058), .ZN(n6073) );
  INV_X1 U5043 ( .A(n6496), .ZN(n10012) );
  NAND2_X1 U5044 ( .A1(n5093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4853) );
  XNOR2_X1 U5045 ( .A(n5891), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6471) );
  XNOR2_X1 U5046 ( .A(n5430), .B(n5429), .ZN(n6990) );
  INV_X1 U5047 ( .A(n4649), .ZN(n6272) );
  OR2_X1 U5048 ( .A1(n4525), .A2(n9870), .ZN(P1_U3517) );
  OR2_X1 U5049 ( .A1(n4524), .A2(n9782), .ZN(P1_U3549) );
  NAND2_X2 U5050 ( .A1(n7766), .A2(n9083), .ZN(n7765) );
  NAND2_X2 U5051 ( .A1(n7679), .A2(n6509), .ZN(n7766) );
  XNOR2_X2 U5052 ( .A(n6641), .B(n6637), .ZN(n8213) );
  OAI21_X2 U5053 ( .B1(n7711), .B2(n4528), .A(n4738), .ZN(n7883) );
  AND2_X1 U5054 ( .A1(n8223), .A2(n8315), .ZN(n4514) );
  NAND2_X4 U5055 ( .A1(n6073), .A2(n6072), .ZN(n9131) );
  NAND4_X2 U5057 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n9354)
         );
  XNOR2_X2 U5058 ( .A(n5907), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5908) );
  AOI21_X2 U5059 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7067), .A(n7972), .ZN(
        n6705) );
  OR2_X1 U5060 ( .A1(n10107), .A2(n7418), .ZN(n4817) );
  OAI21_X2 U5061 ( .B1(n5002), .B2(P2_RD_REG_SCAN_IN), .A(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U5062 ( .A1(n9044), .A2(n9043), .ZN(n9042) );
  OAI21_X1 U5063 ( .B1(n8690), .B2(n4888), .A(n4615), .ZN(n8673) );
  AND2_X1 U5064 ( .A1(n9047), .A2(n4598), .ZN(n4732) );
  OAI21_X1 U5065 ( .B1(n8444), .B2(n8502), .A(n8727), .ZN(n8715) );
  NAND2_X1 U5066 ( .A1(n9692), .A2(n9695), .ZN(n9691) );
  NAND2_X1 U5067 ( .A1(n7984), .A2(n6555), .ZN(n9725) );
  NAND2_X1 U5068 ( .A1(n4944), .A2(n4943), .ZN(n8114) );
  NAND2_X1 U5069 ( .A1(n6505), .A2(n6504), .ZN(n7392) );
  NAND2_X1 U5070 ( .A1(n5689), .A2(n5688), .ZN(n8648) );
  NOR2_X2 U5071 ( .A1(n5687), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5704) );
  NOR2_X1 U5072 ( .A1(n7566), .A2(n7820), .ZN(n7565) );
  OR2_X2 U5073 ( .A1(n5619), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5631) );
  INV_X1 U5074 ( .A(n10131), .ZN(n10157) );
  INV_X1 U5075 ( .A(n10029), .ZN(n9971) );
  NAND2_X1 U5076 ( .A1(n6547), .A2(n7577), .ZN(n9064) );
  INV_X1 U5077 ( .A(n9355), .ZN(n7579) );
  CLKBUF_X3 U5078 ( .A(n5970), .Z(n5987) );
  INV_X1 U5079 ( .A(n8513), .ZN(n7500) );
  INV_X1 U5080 ( .A(n7422), .ZN(n7620) );
  INV_X1 U5081 ( .A(n6881), .ZN(n5775) );
  INV_X1 U5082 ( .A(n6218), .ZN(n4516) );
  XNOR2_X1 U5083 ( .A(n5324), .B(n5323), .ZN(n6685) );
  INV_X2 U5084 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OAI21_X1 U5085 ( .B1(n9590), .B2(n9589), .A(n4990), .ZN(n9577) );
  NOR2_X1 U5086 ( .A1(n8615), .A2(n4518), .ZN(n4572) );
  NAND2_X1 U5087 ( .A1(n6526), .A2(n5166), .ZN(n4989) );
  MUX2_X1 U5088 ( .A(n8854), .B(n8853), .S(n10196), .Z(n8855) );
  MUX2_X1 U5089 ( .A(n8796), .B(n8853), .S(n10213), .Z(n8797) );
  AOI22_X1 U5090 ( .A1(n8631), .A2(n5712), .B1(n8646), .B2(n8843), .ZN(n5725)
         );
  CLKBUF_X1 U5091 ( .A(n9696), .Z(n4636) );
  OAI22_X1 U5092 ( .A1(n9705), .A2(n6521), .B1(n9737), .B2(n9720), .ZN(n9696)
         );
  NAND2_X1 U5093 ( .A1(n4733), .A2(n4570), .ZN(n9015) );
  NAND2_X1 U5094 ( .A1(n9042), .A2(n4732), .ZN(n4733) );
  NAND2_X1 U5095 ( .A1(n9691), .A2(n5049), .ZN(n9674) );
  NAND2_X1 U5096 ( .A1(n4786), .A2(n4791), .ZN(n4785) );
  NAND2_X1 U5097 ( .A1(n6888), .A2(n6854), .ZN(n6916) );
  NAND2_X1 U5098 ( .A1(n9725), .A2(n6557), .ZN(n9726) );
  AOI21_X1 U5099 ( .B1(n6839), .B2(n6840), .A(n4788), .ZN(n4787) );
  NAND2_X1 U5100 ( .A1(n5092), .A2(n5091), .ZN(n5090) );
  OR2_X1 U5101 ( .A1(n8106), .A2(n8105), .ZN(n5092) );
  OR2_X1 U5102 ( .A1(n6836), .A2(n8664), .ZN(n6838) );
  OR2_X1 U5103 ( .A1(n8009), .A2(n4945), .ZN(n4944) );
  OR2_X1 U5104 ( .A1(n7841), .A2(n9927), .ZN(n7912) );
  AND2_X1 U5105 ( .A1(n5710), .A2(n5709), .ZN(n5766) );
  NAND2_X1 U5106 ( .A1(n6233), .A2(n6232), .ZN(n8964) );
  AND2_X1 U5107 ( .A1(n5704), .A2(n8335), .ZN(n8620) );
  NAND2_X2 U5108 ( .A1(n5462), .A2(n5461), .ZN(n8237) );
  NAND2_X1 U5109 ( .A1(n5543), .A2(n5542), .ZN(n8244) );
  NAND2_X1 U5110 ( .A1(n6151), .A2(n6150), .ZN(n7791) );
  NOR2_X1 U5111 ( .A1(n7565), .A2(n6699), .ZN(n7721) );
  XNOR2_X1 U5112 ( .A(n5456), .B(n5455), .ZN(n7101) );
  NAND2_X1 U5113 ( .A1(n6134), .A2(n6133), .ZN(n7543) );
  NAND2_X1 U5114 ( .A1(n6113), .A2(n6112), .ZN(n7870) );
  NOR2_X2 U5115 ( .A1(n5631), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5651) );
  AND2_X1 U5116 ( .A1(n5433), .A2(n5432), .ZN(n7861) );
  NOR2_X1 U5117 ( .A1(n7367), .A2(n6697), .ZN(n6698) );
  NAND2_X1 U5118 ( .A1(n6094), .A2(n6093), .ZN(n7442) );
  NAND2_X1 U5119 ( .A1(n10076), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n4640) );
  NAND4_X1 U5120 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n10029)
         );
  OR2_X1 U5121 ( .A1(n6980), .A2(n6535), .ZN(n6030) );
  OAI211_X1 U5122 ( .C1(n6678), .C2(n6685), .A(n5330), .B(n5329), .ZN(n7345)
         );
  INV_X1 U5123 ( .A(n6239), .ZN(n6413) );
  AND2_X2 U5124 ( .A1(n7020), .A2(n6962), .ZN(P1_U3973) );
  INV_X2 U5125 ( .A(n5328), .ZN(n6875) );
  AOI21_X1 U5126 ( .B1(n4588), .B2(n5021), .A(n5522), .ZN(n4703) );
  NAND2_X2 U5127 ( .A1(n5286), .A2(n5285), .ZN(n6881) );
  NAND2_X2 U5128 ( .A1(n5286), .A2(n5287), .ZN(n5562) );
  NAND2_X2 U5129 ( .A1(n6678), .A2(n4637), .ZN(n6873) );
  NAND2_X1 U5130 ( .A1(n6678), .A2(n5176), .ZN(n5328) );
  NAND2_X1 U5131 ( .A1(n5190), .A2(n5189), .ZN(n5392) );
  AND2_X1 U5132 ( .A1(n5021), .A2(n4706), .ZN(n4705) );
  INV_X1 U5133 ( .A(n5773), .ZN(n6925) );
  NAND2_X2 U5134 ( .A1(n5772), .A2(n5773), .ZN(n6678) );
  CLKBUF_X1 U5135 ( .A(n6190), .Z(n9060) );
  INV_X1 U5136 ( .A(n6190), .ZN(n6172) );
  CLKBUF_X3 U5137 ( .A(n6272), .Z(n4526) );
  AOI21_X1 U5138 ( .B1(n5010), .B2(n5008), .A(n5007), .ZN(n5006) );
  NAND2_X1 U5139 ( .A1(n9906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U5140 ( .A(n5483), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U5141 ( .A1(n6450), .A2(n5883), .ZN(n7018) );
  XNOR2_X1 U5142 ( .A(n5855), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9249) );
  NOR2_X1 U5143 ( .A1(n5788), .A2(n5269), .ZN(n5797) );
  NAND2_X1 U5144 ( .A1(n4728), .A2(n5879), .ZN(n7982) );
  NAND2_X1 U5145 ( .A1(n5854), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5855) );
  INV_X2 U5146 ( .A(n7295), .ZN(n4517) );
  OAI21_X1 U5147 ( .B1(n4727), .B2(n6130), .A(n4587), .ZN(n5879) );
  XNOR2_X1 U5148 ( .A(n5195), .B(n10454), .ZN(n5412) );
  NAND2_X1 U5149 ( .A1(n5393), .A2(n5260), .ZN(n5409) );
  NOR2_X1 U5150 ( .A1(n5265), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5130) );
  AND2_X1 U5151 ( .A1(n6026), .A2(n5867), .ZN(n6052) );
  AND3_X1 U5152 ( .A1(n4856), .A2(n4855), .A3(n4854), .ZN(n5264) );
  INV_X1 U5153 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10606) );
  INV_X1 U5154 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5867) );
  INV_X1 U5155 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5346) );
  INV_X1 U5156 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5323) );
  INV_X2 U5157 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5158 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4856) );
  INV_X1 U5159 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4855) );
  INV_X1 U5160 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4854) );
  INV_X2 U5161 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5861) );
  NOR2_X1 U5162 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5837) );
  INV_X1 U5163 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6206) );
  INV_X1 U5164 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U5165 ( .A1(n6841), .A2(n4784), .ZN(n4783) );
  AND2_X1 U5166 ( .A1(n4791), .A2(n6839), .ZN(n4784) );
  NAND2_X1 U5167 ( .A1(n4519), .A2(n4958), .ZN(n4518) );
  NAND2_X1 U5168 ( .A1(n8616), .A2(n8617), .ZN(n4519) );
  NOR2_X2 U5169 ( .A1(n8612), .A2(n6714), .ZN(n6717) );
  NAND2_X1 U5170 ( .A1(n4986), .A2(n4523), .ZN(n4520) );
  AND2_X2 U5171 ( .A1(n4520), .A2(n4521), .ZN(n9647) );
  OR2_X1 U5172 ( .A1(n4522), .A2(n6524), .ZN(n4521) );
  INV_X1 U5173 ( .A(n6525), .ZN(n4522) );
  AND2_X1 U5174 ( .A1(n4983), .A2(n6525), .ZN(n4523) );
  NAND2_X1 U5175 ( .A1(n10103), .A2(n10102), .ZN(n10101) );
  AND2_X1 U5177 ( .A1(n9798), .A2(n9871), .ZN(n4524) );
  MUX2_X1 U5178 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9869), .S(n10094), .Z(n9782) );
  NOR2_X1 U5179 ( .A1(n5500), .A2(n5499), .ZN(n5161) );
  AOI21_X2 U5180 ( .B1(n4693), .B2(n4695), .A(n4581), .ZN(n4691) );
  AOI22_X2 U5181 ( .A1(n8715), .A2(n6895), .B1(n8708), .B2(n8881), .ZN(n8704)
         );
  AND2_X1 U5182 ( .A1(n9879), .A2(n9871), .ZN(n4525) );
  MUX2_X1 U5183 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9869), .S(n10078), .Z(n9870) );
  NOR2_X1 U5184 ( .A1(n5596), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5311) );
  OR2_X2 U5185 ( .A1(n5663), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5687) );
  NOR2_X2 U5186 ( .A1(n5544), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5559) );
  OR2_X1 U5187 ( .A1(n9750), .A2(n5919), .ZN(n6494) );
  INV_X1 U5188 ( .A(n9750), .ZN(n7125) );
  NAND2_X2 U5189 ( .A1(n5895), .A2(n5832), .ZN(n5951) );
  XNOR2_X2 U5190 ( .A(n8849), .B(n8633), .ZN(n8644) );
  NAND2_X4 U5191 ( .A1(n5694), .A2(n5693), .ZN(n8633) );
  OAI221_X1 U5192 ( .B1(n10390), .B2(keyinput_g39), .C1(n5868), .C2(
        keyinput_g111), .A(n10389), .ZN(n10400) );
  INV_X2 U5193 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5868) );
  NOR2_X4 U5194 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5895) );
  XNOR2_X2 U5195 ( .A(n6539), .B(n9096), .ZN(n8312) );
  INV_X2 U5196 ( .A(n5909), .ZN(n8223) );
  AND2_X4 U5197 ( .A1(n5908), .A2(n8223), .ZN(n5991) );
  NAND2_X1 U5198 ( .A1(n5909), .A2(n5908), .ZN(n6239) );
  NAND2_X2 U5199 ( .A1(n6471), .A2(n9300), .ZN(n4649) );
  INV_X1 U5200 ( .A(n6218), .ZN(n4527) );
  NAND2_X1 U5201 ( .A1(n5909), .A2(n8315), .ZN(n6218) );
  AOI21_X1 U5202 ( .B1(n5025), .B2(n5026), .A(n5455), .ZN(n5023) );
  NOR2_X1 U5203 ( .A1(n5429), .A2(n5011), .ZN(n5010) );
  INV_X1 U5204 ( .A(n5197), .ZN(n5011) );
  AND2_X1 U5205 ( .A1(n10125), .A2(n6751), .ZN(n6749) );
  NAND2_X1 U5206 ( .A1(n7700), .A2(n7547), .ZN(n7216) );
  OR2_X1 U5207 ( .A1(n8756), .A2(n5602), .ZN(n4878) );
  AND2_X1 U5208 ( .A1(n5345), .A2(n4593), .ZN(n5393) );
  INV_X1 U5209 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5126) );
  AND2_X1 U5210 ( .A1(n5035), .A2(n5256), .ZN(n5034) );
  NAND2_X1 U5211 ( .A1(n5613), .A2(n5252), .ZN(n5035) );
  OAI211_X1 U5212 ( .C1(n5000), .C2(n6948), .A(n4998), .B(n4999), .ZN(n4792)
         );
  NOR2_X1 U5213 ( .A1(n6889), .A2(n6946), .ZN(n4999) );
  NAND2_X1 U5214 ( .A1(n5000), .A2(n6864), .ZN(n4998) );
  INV_X1 U5215 ( .A(n5562), .ZN(n5719) );
  NAND2_X1 U5216 ( .A1(n6706), .A2(n4948), .ZN(n4943) );
  NAND2_X1 U5217 ( .A1(n4948), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4945) );
  INV_X1 U5218 ( .A(n6916), .ZN(n6846) );
  NAND2_X1 U5219 ( .A1(n4649), .A2(n5176), .ZN(n6190) );
  INV_X1 U5220 ( .A(n6789), .ZN(n4802) );
  NOR2_X1 U5221 ( .A1(n6916), .A2(n6845), .ZN(n4791) );
  NAND2_X1 U5222 ( .A1(n5584), .A2(n5236), .ZN(n5039) );
  INV_X1 U5223 ( .A(n9218), .ZN(n4675) );
  NOR2_X1 U5224 ( .A1(n4720), .A2(n5039), .ZN(n4719) );
  INV_X1 U5225 ( .A(n4721), .ZN(n4720) );
  NAND2_X1 U5226 ( .A1(n5023), .A2(n4707), .ZN(n4706) );
  INV_X1 U5227 ( .A(n5211), .ZN(n4707) );
  AOI21_X1 U5228 ( .B1(n5023), .B2(n5024), .A(n4582), .ZN(n5021) );
  INV_X1 U5229 ( .A(n5025), .ZN(n5024) );
  NAND2_X1 U5230 ( .A1(n5199), .A2(n10632), .ZN(n5202) );
  INV_X1 U5231 ( .A(n4928), .ZN(n4926) );
  AOI21_X1 U5232 ( .B1(n8383), .B2(n4906), .A(n4542), .ZN(n4905) );
  OR2_X1 U5233 ( .A1(n8098), .A2(n8127), .ZN(n6772) );
  OR2_X1 U5234 ( .A1(n8294), .A2(n8293), .ZN(n8295) );
  INV_X1 U5235 ( .A(n8629), .ZN(n4698) );
  INV_X1 U5236 ( .A(n8318), .ZN(n5286) );
  NOR2_X1 U5237 ( .A1(n6690), .A2(n7488), .ZN(n6691) );
  NOR2_X1 U5238 ( .A1(n6690), .A2(n6585), .ZN(n6586) );
  NOR2_X1 U5239 ( .A1(n6692), .A2(n6971), .ZN(n6694) );
  NOR2_X1 U5240 ( .A1(n6587), .A2(n6971), .ZN(n6588) );
  NOR2_X1 U5241 ( .A1(n8568), .A2(n4632), .ZN(n6605) );
  NOR2_X1 U5242 ( .A1(n8582), .A2(n8171), .ZN(n4632) );
  NOR2_X1 U5243 ( .A1(n10131), .A2(n8512), .ZN(n4885) );
  NAND2_X1 U5244 ( .A1(n5369), .A2(n5368), .ZN(n4869) );
  INV_X1 U5245 ( .A(n8856), .ZN(n6836) );
  OR2_X1 U5246 ( .A1(n8866), .A2(n8692), .ZN(n6826) );
  NOR2_X1 U5247 ( .A1(n6893), .A2(n5761), .ZN(n5762) );
  AND2_X1 U5248 ( .A1(n8686), .A2(n6827), .ZN(n5761) );
  NOR2_X1 U5249 ( .A1(n5756), .A2(n6819), .ZN(n5757) );
  OR2_X1 U5250 ( .A1(n8444), .A2(n8745), .ZN(n8699) );
  OR2_X1 U5251 ( .A1(n8892), .A2(n8759), .ZN(n6801) );
  NAND2_X1 U5252 ( .A1(n8932), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U5253 ( .A1(n5157), .A2(n5920), .ZN(n5922) );
  XNOR2_X1 U5254 ( .A(n5917), .B(n6438), .ZN(n5924) );
  NAND2_X1 U5255 ( .A1(n5916), .A2(n5915), .ZN(n5917) );
  OR2_X1 U5256 ( .A1(n9871), .A2(n9608), .ZN(n9223) );
  NAND2_X1 U5257 ( .A1(n6850), .A2(n6849), .ZN(n6867) );
  NAND2_X1 U5258 ( .A1(n5017), .A2(SI_29_), .ZN(n6850) );
  XNOR2_X1 U5259 ( .A(n6848), .B(n6847), .ZN(n5017) );
  NAND2_X1 U5260 ( .A1(n5681), .A2(n5680), .ZN(n5697) );
  AOI21_X1 U5261 ( .B1(n5614), .B2(n5032), .A(n5030), .ZN(n5675) );
  AND2_X1 U5262 ( .A1(n5642), .A2(n5252), .ZN(n5032) );
  OAI21_X1 U5263 ( .B1(n5034), .B2(n5031), .A(n5644), .ZN(n5030) );
  INV_X1 U5264 ( .A(n5642), .ZN(n5031) );
  AND2_X1 U5265 ( .A1(n4713), .A2(n4619), .ZN(n4711) );
  NAND2_X1 U5266 ( .A1(n5086), .A2(n5087), .ZN(n6189) );
  AND2_X1 U5267 ( .A1(n5088), .A2(n5870), .ZN(n5087) );
  NOR2_X1 U5268 ( .A1(n5836), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5088) );
  INV_X1 U5269 ( .A(n5023), .ZN(n4708) );
  NAND2_X1 U5270 ( .A1(n5005), .A2(n5003), .ZN(n5502) );
  AOI21_X1 U5271 ( .B1(n5006), .B2(n5009), .A(n5004), .ZN(n5003) );
  INV_X1 U5272 ( .A(n5165), .ZN(n5004) );
  OAI21_X1 U5273 ( .B1(n5391), .B2(n4695), .A(n5412), .ZN(n4694) );
  INV_X1 U5274 ( .A(n5194), .ZN(n4695) );
  AND2_X1 U5275 ( .A1(n4555), .A2(n7218), .ZN(n8281) );
  NAND2_X1 U5276 ( .A1(n8373), .A2(n8434), .ZN(n8300) );
  AND2_X1 U5277 ( .A1(n6772), .A2(n6774), .ZN(n8077) );
  OR2_X1 U5278 ( .A1(n5339), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U5279 ( .A1(n6692), .A2(n6971), .ZN(n6693) );
  AND2_X1 U5280 ( .A1(n4824), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U5281 ( .A1(n7148), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U5282 ( .A1(n4832), .A2(n4831), .ZN(n4952) );
  INV_X1 U5283 ( .A(n8577), .ZN(n4831) );
  AOI21_X1 U5284 ( .B1(n8662), .B2(n8667), .A(n4612), .ZN(n8651) );
  NAND2_X1 U5285 ( .A1(n5583), .A2(n5582), .ZN(n8756) );
  NOR2_X1 U5286 ( .A1(n7814), .A2(n6745), .ZN(n5110) );
  NAND2_X1 U5287 ( .A1(n4887), .A2(n4553), .ZN(n4886) );
  INV_X1 U5288 ( .A(n10117), .ZN(n4887) );
  INV_X1 U5289 ( .A(n10118), .ZN(n8762) );
  OR2_X1 U5290 ( .A1(n8767), .A2(n8744), .ZN(n6805) );
  XNOR2_X1 U5291 ( .A(n5284), .B(n8903), .ZN(n5285) );
  NAND2_X1 U5292 ( .A1(n8905), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5284) );
  INV_X1 U5293 ( .A(n5130), .ZN(n5128) );
  INV_X1 U5294 ( .A(n8932), .ZN(n4759) );
  AND2_X1 U5295 ( .A1(n9056), .A2(n9559), .ZN(n9296) );
  NOR2_X1 U5296 ( .A1(n4772), .A2(n4771), .ZN(n9431) );
  INV_X1 U5297 ( .A(n9434), .ZN(n4771) );
  INV_X1 U5298 ( .A(n4965), .ZN(n4964) );
  NAND2_X1 U5299 ( .A1(n9674), .A2(n9186), .ZN(n9660) );
  NAND2_X1 U5300 ( .A1(n6515), .A2(n6514), .ZN(n7916) );
  AND2_X1 U5301 ( .A1(n9085), .A2(n9276), .ZN(n5062) );
  NAND2_X1 U5302 ( .A1(n6537), .A2(n6536), .ZN(n8307) );
  OR2_X1 U5303 ( .A1(n8319), .A2(n6535), .ZN(n6537) );
  NAND2_X1 U5304 ( .A1(n5029), .A2(n5034), .ZN(n5643) );
  NAND2_X1 U5305 ( .A1(n5036), .A2(n5236), .ZN(n5585) );
  NAND2_X1 U5306 ( .A1(n5231), .A2(n5040), .ZN(n5036) );
  OAI21_X1 U5307 ( .B1(n5426), .B2(n5009), .A(n5006), .ZN(n5441) );
  INV_X1 U5308 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5002) );
  INV_X1 U5309 ( .A(n8849), .ZN(n8360) );
  OR2_X1 U5310 ( .A1(n8009), .A2(n5487), .ZN(n4947) );
  XNOR2_X1 U5311 ( .A(n6705), .B(n8020), .ZN(n8009) );
  OAI21_X1 U5312 ( .B1(n8611), .B2(n10267), .A(n8595), .ZN(n5104) );
  INV_X1 U5313 ( .A(n8613), .ZN(n4818) );
  AOI21_X1 U5314 ( .B1(n5785), .B2(n10123), .A(n5784), .ZN(n8350) );
  NAND2_X1 U5315 ( .A1(n4810), .A2(n4809), .ZN(n4808) );
  INV_X1 U5316 ( .A(n7341), .ZN(n4810) );
  AOI21_X1 U5317 ( .B1(n6746), .B2(n6749), .A(n6745), .ZN(n4806) );
  OR2_X1 U5318 ( .A1(n4531), .A2(n4595), .ZN(n4797) );
  NOR2_X1 U5319 ( .A1(n8149), .A2(n4801), .ZN(n4800) );
  INV_X1 U5320 ( .A(n6786), .ZN(n4801) );
  OAI21_X1 U5321 ( .B1(n4645), .B2(n4644), .A(n4642), .ZN(n9157) );
  NAND2_X1 U5322 ( .A1(n9154), .A2(n9263), .ZN(n4644) );
  NOR2_X1 U5323 ( .A1(n5057), .A2(n4643), .ZN(n4642) );
  AOI21_X1 U5324 ( .B1(n9152), .B2(n9151), .A(n4646), .ZN(n4645) );
  OR2_X1 U5325 ( .A1(n4659), .A2(n4657), .ZN(n4656) );
  NOR2_X1 U5326 ( .A1(n4666), .A2(n4658), .ZN(n4657) );
  INV_X1 U5327 ( .A(n9270), .ZN(n4658) );
  AND2_X1 U5328 ( .A1(n4663), .A2(n4660), .ZN(n4659) );
  AND2_X1 U5329 ( .A1(n9162), .A2(n9277), .ZN(n4663) );
  NAND2_X1 U5330 ( .A1(n4664), .A2(n4661), .ZN(n4660) );
  INV_X1 U5331 ( .A(n9274), .ZN(n4661) );
  NAND2_X1 U5332 ( .A1(n9165), .A2(n9278), .ZN(n4662) );
  NOR2_X1 U5333 ( .A1(n8149), .A2(n5495), .ZN(n4799) );
  AND2_X1 U5334 ( .A1(n4797), .A2(n4798), .ZN(n4796) );
  OR2_X1 U5335 ( .A1(n4531), .A2(n6783), .ZN(n4798) );
  INV_X1 U5336 ( .A(n4797), .ZN(n4794) );
  AOI21_X1 U5337 ( .B1(n9188), .B2(n9187), .A(n4684), .ZN(n4683) );
  INV_X1 U5338 ( .A(n9661), .ZN(n4684) );
  AND2_X1 U5339 ( .A1(n4686), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U5340 ( .A1(n4683), .A2(n4681), .ZN(n4680) );
  INV_X1 U5341 ( .A(n9192), .ZN(n4686) );
  INV_X1 U5342 ( .A(n9187), .ZN(n4681) );
  INV_X1 U5343 ( .A(n4683), .ZN(n4682) );
  AND2_X1 U5344 ( .A1(n8396), .A2(n8457), .ZN(n8272) );
  INV_X1 U5345 ( .A(n4787), .ZN(n4786) );
  OR2_X1 U5346 ( .A1(n8291), .A2(n8290), .ZN(n8296) );
  XNOR2_X1 U5347 ( .A(n8856), .B(n7421), .ZN(n8324) );
  OR2_X1 U5348 ( .A1(n8838), .A2(n6855), .ZN(n6918) );
  NAND2_X1 U5349 ( .A1(n6888), .A2(n4701), .ZN(n4700) );
  NOR2_X1 U5350 ( .A1(n4702), .A2(n8630), .ZN(n4701) );
  INV_X1 U5351 ( .A(n5767), .ZN(n4702) );
  INV_X1 U5352 ( .A(n5089), .ZN(n6592) );
  NAND2_X1 U5353 ( .A1(n7718), .A2(n6702), .ZN(n4954) );
  AOI21_X1 U5354 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7148), .A(n8535), .ZN(
        n6602) );
  INV_X1 U5355 ( .A(n5117), .ZN(n5115) );
  AOI21_X1 U5356 ( .B1(n6791), .B2(n6790), .A(n5118), .ZN(n5117) );
  INV_X1 U5357 ( .A(n6728), .ZN(n5118) );
  OR2_X1 U5358 ( .A1(n8830), .A2(n8761), .ZN(n6799) );
  OR2_X1 U5359 ( .A1(n10176), .A2(n8024), .ZN(n8073) );
  INV_X1 U5360 ( .A(n4553), .ZN(n4882) );
  NAND2_X1 U5361 ( .A1(n10137), .A2(n8515), .ZN(n6732) );
  NAND2_X1 U5362 ( .A1(n7271), .A2(n7345), .ZN(n5739) );
  OR2_X1 U5363 ( .A1(n8860), .A2(n8653), .ZN(n6834) );
  NAND2_X1 U5364 ( .A1(n8809), .A2(n8717), .ZN(n6818) );
  OR2_X1 U5365 ( .A1(n8809), .A2(n8717), .ZN(n5760) );
  NOR2_X1 U5366 ( .A1(n8739), .A2(n4877), .ZN(n4876) );
  INV_X1 U5367 ( .A(n5601), .ZN(n4877) );
  NAND2_X1 U5368 ( .A1(n4858), .A2(n4857), .ZN(n8136) );
  AOI21_X1 U5369 ( .B1(n5162), .B2(n4559), .A(n4860), .ZN(n4858) );
  NOR2_X1 U5370 ( .A1(n8372), .A2(n5749), .ZN(n4860) );
  NAND2_X1 U5371 ( .A1(n4597), .A2(n4631), .ZN(n5518) );
  NAND2_X1 U5372 ( .A1(n4586), .A2(n5748), .ZN(n5137) );
  NOR2_X1 U5373 ( .A1(n8124), .A2(n5140), .ZN(n5139) );
  OR2_X1 U5374 ( .A1(n8989), .A2(n4621), .ZN(n4753) );
  OAI21_X1 U5375 ( .B1(n4753), .B2(n4754), .A(n4606), .ZN(n4749) );
  NOR2_X1 U5376 ( .A1(n4560), .A2(n4743), .ZN(n4742) );
  INV_X1 U5377 ( .A(n6109), .ZN(n4743) );
  INV_X1 U5378 ( .A(n8958), .ZN(n5077) );
  NOR2_X1 U5379 ( .A1(n5079), .A2(n4540), .ZN(n5078) );
  INV_X1 U5380 ( .A(n6006), .ZN(n4726) );
  NOR2_X1 U5381 ( .A1(n8307), .A2(n9867), .ZN(n4965) );
  NOR2_X1 U5382 ( .A1(n4971), .A2(n9636), .ZN(n4970) );
  INV_X1 U5383 ( .A(n4972), .ZN(n4971) );
  NOR2_X1 U5384 ( .A1(n7791), .A2(n7543), .ZN(n4975) );
  NAND2_X1 U5385 ( .A1(n4718), .A2(n4578), .ZN(n5303) );
  NAND2_X1 U5386 ( .A1(n5537), .A2(n4719), .ZN(n4718) );
  NAND2_X1 U5387 ( .A1(n4717), .A2(n4564), .ZN(n4716) );
  INV_X1 U5388 ( .A(n5217), .ZN(n5028) );
  INV_X1 U5389 ( .A(n5469), .ZN(n5220) );
  XNOR2_X1 U5390 ( .A(n5219), .B(n5218), .ZN(n5469) );
  NAND2_X1 U5391 ( .A1(n5214), .A2(n10408), .ZN(n5217) );
  NAND2_X1 U5392 ( .A1(n5202), .A2(n5201), .ZN(n5429) );
  INV_X1 U5393 ( .A(SI_7_), .ZN(n10365) );
  INV_X1 U5394 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U5395 ( .A1(n4931), .A2(n4929), .ZN(n8361) );
  AOI21_X1 U5396 ( .B1(n4932), .B2(n4934), .A(n4930), .ZN(n4929) );
  INV_X1 U5397 ( .A(n8362), .ZN(n4930) );
  AND2_X1 U5398 ( .A1(n8445), .A2(n8260), .ZN(n8383) );
  INV_X1 U5399 ( .A(n8516), .ZN(n7227) );
  AND2_X1 U5400 ( .A1(n8092), .A2(n8070), .ZN(n8071) );
  AND2_X1 U5401 ( .A1(n8290), .A2(n8287), .ZN(n8405) );
  NAND2_X1 U5402 ( .A1(n4910), .A2(n4908), .ZN(n8427) );
  AOI21_X1 U5403 ( .B1(n4911), .B2(n4912), .A(n4909), .ZN(n4908) );
  INV_X1 U5404 ( .A(n8425), .ZN(n4909) );
  AND2_X1 U5405 ( .A1(n8404), .A2(n8284), .ZN(n8435) );
  NAND2_X1 U5406 ( .A1(n4922), .A2(n4565), .ZN(n8062) );
  INV_X1 U5407 ( .A(n8034), .ZN(n4927) );
  NAND2_X1 U5408 ( .A1(n8229), .A2(n4939), .ZN(n4937) );
  AND2_X1 U5409 ( .A1(n8299), .A2(n8707), .ZN(n4915) );
  AND2_X1 U5410 ( .A1(n8435), .A2(n8295), .ZN(n8299) );
  NAND2_X1 U5411 ( .A1(n8279), .A2(n8278), .ZN(n8434) );
  NAND2_X1 U5412 ( .A1(n7115), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n8212) );
  INV_X1 U5413 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4942) );
  OAI21_X1 U5414 ( .B1(n6685), .B2(n6684), .A(n6686), .ZN(n8208) );
  NOR2_X1 U5415 ( .A1(n6683), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U5416 ( .A1(n4817), .A2(n4816), .ZN(n10103) );
  NAND2_X1 U5417 ( .A1(n10107), .A2(n7418), .ZN(n4816) );
  NAND2_X1 U5418 ( .A1(n7237), .A2(n4834), .ZN(n7140) );
  NAND2_X1 U5419 ( .A1(n4634), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7235) );
  INV_X1 U5420 ( .A(n7140), .ZN(n4634) );
  INV_X1 U5421 ( .A(n6694), .ZN(n4957) );
  NAND2_X1 U5422 ( .A1(n6693), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4956) );
  NAND2_X1 U5423 ( .A1(n6693), .A2(n4829), .ZN(n4827) );
  INV_X1 U5424 ( .A(n7368), .ZN(n4830) );
  INV_X1 U5425 ( .A(n7563), .ZN(n4633) );
  INV_X1 U5426 ( .A(n7727), .ZN(n4845) );
  NAND2_X1 U5427 ( .A1(n4847), .A2(n4551), .ZN(n4846) );
  OR2_X1 U5428 ( .A1(n7721), .A2(n7720), .ZN(n7718) );
  XNOR2_X1 U5429 ( .A(n4954), .B(n4953), .ZN(n7901) );
  INV_X1 U5430 ( .A(n7905), .ZN(n4953) );
  NAND2_X1 U5431 ( .A1(n7096), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5091) );
  AND2_X1 U5432 ( .A1(n4826), .A2(n4556), .ZN(n8545) );
  OR2_X1 U5433 ( .A1(n8552), .A2(n6710), .ZN(n4832) );
  XNOR2_X1 U5434 ( .A(n6602), .B(n6708), .ZN(n8560) );
  NOR2_X1 U5435 ( .A1(n6708), .A2(n6602), .ZN(n6603) );
  AND2_X1 U5436 ( .A1(n4952), .A2(n4951), .ZN(n6711) );
  NAND2_X1 U5437 ( .A1(n7265), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4951) );
  AOI21_X1 U5438 ( .B1(n4876), .B2(n5602), .A(n4879), .ZN(n4875) );
  AND2_X1 U5439 ( .A1(n8892), .A2(n8728), .ZN(n4879) );
  AND2_X1 U5440 ( .A1(n6805), .A2(n6804), .ZN(n8755) );
  INV_X1 U5441 ( .A(n6774), .ZN(n5140) );
  AOI21_X1 U5442 ( .B1(n4529), .B2(n6902), .A(n5133), .ZN(n5132) );
  OR2_X1 U5443 ( .A1(n7920), .A2(n6902), .ZN(n5134) );
  NAND2_X1 U5444 ( .A1(n5134), .A2(n4529), .ZN(n8049) );
  AND4_X1 U5445 ( .A1(n5453), .A2(n5452), .A3(n5451), .A4(n5450), .ZN(n8059)
         );
  AND4_X1 U5446 ( .A1(n5493), .A2(n5492), .A3(n5491), .A4(n5490), .ZN(n8127)
         );
  INV_X1 U5447 ( .A(n4885), .ZN(n4883) );
  NAND2_X1 U5448 ( .A1(n4865), .A2(n4864), .ZN(n4863) );
  NAND2_X1 U5449 ( .A1(n8516), .A2(n7191), .ZN(n6896) );
  INV_X1 U5450 ( .A(n5124), .ZN(n5123) );
  XNOR2_X1 U5451 ( .A(n8843), .B(n8646), .ZN(n8630) );
  NAND2_X1 U5452 ( .A1(n5764), .A2(n6834), .ZN(n8655) );
  AOI21_X1 U5453 ( .B1(n8651), .B2(n5671), .A(n5670), .ZN(n8643) );
  AND2_X1 U5454 ( .A1(n6836), .A2(n8645), .ZN(n5670) );
  NOR2_X1 U5455 ( .A1(n8872), .A2(n8677), .ZN(n4888) );
  NOR2_X1 U5456 ( .A1(n5762), .A2(n5141), .ZN(n5147) );
  INV_X1 U5457 ( .A(n5148), .ZN(n5141) );
  OR2_X1 U5458 ( .A1(n5762), .A2(n5763), .ZN(n5146) );
  OR2_X1 U5459 ( .A1(n6822), .A2(n6825), .ZN(n8674) );
  OR2_X1 U5460 ( .A1(n8719), .A2(n8708), .ZN(n8701) );
  NAND2_X1 U5461 ( .A1(n5297), .A2(n5296), .ZN(n8444) );
  NAND2_X1 U5462 ( .A1(n4878), .A2(n5601), .ZN(n8740) );
  AND2_X1 U5463 ( .A1(n4878), .A2(n4876), .ZN(n8743) );
  INV_X1 U5464 ( .A(n5162), .ZN(n4862) );
  INV_X1 U5465 ( .A(n8760), .ZN(n10120) );
  AND2_X1 U5466 ( .A1(n5774), .A2(n6952), .ZN(n10118) );
  NAND2_X1 U5467 ( .A1(n8051), .A2(n5139), .ZN(n8122) );
  NOR2_X1 U5468 ( .A1(n5150), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4814) );
  NAND2_X1 U5469 ( .A1(n5152), .A2(n5151), .ZN(n5150) );
  AND2_X1 U5470 ( .A1(n5270), .A2(n5273), .ZN(n5152) );
  INV_X1 U5471 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5790) );
  INV_X1 U5472 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5792) );
  AND2_X1 U5473 ( .A1(n5727), .A2(n5726), .ZN(n5730) );
  XNOR2_X1 U5474 ( .A(n5394), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U5475 ( .A1(n5127), .A2(n5259), .ZN(n5378) );
  INV_X1 U5476 ( .A(n5360), .ZN(n5127) );
  OR2_X1 U5477 ( .A1(n6932), .A2(n6931), .ZN(n5085) );
  NOR2_X1 U5478 ( .A1(n8931), .A2(n4755), .ZN(n4754) );
  INV_X1 U5479 ( .A(n4753), .ZN(n4751) );
  NAND2_X1 U5480 ( .A1(n5068), .A2(n4554), .ZN(n8921) );
  NAND2_X1 U5481 ( .A1(n8999), .A2(n5073), .ZN(n5068) );
  INV_X1 U5482 ( .A(n5065), .ZN(n8983) );
  NAND2_X1 U5483 ( .A1(n4530), .A2(n4606), .ZN(n5067) );
  NOR2_X1 U5484 ( .A1(n5069), .A2(n4536), .ZN(n5066) );
  NOR2_X1 U5485 ( .A1(n9023), .A2(n6405), .ZN(n6930) );
  NAND2_X1 U5486 ( .A1(n4667), .A2(n4669), .ZN(n9332) );
  AND2_X1 U5487 ( .A1(n4601), .A2(n4670), .ZN(n4669) );
  NAND2_X1 U5488 ( .A1(n4770), .A2(n4769), .ZN(n4768) );
  NAND2_X1 U5489 ( .A1(n9408), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4769) );
  NOR2_X1 U5490 ( .A1(n7321), .A2(n4622), .ZN(n4772) );
  NOR2_X1 U5491 ( .A1(n9056), .A2(n4547), .ZN(n4962) );
  INV_X1 U5492 ( .A(n5054), .ZN(n5053) );
  AOI21_X1 U5493 ( .B1(n5054), .B2(n5052), .A(n5051), .ZN(n5050) );
  AND2_X1 U5494 ( .A1(n9205), .A2(n9576), .ZN(n5054) );
  NAND2_X1 U5495 ( .A1(n5055), .A2(n9205), .ZN(n9570) );
  OR2_X1 U5496 ( .A1(n9871), .A2(n9783), .ZN(n4990) );
  AND4_X1 U5497 ( .A1(n6435), .A2(n6434), .A3(n6433), .A4(n6432), .ZN(n9597)
         );
  INV_X1 U5498 ( .A(n5046), .ZN(n5045) );
  AOI21_X1 U5499 ( .B1(n5046), .B2(n5044), .A(n5043), .ZN(n5042) );
  INV_X1 U5500 ( .A(n9227), .ZN(n5043) );
  NAND2_X1 U5501 ( .A1(n4986), .A2(n4983), .ZN(n9662) );
  INV_X1 U5502 ( .A(n4984), .ZN(n4983) );
  OAI22_X1 U5503 ( .A1(n6523), .A2(n4985), .B1(n9184), .B2(n9896), .ZN(n4984)
         );
  AND2_X1 U5504 ( .A1(n9677), .A2(n9185), .ZN(n5049) );
  AND2_X1 U5505 ( .A1(n9185), .A2(n9183), .ZN(n9695) );
  INV_X1 U5506 ( .A(n4994), .ZN(n4993) );
  AOI21_X1 U5507 ( .B1(n4994), .B2(n4992), .A(n4573), .ZN(n4991) );
  AND2_X1 U5508 ( .A1(n4995), .A2(n6517), .ZN(n4994) );
  AND2_X1 U5509 ( .A1(n9277), .A2(n9280), .ZN(n9085) );
  NAND2_X1 U5510 ( .A1(n7778), .A2(n5063), .ZN(n7838) );
  AND2_X1 U5511 ( .A1(n4552), .A2(n9163), .ZN(n5063) );
  AND2_X1 U5512 ( .A1(n9081), .A2(n9154), .ZN(n5058) );
  NAND2_X1 U5513 ( .A1(n5060), .A2(n5059), .ZN(n7524) );
  INV_X1 U5514 ( .A(n7523), .ZN(n5060) );
  NAND2_X1 U5515 ( .A1(n9062), .A2(n9061), .ZN(n9564) );
  XNOR2_X1 U5516 ( .A(n6871), .B(n6870), .ZN(n9053) );
  OAI22_X1 U5517 ( .A1(n6867), .A2(n6866), .B1(SI_30_), .B2(n6865), .ZN(n6871)
         );
  XNOR2_X1 U5518 ( .A(n6867), .B(n6866), .ZN(n9059) );
  XNOR2_X1 U5519 ( .A(n5660), .B(n5672), .ZN(n8038) );
  NAND2_X1 U5520 ( .A1(n5656), .A2(n5676), .ZN(n5660) );
  NAND2_X1 U5521 ( .A1(n5675), .A2(n5673), .ZN(n5656) );
  INV_X1 U5522 ( .A(n5880), .ZN(n4727) );
  XNOR2_X1 U5523 ( .A(n5675), .B(n5673), .ZN(n7961) );
  XNOR2_X1 U5524 ( .A(n5628), .B(n5627), .ZN(n7930) );
  NAND2_X1 U5525 ( .A1(n4710), .A2(n4709), .ZN(n5614) );
  AOI21_X1 U5526 ( .B1(n4711), .B2(n4715), .A(n4616), .ZN(n4709) );
  NAND2_X1 U5527 ( .A1(n4996), .A2(n4711), .ZN(n4710) );
  NAND2_X1 U5528 ( .A1(n4712), .A2(n4713), .ZN(n5605) );
  OR2_X1 U5529 ( .A1(n4996), .A2(n4715), .ZN(n4712) );
  NAND2_X1 U5530 ( .A1(n5845), .A2(n5844), .ZN(n6286) );
  NAND2_X1 U5531 ( .A1(n5231), .A2(n5230), .ZN(n5570) );
  NAND2_X1 U5532 ( .A1(n4723), .A2(n5227), .ZN(n5553) );
  OAI21_X1 U5533 ( .B1(n5212), .B2(n4708), .A(n4705), .ZN(n5523) );
  INV_X1 U5534 ( .A(n4694), .ZN(n4693) );
  XNOR2_X1 U5535 ( .A(n5188), .B(n5187), .ZN(n5376) );
  AND3_X1 U5536 ( .A1(n5301), .A2(n5300), .A3(n5299), .ZN(n8745) );
  AND2_X1 U5537 ( .A1(n5638), .A2(n5637), .ZN(n8692) );
  OR2_X1 U5538 ( .A1(n5328), .A2(n8221), .ZN(n5350) );
  AND4_X1 U5539 ( .A1(n5390), .A2(n5389), .A3(n5388), .A4(n5387), .ZN(n7693)
         );
  NAND2_X1 U5540 ( .A1(n4689), .A2(n4534), .ZN(n4688) );
  NAND2_X1 U5541 ( .A1(n6924), .A2(n6923), .ZN(n4689) );
  NAND4_X1 U5542 ( .A1(n5440), .A2(n5439), .A3(n5438), .A4(n5437), .ZN(n8511)
         );
  OR2_X1 U5543 ( .A1(n5343), .A2(n5436), .ZN(n5437) );
  NAND4_X1 U5544 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n8512)
         );
  INV_X1 U5545 ( .A(n7693), .ZN(n10119) );
  NAND4_X1 U5546 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .ZN(n8513)
         );
  INV_X1 U5547 ( .A(n6706), .ZN(n4946) );
  NOR2_X1 U5548 ( .A1(n8553), .A2(n6614), .ZN(n8552) );
  NOR2_X1 U5549 ( .A1(n8586), .A2(n8778), .ZN(n8585) );
  NAND2_X1 U5550 ( .A1(n8594), .A2(n10095), .ZN(n5105) );
  OAI21_X1 U5551 ( .B1(n8593), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8592), .ZN(
        n5106) );
  INV_X1 U5552 ( .A(n4819), .ZN(n8614) );
  OR2_X1 U5553 ( .A1(n8619), .A2(n8618), .ZN(n4958) );
  NOR2_X1 U5554 ( .A1(n8591), .A2(n6606), .ZN(n8602) );
  NOR2_X1 U5555 ( .A1(n8600), .A2(n6608), .ZN(n6609) );
  NAND2_X1 U5556 ( .A1(n5593), .A2(n5592), .ZN(n8767) );
  NAND2_X1 U5557 ( .A1(n5111), .A2(n6744), .ZN(n7812) );
  INV_X1 U5558 ( .A(n10133), .ZN(n8776) );
  INV_X1 U5559 ( .A(n8860), .ZN(n8798) );
  NAND2_X1 U5560 ( .A1(n5786), .A2(n10181), .ZN(n5787) );
  NAND2_X1 U5561 ( .A1(n5686), .A2(n5685), .ZN(n8849) );
  NAND2_X1 U5562 ( .A1(n8220), .A2(n6875), .ZN(n5686) );
  XNOR2_X1 U5563 ( .A(n4901), .B(n5308), .ZN(n7547) );
  NAND2_X1 U5564 ( .A1(n5589), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U5565 ( .A1(n5304), .A2(n5305), .ZN(n5571) );
  NAND2_X1 U5566 ( .A1(n6266), .A2(n9012), .ZN(n4761) );
  NOR2_X1 U5567 ( .A1(n6930), .A2(n5085), .ZN(n6935) );
  AND2_X1 U5568 ( .A1(n6468), .A2(n9025), .ZN(n6467) );
  AOI21_X1 U5569 ( .B1(n9023), .B2(n5084), .A(n5082), .ZN(n5081) );
  INV_X1 U5570 ( .A(n5085), .ZN(n5084) );
  OAI21_X1 U5571 ( .B1(n5085), .B2(n5083), .A(n4609), .ZN(n5082) );
  INV_X1 U5572 ( .A(n6405), .ZN(n5083) );
  OR2_X1 U5573 ( .A1(n4649), .A2(n7028), .ZN(n4648) );
  NOR2_X1 U5574 ( .A1(n8950), .A2(n8949), .ZN(n9023) );
  NAND2_X1 U5575 ( .A1(n6210), .A2(n6209), .ZN(n9927) );
  NOR2_X1 U5576 ( .A1(n7042), .A2(n4767), .ZN(n7047) );
  AND2_X1 U5577 ( .A1(n7043), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4767) );
  NAND2_X1 U5578 ( .A1(n6346), .A2(n6345), .ZN(n9656) );
  NAND2_X1 U5579 ( .A1(n6568), .A2(n5168), .ZN(n6725) );
  AND2_X1 U5580 ( .A1(n8307), .A2(n9879), .ZN(n6727) );
  OAI21_X1 U5581 ( .B1(n6848), .B2(n5015), .A(n5013), .ZN(n8319) );
  AOI22_X1 U5582 ( .A1(n5016), .A2(SI_29_), .B1(n6847), .B2(n5717), .ZN(n5015)
         );
  OAI22_X1 U5583 ( .A1(n5016), .A2(n5717), .B1(n6847), .B2(SI_29_), .ZN(n5014)
         );
  INV_X1 U5584 ( .A(n4813), .ZN(n4812) );
  OAI22_X1 U5585 ( .A1(n5739), .A2(n6948), .B1(n6732), .B2(n6952), .ZN(n4813)
         );
  NAND2_X1 U5586 ( .A1(n4811), .A2(n4568), .ZN(n4807) );
  NAND2_X1 U5587 ( .A1(n6731), .A2(n6730), .ZN(n4811) );
  INV_X1 U5588 ( .A(n9153), .ZN(n4646) );
  INV_X1 U5589 ( .A(n9155), .ZN(n4643) );
  NAND2_X1 U5590 ( .A1(n9280), .A2(n9207), .ZN(n4666) );
  AND2_X1 U5591 ( .A1(n4656), .A2(n4662), .ZN(n4651) );
  NAND2_X1 U5592 ( .A1(n4653), .A2(n4662), .ZN(n4652) );
  INV_X1 U5593 ( .A(n4654), .ZN(n4653) );
  AOI21_X1 U5594 ( .B1(n4659), .B2(n4665), .A(n4655), .ZN(n4654) );
  NOR2_X1 U5595 ( .A1(n4666), .A2(n4561), .ZN(n4655) );
  NAND2_X1 U5596 ( .A1(n4794), .A2(n4577), .ZN(n4793) );
  NAND2_X1 U5597 ( .A1(n4783), .A2(n4537), .ZN(n4790) );
  NAND2_X1 U5598 ( .A1(n4685), .A2(n9193), .ZN(n9198) );
  AOI21_X1 U5599 ( .B1(n4679), .B2(n4682), .A(n4591), .ZN(n4678) );
  AND2_X1 U5600 ( .A1(n8267), .A2(n4563), .ZN(n8268) );
  OR2_X1 U5601 ( .A1(n8265), .A2(n8394), .ZN(n8267) );
  INV_X1 U5602 ( .A(n6838), .ZN(n5125) );
  AND2_X1 U5603 ( .A1(n5521), .A2(n4559), .ZN(n4859) );
  AND2_X1 U5604 ( .A1(n7654), .A2(n7611), .ZN(n4980) );
  INV_X1 U5605 ( .A(n6503), .ZN(n4981) );
  INV_X1 U5606 ( .A(n5039), .ZN(n4717) );
  INV_X1 U5607 ( .A(n5038), .ZN(n5037) );
  OAI21_X1 U5608 ( .B1(n5040), .B2(n5039), .A(n5239), .ZN(n5038) );
  NOR2_X1 U5609 ( .A1(n4567), .A2(n4722), .ZN(n4721) );
  INV_X1 U5610 ( .A(n5227), .ZN(n4722) );
  INV_X1 U5611 ( .A(n5535), .ZN(n5226) );
  INV_X1 U5612 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10440) );
  AOI21_X1 U5613 ( .B1(n4935), .B2(n4933), .A(n8363), .ZN(n4932) );
  INV_X1 U5614 ( .A(n4939), .ZN(n4933) );
  INV_X1 U5615 ( .A(n4935), .ZN(n4934) );
  AOI21_X1 U5616 ( .B1(n8250), .B2(n8483), .A(n8426), .ZN(n4911) );
  INV_X1 U5617 ( .A(n8250), .ZN(n4912) );
  OR2_X1 U5618 ( .A1(n8228), .A2(n8507), .ZN(n4939) );
  INV_X1 U5619 ( .A(n7551), .ZN(n4921) );
  NAND2_X1 U5620 ( .A1(n4783), .A2(n4785), .ZN(n6860) );
  NAND2_X1 U5621 ( .A1(n4837), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4836) );
  NAND2_X1 U5622 ( .A1(n10101), .A2(n6687), .ZN(n6688) );
  NOR2_X1 U5623 ( .A1(n7368), .A2(n7670), .ZN(n4829) );
  OR2_X1 U5624 ( .A1(n7364), .A2(n6591), .ZN(n5089) );
  INV_X1 U5625 ( .A(n8115), .ZN(n4948) );
  INV_X1 U5626 ( .A(n8048), .ZN(n5133) );
  NAND2_X1 U5627 ( .A1(n4585), .A2(n4869), .ZN(n4864) );
  NAND2_X1 U5628 ( .A1(n4871), .A2(n5398), .ZN(n4865) );
  NAND2_X1 U5629 ( .A1(n7333), .A2(n4867), .ZN(n4866) );
  INV_X1 U5630 ( .A(n5368), .ZN(n4868) );
  OAI21_X1 U5631 ( .B1(n6897), .B2(n7341), .A(n5739), .ZN(n7410) );
  NAND2_X1 U5632 ( .A1(n7410), .A2(n7411), .ZN(n7409) );
  OAI21_X1 U5633 ( .B1(n5803), .B2(P2_D_REG_0__SCAN_IN), .A(n6992), .ZN(n7215)
         );
  NOR2_X1 U5634 ( .A1(n5125), .A2(n5121), .ZN(n5120) );
  INV_X1 U5635 ( .A(n6834), .ZN(n5121) );
  OAI21_X1 U5636 ( .B1(n8656), .B2(n5125), .A(n8644), .ZN(n5124) );
  NOR2_X1 U5637 ( .A1(n5754), .A2(n5149), .ZN(n5148) );
  INV_X1 U5638 ( .A(n6805), .ZN(n5149) );
  OR2_X1 U5639 ( .A1(n6949), .A2(n5824), .ZN(n7303) );
  INV_X1 U5640 ( .A(n5269), .ZN(n5151) );
  INV_X1 U5641 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U5642 ( .A1(n5304), .A2(n4917), .ZN(n5307) );
  NOR2_X1 U5643 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4917) );
  INV_X1 U5644 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U5645 ( .A1(n8998), .A2(n9003), .ZN(n5072) );
  OR2_X1 U5646 ( .A1(n8998), .A2(n9003), .ZN(n5073) );
  OAI21_X1 U5647 ( .B1(n4554), .B2(n5071), .A(n5070), .ZN(n5069) );
  INV_X1 U5648 ( .A(n8981), .ZN(n5070) );
  INV_X1 U5649 ( .A(n8982), .ZN(n5071) );
  NAND2_X1 U5650 ( .A1(n7353), .A2(n6070), .ZN(n6088) );
  NOR2_X1 U5651 ( .A1(n6095), .A2(n7714), .ZN(n6115) );
  AND2_X1 U5652 ( .A1(n6440), .A2(n9748), .ZN(n5941) );
  AND2_X1 U5653 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6013) );
  NAND2_X1 U5654 ( .A1(n9218), .A2(n4674), .ZN(n4673) );
  INV_X1 U5655 ( .A(n9211), .ZN(n4674) );
  NOR2_X1 U5656 ( .A1(n9217), .A2(n9296), .ZN(n4676) );
  NOR2_X1 U5657 ( .A1(n4672), .A2(n5051), .ZN(n4668) );
  OR2_X1 U5658 ( .A1(n4675), .A2(n9212), .ZN(n4672) );
  OR2_X1 U5659 ( .A1(n4675), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U5660 ( .A1(n9096), .A2(n4608), .ZN(n4671) );
  AND2_X1 U5661 ( .A1(n9479), .A2(n4764), .ZN(n9495) );
  NAND2_X1 U5662 ( .A1(n9480), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4764) );
  INV_X1 U5663 ( .A(n9646), .ZN(n5044) );
  OR2_X1 U5664 ( .A1(n9878), .A2(n9030), .ZN(n9245) );
  AND2_X1 U5665 ( .A1(n5047), .A2(n9224), .ZN(n5046) );
  NOR2_X1 U5666 ( .A1(n9656), .A2(n9670), .ZN(n4972) );
  NAND2_X1 U5667 ( .A1(n4557), .A2(n6522), .ZN(n4985) );
  NOR2_X1 U5668 ( .A1(n6523), .A2(n4988), .ZN(n4987) );
  INV_X1 U5669 ( .A(n6522), .ZN(n4988) );
  NAND2_X1 U5670 ( .A1(n4967), .A2(n4966), .ZN(n9683) );
  NAND2_X1 U5671 ( .A1(n9085), .A2(n6516), .ZN(n4995) );
  INV_X1 U5672 ( .A(n6516), .ZN(n4992) );
  AND2_X1 U5673 ( .A1(n6115), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6135) );
  OR2_X1 U5674 ( .A1(n7442), .A2(n7866), .ZN(n9151) );
  NOR2_X1 U5675 ( .A1(n6032), .A2(n6031), .ZN(n6056) );
  NAND2_X1 U5676 ( .A1(n9684), .A2(n9892), .ZN(n9667) );
  NAND2_X1 U5677 ( .A1(n9740), .A2(n9905), .ZN(n9739) );
  NAND2_X1 U5678 ( .A1(n6286), .A2(n9335), .ZN(n6542) );
  NAND2_X1 U5679 ( .A1(n4997), .A2(n5698), .ZN(n5714) );
  NAND2_X1 U5680 ( .A1(n5697), .A2(n5696), .ZN(n4997) );
  AND2_X1 U5681 ( .A1(n5887), .A2(n5881), .ZN(n5888) );
  NAND2_X1 U5682 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n4731) );
  INV_X2 U5683 ( .A(n5176), .ZN(n5186) );
  AOI21_X1 U5684 ( .B1(n4618), .B2(n5246), .A(n4714), .ZN(n4713) );
  NOR2_X1 U5685 ( .A1(n5245), .A2(SI_20_), .ZN(n4714) );
  NOR2_X1 U5686 ( .A1(n5246), .A2(n10599), .ZN(n4715) );
  NOR2_X1 U5687 ( .A1(n5569), .A2(n5041), .ZN(n5040) );
  INV_X1 U5688 ( .A(n5230), .ZN(n5041) );
  NAND2_X1 U5689 ( .A1(n4723), .A2(n4721), .ZN(n5231) );
  OR2_X1 U5690 ( .A1(n5537), .A2(n5228), .ZN(n4723) );
  AOI21_X1 U5691 ( .B1(n5480), .B2(n5027), .A(n4583), .ZN(n5025) );
  NOR2_X1 U5692 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5834) );
  NAND2_X1 U5693 ( .A1(n5205), .A2(n10618), .ZN(n5501) );
  XNOR2_X1 U5694 ( .A(n5210), .B(n5208), .ZN(n5503) );
  INV_X1 U5695 ( .A(n5202), .ZN(n5007) );
  INV_X1 U5696 ( .A(n5425), .ZN(n5008) );
  INV_X1 U5697 ( .A(n5010), .ZN(n5009) );
  INV_X1 U5698 ( .A(SI_6_), .ZN(n10454) );
  NAND2_X1 U5699 ( .A1(n5018), .A2(SI_3_), .ZN(n5182) );
  OAI21_X1 U5700 ( .B1(n5186), .B2(n5020), .A(n5019), .ZN(n5018) );
  NAND2_X1 U5701 ( .A1(n5186), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5019) );
  INV_X1 U5702 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4687) );
  XNOR2_X1 U5703 ( .A(n5274), .B(n5273), .ZN(n5773) );
  NAND2_X1 U5704 ( .A1(n5272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U5705 ( .A1(n4904), .A2(n8383), .ZN(n8391) );
  NAND2_X1 U5706 ( .A1(n8381), .A2(n8382), .ZN(n4904) );
  AND2_X1 U5707 ( .A1(n8415), .A2(n8416), .ZN(n8250) );
  INV_X1 U5708 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U5709 ( .A1(n4921), .A2(n7549), .ZN(n4920) );
  AND2_X1 U5710 ( .A1(n8468), .A2(n8253), .ZN(n8425) );
  NAND2_X1 U5711 ( .A1(n7498), .A2(n7497), .ZN(n7552) );
  AOI21_X1 U5712 ( .B1(n4925), .B2(n4928), .A(n4541), .ZN(n4924) );
  NAND2_X1 U5713 ( .A1(n4923), .A2(n4925), .ZN(n4922) );
  INV_X1 U5714 ( .A(n7802), .ZN(n4923) );
  NOR2_X1 U5715 ( .A1(n8231), .A2(n4936), .ZN(n4935) );
  INV_X1 U5716 ( .A(n4938), .ZN(n4936) );
  NAND2_X1 U5717 ( .A1(n8228), .A2(n8507), .ZN(n4938) );
  AOI21_X1 U5718 ( .B1(n4905), .B2(n4907), .A(n4579), .ZN(n4903) );
  INV_X1 U5719 ( .A(n8383), .ZN(n4907) );
  OR2_X1 U5720 ( .A1(n5511), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U5721 ( .A1(n5575), .A2(n10452), .ZN(n5594) );
  INV_X1 U5722 ( .A(n10121), .ZN(n7830) );
  AOI21_X1 U5723 ( .B1(n6863), .B2(n8834), .A(n4809), .ZN(n6891) );
  AOI21_X1 U5724 ( .B1(n4698), .B2(n4548), .A(n4589), .ZN(n6890) );
  AND2_X1 U5725 ( .A1(n6884), .A2(n5724), .ZN(n8499) );
  NAND2_X1 U5726 ( .A1(n6876), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U5727 ( .A1(n4940), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U5728 ( .A1(n8206), .A2(n6686), .ZN(n10102) );
  NAND2_X1 U5729 ( .A1(n4849), .A2(n4848), .ZN(n7287) );
  NAND2_X1 U5730 ( .A1(n6587), .A2(n6971), .ZN(n4848) );
  NOR2_X1 U5731 ( .A1(n7286), .A2(n6588), .ZN(n7366) );
  XNOR2_X1 U5732 ( .A(n5089), .B(n6983), .ZN(n7563) );
  OR2_X1 U5733 ( .A1(n4562), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5442) );
  OR2_X1 U5734 ( .A1(n4845), .A2(n4843), .ZN(n4842) );
  INV_X1 U5735 ( .A(n6595), .ZN(n4843) );
  INV_X1 U5736 ( .A(n4954), .ZN(n6703) );
  NAND2_X1 U5737 ( .A1(n4544), .A2(n7964), .ZN(n5100) );
  NAND2_X1 U5738 ( .A1(n5101), .A2(n4544), .ZN(n5099) );
  INV_X1 U5739 ( .A(n8536), .ZN(n4841) );
  XNOR2_X1 U5740 ( .A(n5090), .B(n4825), .ZN(n8520) );
  OAI21_X1 U5741 ( .B1(n8590), .B2(n4851), .A(n4850), .ZN(n8600) );
  NAND2_X1 U5742 ( .A1(n4852), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4851) );
  AND3_X1 U5743 ( .A1(n5612), .A2(n5611), .A3(n5610), .ZN(n8708) );
  NAND2_X1 U5744 ( .A1(n4874), .A2(n4533), .ZN(n8727) );
  AOI21_X1 U5745 ( .B1(n5117), .B2(n5114), .A(n6793), .ZN(n5113) );
  INV_X1 U5746 ( .A(n6791), .ZN(n5114) );
  NAND2_X1 U5747 ( .A1(n6799), .A2(n6803), .ZN(n8781) );
  AND2_X1 U5748 ( .A1(n5559), .A2(n5558), .ZN(n5575) );
  OR2_X1 U5749 ( .A1(n5529), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5544) );
  NOR2_X1 U5750 ( .A1(n5489), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5475) );
  OR2_X1 U5751 ( .A1(n5513), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U5752 ( .A1(n5448), .A2(n5447), .ZN(n5511) );
  INV_X1 U5753 ( .A(n8509), .ZN(n8024) );
  AND2_X1 U5754 ( .A1(n5434), .A2(n10566), .ZN(n5448) );
  INV_X1 U5755 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10566) );
  INV_X1 U5756 ( .A(n4881), .ZN(n4880) );
  AOI21_X1 U5757 ( .B1(n4884), .B2(n4882), .A(n4590), .ZN(n4881) );
  NAND2_X1 U5758 ( .A1(n10127), .A2(n6749), .ZN(n5111) );
  NOR2_X1 U5759 ( .A1(n5416), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5434) );
  OR2_X1 U5760 ( .A1(n5402), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U5761 ( .A1(n7478), .A2(n6742), .ZN(n10127) );
  INV_X1 U5762 ( .A(n4870), .ZN(n7665) );
  AOI21_X1 U5763 ( .B1(n4873), .B2(n4626), .A(n4871), .ZN(n4870) );
  NAND2_X1 U5764 ( .A1(n7333), .A2(n5368), .ZN(n4873) );
  AND2_X1 U5765 ( .A1(n6747), .A2(n6741), .ZN(n7332) );
  INV_X1 U5766 ( .A(n6898), .ZN(n7411) );
  NAND2_X1 U5767 ( .A1(n7227), .A2(n7308), .ZN(n7341) );
  NAND2_X1 U5768 ( .A1(n8646), .A2(n10120), .ZN(n4895) );
  OAI211_X1 U5769 ( .C1(n8753), .C2(n5144), .A(n5143), .B(n6826), .ZN(n8668)
         );
  NAND2_X1 U5770 ( .A1(n5146), .A2(n6824), .ZN(n5144) );
  INV_X1 U5771 ( .A(n5147), .ZN(n5142) );
  NAND2_X1 U5772 ( .A1(n6834), .A2(n6833), .ZN(n8667) );
  NAND2_X1 U5773 ( .A1(n5758), .A2(n4696), .ZN(n8686) );
  NAND2_X1 U5774 ( .A1(n5759), .A2(n4697), .ZN(n4696) );
  AND2_X1 U5775 ( .A1(n8697), .A2(n5758), .ZN(n8685) );
  NAND2_X1 U5776 ( .A1(n8753), .A2(n5148), .ZN(n8698) );
  AND2_X1 U5777 ( .A1(n5760), .A2(n6818), .ZN(n8705) );
  AND2_X1 U5778 ( .A1(n5624), .A2(n5623), .ZN(n8717) );
  NAND2_X1 U5779 ( .A1(n8133), .A2(n8134), .ZN(n8166) );
  INV_X1 U5780 ( .A(n5136), .ZN(n5135) );
  OAI21_X1 U5781 ( .B1(n5139), .B2(n5137), .A(n5160), .ZN(n5136) );
  INV_X1 U5782 ( .A(n7345), .ZN(n10137) );
  NAND2_X1 U5783 ( .A1(n4815), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U5784 ( .A1(n5587), .A2(n5586), .ZN(n5589) );
  INV_X1 U5785 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U5786 ( .A1(n5345), .A2(n5346), .ZN(n5360) );
  NAND2_X1 U5787 ( .A1(n7998), .A2(n4575), .ZN(n8911) );
  NAND2_X1 U5788 ( .A1(n4745), .A2(n6126), .ZN(n6127) );
  XNOR2_X1 U5789 ( .A(n6088), .B(n6086), .ZN(n7591) );
  INV_X1 U5790 ( .A(n9775), .ZN(n9195) );
  OR2_X1 U5791 ( .A1(n6235), .A2(n6234), .ZN(n8971) );
  AND2_X1 U5792 ( .A1(n8982), .A2(n8981), .ZN(n4737) );
  OR2_X1 U5793 ( .A1(n7579), .A2(n6400), .ZN(n5982) );
  OR2_X1 U5794 ( .A1(n6076), .A2(n6075), .ZN(n6095) );
  OR2_X1 U5795 ( .A1(n6175), .A2(n8002), .ZN(n6195) );
  NAND2_X1 U5796 ( .A1(n4750), .A2(n4748), .ZN(n4760) );
  INV_X1 U5797 ( .A(n4749), .ZN(n4748) );
  NAND2_X1 U5798 ( .A1(n8999), .A2(n8998), .ZN(n9002) );
  NAND2_X1 U5799 ( .A1(n4744), .A2(n4740), .ZN(n7880) );
  INV_X1 U5800 ( .A(n4745), .ZN(n4744) );
  INV_X1 U5801 ( .A(n4739), .ZN(n4738) );
  OAI21_X1 U5802 ( .B1(n4528), .B2(n4742), .A(n7881), .ZN(n4739) );
  INV_X1 U5803 ( .A(n6265), .ZN(n5076) );
  NOR2_X1 U5804 ( .A1(n8971), .A2(n6275), .ZN(n6276) );
  OAI21_X1 U5805 ( .B1(n6002), .B2(n4726), .A(n6025), .ZN(n4725) );
  NOR2_X1 U5806 ( .A1(n6003), .A2(n4726), .ZN(n4724) );
  INV_X1 U5807 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6031) );
  NOR2_X1 U5808 ( .A1(n7201), .A2(n4766), .ZN(n9414) );
  AND2_X1 U5809 ( .A1(n7202), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U5810 ( .A1(n9414), .A2(n9415), .ZN(n9413) );
  NOR2_X1 U5811 ( .A1(n6110), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6131) );
  NOR2_X1 U5812 ( .A1(n9431), .A2(n4623), .ZN(n7325) );
  NAND2_X1 U5813 ( .A1(n6986), .A2(n4649), .ZN(n7022) );
  NAND2_X1 U5814 ( .A1(n6533), .A2(n9569), .ZN(n9579) );
  INV_X1 U5815 ( .A(n9577), .ZN(n6533) );
  AND2_X1 U5816 ( .A1(n6477), .A2(n6431), .ZN(n9582) );
  NAND2_X1 U5817 ( .A1(n9645), .A2(n9646), .ZN(n5048) );
  NAND2_X1 U5818 ( .A1(n5048), .A2(n5046), .ZN(n9633) );
  NAND2_X1 U5819 ( .A1(n9684), .A2(n4972), .ZN(n9652) );
  AND2_X1 U5820 ( .A1(n4539), .A2(n10069), .ZN(n4973) );
  NAND2_X1 U5821 ( .A1(n7530), .A2(n4975), .ZN(n7767) );
  NAND2_X1 U5822 ( .A1(n5059), .A2(n9269), .ZN(n5056) );
  NAND2_X1 U5823 ( .A1(n7530), .A2(n7891), .ZN(n7682) );
  AND2_X1 U5824 ( .A1(n7468), .A2(n7472), .ZN(n7530) );
  NOR2_X1 U5825 ( .A1(n7436), .A2(n7442), .ZN(n7468) );
  AND2_X1 U5826 ( .A1(n9151), .A2(n9148), .ZN(n9077) );
  NAND2_X1 U5827 ( .A1(n4969), .A2(n4968), .ZN(n7436) );
  INV_X1 U5828 ( .A(n9984), .ZN(n4969) );
  NAND2_X1 U5829 ( .A1(n9985), .A2(n10049), .ZN(n9984) );
  NOR2_X1 U5830 ( .A1(n7657), .A2(n10041), .ZN(n9985) );
  OR2_X1 U5831 ( .A1(n7604), .A2(n10031), .ZN(n7657) );
  OR2_X1 U5832 ( .A1(n7627), .A2(n7583), .ZN(n7604) );
  NAND2_X1 U5833 ( .A1(n7742), .A2(n10019), .ZN(n7627) );
  AND2_X1 U5834 ( .A1(n7744), .A2(n10012), .ZN(n7742) );
  AND2_X1 U5835 ( .A1(n6546), .A2(n6545), .ZN(n7737) );
  NOR2_X1 U5836 ( .A1(n5919), .A2(n9748), .ZN(n7744) );
  NAND2_X1 U5837 ( .A1(n4514), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U5838 ( .A1(n5716), .A2(n5715), .ZN(n6848) );
  NAND2_X1 U5839 ( .A1(n5714), .A2(n5713), .ZN(n5716) );
  XNOR2_X1 U5840 ( .A(n5714), .B(n5713), .ZN(n8101) );
  NAND2_X1 U5841 ( .A1(n5879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U5842 ( .A1(n4996), .A2(n5245), .ZN(n5295) );
  OAI21_X1 U5843 ( .B1(n5481), .B2(n5480), .A(n5217), .ZN(n5470) );
  NAND2_X1 U5844 ( .A1(n5012), .A2(n5197), .ZN(n5430) );
  NAND2_X1 U5845 ( .A1(n5426), .A2(n5425), .ZN(n5012) );
  NAND2_X1 U5846 ( .A1(n5193), .A2(SI_5_), .ZN(n5194) );
  INV_X1 U5847 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5833) );
  NOR2_X1 U5848 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5064) );
  XNOR2_X1 U5849 ( .A(n5018), .B(n10570), .ZN(n5364) );
  NOR2_X1 U5850 ( .A1(n7802), .A2(n7803), .ZN(n7826) );
  NAND2_X1 U5851 ( .A1(n8280), .A2(n8434), .ZN(n8374) );
  NOR2_X1 U5852 ( .A1(n7426), .A2(n7427), .ZN(n7494) );
  NOR2_X1 U5853 ( .A1(n7826), .A2(n4928), .ZN(n8031) );
  AND2_X1 U5854 ( .A1(n8397), .A2(n8396), .ZN(n8459) );
  NAND2_X1 U5855 ( .A1(n8082), .A2(n8081), .ZN(n8229) );
  OR2_X1 U5856 ( .A1(n8080), .A2(n8079), .ZN(n8081) );
  AND2_X1 U5857 ( .A1(n8288), .A2(n8405), .ZN(n8407) );
  AND4_X1 U5858 ( .A1(n5375), .A2(n5374), .A3(n5373), .A4(n5372), .ZN(n7554)
         );
  AND3_X1 U5859 ( .A1(n5397), .A2(n5396), .A3(n5395), .ZN(n7555) );
  NAND2_X1 U5860 ( .A1(n4919), .A2(n4920), .ZN(n7689) );
  AND3_X1 U5861 ( .A1(n5382), .A2(n5381), .A3(n5380), .ZN(n10147) );
  NAND2_X1 U5862 ( .A1(n4922), .A2(n4924), .ZN(n8033) );
  AND3_X1 U5863 ( .A1(n5317), .A2(n5316), .A3(n5315), .ZN(n8759) );
  AND2_X1 U5864 ( .A1(n4937), .A2(n4935), .ZN(n8364) );
  NAND2_X1 U5865 ( .A1(n4937), .A2(n4938), .ZN(n8230) );
  AND4_X1 U5866 ( .A1(n5581), .A2(n5580), .A3(n5579), .A4(n5578), .ZN(n8761)
         );
  NAND2_X1 U5867 ( .A1(n4919), .A2(n4918), .ZN(n7800) );
  AND2_X1 U5868 ( .A1(n4532), .A2(n7691), .ZN(n4918) );
  AND2_X1 U5869 ( .A1(n4919), .A2(n4532), .ZN(n7692) );
  AOI21_X1 U5870 ( .B1(n8666), .B2(n5719), .A(n5655), .ZN(n8653) );
  INV_X1 U5871 ( .A(n8299), .ZN(n4916) );
  INV_X1 U5872 ( .A(n8482), .ZN(n8472) );
  INV_X1 U5873 ( .A(n8490), .ZN(n8479) );
  INV_X1 U5874 ( .A(n8378), .ZN(n8496) );
  NAND2_X1 U5875 ( .A1(n8246), .A2(n8245), .ZN(n8485) );
  INV_X1 U5876 ( .A(n8717), .ZN(n8501) );
  INV_X1 U5877 ( .A(n7554), .ZN(n7666) );
  NAND2_X1 U5878 ( .A1(n5344), .A2(n5107), .ZN(n8514) );
  INV_X1 U5879 ( .A(n5108), .ZN(n5107) );
  AND2_X1 U5880 ( .A1(n5341), .A2(n5340), .ZN(n5344) );
  OAI21_X1 U5881 ( .B1(n6881), .B2(n10200), .A(n5109), .ZN(n5108) );
  OR2_X1 U5882 ( .A1(n5562), .A2(n8209), .ZN(n5321) );
  OR2_X1 U5883 ( .A1(n6881), .A2(n5318), .ZN(n5322) );
  NAND2_X1 U5884 ( .A1(n5153), .A2(n4781), .ZN(n8516) );
  INV_X1 U5885 ( .A(n4782), .ZN(n4781) );
  OAI22_X1 U5886 ( .A1(n6582), .A2(n6881), .B1(n5562), .B2(n10630), .ZN(n4782)
         );
  OR2_X1 U5887 ( .A1(n7176), .A2(n7174), .ZN(n8606) );
  OAI21_X1 U5888 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7115), .A(n8212), .ZN(n7116) );
  NAND2_X1 U5889 ( .A1(n6637), .A2(n4941), .ZN(n6583) );
  NAND2_X1 U5890 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n4942), .ZN(n4941) );
  OAI21_X1 U5891 ( .B1(n8205), .B2(n5318), .A(n6584), .ZN(n10111) );
  INV_X1 U5892 ( .A(n7235), .ZN(n7139) );
  NAND2_X1 U5893 ( .A1(n4957), .A2(n6693), .ZN(n7283) );
  INV_X1 U5894 ( .A(n4956), .ZN(n4955) );
  AND2_X1 U5895 ( .A1(n4957), .A2(n4956), .ZN(n7369) );
  NAND2_X1 U5896 ( .A1(n4846), .A2(n4845), .ZN(n7730) );
  INV_X1 U5897 ( .A(n4846), .ZN(n7728) );
  NOR2_X1 U5898 ( .A1(n7893), .A2(n5445), .ZN(n7892) );
  NOR2_X1 U5899 ( .A1(n7892), .A2(n6597), .ZN(n7965) );
  NAND2_X1 U5900 ( .A1(n4823), .A2(n4549), .ZN(n4822) );
  INV_X1 U5901 ( .A(n8114), .ZN(n4823) );
  NAND2_X1 U5902 ( .A1(n8114), .A2(n4825), .ZN(n4820) );
  NAND2_X1 U5903 ( .A1(n4545), .A2(n4825), .ZN(n4824) );
  INV_X1 U5904 ( .A(n5090), .ZN(n6600) );
  NOR2_X1 U5905 ( .A1(n8520), .A2(n8190), .ZN(n8521) );
  INV_X1 U5906 ( .A(n4950), .ZN(n8543) );
  NAND2_X1 U5907 ( .A1(n4840), .A2(n4838), .ZN(n8535) );
  NAND2_X1 U5908 ( .A1(n6601), .A2(n4841), .ZN(n4840) );
  OR2_X1 U5909 ( .A1(n8520), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U5910 ( .A1(n4841), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4839) );
  INV_X1 U5911 ( .A(n5097), .ZN(n8558) );
  OR2_X1 U5912 ( .A1(n8560), .A2(n8559), .ZN(n5097) );
  INV_X1 U5913 ( .A(n6603), .ZN(n5096) );
  INV_X1 U5914 ( .A(n4832), .ZN(n8578) );
  INV_X1 U5915 ( .A(n4952), .ZN(n8576) );
  NAND2_X1 U5916 ( .A1(n5098), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U5917 ( .A1(n6603), .A2(n5098), .ZN(n5094) );
  INV_X1 U5918 ( .A(n8569), .ZN(n5098) );
  AOI21_X1 U5919 ( .B1(n9053), .B2(n6875), .A(n6874), .ZN(n8625) );
  XNOR2_X1 U5920 ( .A(n6886), .B(n6846), .ZN(n8347) );
  NAND2_X1 U5921 ( .A1(n4699), .A2(n5767), .ZN(n6886) );
  OR2_X1 U5922 ( .A1(n8620), .A2(n5705), .ZN(n8639) );
  AND2_X1 U5923 ( .A1(n5630), .A2(n5629), .ZN(n8680) );
  NAND2_X1 U5924 ( .A1(n5616), .A2(n5615), .ZN(n8809) );
  NAND2_X1 U5925 ( .A1(n5607), .A2(n5606), .ZN(n8719) );
  NAND2_X1 U5926 ( .A1(n5574), .A2(n5573), .ZN(n8830) );
  NOR2_X1 U5927 ( .A1(n5138), .A2(n5140), .ZN(n5172) );
  INV_X1 U5928 ( .A(n8051), .ZN(n5138) );
  AND2_X1 U5929 ( .A1(n5134), .A2(n6759), .ZN(n7949) );
  NAND2_X1 U5930 ( .A1(n5444), .A2(n5443), .ZN(n10171) );
  NAND2_X1 U5931 ( .A1(n4886), .A2(n4883), .ZN(n7815) );
  NAND2_X1 U5932 ( .A1(n4872), .A2(n5368), .ZN(n7486) );
  OR2_X1 U5933 ( .A1(n7333), .A2(n5369), .ZN(n4872) );
  INV_X1 U5934 ( .A(n8770), .ZN(n10132) );
  INV_X1 U5935 ( .A(n7273), .ZN(n10142) );
  AND3_X1 U5936 ( .A1(n10181), .A2(n7177), .A3(n7176), .ZN(n10133) );
  NOR2_X1 U5937 ( .A1(n10213), .A2(n8793), .ZN(n4892) );
  NAND2_X1 U5938 ( .A1(n6853), .A2(n6852), .ZN(n8838) );
  NAND2_X1 U5939 ( .A1(n8635), .A2(n8634), .ZN(n8636) );
  NAND2_X1 U5940 ( .A1(n8633), .A2(n10118), .ZN(n8634) );
  NAND2_X1 U5941 ( .A1(n5122), .A2(n6838), .ZN(n8642) );
  NAND2_X1 U5942 ( .A1(n8655), .A2(n8656), .ZN(n5122) );
  AOI21_X1 U5943 ( .B1(n4896), .B2(n10123), .A(n4893), .ZN(n8847) );
  NAND2_X1 U5944 ( .A1(n4895), .A2(n4894), .ZN(n4893) );
  XNOR2_X1 U5945 ( .A(n8643), .B(n4788), .ZN(n4896) );
  NAND2_X1 U5946 ( .A1(n8645), .A2(n10118), .ZN(n4894) );
  AND2_X1 U5947 ( .A1(n5662), .A2(n5661), .ZN(n8856) );
  NAND2_X1 U5948 ( .A1(n5650), .A2(n5649), .ZN(n8860) );
  INV_X1 U5949 ( .A(n8680), .ZN(n8866) );
  NAND2_X1 U5950 ( .A1(n8753), .A2(n5147), .ZN(n5145) );
  NAND2_X1 U5951 ( .A1(n5310), .A2(n5309), .ZN(n8892) );
  AND2_X1 U5952 ( .A1(n8748), .A2(n8747), .ZN(n8890) );
  NAND2_X1 U5953 ( .A1(n8753), .A2(n6805), .ZN(n8738) );
  NAND2_X1 U5954 ( .A1(n5557), .A2(n5556), .ZN(n8414) );
  NAND2_X1 U5955 ( .A1(n5116), .A2(n6791), .ZN(n8164) );
  OR2_X1 U5956 ( .A1(n8142), .A2(n6790), .ZN(n5116) );
  NAND2_X1 U5957 ( .A1(n5528), .A2(n5527), .ZN(n8240) );
  AND2_X1 U5958 ( .A1(n4862), .A2(n4861), .ZN(n8150) );
  NAND2_X1 U5959 ( .A1(n7921), .A2(n5521), .ZN(n4861) );
  INV_X1 U5960 ( .A(n8900), .ZN(n8891) );
  NAND2_X1 U5961 ( .A1(n8122), .A2(n5748), .ZN(n8179) );
  XNOR2_X1 U5962 ( .A(n5791), .B(n5790), .ZN(n7963) );
  NAND2_X1 U5963 ( .A1(n5795), .A2(n5794), .ZN(n7932) );
  MUX2_X1 U5964 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5732), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5734) );
  XNOR2_X1 U5965 ( .A(n5506), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7905) );
  INV_X1 U5966 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6972) );
  INV_X1 U5967 ( .A(n5345), .ZN(n5093) );
  NAND2_X1 U5968 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5324) );
  NAND2_X1 U5969 ( .A1(n7880), .A2(n6127), .ZN(n7864) );
  NAND2_X1 U5970 ( .A1(n6289), .A2(n6288), .ZN(n9843) );
  OAI22_X1 U5971 ( .A1(n9060), .A2(n8342), .B1(n9340), .B2(n4649), .ZN(n6287)
         );
  OR2_X1 U5972 ( .A1(n5944), .A2(n6387), .ZN(n5945) );
  INV_X1 U5973 ( .A(n4746), .ZN(n8941) );
  INV_X1 U5974 ( .A(n4754), .ZN(n4747) );
  NAND2_X1 U5975 ( .A1(n9042), .A2(n9047), .ZN(n8960) );
  NAND2_X1 U5976 ( .A1(n5080), .A2(n8957), .ZN(n8970) );
  OR2_X1 U5977 ( .A1(n8960), .A2(n8958), .ZN(n5080) );
  NAND2_X1 U5978 ( .A1(n6252), .A2(n6251), .ZN(n8977) );
  NAND2_X1 U5979 ( .A1(n6361), .A2(n6360), .ZN(n9636) );
  NAND2_X1 U5980 ( .A1(n4734), .A2(n9025), .ZN(n8987) );
  NAND2_X1 U5981 ( .A1(n4736), .A2(n4735), .ZN(n4734) );
  INV_X1 U5982 ( .A(n8983), .ZN(n4735) );
  NAND2_X1 U5983 ( .A1(n8921), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U5984 ( .A1(n4752), .A2(n4756), .ZN(n8991) );
  NAND2_X1 U5985 ( .A1(n4759), .A2(n4758), .ZN(n4752) );
  OAI21_X1 U5986 ( .B1(n7107), .B2(n7108), .A(n5947), .ZN(n7123) );
  OR2_X1 U5987 ( .A1(n6476), .A2(n6475), .ZN(n9028) );
  INV_X1 U5988 ( .A(n9046), .ZN(n9025) );
  INV_X1 U5989 ( .A(n9332), .ZN(n9331) );
  AND2_X1 U5990 ( .A1(n4768), .A2(n7017), .ZN(n7042) );
  INV_X1 U5991 ( .A(n4768), .ZN(n7025) );
  NOR2_X1 U5992 ( .A1(n7072), .A2(n4605), .ZN(n7076) );
  NOR2_X1 U5993 ( .A1(n7076), .A2(n7075), .ZN(n7201) );
  INV_X1 U5994 ( .A(n4772), .ZN(n9433) );
  OR2_X1 U5995 ( .A1(n9463), .A2(n4765), .ZN(n9479) );
  INV_X1 U5996 ( .A(n9465), .ZN(n4765) );
  INV_X1 U5997 ( .A(n9463), .ZN(n9464) );
  NAND2_X1 U5998 ( .A1(n9946), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4776) );
  INV_X1 U5999 ( .A(n9556), .ZN(n4775) );
  OAI21_X1 U6000 ( .B1(n9554), .B2(n9962), .A(n9553), .ZN(n4780) );
  OAI21_X1 U6001 ( .B1(n9550), .B2(n9962), .A(n4778), .ZN(n4777) );
  OR2_X1 U6002 ( .A1(n9552), .A2(n9957), .ZN(n4778) );
  NOR2_X1 U6003 ( .A1(n9557), .A2(n9715), .ZN(n9762) );
  NAND2_X1 U6004 ( .A1(n9056), .A2(n4547), .ZN(n4960) );
  NAND2_X1 U6005 ( .A1(n9593), .A2(n4962), .ZN(n4961) );
  NOR2_X1 U6006 ( .A1(n9565), .A2(n9715), .ZN(n9766) );
  AOI21_X1 U6007 ( .B1(n6565), .B2(n10075), .A(n6564), .ZN(n8314) );
  NAND2_X1 U6008 ( .A1(n5055), .A2(n5054), .ZN(n9572) );
  INV_X1 U6009 ( .A(n9783), .ZN(n9608) );
  NAND2_X1 U6010 ( .A1(n6390), .A2(n6389), .ZN(n9613) );
  NAND2_X1 U6011 ( .A1(n4989), .A2(n6527), .ZN(n9641) );
  AND2_X1 U6012 ( .A1(n9691), .A2(n9185), .ZN(n9675) );
  OAI21_X1 U6013 ( .B1(n4636), .B2(n4557), .A(n6522), .ZN(n9678) );
  NAND2_X1 U6014 ( .A1(n6315), .A2(n6314), .ZN(n9688) );
  NAND2_X1 U6015 ( .A1(n6274), .A2(n6273), .ZN(n9744) );
  NAND2_X1 U6016 ( .A1(n9923), .A2(n6516), .ZN(n7983) );
  OR2_X1 U6017 ( .A1(n7916), .A2(n9085), .ZN(n9923) );
  AND2_X1 U6018 ( .A1(n7838), .A2(n9276), .ZN(n7908) );
  AND2_X1 U6019 ( .A1(n7778), .A2(n9163), .ZN(n5171) );
  NAND2_X1 U6020 ( .A1(n7765), .A2(n6510), .ZN(n7777) );
  AND2_X1 U6021 ( .A1(n7524), .A2(n9154), .ZN(n7677) );
  NAND2_X1 U6022 ( .A1(n5058), .A2(n7524), .ZN(n7676) );
  NAND2_X1 U6023 ( .A1(n6034), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U6024 ( .A1(n6411), .A2(n6410), .ZN(n9871) );
  AND2_X1 U6025 ( .A1(n7020), .A2(n6987), .ZN(n9995) );
  OR2_X1 U6026 ( .A1(n4730), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U6027 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n4729) );
  NOR2_X1 U6028 ( .A1(n5880), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4730) );
  NAND2_X1 U6029 ( .A1(n5033), .A2(n5252), .ZN(n5257) );
  CLKBUF_X1 U6030 ( .A(n6286), .Z(n9340) );
  INV_X1 U6031 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U6032 ( .A1(n5896), .A2(n4763), .ZN(n7028) );
  XNOR2_X1 U6033 ( .A(n4688), .B(n7547), .ZN(n6929) );
  NAND2_X1 U6034 ( .A1(n8596), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7119) );
  INV_X1 U6035 ( .A(n4947), .ZN(n8008) );
  INV_X1 U6036 ( .A(n5092), .ZN(n8104) );
  AOI21_X1 U6037 ( .B1(n5106), .B2(n10114), .A(n5102), .ZN(n8598) );
  NAND2_X1 U6038 ( .A1(n5105), .A2(n5103), .ZN(n5102) );
  OAI21_X1 U6039 ( .B1(n8612), .B2(n4535), .A(n6720), .ZN(n4959) );
  OR2_X1 U6040 ( .A1(n6611), .A2(n8618), .ZN(n6723) );
  AOI21_X1 U6041 ( .B1(n5828), .B2(n6959), .A(n6958), .ZN(n6960) );
  OAI21_X1 U6042 ( .B1(n8847), .B2(n10211), .A(n4889), .ZN(P2_U3486) );
  INV_X1 U6043 ( .A(n4890), .ZN(n4889) );
  OAI21_X1 U6044 ( .B1(n8852), .B2(n8823), .A(n4891), .ZN(n4890) );
  NOR2_X1 U6045 ( .A1(n4624), .A2(n4892), .ZN(n4891) );
  NOR2_X1 U6046 ( .A1(n5081), .A2(n6490), .ZN(n6491) );
  NAND2_X1 U6047 ( .A1(n4779), .A2(n4773), .ZN(P1_U3262) );
  AOI21_X1 U6048 ( .B1(n4777), .B2(n9340), .A(n4774), .ZN(n4773) );
  NAND2_X1 U6049 ( .A1(n4780), .A2(n9555), .ZN(n4779) );
  NAND2_X1 U6050 ( .A1(n4776), .A2(n4775), .ZN(n4774) );
  NOR2_X1 U6051 ( .A1(n6577), .A2(n5169), .ZN(n6578) );
  NOR2_X1 U6052 ( .A1(n6727), .A2(n4627), .ZN(n4976) );
  NAND2_X1 U6053 ( .A1(n6725), .A2(n10078), .ZN(n4977) );
  INV_X1 U6054 ( .A(n5991), .ZN(n6114) );
  INV_X2 U6055 ( .A(n6114), .ZN(n6074) );
  AND2_X1 U6056 ( .A1(n4741), .A2(n4740), .ZN(n4528) );
  INV_X1 U6057 ( .A(n6847), .ZN(n5016) );
  NAND2_X2 U6058 ( .A1(n5287), .A2(n8318), .ZN(n5339) );
  AND2_X1 U6059 ( .A1(n7951), .A2(n6759), .ZN(n4529) );
  AND2_X1 U6060 ( .A1(n5073), .A2(n8982), .ZN(n4530) );
  AND2_X1 U6061 ( .A1(n8141), .A2(n4802), .ZN(n4531) );
  AND2_X1 U6062 ( .A1(n4920), .A2(n4584), .ZN(n4532) );
  INV_X1 U6063 ( .A(n5740), .ZN(n4871) );
  AND2_X1 U6064 ( .A1(n4875), .A2(n8731), .ZN(n4533) );
  AND2_X1 U6065 ( .A1(n4792), .A2(n4614), .ZN(n4534) );
  AND2_X1 U6066 ( .A1(n8614), .A2(n8613), .ZN(n4535) );
  AND2_X1 U6067 ( .A1(n4530), .A2(n5075), .ZN(n4536) );
  AND2_X1 U6068 ( .A1(n4785), .A2(n4580), .ZN(n4537) );
  AND2_X1 U6069 ( .A1(n7497), .A2(n4921), .ZN(n4538) );
  AND2_X1 U6070 ( .A1(n4975), .A2(n4974), .ZN(n4539) );
  AND2_X1 U6071 ( .A1(n8968), .A2(n8967), .ZN(n4540) );
  AND2_X1 U6072 ( .A1(n8029), .A2(n8028), .ZN(n4541) );
  NAND2_X1 U6073 ( .A1(n8445), .A2(n8268), .ZN(n4542) );
  AND2_X1 U6074 ( .A1(n4836), .A2(n4833), .ZN(n4543) );
  OR2_X1 U6075 ( .A1(n7978), .A2(n10208), .ZN(n4544) );
  AND2_X1 U6076 ( .A1(n7096), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4545) );
  AND2_X1 U6077 ( .A1(n4617), .A2(n7880), .ZN(n4546) );
  OR2_X1 U6078 ( .A1(n9564), .A2(n4964), .ZN(n4547) );
  AND2_X1 U6079 ( .A1(n9291), .A2(n9316), .ZN(n9096) );
  INV_X1 U6080 ( .A(n8931), .ZN(n4758) );
  AND2_X1 U6081 ( .A1(n6888), .A2(n5767), .ZN(n4548) );
  AND2_X1 U6082 ( .A1(n5277), .A2(n5276), .ZN(n8805) );
  INV_X1 U6083 ( .A(n8805), .ZN(n8872) );
  NOR2_X1 U6084 ( .A1(n4545), .A2(n4825), .ZN(n4549) );
  AND2_X1 U6085 ( .A1(n4970), .A2(n9626), .ZN(n4550) );
  NAND2_X1 U6086 ( .A1(n4633), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4847) );
  INV_X1 U6087 ( .A(n7865), .ZN(n4741) );
  XNOR2_X1 U6088 ( .A(n5280), .B(n5271), .ZN(n5772) );
  INV_X2 U6089 ( .A(n5943), .ZN(n6438) );
  NAND2_X1 U6090 ( .A1(n4760), .A2(n5074), .ZN(n8999) );
  INV_X1 U6091 ( .A(n6902), .ZN(n5745) );
  OR2_X1 U6092 ( .A1(n7570), .A2(n6592), .ZN(n4551) );
  AND2_X1 U6093 ( .A1(n9276), .A2(n9164), .ZN(n4552) );
  OAI21_X1 U6094 ( .B1(n8999), .B2(n8998), .A(n9003), .ZN(n8922) );
  OR2_X1 U6095 ( .A1(n7805), .A2(n10157), .ZN(n4553) );
  AND2_X1 U6096 ( .A1(n8923), .A2(n5072), .ZN(n4554) );
  OR2_X1 U6097 ( .A1(n7215), .A2(n7214), .ZN(n4555) );
  OR2_X1 U6098 ( .A1(n8532), .A2(n6707), .ZN(n4556) );
  AND2_X1 U6099 ( .A1(n9698), .A2(n9828), .ZN(n4557) );
  OR2_X1 U6100 ( .A1(n5828), .A2(n8499), .ZN(n6888) );
  AND2_X1 U6101 ( .A1(n9684), .A2(n4970), .ZN(n4558) );
  OR2_X1 U6102 ( .A1(n8240), .A2(n8505), .ZN(n4559) );
  INV_X1 U6103 ( .A(n9269), .ZN(n5057) );
  INV_X1 U6104 ( .A(n8514), .ZN(n5351) );
  OR2_X1 U6105 ( .A1(n10171), .A2(n8059), .ZN(n6759) );
  NAND2_X1 U6106 ( .A1(n5739), .A2(n6732), .ZN(n6897) );
  AND2_X1 U6107 ( .A1(n6126), .A2(n7865), .ZN(n4560) );
  NAND4_X1 U6108 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n8515)
         );
  INV_X1 U6109 ( .A(n8515), .ZN(n7271) );
  AND2_X1 U6110 ( .A1(n9274), .A2(n9161), .ZN(n4561) );
  OR2_X1 U6111 ( .A1(n5409), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n4562) );
  INV_X1 U6112 ( .A(n7029), .ZN(n4647) );
  NAND2_X1 U6113 ( .A1(n6332), .A2(n6331), .ZN(n9670) );
  INV_X1 U6114 ( .A(n6690), .ZN(n7254) );
  XNOR2_X1 U6115 ( .A(n5379), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6690) );
  AND4_X1 U6116 ( .A1(n5895), .A2(n5064), .A3(n5832), .A4(n5833), .ZN(n6026)
         );
  AOI21_X1 U6117 ( .B1(n4926), .B2(n7803), .A(n8030), .ZN(n4925) );
  OR2_X1 U6118 ( .A1(n8266), .A2(n8456), .ZN(n4563) );
  AND2_X1 U6119 ( .A1(n4721), .A2(n5228), .ZN(n4564) );
  AND2_X1 U6120 ( .A1(n4924), .A2(n4927), .ZN(n4565) );
  NOR2_X1 U6121 ( .A1(n10121), .A2(n7823), .ZN(n4566) );
  NAND2_X1 U6122 ( .A1(n6131), .A2(n5860), .ZN(n6149) );
  NOR2_X1 U6123 ( .A1(n5229), .A2(SI_16_), .ZN(n4567) );
  AND2_X1 U6124 ( .A1(n5739), .A2(n4808), .ZN(n4568) );
  INV_X1 U6125 ( .A(n4665), .ZN(n4664) );
  AND2_X1 U6126 ( .A1(n8866), .A2(n8692), .ZN(n6825) );
  NAND2_X1 U6127 ( .A1(n6193), .A2(n6192), .ZN(n9111) );
  NAND2_X1 U6128 ( .A1(n9927), .A2(n10065), .ZN(n4569) );
  OR2_X1 U6129 ( .A1(n5078), .A2(n5076), .ZN(n4570) );
  NAND2_X1 U6130 ( .A1(n9744), .A2(n9711), .ZN(n4571) );
  AND2_X1 U6131 ( .A1(n8977), .A2(n9918), .ZN(n4573) );
  AND2_X1 U6132 ( .A1(n5097), .A2(n5096), .ZN(n4574) );
  AND2_X1 U6133 ( .A1(n6202), .A2(n6188), .ZN(n4575) );
  AND2_X1 U6134 ( .A1(n5048), .A2(n9224), .ZN(n4576) );
  NAND2_X1 U6135 ( .A1(n4897), .A2(n7271), .ZN(n4898) );
  NAND2_X1 U6136 ( .A1(n8141), .A2(n4799), .ZN(n4577) );
  AND2_X1 U6137 ( .A1(n5037), .A2(n4716), .ZN(n4578) );
  INV_X1 U6138 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5259) );
  NOR2_X1 U6139 ( .A1(n8274), .A2(n8273), .ZN(n4579) );
  NAND2_X1 U6140 ( .A1(n6846), .A2(n6859), .ZN(n4580) );
  AND2_X1 U6141 ( .A1(n5195), .A2(SI_6_), .ZN(n4581) );
  AND2_X1 U6142 ( .A1(n5221), .A2(SI_13_), .ZN(n4582) );
  AND2_X1 U6143 ( .A1(n5219), .A2(SI_12_), .ZN(n4583) );
  NAND2_X1 U6144 ( .A1(n7690), .A2(n7693), .ZN(n4584) );
  AND2_X1 U6145 ( .A1(n5741), .A2(n5398), .ZN(n4585) );
  OR2_X1 U6146 ( .A1(n8237), .A2(n8226), .ZN(n4586) );
  AND2_X1 U6147 ( .A1(n5877), .A2(n4731), .ZN(n4587) );
  INV_X1 U6148 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5860) );
  XNOR2_X1 U6149 ( .A(n5221), .B(SI_13_), .ZN(n5455) );
  INV_X1 U6150 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6130) );
  AND2_X1 U6151 ( .A1(n4706), .A2(n4708), .ZN(n4588) );
  NAND2_X1 U6152 ( .A1(n6887), .A2(n4700), .ZN(n4589) );
  AND2_X1 U6153 ( .A1(n10121), .A2(n7823), .ZN(n4590) );
  NAND2_X1 U6154 ( .A1(n9191), .A2(n5047), .ZN(n4591) );
  OR2_X1 U6155 ( .A1(n9111), .A2(n9346), .ZN(n4592) );
  AND3_X1 U6156 ( .A1(n5346), .A2(n5259), .A3(n5126), .ZN(n4593) );
  AND2_X1 U6157 ( .A1(n6753), .A2(n6952), .ZN(n4594) );
  AND2_X1 U6158 ( .A1(n8141), .A2(n4800), .ZN(n4595) );
  AND2_X1 U6159 ( .A1(n8237), .A2(n8506), .ZN(n6785) );
  NOR2_X1 U6160 ( .A1(n10041), .A2(n10029), .ZN(n4596) );
  NAND2_X1 U6161 ( .A1(n6783), .A2(n5497), .ZN(n4597) );
  AND2_X1 U6162 ( .A1(n6265), .A2(n5077), .ZN(n4598) );
  INV_X1 U6163 ( .A(n5027), .ZN(n5026) );
  NOR2_X1 U6164 ( .A1(n5220), .A2(n5028), .ZN(n5027) );
  NOR2_X1 U6165 ( .A1(n4566), .A2(n4885), .ZN(n4884) );
  AND2_X1 U6166 ( .A1(n6545), .A2(n6547), .ZN(n4599) );
  AND2_X1 U6167 ( .A1(n4592), .A2(n6510), .ZN(n4600) );
  INV_X1 U6168 ( .A(n9576), .ZN(n9569) );
  AND2_X1 U6169 ( .A1(n9290), .A2(n9206), .ZN(n9576) );
  AND2_X1 U6170 ( .A1(n4673), .A2(n4676), .ZN(n4601) );
  AND2_X1 U6171 ( .A1(n6918), .A2(n6888), .ZN(n4602) );
  OR2_X1 U6172 ( .A1(n8298), .A2(n8297), .ZN(n4603) );
  INV_X1 U6173 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5554) );
  INV_X1 U6174 ( .A(n5918), .ZN(n6042) );
  NAND2_X1 U6175 ( .A1(n7711), .A2(n6109), .ZN(n4745) );
  XNOR2_X1 U6176 ( .A(n5361), .B(n5259), .ZN(n6963) );
  INV_X1 U6177 ( .A(n6963), .ZN(n4833) );
  AND2_X1 U6178 ( .A1(n8485), .A2(n8250), .ZN(n4604) );
  NAND2_X1 U6179 ( .A1(n5454), .A2(n6902), .ZN(n7921) );
  INV_X1 U6180 ( .A(n8511), .ZN(n8028) );
  INV_X1 U6181 ( .A(n8644), .ZN(n4788) );
  INV_X1 U6182 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5020) );
  AND2_X1 U6183 ( .A1(n7077), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4605) );
  OR2_X1 U6184 ( .A1(n8939), .A2(n8938), .ZN(n4606) );
  AND2_X1 U6185 ( .A1(n7530), .A2(n4539), .ZN(n4607) );
  OAI21_X1 U6186 ( .B1(n8319), .B2(n5328), .A(n5718), .ZN(n5828) );
  INV_X1 U6187 ( .A(n9063), .ZN(n5059) );
  AND2_X1 U6188 ( .A1(n9209), .A2(n9215), .ZN(n4608) );
  XNOR2_X1 U6189 ( .A(n5878), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6450) );
  INV_X1 U6190 ( .A(n8507), .ZN(n8232) );
  INV_X1 U6191 ( .A(n8149), .ZN(n4803) );
  AND3_X1 U6192 ( .A1(n6486), .A2(n9025), .A3(n6485), .ZN(n4609) );
  AND2_X1 U6193 ( .A1(n9223), .A2(n9205), .ZN(n9589) );
  INV_X1 U6194 ( .A(n9589), .ZN(n5052) );
  NOR2_X1 U6195 ( .A1(n6601), .A2(n8521), .ZN(n4610) );
  AND2_X1 U6196 ( .A1(n4874), .A2(n4875), .ZN(n4611) );
  NAND2_X1 U6197 ( .A1(n6426), .A2(n6425), .ZN(n9867) );
  INV_X1 U6198 ( .A(n4967), .ZN(n9714) );
  NOR2_X1 U6199 ( .A1(n9739), .A2(n9843), .ZN(n4967) );
  AND2_X1 U6200 ( .A1(n8798), .A2(n8653), .ZN(n4612) );
  OR2_X1 U6201 ( .A1(n9867), .A2(n9597), .ZN(n9290) );
  INV_X1 U6202 ( .A(n9290), .ZN(n5051) );
  INV_X1 U6203 ( .A(n5075), .ZN(n5074) );
  NOR2_X1 U6204 ( .A1(n6330), .A2(n6329), .ZN(n5075) );
  AND2_X1 U6205 ( .A1(n4947), .A2(n4946), .ZN(n4613) );
  AND2_X1 U6206 ( .A1(n5292), .A2(n5291), .ZN(n8707) );
  INV_X1 U6207 ( .A(n8707), .ZN(n8677) );
  NAND2_X1 U6208 ( .A1(n6378), .A2(n6377), .ZN(n9878) );
  NAND2_X1 U6209 ( .A1(n8834), .A2(n6885), .ZN(n4614) );
  OR2_X1 U6210 ( .A1(n8414), .A2(n8487), .ZN(n6792) );
  NAND2_X1 U6211 ( .A1(n8872), .A2(n8677), .ZN(n4615) );
  AND2_X1 U6212 ( .A1(n5247), .A2(SI_21_), .ZN(n4616) );
  AND2_X1 U6213 ( .A1(n6127), .A2(n4741), .ZN(n4617) );
  NAND2_X1 U6214 ( .A1(n5245), .A2(SI_20_), .ZN(n4618) );
  INV_X1 U6215 ( .A(n4757), .ZN(n4756) );
  NOR2_X1 U6216 ( .A1(n6302), .A2(n6303), .ZN(n4757) );
  OR2_X1 U6217 ( .A1(n5247), .A2(SI_21_), .ZN(n4619) );
  AND2_X1 U6218 ( .A1(n6527), .A2(n5170), .ZN(n4620) );
  AND2_X1 U6219 ( .A1(n4757), .A2(n8988), .ZN(n4621) );
  INV_X1 U6220 ( .A(n5711), .ZN(n8843) );
  AND2_X1 U6221 ( .A1(n5703), .A2(n5702), .ZN(n5711) );
  INV_X1 U6222 ( .A(n9096), .ZN(n9212) );
  AND2_X1 U6223 ( .A1(n9055), .A2(n9054), .ZN(n9860) );
  XNOR2_X1 U6224 ( .A(n5729), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7175) );
  INV_X1 U6225 ( .A(n7175), .ZN(n4809) );
  INV_X1 U6226 ( .A(n8532), .ZN(n4825) );
  NAND2_X1 U6227 ( .A1(n6306), .A2(n6305), .ZN(n9698) );
  INV_X1 U6228 ( .A(n9698), .ZN(n4966) );
  INV_X1 U6229 ( .A(n6126), .ZN(n4740) );
  NAND2_X1 U6230 ( .A1(n5800), .A2(n5801), .ZN(n5803) );
  AND2_X1 U6231 ( .A1(n7322), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4622) );
  AND2_X1 U6232 ( .A1(n9436), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U6233 ( .A1(n4982), .A2(n6503), .ZN(n7653) );
  INV_X1 U6234 ( .A(n8382), .ZN(n4906) );
  INV_X1 U6235 ( .A(n8957), .ZN(n5079) );
  INV_X1 U6236 ( .A(n8988), .ZN(n4755) );
  AND2_X1 U6237 ( .A1(n8849), .A2(n6959), .ZN(n4624) );
  AND2_X1 U6238 ( .A1(n7257), .A2(n6006), .ZN(n4625) );
  AND2_X1 U6239 ( .A1(n4869), .A2(n5741), .ZN(n4626) );
  NOR2_X1 U6240 ( .A1(n10078), .A2(n6726), .ZN(n4627) );
  NOR2_X1 U6241 ( .A1(n7965), .A2(n7964), .ZN(n4628) );
  OAI21_X1 U6242 ( .B1(n4725), .B2(n4724), .A(n6050), .ZN(n7454) );
  INV_X1 U6243 ( .A(n9131), .ZN(n4968) );
  NAND2_X1 U6244 ( .A1(n6174), .A2(n6173), .ZN(n7997) );
  INV_X1 U6245 ( .A(n7997), .ZN(n4974) );
  NOR2_X1 U6246 ( .A1(n7107), .A2(n7108), .ZN(n4629) );
  AND2_X1 U6247 ( .A1(n4955), .A2(n4957), .ZN(n4630) );
  NAND2_X1 U6248 ( .A1(n5734), .A2(n5733), .ZN(n7700) );
  NAND2_X1 U6249 ( .A1(n9400), .A2(n9401), .ZN(n4770) );
  AOI21_X1 U6250 ( .B1(n8596), .B2(n8597), .A(n5104), .ZN(n5103) );
  XNOR2_X1 U6251 ( .A(n6605), .B(n8597), .ZN(n8590) );
  XNOR2_X1 U6252 ( .A(n6711), .B(n8597), .ZN(n8586) );
  NAND2_X1 U6253 ( .A1(n10092), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4638) );
  NOR2_X4 U6254 ( .A1(n9991), .A2(n7518), .ZN(n9731) );
  OAI21_X1 U6255 ( .B1(P1_RD_REG_SCAN_IN), .B2(P1_ADDR_REG_19__SCAN_IN), .A(
        n4687), .ZN(n5173) );
  OAI22_X1 U6256 ( .A1(n8704), .A2(n8705), .B1(n8501), .B2(n8809), .ZN(n8690)
         );
  OAI22_X1 U6257 ( .A1(n8673), .A2(n5639), .B1(n8866), .B2(n8500), .ZN(n8662)
         );
  AOI21_X1 U6258 ( .B1(n8637), .B2(n10123), .A(n8636), .ZN(n8841) );
  NAND2_X1 U6259 ( .A1(n5161), .A2(n8042), .ZN(n4631) );
  NAND2_X1 U6260 ( .A1(n5481), .A2(n5027), .ZN(n5022) );
  NAND2_X1 U6261 ( .A1(n5022), .A2(n5025), .ZN(n5456) );
  OAI21_X2 U6262 ( .B1(n7916), .B2(n4993), .A(n4991), .ZN(n9730) );
  OR2_X1 U6263 ( .A1(n10041), .A2(n9971), .ZN(n9119) );
  OR2_X1 U6264 ( .A1(n10031), .A2(n7580), .ZN(n9258) );
  INV_X4 U6265 ( .A(n6239), .ZN(n6478) );
  NAND2_X1 U6266 ( .A1(n4977), .A2(n4976), .ZN(P1_U3519) );
  NAND2_X1 U6267 ( .A1(n4844), .A2(n4842), .ZN(n6596) );
  NOR2_X1 U6268 ( .A1(n7287), .A2(n5383), .ZN(n7286) );
  INV_X1 U6269 ( .A(n6588), .ZN(n4849) );
  NAND2_X1 U6270 ( .A1(n10110), .A2(n4836), .ZN(n4835) );
  NAND2_X1 U6271 ( .A1(n4692), .A2(n5194), .ZN(n5413) );
  NAND2_X1 U6272 ( .A1(n4635), .A2(n5179), .ZN(n5348) );
  NAND2_X1 U6273 ( .A1(n5326), .A2(n5327), .ZN(n4635) );
  NAND2_X1 U6274 ( .A1(n4639), .A2(n4638), .ZN(n9772) );
  NAND2_X1 U6275 ( .A1(n9865), .A2(n10094), .ZN(n4639) );
  NAND2_X1 U6276 ( .A1(n4641), .A2(n4640), .ZN(n9866) );
  NAND2_X1 U6277 ( .A1(n9865), .A2(n10078), .ZN(n4641) );
  NAND3_X1 U6278 ( .A1(n5897), .A2(n4648), .A3(n5898), .ZN(n5919) );
  NAND2_X1 U6279 ( .A1(n4649), .A2(n4637), .ZN(n5948) );
  NAND2_X1 U6280 ( .A1(n4526), .A2(n4647), .ZN(n5953) );
  MUX2_X1 U6281 ( .A(n9912), .B(P1_IR_REG_0__SCAN_IN), .S(n6272), .Z(n9748) );
  NAND2_X1 U6282 ( .A1(n9160), .A2(n4651), .ZN(n4650) );
  NAND2_X1 U6283 ( .A1(n4650), .A2(n4652), .ZN(n9167) );
  NAND2_X1 U6284 ( .A1(n9161), .A2(n9270), .ZN(n4665) );
  INV_X1 U6285 ( .A(n7649), .ZN(n9065) );
  XNOR2_X2 U6286 ( .A(n10001), .B(n6493), .ZN(n7649) );
  NAND2_X1 U6287 ( .A1(n9065), .A2(n7638), .ZN(n6546) );
  NAND2_X1 U6288 ( .A1(n9210), .A2(n4668), .ZN(n4667) );
  NAND2_X1 U6289 ( .A1(n4677), .A2(n4678), .ZN(n4685) );
  NAND2_X1 U6290 ( .A1(n9189), .A2(n4679), .ZN(n4677) );
  NAND2_X1 U6291 ( .A1(n5392), .A2(n4693), .ZN(n4690) );
  NAND2_X1 U6292 ( .A1(n5392), .A2(n5391), .ZN(n4692) );
  NAND2_X2 U6293 ( .A1(n4690), .A2(n4691), .ZN(n5426) );
  AND2_X1 U6294 ( .A1(n5760), .A2(n8699), .ZN(n4697) );
  NAND2_X1 U6295 ( .A1(n5757), .A2(n5759), .ZN(n5758) );
  NAND2_X1 U6296 ( .A1(n8629), .A2(n8630), .ZN(n4699) );
  NAND2_X1 U6297 ( .A1(n5212), .A2(n4705), .ZN(n4704) );
  NAND2_X1 U6298 ( .A1(n4704), .A2(n4703), .ZN(n5224) );
  NAND2_X1 U6299 ( .A1(n5212), .A2(n5211), .ZN(n5481) );
  NAND2_X1 U6300 ( .A1(n6003), .A2(n6002), .ZN(n7257) );
  OAI21_X2 U6301 ( .B1(n8932), .B2(n4747), .A(n4751), .ZN(n4746) );
  INV_X1 U6302 ( .A(n6285), .ZN(n4762) );
  AND2_X2 U6303 ( .A1(n4762), .A2(n4761), .ZN(n8932) );
  MUX2_X1 U6304 ( .A(n7641), .B(P1_REG2_REG_1__SCAN_IN), .S(n7028), .Z(n9356)
         );
  MUX2_X1 U6305 ( .A(n5894), .B(P1_IR_REG_31__SCAN_IN), .S(n5893), .Z(n4763)
         );
  AND2_X2 U6306 ( .A1(n4942), .A2(n5323), .ZN(n5345) );
  INV_X1 U6307 ( .A(n4790), .ZN(n6856) );
  NAND2_X1 U6308 ( .A1(n4789), .A2(n4602), .ZN(n6857) );
  NAND2_X1 U6309 ( .A1(n4790), .A2(n5711), .ZN(n4789) );
  NAND2_X1 U6310 ( .A1(n4795), .A2(n4793), .ZN(n6795) );
  OR2_X1 U6311 ( .A1(n6784), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U6312 ( .A1(n6769), .A2(n4804), .ZN(n6771) );
  OAI211_X1 U6313 ( .C1(n4806), .C2(n6952), .A(n6758), .B(n4805), .ZN(n4804)
         );
  NAND3_X1 U6314 ( .A1(n6754), .A2(n6752), .A3(n4594), .ZN(n4805) );
  NAND3_X1 U6315 ( .A1(n7411), .A2(n4812), .A3(n4807), .ZN(n6739) );
  NAND2_X1 U6316 ( .A1(n5735), .A2(n4814), .ZN(n4815) );
  NAND2_X1 U6317 ( .A1(n5735), .A2(n5268), .ZN(n5788) );
  INV_X1 U6318 ( .A(n4815), .ZN(n5283) );
  NAND2_X1 U6319 ( .A1(n6688), .A2(n6963), .ZN(n7241) );
  AND2_X2 U6320 ( .A1(n4819), .A2(n4818), .ZN(n8612) );
  OR2_X2 U6321 ( .A1(n8585), .A2(n6712), .ZN(n4819) );
  NOR2_X1 U6322 ( .A1(n8114), .A2(n4545), .ZN(n6707) );
  NAND3_X1 U6323 ( .A1(n4822), .A2(n4824), .A3(n4820), .ZN(n8518) );
  NAND3_X1 U6324 ( .A1(n4822), .A2(n4821), .A3(n4820), .ZN(n4826) );
  INV_X1 U6325 ( .A(n4826), .ZN(n8517) );
  NAND2_X1 U6326 ( .A1(n4828), .A2(n4827), .ZN(n7367) );
  NAND2_X1 U6327 ( .A1(n6694), .A2(n4830), .ZN(n4828) );
  NAND2_X1 U6328 ( .A1(n10110), .A2(n4543), .ZN(n4834) );
  NAND2_X1 U6329 ( .A1(n4835), .A2(n6963), .ZN(n7237) );
  INV_X1 U6330 ( .A(n6645), .ZN(n4837) );
  NAND3_X1 U6331 ( .A1(n4847), .A2(n4551), .A3(n6595), .ZN(n4844) );
  INV_X1 U6332 ( .A(n4847), .ZN(n7562) );
  NAND2_X1 U6333 ( .A1(n6606), .A2(n4852), .ZN(n4850) );
  NOR2_X1 U6334 ( .A1(n8590), .A2(n6604), .ZN(n8591) );
  INV_X1 U6335 ( .A(n8601), .ZN(n4852) );
  MUX2_X1 U6336 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10200), .S(n10107), .Z(
        n10112) );
  XNOR2_X2 U6337 ( .A(n4853), .B(n5346), .ZN(n10107) );
  NAND2_X1 U6338 ( .A1(n8136), .A2(n5550), .ZN(n8133) );
  NAND2_X1 U6339 ( .A1(n4859), .A2(n7921), .ZN(n4857) );
  NAND2_X1 U6340 ( .A1(n4866), .A2(n4863), .ZN(n5400) );
  NOR2_X1 U6341 ( .A1(n4871), .A2(n4868), .ZN(n4867) );
  NAND2_X1 U6342 ( .A1(n8756), .A2(n4876), .ZN(n4874) );
  AOI21_X1 U6343 ( .B1(n10117), .B2(n4884), .A(n4880), .ZN(n7854) );
  NAND2_X1 U6344 ( .A1(n5797), .A2(n5270), .ZN(n5272) );
  AOI22_X2 U6345 ( .A1(n8643), .A2(n5695), .B1(n8654), .B2(n8360), .ZN(n8631)
         );
  OAI21_X1 U6346 ( .B1(n7892), .B2(n5099), .A(n5100), .ZN(n6598) );
  NOR2_X1 U6347 ( .A1(n7366), .A2(n7365), .ZN(n7364) );
  NOR2_X1 U6348 ( .A1(n8010), .A2(n6599), .ZN(n8106) );
  NAND2_X1 U6349 ( .A1(n4959), .A2(n4572), .ZN(P2_U3200) );
  INV_X1 U6350 ( .A(n6597), .ZN(n5101) );
  NAND2_X1 U6351 ( .A1(n5568), .A2(n5567), .ZN(n8771) );
  NAND2_X1 U6352 ( .A1(n5400), .A2(n5399), .ZN(n10117) );
  NAND2_X1 U6353 ( .A1(n6734), .A2(n6733), .ZN(n6898) );
  NAND2_X1 U6354 ( .A1(n5338), .A2(n5337), .ZN(n7412) );
  NAND2_X1 U6355 ( .A1(n5130), .A2(n5156), .ZN(n5129) );
  NAND3_X1 U6356 ( .A1(n4898), .A2(n7220), .A3(n4900), .ZN(n7267) );
  NAND2_X1 U6357 ( .A1(n7219), .A2(n8515), .ZN(n4900) );
  INV_X1 U6358 ( .A(n7219), .ZN(n4897) );
  INV_X1 U6359 ( .A(n4898), .ZN(n7266) );
  NOR2_X1 U6360 ( .A1(n7266), .A2(n4899), .ZN(n7221) );
  NAND2_X1 U6361 ( .A1(n7267), .A2(n4898), .ZN(n7268) );
  INV_X1 U6362 ( .A(n4900), .ZN(n4899) );
  NAND2_X1 U6363 ( .A1(n8381), .A2(n4905), .ZN(n4902) );
  NAND2_X1 U6364 ( .A1(n4902), .A2(n4903), .ZN(n8460) );
  NAND2_X1 U6365 ( .A1(n8246), .A2(n4911), .ZN(n4910) );
  OAI211_X1 U6366 ( .C1(n8434), .C2(n4916), .A(n4913), .B(n4603), .ZN(n4914)
         );
  NAND2_X1 U6367 ( .A1(n8280), .A2(n4915), .ZN(n4913) );
  INV_X1 U6368 ( .A(n4914), .ZN(n8327) );
  NAND3_X1 U6369 ( .A1(n8280), .A2(n8434), .A3(n8707), .ZN(n8373) );
  INV_X1 U6370 ( .A(n5307), .ZN(n5727) );
  NAND2_X1 U6371 ( .A1(n7498), .A2(n4538), .ZN(n4919) );
  AND2_X1 U6372 ( .A1(n7827), .A2(n7830), .ZN(n4928) );
  NAND2_X1 U6373 ( .A1(n8229), .A2(n4932), .ZN(n4931) );
  INV_X1 U6374 ( .A(n8208), .ZN(n4940) );
  MUX2_X1 U6375 ( .A(n8909), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6376 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8909), .S(n6678), .Z(n7308) );
  XNOR2_X2 U6377 ( .A(n6709), .B(n6708), .ZN(n8553) );
  AND2_X2 U6378 ( .A1(n4950), .A2(n4949), .ZN(n6709) );
  OR2_X2 U6379 ( .A1(n8545), .A2(n8544), .ZN(n4950) );
  OR2_X1 U6380 ( .A1(n9593), .A2(n9860), .ZN(n4963) );
  NAND2_X1 U6381 ( .A1(n9593), .A2(n4965), .ZN(n9563) );
  NAND2_X1 U6382 ( .A1(n9593), .A2(n9581), .ZN(n9580) );
  NAND3_X1 U6383 ( .A1(n4963), .A2(n4961), .A3(n4960), .ZN(n9557) );
  NOR2_X2 U6384 ( .A1(n7988), .A2(n8977), .ZN(n9740) );
  NAND2_X1 U6385 ( .A1(n9684), .A2(n4550), .ZN(n9623) );
  NAND2_X1 U6386 ( .A1(n7530), .A2(n4973), .ZN(n7841) );
  NAND2_X1 U6387 ( .A1(n4979), .A2(n4978), .ZN(n9972) );
  AOI21_X1 U6388 ( .B1(n7654), .B2(n4981), .A(n4596), .ZN(n4978) );
  NAND2_X1 U6389 ( .A1(n7603), .A2(n4980), .ZN(n4979) );
  NAND2_X1 U6390 ( .A1(n7603), .A2(n7611), .ZN(n4982) );
  NAND2_X1 U6391 ( .A1(n7765), .A2(n4600), .ZN(n6512) );
  NAND2_X1 U6392 ( .A1(n9696), .A2(n4987), .ZN(n4986) );
  NAND2_X1 U6393 ( .A1(n4989), .A2(n4620), .ZN(n6529) );
  OAI21_X2 U6394 ( .B1(n7438), .B2(n9077), .A(n6506), .ZN(n7462) );
  OAI21_X2 U6395 ( .B1(n7392), .B2(n7391), .A(n7389), .ZN(n7438) );
  OAI21_X2 U6396 ( .B1(n9615), .B2(n6531), .A(n6532), .ZN(n9590) );
  NAND2_X1 U6397 ( .A1(n5244), .A2(n5243), .ZN(n4996) );
  OR2_X2 U6398 ( .A1(n6862), .A2(n6861), .ZN(n5000) );
  NAND2_X2 U6399 ( .A1(n5173), .A2(n5001), .ZN(n5176) );
  NAND2_X1 U6400 ( .A1(n5426), .A2(n5006), .ZN(n5005) );
  NAND2_X1 U6401 ( .A1(n6848), .A2(n5014), .ZN(n5013) );
  NAND2_X1 U6402 ( .A1(n5614), .A2(n5252), .ZN(n5029) );
  OR2_X1 U6403 ( .A1(n5614), .A2(n5613), .ZN(n5033) );
  OAI21_X1 U6404 ( .B1(n9645), .B2(n5045), .A(n5042), .ZN(n9619) );
  INV_X1 U6405 ( .A(n9640), .ZN(n5047) );
  OAI21_X1 U6406 ( .B1(n9588), .B2(n5053), .A(n5050), .ZN(n6559) );
  NAND2_X1 U6407 ( .A1(n9588), .A2(n9589), .ZN(n5055) );
  OAI22_X2 U6408 ( .A1(n5058), .A2(n5057), .B1(n7523), .B2(n5056), .ZN(n7762)
         );
  NAND2_X1 U6409 ( .A1(n6546), .A2(n4599), .ZN(n9253) );
  AOI21_X1 U6410 ( .B1(n5061), .B2(n6548), .A(n9254), .ZN(n9118) );
  NAND2_X1 U6411 ( .A1(n9253), .A2(n9251), .ZN(n5061) );
  NAND2_X2 U6412 ( .A1(n7838), .A2(n5062), .ZN(n7984) );
  OAI21_X2 U6413 ( .B1(n8941), .B2(n5067), .A(n5066), .ZN(n5065) );
  INV_X1 U6414 ( .A(n9015), .ZN(n6266) );
  AOI21_X1 U6415 ( .B1(n9015), .B2(n6284), .A(n9013), .ZN(n6285) );
  NAND2_X1 U6416 ( .A1(n7998), .A2(n6188), .ZN(n6205) );
  INV_X1 U6417 ( .A(n6110), .ZN(n5086) );
  INV_X1 U6418 ( .A(n6189), .ZN(n5843) );
  OAI21_X1 U6419 ( .B1(n8560), .B2(n5095), .A(n5094), .ZN(n8568) );
  XNOR2_X1 U6420 ( .A(n6598), .B(n8020), .ZN(n8011) );
  NAND2_X1 U6421 ( .A1(n7409), .A2(n6734), .ZN(n7331) );
  NAND2_X1 U6422 ( .A1(n5111), .A2(n5110), .ZN(n7811) );
  OR2_X1 U6423 ( .A1(n8142), .A2(n5115), .ZN(n5112) );
  NAND2_X1 U6424 ( .A1(n5112), .A2(n5113), .ZN(n8782) );
  NAND2_X1 U6425 ( .A1(n5119), .A2(n5123), .ZN(n5765) );
  NAND2_X1 U6426 ( .A1(n5764), .A2(n5120), .ZN(n5119) );
  NOR2_X1 U6427 ( .A1(n5409), .A2(n5128), .ZN(n5304) );
  NOR2_X2 U6428 ( .A1(n5129), .A2(n5409), .ZN(n5735) );
  NAND2_X1 U6429 ( .A1(n7920), .A2(n4529), .ZN(n5131) );
  NAND2_X1 U6430 ( .A1(n5131), .A2(n5132), .ZN(n5746) );
  OAI21_X1 U6431 ( .B1(n8051), .B2(n5137), .A(n5135), .ZN(n8148) );
  NAND3_X1 U6432 ( .A1(n5142), .A2(n6824), .A3(n5146), .ZN(n5143) );
  NAND2_X1 U6433 ( .A1(n5145), .A2(n5146), .ZN(n8672) );
  AND2_X1 U6434 ( .A1(n9141), .A2(n9140), .ZN(n9074) );
  OR2_X1 U6435 ( .A1(n6688), .A2(n6963), .ZN(n6689) );
  OR2_X1 U6436 ( .A1(n9266), .A2(n6552), .ZN(n9264) );
  XNOR2_X1 U6437 ( .A(n5178), .B(n5174), .ZN(n5327) );
  NAND2_X1 U6438 ( .A1(n8300), .A2(n8435), .ZN(n8403) );
  NAND2_X1 U6439 ( .A1(n7465), .A2(n7464), .ZN(n7463) );
  XNOR2_X1 U6440 ( .A(n8631), .B(n8630), .ZN(n8637) );
  CLKBUF_X1 U6441 ( .A(n6471), .Z(n9378) );
  INV_X1 U6442 ( .A(n8347), .ZN(n5786) );
  OR2_X1 U6443 ( .A1(n7646), .A2(n5918), .ZN(n5963) );
  NAND2_X1 U6444 ( .A1(n6725), .A2(n10094), .ZN(n6579) );
  XNOR2_X1 U6445 ( .A(n5181), .B(n5180), .ZN(n5347) );
  NAND4_X2 U6446 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n9998)
         );
  NAND4_X2 U6447 ( .A1(n5913), .A2(n5912), .A3(n5910), .A4(n5911), .ZN(n6493)
         );
  NAND2_X1 U6448 ( .A1(n8277), .A2(n8276), .ZN(n8280) );
  INV_X1 U6449 ( .A(n6246), .ZN(n5849) );
  BUF_X2 U6450 ( .A(n6493), .Z(n9750) );
  INV_X1 U6451 ( .A(n5919), .ZN(n10001) );
  AND2_X4 U6452 ( .A1(n8223), .A2(n8315), .ZN(n6034) );
  XNOR2_X2 U6453 ( .A(n5892), .B(n5903), .ZN(n9300) );
  NAND2_X2 U6454 ( .A1(n5899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5892) );
  XNOR2_X1 U6455 ( .A(n8642), .B(n8644), .ZN(n8852) );
  XNOR2_X1 U6456 ( .A(n8629), .B(n8630), .ZN(n8846) );
  NAND2_X1 U6457 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  NAND2_X1 U6458 ( .A1(n5351), .A2(n7273), .ZN(n6734) );
  INV_X1 U6459 ( .A(n7570), .ZN(n6983) );
  AND2_X1 U6460 ( .A1(n5332), .A2(n5331), .ZN(n5153) );
  INV_X1 U6461 ( .A(n8596), .ZN(n6680) );
  AND2_X1 U6462 ( .A1(n5489), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5154) );
  AND2_X1 U6463 ( .A1(n5903), .A2(n5902), .ZN(n5155) );
  AND4_X1 U6464 ( .A1(n5267), .A2(n5266), .A3(n5586), .A4(n5306), .ZN(n5156)
         );
  NAND2_X1 U6465 ( .A1(n9750), .A2(n6042), .ZN(n5157) );
  NAND2_X1 U6466 ( .A1(n6721), .A2(n6720), .ZN(n5158) );
  NAND2_X1 U6467 ( .A1(n9998), .A2(n6042), .ZN(n5159) );
  OR2_X1 U6468 ( .A1(n8194), .A2(n8506), .ZN(n5160) );
  NOR2_X1 U6469 ( .A1(n5520), .A2(n5519), .ZN(n5162) );
  NOR2_X1 U6470 ( .A1(n6956), .A2(n8900), .ZN(n5163) );
  AND3_X1 U6471 ( .A1(n5838), .A2(n5861), .A3(n5858), .ZN(n5164) );
  INV_X1 U6472 ( .A(n9734), .ZN(n9757) );
  AND2_X1 U6473 ( .A1(n5501), .A2(n5207), .ZN(n5165) );
  NAND2_X1 U6474 ( .A1(n6264), .A2(n6263), .ZN(n6265) );
  NAND2_X1 U6475 ( .A1(n9656), .A2(n9816), .ZN(n5166) );
  OR2_X1 U6476 ( .A1(n7018), .A2(n5937), .ZN(n5167) );
  INV_X1 U6477 ( .A(n8625), .ZN(n8834) );
  AND2_X1 U6478 ( .A1(n8314), .A2(n8310), .ZN(n5168) );
  AND2_X1 U6479 ( .A1(n8307), .A2(n9798), .ZN(n5169) );
  OR2_X1 U6480 ( .A1(n9636), .A2(n9806), .ZN(n5170) );
  INV_X1 U6481 ( .A(n8701), .ZN(n5755) );
  NAND2_X1 U6482 ( .A1(n6818), .A2(n5755), .ZN(n5759) );
  AND2_X1 U6483 ( .A1(n5914), .A2(n7018), .ZN(n5885) );
  NOR2_X1 U6484 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5872) );
  AND2_X1 U6485 ( .A1(n8446), .A2(n8272), .ZN(n8273) );
  INV_X1 U6486 ( .A(n6685), .ZN(n6637) );
  OR2_X1 U6487 ( .A1(n8843), .A2(n5766), .ZN(n5767) );
  NOR2_X1 U6488 ( .A1(n8680), .A2(n8692), .ZN(n5639) );
  AND2_X1 U6489 ( .A1(n7710), .A2(n7712), .ZN(n6105) );
  AND4_X1 U6490 ( .A1(n5872), .A2(n5871), .A3(n10606), .A4(n5870), .ZN(n5874)
         );
  INV_X1 U6491 ( .A(n5551), .ZN(n5229) );
  AND2_X1 U6492 ( .A1(n5503), .A2(n5501), .ZN(n5209) );
  NAND2_X1 U6493 ( .A1(n8325), .A2(n8664), .ZN(n8326) );
  NAND2_X1 U6494 ( .A1(n7241), .A2(n6689), .ZN(n7136) );
  INV_X1 U6495 ( .A(n8673), .ZN(n8675) );
  NAND2_X1 U6496 ( .A1(n7921), .A2(n7950), .ZN(n8041) );
  INV_X1 U6497 ( .A(n6204), .ZN(n6202) );
  NOR2_X1 U6498 ( .A1(n6318), .A2(n6317), .ZN(n6333) );
  AND2_X1 U6499 ( .A1(n6333), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6347) );
  OR2_X1 U6500 ( .A1(n9021), .A2(n9022), .ZN(n6405) );
  NOR2_X1 U6501 ( .A1(n6195), .A2(n6194), .ZN(n6211) );
  NAND2_X1 U6502 ( .A1(n6513), .A2(n4569), .ZN(n6515) );
  OR2_X1 U6503 ( .A1(n6848), .A2(n5016), .ZN(n6849) );
  NAND2_X1 U6504 ( .A1(n5675), .A2(n5674), .ZN(n5681) );
  INV_X1 U6505 ( .A(n5841), .ZN(n5842) );
  NAND2_X1 U6506 ( .A1(n5502), .A2(n5209), .ZN(n5212) );
  INV_X1 U6507 ( .A(n8351), .ZN(n8328) );
  AND2_X1 U6508 ( .A1(n8456), .A2(n8263), .ZN(n8396) );
  AND2_X1 U6509 ( .A1(n5311), .A2(n8451), .ZN(n5608) );
  AND2_X1 U6510 ( .A1(n8394), .A2(n8271), .ZN(n8446) );
  OR2_X1 U6511 ( .A1(n5594), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5596) );
  INV_X1 U6512 ( .A(n10107), .ZN(n6645) );
  NOR2_X1 U6513 ( .A1(n7905), .A2(n6596), .ZN(n6597) );
  INV_X1 U6514 ( .A(n10100), .ZN(n6720) );
  NAND2_X1 U6515 ( .A1(n5651), .A2(n8409), .ZN(n5663) );
  NAND2_X1 U6516 ( .A1(n5608), .A2(n10441), .ZN(n5617) );
  INV_X1 U6517 ( .A(n6803), .ZN(n5751) );
  INV_X1 U6518 ( .A(n8124), .ZN(n5747) );
  AND2_X1 U6519 ( .A1(n8073), .A2(n8048), .ZN(n7951) );
  AND2_X1 U6520 ( .A1(n8982), .A2(n6359), .ZN(n8923) );
  NAND2_X1 U6521 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(n6292), .ZN(n6318) );
  AND2_X1 U6522 ( .A1(n6409), .A2(n6408), .ZN(n6931) );
  OR2_X1 U6523 ( .A1(n6153), .A2(n6152), .ZN(n6175) );
  NOR2_X1 U6524 ( .A1(n6362), .A2(n6363), .ZN(n6379) );
  NOR2_X1 U6525 ( .A1(n6404), .A2(n6403), .ZN(n9022) );
  AND2_X1 U6526 ( .A1(n9245), .A2(n9237), .ZN(n9628) );
  AND2_X1 U6527 ( .A1(n9190), .A2(n9224), .ZN(n9646) );
  NAND2_X1 U6528 ( .A1(n6518), .A2(n4571), .ZN(n6520) );
  OR2_X1 U6529 ( .A1(n9340), .A2(n9335), .ZN(n9215) );
  NAND2_X1 U6530 ( .A1(n5217), .A2(n5216), .ZN(n5480) );
  NOR2_X1 U6531 ( .A1(n5183), .A2(n5364), .ZN(n5184) );
  INV_X1 U6532 ( .A(SI_3_), .ZN(n10570) );
  XNOR2_X1 U6533 ( .A(n8630), .B(n7421), .ZN(n8333) );
  INV_X1 U6534 ( .A(n7861), .ZN(n10167) );
  INV_X1 U6535 ( .A(n8403), .ZN(n8438) );
  AND2_X1 U6536 ( .A1(n5669), .A2(n5668), .ZN(n8664) );
  AND4_X1 U6537 ( .A1(n5566), .A2(n5565), .A3(n5564), .A4(n5563), .ZN(n8487)
         );
  OR2_X1 U6538 ( .A1(n5343), .A2(n5401), .ZN(n5407) );
  INV_X1 U6539 ( .A(n7378), .ZN(n10095) );
  NAND2_X1 U6540 ( .A1(n5510), .A2(n5509), .ZN(n10176) );
  INV_X1 U6541 ( .A(n10147), .ZN(n7490) );
  INV_X1 U6542 ( .A(n8829), .ZN(n6959) );
  NOR2_X1 U6543 ( .A1(n10196), .A2(n5722), .ZN(n5829) );
  NAND2_X1 U6544 ( .A1(n8038), .A2(n6875), .ZN(n5662) );
  AND2_X1 U6545 ( .A1(n6801), .A2(n8697), .ZN(n8739) );
  INV_X1 U6546 ( .A(n10183), .ZN(n10195) );
  NOR2_X1 U6547 ( .A1(n8983), .A2(n6376), .ZN(n8950) );
  INV_X1 U6548 ( .A(n9041), .ZN(n9033) );
  INV_X1 U6549 ( .A(n9036), .ZN(n9051) );
  OR2_X1 U6550 ( .A1(n6573), .A2(n6469), .ZN(n9753) );
  INV_X1 U6551 ( .A(n9849), .ZN(n10075) );
  XNOR2_X1 U6552 ( .A(n5196), .B(n10365), .ZN(n5425) );
  INV_X1 U6553 ( .A(n8719), .ZN(n8881) );
  AND2_X1 U6554 ( .A1(n7172), .A2(n7171), .ZN(n8482) );
  AND2_X1 U6555 ( .A1(n7166), .A2(n7165), .ZN(n8490) );
  INV_X1 U6556 ( .A(n5766), .ZN(n8646) );
  INV_X1 U6557 ( .A(n8692), .ZN(n8500) );
  INV_X1 U6558 ( .A(n8487), .ZN(n8773) );
  OR2_X1 U6559 ( .A1(n6719), .A2(n6718), .ZN(n10100) );
  INV_X1 U6560 ( .A(n10213), .ZN(n10211) );
  NOR2_X1 U6561 ( .A1(n5163), .A2(n5829), .ZN(n5830) );
  AND2_X1 U6562 ( .A1(n5827), .A2(n5826), .ZN(n10198) );
  AND2_X1 U6563 ( .A1(n6673), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6997) );
  INV_X1 U6564 ( .A(n7978), .ZN(n7067) );
  INV_X1 U6565 ( .A(n6942), .ZN(n6943) );
  NAND2_X1 U6566 ( .A1(n6935), .A2(n6467), .ZN(n6492) );
  OR2_X1 U6567 ( .A1(n6476), .A2(n6466), .ZN(n9046) );
  AND2_X1 U6568 ( .A1(n9753), .A2(n6470), .ZN(n9036) );
  INV_X1 U6569 ( .A(n4511), .ZN(n9719) );
  AND2_X1 U6570 ( .A1(n9753), .A2(n7510), .ZN(n9734) );
  OR2_X1 U6571 ( .A1(n6724), .A2(n6575), .ZN(n10092) );
  OR2_X1 U6572 ( .A1(n6724), .A2(n7507), .ZN(n10076) );
  INV_X1 U6573 ( .A(n9993), .ZN(n9992) );
  INV_X1 U6574 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10457) );
  INV_X1 U6575 ( .A(n8606), .ZN(P2_U3893) );
  NAND2_X1 U6576 ( .A1(n6579), .A2(n6578), .ZN(P1_U3551) );
  MUX2_X1 U6577 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5176), .Z(n5178) );
  INV_X1 U6578 ( .A(SI_1_), .ZN(n5174) );
  AND2_X1 U6579 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5175) );
  NAND2_X1 U6580 ( .A1(n6965), .A2(n5175), .ZN(n5933) );
  AND2_X1 U6581 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6582 ( .A1(n5176), .A2(n5177), .ZN(n5335) );
  NAND2_X1 U6583 ( .A1(n5933), .A2(n5335), .ZN(n5326) );
  NAND2_X1 U6584 ( .A1(n5178), .A2(SI_1_), .ZN(n5179) );
  MUX2_X1 U6585 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5186), .Z(n5181) );
  INV_X1 U6586 ( .A(SI_2_), .ZN(n5180) );
  NAND2_X1 U6587 ( .A1(n5348), .A2(n5347), .ZN(n5363) );
  NAND2_X1 U6588 ( .A1(n5181), .A2(SI_2_), .ZN(n5362) );
  AND2_X1 U6589 ( .A1(n5362), .A2(n5182), .ZN(n5185) );
  INV_X1 U6590 ( .A(n5182), .ZN(n5183) );
  AOI21_X2 U6591 ( .B1(n5363), .B2(n5185), .A(n5184), .ZN(n5377) );
  BUF_X8 U6592 ( .A(n5186), .Z(n6965) );
  MUX2_X1 U6593 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6965), .Z(n5188) );
  INV_X1 U6594 ( .A(SI_4_), .ZN(n5187) );
  NAND2_X1 U6595 ( .A1(n5377), .A2(n5376), .ZN(n5190) );
  NAND2_X1 U6596 ( .A1(n5188), .A2(SI_4_), .ZN(n5189) );
  INV_X1 U6597 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5191) );
  MUX2_X1 U6598 ( .A(n6972), .B(n5191), .S(n6965), .Z(n5192) );
  XNOR2_X2 U6599 ( .A(n5192), .B(SI_5_), .ZN(n5391) );
  INV_X1 U6600 ( .A(n5192), .ZN(n5193) );
  MUX2_X1 U6601 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6965), .Z(n5195) );
  MUX2_X1 U6602 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6965), .Z(n5196) );
  NAND2_X1 U6603 ( .A1(n5196), .A2(SI_7_), .ZN(n5197) );
  INV_X1 U6604 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7009) );
  INV_X1 U6605 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5198) );
  MUX2_X1 U6606 ( .A(n7009), .B(n5198), .S(n6965), .Z(n5199) );
  INV_X1 U6607 ( .A(SI_8_), .ZN(n10632) );
  INV_X1 U6608 ( .A(n5199), .ZN(n5200) );
  NAND2_X1 U6609 ( .A1(n5200), .A2(SI_8_), .ZN(n5201) );
  INV_X1 U6610 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5204) );
  INV_X1 U6611 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5203) );
  MUX2_X1 U6612 ( .A(n5204), .B(n5203), .S(n6965), .Z(n5205) );
  INV_X1 U6613 ( .A(SI_9_), .ZN(n10618) );
  INV_X1 U6614 ( .A(n5205), .ZN(n5206) );
  NAND2_X1 U6615 ( .A1(n5206), .A2(SI_9_), .ZN(n5207) );
  MUX2_X1 U6616 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6965), .Z(n5210) );
  INV_X1 U6617 ( .A(SI_10_), .ZN(n5208) );
  NAND2_X1 U6618 ( .A1(n5210), .A2(SI_10_), .ZN(n5211) );
  INV_X1 U6619 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5213) );
  MUX2_X1 U6620 ( .A(n5213), .B(n10457), .S(n6965), .Z(n5214) );
  INV_X1 U6621 ( .A(SI_11_), .ZN(n10408) );
  INV_X1 U6622 ( .A(n5214), .ZN(n5215) );
  NAND2_X1 U6623 ( .A1(n5215), .A2(SI_11_), .ZN(n5216) );
  MUX2_X1 U6624 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6965), .Z(n5219) );
  INV_X1 U6625 ( .A(SI_12_), .ZN(n5218) );
  MUX2_X1 U6626 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6965), .Z(n5221) );
  MUX2_X1 U6627 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6965), .Z(n5222) );
  XNOR2_X1 U6628 ( .A(n5222), .B(SI_14_), .ZN(n5522) );
  NAND2_X1 U6629 ( .A1(n5222), .A2(SI_14_), .ZN(n5223) );
  NAND2_X1 U6630 ( .A1(n5224), .A2(n5223), .ZN(n5537) );
  MUX2_X1 U6631 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6965), .Z(n5535) );
  INV_X1 U6632 ( .A(SI_15_), .ZN(n5225) );
  NOR2_X1 U6633 ( .A1(n5226), .A2(n5225), .ZN(n5228) );
  NAND2_X1 U6634 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  INV_X1 U6635 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7264) );
  INV_X1 U6636 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10374) );
  MUX2_X1 U6637 ( .A(n7264), .B(n10374), .S(n4637), .Z(n5551) );
  NAND2_X1 U6638 ( .A1(n5229), .A2(SI_16_), .ZN(n5230) );
  INV_X1 U6639 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5232) );
  INV_X1 U6640 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10366) );
  MUX2_X1 U6641 ( .A(n5232), .B(n10366), .S(n6965), .Z(n5233) );
  INV_X1 U6642 ( .A(SI_17_), .ZN(n10568) );
  NAND2_X1 U6643 ( .A1(n5233), .A2(n10568), .ZN(n5236) );
  INV_X1 U6644 ( .A(n5233), .ZN(n5234) );
  NAND2_X1 U6645 ( .A1(n5234), .A2(SI_17_), .ZN(n5235) );
  NAND2_X1 U6646 ( .A1(n5236), .A2(n5235), .ZN(n5569) );
  MUX2_X1 U6647 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4637), .Z(n5238) );
  INV_X1 U6648 ( .A(SI_18_), .ZN(n5237) );
  XNOR2_X1 U6649 ( .A(n5238), .B(n5237), .ZN(n5584) );
  NAND2_X1 U6650 ( .A1(n5238), .A2(SI_18_), .ZN(n5239) );
  INV_X1 U6651 ( .A(n5303), .ZN(n5244) );
  INV_X1 U6652 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7548) );
  INV_X1 U6653 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8342) );
  MUX2_X1 U6654 ( .A(n7548), .B(n8342), .S(n6965), .Z(n5240) );
  INV_X1 U6655 ( .A(SI_19_), .ZN(n10575) );
  NAND2_X1 U6656 ( .A1(n5240), .A2(n10575), .ZN(n5245) );
  INV_X1 U6657 ( .A(n5240), .ZN(n5241) );
  NAND2_X1 U6658 ( .A1(n5241), .A2(SI_19_), .ZN(n5242) );
  NAND2_X1 U6659 ( .A1(n5245), .A2(n5242), .ZN(n5302) );
  INV_X1 U6660 ( .A(n5302), .ZN(n5243) );
  INV_X1 U6661 ( .A(SI_20_), .ZN(n10599) );
  MUX2_X1 U6662 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4637), .Z(n5293) );
  INV_X1 U6663 ( .A(n5293), .ZN(n5246) );
  INV_X1 U6664 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7776) );
  INV_X1 U6665 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7789) );
  MUX2_X1 U6666 ( .A(n7776), .B(n7789), .S(n6965), .Z(n5603) );
  INV_X1 U6667 ( .A(n5603), .ZN(n5247) );
  INV_X1 U6668 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7852) );
  INV_X1 U6669 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10642) );
  MUX2_X1 U6670 ( .A(n7852), .B(n10642), .S(n4637), .Z(n5249) );
  INV_X1 U6671 ( .A(SI_22_), .ZN(n5248) );
  NAND2_X1 U6672 ( .A1(n5249), .A2(n5248), .ZN(n5252) );
  INV_X1 U6673 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6674 ( .A1(n5250), .A2(SI_22_), .ZN(n5251) );
  NAND2_X1 U6675 ( .A1(n5252), .A2(n5251), .ZN(n5613) );
  INV_X1 U6676 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5275) );
  INV_X1 U6677 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6344) );
  MUX2_X1 U6678 ( .A(n5275), .B(n6344), .S(n4637), .Z(n5253) );
  INV_X1 U6679 ( .A(SI_23_), .ZN(n10585) );
  NAND2_X1 U6680 ( .A1(n5253), .A2(n10585), .ZN(n5641) );
  INV_X1 U6681 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U6682 ( .A1(n5254), .A2(SI_23_), .ZN(n5255) );
  AND2_X1 U6683 ( .A1(n5641), .A2(n5255), .ZN(n5256) );
  OR2_X1 U6684 ( .A1(n5257), .A2(n5256), .ZN(n5258) );
  NAND2_X1 U6685 ( .A1(n5643), .A2(n5258), .ZN(n7877) );
  NOR2_X1 U6686 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5263) );
  NOR2_X1 U6687 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5262) );
  NOR2_X1 U6688 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5261) );
  NAND4_X1 U6689 ( .A1(n5264), .A2(n5263), .A3(n5262), .A4(n5261), .ZN(n5265)
         );
  NOR2_X1 U6690 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5267) );
  NOR2_X1 U6691 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5266) );
  INV_X1 U6692 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5306) );
  INV_X1 U6693 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5268) );
  NAND3_X1 U6694 ( .A1(n5792), .A2(n5818), .A3(n5790), .ZN(n5269) );
  INV_X1 U6695 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5270) );
  INV_X1 U6696 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5273) );
  INV_X1 U6697 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6698 ( .A1(n7877), .A2(n6875), .ZN(n5277) );
  OR2_X1 U6699 ( .A1(n6873), .A2(n5275), .ZN(n5276) );
  NOR2_X2 U6700 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5384) );
  NAND2_X1 U6701 ( .A1(n5384), .A2(n5385), .ZN(n5402) );
  INV_X1 U6702 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5447) );
  INV_X1 U6703 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6704 ( .A1(n5475), .A2(n5463), .ZN(n5529) );
  INV_X1 U6705 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5558) );
  INV_X1 U6706 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10452) );
  INV_X1 U6707 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8451) );
  INV_X1 U6708 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10441) );
  OR2_X2 U6709 ( .A1(n5617), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U6710 ( .A1(n5619), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6711 ( .A1(n5631), .A2(n5278), .ZN(n8694) );
  NAND2_X1 U6712 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5279) );
  NOR2_X1 U6713 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5282) );
  NAND2_X1 U6714 ( .A1(n5283), .A2(n5282), .ZN(n8905) );
  INV_X1 U6715 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U6716 ( .A1(n8694), .A2(n5719), .ZN(n5292) );
  INV_X1 U6717 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U6718 ( .A1(n5775), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6719 ( .A1(n5776), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5288) );
  OAI211_X1 U6720 ( .C1(n8871), .C2(n5343), .A(n5289), .B(n5288), .ZN(n5290)
         );
  INV_X1 U6721 ( .A(n5290), .ZN(n5291) );
  XNOR2_X1 U6722 ( .A(n5293), .B(n10599), .ZN(n5294) );
  XNOR2_X1 U6723 ( .A(n5295), .B(n5294), .ZN(n7600) );
  NAND2_X1 U6724 ( .A1(n7600), .A2(n6875), .ZN(n5297) );
  INV_X1 U6725 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7699) );
  OR2_X1 U6726 ( .A1(n6873), .A2(n7699), .ZN(n5296) );
  NOR2_X1 U6727 ( .A1(n5311), .A2(n8451), .ZN(n5298) );
  OR2_X1 U6728 ( .A1(n5608), .A2(n5298), .ZN(n8733) );
  NAND2_X1 U6729 ( .A1(n8733), .A2(n5719), .ZN(n5301) );
  AOI22_X1 U6730 ( .A1(n5775), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5776), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6731 ( .A1(n6876), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5299) );
  INV_X1 U6732 ( .A(n8745), .ZN(n8502) );
  XNOR2_X1 U6733 ( .A(n5303), .B(n5302), .ZN(n7546) );
  NAND2_X1 U6734 ( .A1(n7546), .A2(n6875), .ZN(n5310) );
  INV_X1 U6735 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6736 ( .A1(n5307), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5587) );
  INV_X1 U6737 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5308) );
  INV_X1 U6738 ( .A(n7547), .ZN(n7346) );
  AOI22_X1 U6739 ( .A1(n5591), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7346), .B2(
        n5590), .ZN(n5309) );
  AND2_X1 U6740 ( .A1(n5596), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5312) );
  OR2_X1 U6741 ( .A1(n5312), .A2(n5311), .ZN(n8750) );
  NAND2_X1 U6742 ( .A1(n8750), .A2(n5719), .ZN(n5317) );
  INV_X1 U6743 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8820) );
  OR2_X1 U6744 ( .A1(n6881), .A2(n8820), .ZN(n5314) );
  INV_X1 U6745 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8749) );
  OR2_X1 U6746 ( .A1(n5339), .A2(n8749), .ZN(n5313) );
  AND2_X1 U6747 ( .A1(n5314), .A2(n5313), .ZN(n5316) );
  NAND2_X1 U6748 ( .A1(n6876), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5315) );
  INV_X1 U6749 ( .A(n8759), .ZN(n8728) );
  INV_X1 U6750 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5318) );
  INV_X1 U6751 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U6752 ( .A1(n6876), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5320) );
  INV_X1 U6753 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6634) );
  OR2_X1 U6754 ( .A1(n5339), .A2(n6634), .ZN(n5319) );
  AND2_X1 U6755 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n4637), .ZN(n5325) );
  NAND2_X1 U6756 ( .A1(n6678), .A2(n5325), .ZN(n5330) );
  XNOR2_X1 U6757 ( .A(n5326), .B(n5327), .ZN(n6982) );
  OR2_X1 U6758 ( .A1(n5328), .A2(n6982), .ZN(n5329) );
  INV_X1 U6759 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6582) );
  INV_X1 U6760 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10630) );
  NAND2_X1 U6761 ( .A1(n6876), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5332) );
  INV_X1 U6762 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6683) );
  OR2_X1 U6763 ( .A1(n5339), .A2(n6683), .ZN(n5331) );
  NAND2_X1 U6764 ( .A1(n5176), .A2(SI_0_), .ZN(n5334) );
  INV_X1 U6765 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6766 ( .A1(n5334), .A2(n5333), .ZN(n5336) );
  AND2_X1 U6767 ( .A1(n5336), .A2(n5335), .ZN(n8909) );
  NAND2_X1 U6768 ( .A1(n8516), .A2(n7308), .ZN(n7340) );
  NAND2_X1 U6769 ( .A1(n6897), .A2(n7340), .ZN(n5338) );
  NAND2_X1 U6770 ( .A1(n7271), .A2(n10137), .ZN(n5337) );
  INV_X1 U6771 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7418) );
  OR2_X1 U6772 ( .A1(n5339), .A2(n7418), .ZN(n5341) );
  INV_X1 U6773 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7276) );
  OR2_X1 U6774 ( .A1(n5562), .A2(n7276), .ZN(n5340) );
  INV_X1 U6775 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5342) );
  XNOR2_X1 U6776 ( .A(n5348), .B(n5347), .ZN(n8221) );
  INV_X1 U6777 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8222) );
  OR2_X1 U6778 ( .A1(n6873), .A2(n8222), .ZN(n5349) );
  OAI211_X1 U6779 ( .C1(n6678), .C2(n10107), .A(n5350), .B(n5349), .ZN(n7273)
         );
  NAND2_X1 U6780 ( .A1(n10142), .A2(n8514), .ZN(n6733) );
  NAND2_X1 U6781 ( .A1(n7412), .A2(n6898), .ZN(n5353) );
  NAND2_X1 U6782 ( .A1(n5351), .A2(n10142), .ZN(n5352) );
  NAND2_X1 U6783 ( .A1(n5353), .A2(n5352), .ZN(n7333) );
  NAND2_X1 U6784 ( .A1(n6876), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5359) );
  INV_X1 U6785 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5354) );
  OR2_X1 U6786 ( .A1(n6881), .A2(n5354), .ZN(n5358) );
  INV_X1 U6787 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5355) );
  OR2_X1 U6788 ( .A1(n5562), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6789 ( .A1(n5360), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6790 ( .A1(n5363), .A2(n5362), .ZN(n5365) );
  XNOR2_X1 U6791 ( .A(n5365), .B(n5364), .ZN(n6968) );
  OR2_X1 U6792 ( .A1(n5328), .A2(n6968), .ZN(n5367) );
  OR2_X1 U6793 ( .A1(n6873), .A2(n5020), .ZN(n5366) );
  OAI211_X1 U6794 ( .C1(n6678), .C2(n6963), .A(n5367), .B(n5366), .ZN(n7422)
         );
  NOR2_X1 U6795 ( .A1(n8513), .A2(n7422), .ZN(n5369) );
  NAND2_X1 U6796 ( .A1(n8513), .A2(n7422), .ZN(n5368) );
  NAND2_X1 U6797 ( .A1(n5775), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5375) );
  INV_X1 U6798 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7488) );
  OR2_X1 U6799 ( .A1(n5339), .A2(n7488), .ZN(n5374) );
  AND2_X1 U6800 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5370) );
  NOR2_X1 U6801 ( .A1(n5384), .A2(n5370), .ZN(n7505) );
  OR2_X1 U6802 ( .A1(n5562), .A2(n7505), .ZN(n5373) );
  INV_X1 U6803 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5371) );
  OR2_X1 U6804 ( .A1(n5343), .A2(n5371), .ZN(n5372) );
  XNOR2_X1 U6805 ( .A(n5377), .B(n5376), .ZN(n6970) );
  OR2_X1 U6806 ( .A1(n5328), .A2(n6970), .ZN(n5382) );
  INV_X1 U6807 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6964) );
  OR2_X1 U6808 ( .A1(n6873), .A2(n6964), .ZN(n5381) );
  NAND2_X1 U6809 ( .A1(n5378), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6810 ( .A1(n5590), .A2(n6690), .ZN(n5380) );
  NAND2_X1 U6811 ( .A1(n7554), .A2(n10147), .ZN(n5741) );
  NAND2_X1 U6812 ( .A1(n7666), .A2(n7490), .ZN(n5740) );
  NAND2_X1 U6813 ( .A1(n6876), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5390) );
  INV_X1 U6814 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7670) );
  OR2_X1 U6815 ( .A1(n5339), .A2(n7670), .ZN(n5389) );
  INV_X1 U6816 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5383) );
  OR2_X1 U6817 ( .A1(n6881), .A2(n5383), .ZN(n5388) );
  OR2_X1 U6818 ( .A1(n5385), .A2(n5384), .ZN(n5386) );
  AND2_X1 U6819 ( .A1(n5402), .A2(n5386), .ZN(n7671) );
  OR2_X1 U6820 ( .A1(n5562), .A2(n7671), .ZN(n5387) );
  XNOR2_X1 U6821 ( .A(n5392), .B(n5391), .ZN(n6977) );
  OR2_X1 U6822 ( .A1(n5328), .A2(n6977), .ZN(n5397) );
  OR2_X1 U6823 ( .A1(n6873), .A2(n6972), .ZN(n5396) );
  OR2_X1 U6824 ( .A1(n5393), .A2(n5554), .ZN(n5394) );
  NAND2_X1 U6825 ( .A1(n5590), .A2(n6971), .ZN(n5395) );
  NAND2_X1 U6826 ( .A1(n7693), .A2(n7555), .ZN(n5398) );
  INV_X1 U6827 ( .A(n7555), .ZN(n10151) );
  NAND2_X1 U6828 ( .A1(n10119), .A2(n10151), .ZN(n5399) );
  NAND2_X1 U6829 ( .A1(n5776), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5408) );
  INV_X1 U6830 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6831 ( .A1(n5402), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5403) );
  AND2_X1 U6832 ( .A1(n5416), .A2(n5403), .ZN(n10124) );
  OR2_X1 U6833 ( .A1(n5562), .A2(n10124), .ZN(n5406) );
  INV_X1 U6834 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5404) );
  OR2_X1 U6835 ( .A1(n6881), .A2(n5404), .ZN(n5405) );
  NAND2_X1 U6836 ( .A1(n5409), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5410) );
  MUX2_X1 U6837 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5410), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5411) );
  NAND2_X1 U6838 ( .A1(n5411), .A2(n4562), .ZN(n6979) );
  XNOR2_X1 U6839 ( .A(n5413), .B(n5412), .ZN(n6980) );
  OR2_X1 U6840 ( .A1(n5328), .A2(n6980), .ZN(n5415) );
  INV_X1 U6841 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6981) );
  OR2_X1 U6842 ( .A1(n6873), .A2(n6981), .ZN(n5414) );
  OAI211_X1 U6843 ( .C1(n6678), .C2(n6979), .A(n5415), .B(n5414), .ZN(n10131)
         );
  NAND2_X1 U6844 ( .A1(n6876), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5422) );
  INV_X1 U6845 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7820) );
  OR2_X1 U6846 ( .A1(n5339), .A2(n7820), .ZN(n5421) );
  AND2_X1 U6847 ( .A1(n5416), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5417) );
  NOR2_X1 U6848 ( .A1(n5434), .A2(n5417), .ZN(n7821) );
  OR2_X1 U6849 ( .A1(n5562), .A2(n7821), .ZN(n5420) );
  INV_X1 U6850 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5418) );
  OR2_X1 U6851 ( .A1(n6881), .A2(n5418), .ZN(n5419) );
  NAND4_X1 U6852 ( .A1(n5422), .A2(n5421), .A3(n5420), .A4(n5419), .ZN(n10121)
         );
  NAND2_X1 U6853 ( .A1(n4562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5423) );
  MUX2_X1 U6854 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5423), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5424) );
  AND2_X1 U6855 ( .A1(n5424), .A2(n5442), .ZN(n7570) );
  XNOR2_X1 U6856 ( .A(n5426), .B(n5425), .ZN(n6985) );
  OR2_X1 U6857 ( .A1(n5328), .A2(n6985), .ZN(n5428) );
  INV_X1 U6858 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6984) );
  OR2_X1 U6859 ( .A1(n6873), .A2(n6984), .ZN(n5427) );
  OAI211_X1 U6860 ( .C1(n6678), .C2(n6983), .A(n5428), .B(n5427), .ZN(n7823)
         );
  NAND2_X1 U6861 ( .A1(n6990), .A2(n6875), .ZN(n5433) );
  NAND2_X1 U6862 ( .A1(n5442), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5431) );
  XNOR2_X1 U6863 ( .A(n5431), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7733) );
  AOI22_X1 U6864 ( .A1(n5591), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5590), .B2(
        n7733), .ZN(n5432) );
  NAND2_X1 U6865 ( .A1(n5776), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5440) );
  INV_X1 U6866 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6593) );
  OR2_X1 U6867 ( .A1(n6881), .A2(n6593), .ZN(n5439) );
  NOR2_X1 U6868 ( .A1(n5434), .A2(n10566), .ZN(n5435) );
  OR2_X1 U6869 ( .A1(n5448), .A2(n5435), .ZN(n7859) );
  INV_X1 U6870 ( .A(n7859), .ZN(n7833) );
  OR2_X1 U6871 ( .A1(n5562), .A2(n7833), .ZN(n5438) );
  INV_X1 U6872 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6873 ( .A1(n7861), .A2(n8511), .ZN(n6755) );
  NAND2_X1 U6874 ( .A1(n8028), .A2(n10167), .ZN(n6762) );
  NAND2_X1 U6875 ( .A1(n6755), .A2(n6762), .ZN(n7857) );
  NAND2_X1 U6876 ( .A1(n7854), .A2(n7857), .ZN(n7853) );
  NAND2_X1 U6877 ( .A1(n7861), .A2(n8028), .ZN(n7922) );
  NAND2_X1 U6878 ( .A1(n7853), .A2(n7922), .ZN(n5454) );
  XNOR2_X1 U6879 ( .A(n5441), .B(n5165), .ZN(n7061) );
  NAND2_X1 U6880 ( .A1(n7061), .A2(n6875), .ZN(n5444) );
  NOR2_X1 U6881 ( .A1(n5442), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5458) );
  OR2_X1 U6882 ( .A1(n5458), .A2(n5554), .ZN(n5506) );
  AOI22_X1 U6883 ( .A1(n5591), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5590), .B2(
        n7905), .ZN(n5443) );
  NAND2_X1 U6884 ( .A1(n6876), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5453) );
  INV_X1 U6885 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5445) );
  OR2_X1 U6886 ( .A1(n6881), .A2(n5445), .ZN(n5452) );
  INV_X1 U6887 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5446) );
  OR2_X1 U6888 ( .A1(n5339), .A2(n5446), .ZN(n5451) );
  OR2_X1 U6889 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  AND2_X1 U6890 ( .A1(n5511), .A2(n5449), .ZN(n8027) );
  OR2_X1 U6891 ( .A1(n5562), .A2(n8027), .ZN(n5450) );
  NAND2_X1 U6892 ( .A1(n10171), .A2(n8059), .ZN(n6763) );
  NAND2_X1 U6893 ( .A1(n6759), .A2(n6763), .ZN(n6902) );
  INV_X1 U6894 ( .A(n8059), .ZN(n8510) );
  OR2_X1 U6895 ( .A1(n10171), .A2(n8510), .ZN(n7950) );
  NAND2_X1 U6896 ( .A1(n7101), .A2(n6875), .ZN(n5462) );
  NOR2_X1 U6897 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5457) );
  AND2_X1 U6898 ( .A1(n5458), .A2(n5457), .ZN(n5482) );
  INV_X1 U6899 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6900 ( .A1(n5482), .A2(n5459), .ZN(n5471) );
  OR2_X1 U6901 ( .A1(n5471), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6902 ( .A1(n5460), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5525) );
  XNOR2_X1 U6903 ( .A(n5525), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8532) );
  AOI22_X1 U6904 ( .A1(n5591), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5590), .B2(
        n8532), .ZN(n5461) );
  NAND2_X1 U6905 ( .A1(n6876), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5468) );
  INV_X1 U6906 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8190) );
  OR2_X1 U6907 ( .A1(n6881), .A2(n8190), .ZN(n5467) );
  INV_X1 U6908 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8519) );
  OR2_X1 U6909 ( .A1(n5339), .A2(n8519), .ZN(n5466) );
  OR2_X1 U6910 ( .A1(n5475), .A2(n5463), .ZN(n5464) );
  AND2_X1 U6911 ( .A1(n5464), .A2(n5529), .ZN(n8235) );
  OR2_X1 U6912 ( .A1(n5562), .A2(n8235), .ZN(n5465) );
  NAND4_X1 U6913 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n8506)
         );
  OR2_X1 U6914 ( .A1(n8237), .A2(n8506), .ZN(n6783) );
  XNOR2_X1 U6915 ( .A(n5470), .B(n5469), .ZN(n7094) );
  NAND2_X1 U6916 ( .A1(n7094), .A2(n6875), .ZN(n5474) );
  NAND2_X1 U6917 ( .A1(n5471), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5472) );
  XNOR2_X1 U6918 ( .A(n5472), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8119) );
  AOI22_X1 U6919 ( .A1(n5591), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5590), .B2(
        n8119), .ZN(n5473) );
  NAND2_X1 U6920 ( .A1(n6876), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5479) );
  INV_X1 U6921 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6624) );
  OR2_X1 U6922 ( .A1(n6881), .A2(n6624), .ZN(n5478) );
  INV_X1 U6923 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8129) );
  OR2_X1 U6924 ( .A1(n5339), .A2(n8129), .ZN(n5477) );
  NOR2_X1 U6925 ( .A1(n5475), .A2(n5154), .ZN(n8128) );
  OR2_X1 U6926 ( .A1(n5562), .A2(n8128), .ZN(n5476) );
  NAND4_X1 U6927 ( .A1(n5479), .A2(n5478), .A3(n5477), .A4(n5476), .ZN(n8507)
         );
  OR2_X1 U6928 ( .A1(n10194), .A2(n8507), .ZN(n8182) );
  NOR2_X1 U6929 ( .A1(n6785), .A2(n8182), .ZN(n5498) );
  XNOR2_X1 U6930 ( .A(n5481), .B(n5480), .ZN(n7070) );
  NAND2_X1 U6931 ( .A1(n7070), .A2(n6875), .ZN(n5485) );
  OR2_X1 U6932 ( .A1(n5482), .A2(n5554), .ZN(n5483) );
  AOI22_X1 U6933 ( .A1(n5591), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5590), .B2(
        n8020), .ZN(n5484) );
  NAND2_X1 U6934 ( .A1(n5485), .A2(n5484), .ZN(n8098) );
  NAND2_X1 U6935 ( .A1(n6876), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5493) );
  INV_X1 U6936 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5486) );
  OR2_X1 U6937 ( .A1(n6881), .A2(n5486), .ZN(n5492) );
  INV_X1 U6938 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5487) );
  OR2_X1 U6939 ( .A1(n5339), .A2(n5487), .ZN(n5491) );
  NAND2_X1 U6940 ( .A1(n5513), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5488) );
  AND2_X1 U6941 ( .A1(n5489), .A2(n5488), .ZN(n8096) );
  OR2_X1 U6942 ( .A1(n5562), .A2(n8096), .ZN(n5490) );
  INV_X1 U6943 ( .A(n8127), .ZN(n8508) );
  NAND2_X1 U6944 ( .A1(n8098), .A2(n8508), .ZN(n8123) );
  NAND2_X1 U6945 ( .A1(n10194), .A2(n8507), .ZN(n5494) );
  AND2_X1 U6946 ( .A1(n8123), .A2(n5494), .ZN(n8180) );
  INV_X1 U6947 ( .A(n6785), .ZN(n5495) );
  AND2_X1 U6948 ( .A1(n8180), .A2(n5495), .ZN(n5496) );
  NOR2_X1 U6949 ( .A1(n5498), .A2(n5496), .ZN(n5497) );
  NAND2_X1 U6950 ( .A1(n8098), .A2(n8127), .ZN(n6774) );
  OR2_X1 U6951 ( .A1(n8077), .A2(n5498), .ZN(n5500) );
  INV_X1 U6952 ( .A(n6783), .ZN(n5499) );
  NAND2_X1 U6953 ( .A1(n5502), .A2(n5501), .ZN(n5504) );
  XNOR2_X1 U6954 ( .A(n5504), .B(n5503), .ZN(n7065) );
  NAND2_X1 U6955 ( .A1(n7065), .A2(n6875), .ZN(n5510) );
  INV_X1 U6956 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U6957 ( .A1(n5506), .A2(n5505), .ZN(n5507) );
  NAND2_X1 U6958 ( .A1(n5507), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5508) );
  XNOR2_X1 U6959 ( .A(n5508), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7978) );
  AOI22_X1 U6960 ( .A1(n5591), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5590), .B2(
        n7978), .ZN(n5509) );
  NAND2_X1 U6961 ( .A1(n6876), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5517) );
  OR2_X1 U6962 ( .A1(n6881), .A2(n10208), .ZN(n5516) );
  INV_X1 U6963 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7956) );
  OR2_X1 U6964 ( .A1(n5339), .A2(n7956), .ZN(n5515) );
  NAND2_X1 U6965 ( .A1(n5511), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5512) );
  AND2_X1 U6966 ( .A1(n5513), .A2(n5512), .ZN(n8066) );
  OR2_X1 U6967 ( .A1(n5562), .A2(n8066), .ZN(n5514) );
  NAND4_X1 U6968 ( .A1(n5517), .A2(n5516), .A3(n5515), .A4(n5514), .ZN(n8509)
         );
  OR2_X1 U6969 ( .A1(n10176), .A2(n8509), .ZN(n8042) );
  AND2_X1 U6970 ( .A1(n7950), .A2(n5518), .ZN(n5521) );
  INV_X1 U6971 ( .A(n5518), .ZN(n5520) );
  NAND2_X1 U6972 ( .A1(n10176), .A2(n8509), .ZN(n8076) );
  AND2_X1 U6973 ( .A1(n8076), .A2(n4597), .ZN(n5519) );
  XNOR2_X1 U6974 ( .A(n5523), .B(n5522), .ZN(n7147) );
  NAND2_X1 U6975 ( .A1(n7147), .A2(n6875), .ZN(n5528) );
  INV_X1 U6976 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6977 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  NAND2_X1 U6978 ( .A1(n5526), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5539) );
  XNOR2_X1 U6979 ( .A(n5539), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8549) );
  AOI22_X1 U6980 ( .A1(n5591), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5590), .B2(
        n8549), .ZN(n5527) );
  NAND2_X1 U6981 ( .A1(n6876), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5534) );
  INV_X1 U6982 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8155) );
  OR2_X1 U6983 ( .A1(n6881), .A2(n8155), .ZN(n5533) );
  INV_X1 U6984 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6618) );
  OR2_X1 U6985 ( .A1(n5339), .A2(n6618), .ZN(n5532) );
  NAND2_X1 U6986 ( .A1(n5529), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5530) );
  AND2_X1 U6987 ( .A1(n5544), .A2(n5530), .ZN(n8367) );
  OR2_X1 U6988 ( .A1(n5562), .A2(n8367), .ZN(n5531) );
  NAND4_X1 U6989 ( .A1(n5534), .A2(n5533), .A3(n5532), .A4(n5531), .ZN(n8505)
         );
  INV_X1 U6990 ( .A(n8240), .ZN(n8372) );
  INV_X1 U6991 ( .A(n8505), .ZN(n5749) );
  XNOR2_X1 U6992 ( .A(n5535), .B(SI_15_), .ZN(n5536) );
  XNOR2_X1 U6993 ( .A(n5537), .B(n5536), .ZN(n7210) );
  NAND2_X1 U6994 ( .A1(n7210), .A2(n6875), .ZN(n5543) );
  INV_X1 U6995 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6996 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  NAND2_X1 U6997 ( .A1(n5540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5541) );
  XNOR2_X1 U6998 ( .A(n5541), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6708) );
  AOI22_X1 U6999 ( .A1(n5591), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5590), .B2(
        n6708), .ZN(n5542) );
  NAND2_X1 U7000 ( .A1(n6876), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5549) );
  INV_X1 U7001 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8559) );
  OR2_X1 U7002 ( .A1(n6881), .A2(n8559), .ZN(n5548) );
  INV_X1 U7003 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6614) );
  OR2_X1 U7004 ( .A1(n5339), .A2(n6614), .ZN(n5547) );
  AND2_X1 U7005 ( .A1(n5544), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5545) );
  NOR2_X1 U7006 ( .A1(n5559), .A2(n5545), .ZN(n8489) );
  OR2_X1 U7007 ( .A1(n5562), .A2(n8489), .ZN(n5546) );
  NAND4_X1 U7008 ( .A1(n5549), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(n8504)
         );
  OR2_X1 U7009 ( .A1(n8244), .A2(n8504), .ZN(n5550) );
  NAND2_X1 U7010 ( .A1(n8244), .A2(n8504), .ZN(n8134) );
  XNOR2_X1 U7011 ( .A(n5551), .B(SI_16_), .ZN(n5552) );
  XNOR2_X1 U7012 ( .A(n5553), .B(n5552), .ZN(n7263) );
  NAND2_X1 U7013 ( .A1(n7263), .A2(n6875), .ZN(n5557) );
  OR2_X1 U7014 ( .A1(n5304), .A2(n5554), .ZN(n5555) );
  XNOR2_X1 U7015 ( .A(n5555), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8582) );
  AOI22_X1 U7016 ( .A1(n5591), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5590), .B2(
        n8582), .ZN(n5556) );
  NAND2_X1 U7017 ( .A1(n6876), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5566) );
  INV_X1 U7018 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8171) );
  OR2_X1 U7019 ( .A1(n6881), .A2(n8171), .ZN(n5565) );
  INV_X1 U7020 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8175) );
  OR2_X1 U7021 ( .A1(n5339), .A2(n8175), .ZN(n5564) );
  NOR2_X1 U7022 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  OR2_X1 U7023 ( .A1(n5575), .A2(n5560), .ZN(n8421) );
  INV_X1 U7024 ( .A(n8421), .ZN(n5561) );
  OR2_X1 U7025 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  NAND2_X1 U7026 ( .A1(n8414), .A2(n8487), .ZN(n6728) );
  NAND2_X1 U7027 ( .A1(n6792), .A2(n6728), .ZN(n6907) );
  NAND2_X1 U7028 ( .A1(n8166), .A2(n6907), .ZN(n5568) );
  NAND2_X1 U7029 ( .A1(n8414), .A2(n8773), .ZN(n5567) );
  XNOR2_X1 U7030 ( .A(n5570), .B(n5569), .ZN(n7294) );
  NAND2_X1 U7031 ( .A1(n7294), .A2(n6875), .ZN(n5574) );
  NAND2_X1 U7032 ( .A1(n5571), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5572) );
  XNOR2_X1 U7033 ( .A(n5572), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8597) );
  AOI22_X1 U7034 ( .A1(n5591), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5590), .B2(
        n8597), .ZN(n5573) );
  OR2_X1 U7035 ( .A1(n5575), .A2(n10452), .ZN(n5576) );
  NAND2_X1 U7036 ( .A1(n5594), .A2(n5576), .ZN(n8775) );
  NAND2_X1 U7037 ( .A1(n5719), .A2(n8775), .ZN(n5581) );
  INV_X1 U7038 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6604) );
  OR2_X1 U7039 ( .A1(n6881), .A2(n6604), .ZN(n5580) );
  INV_X1 U7040 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8778) );
  OR2_X1 U7041 ( .A1(n5339), .A2(n8778), .ZN(n5579) );
  INV_X1 U7042 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5577) );
  OR2_X1 U7043 ( .A1(n5343), .A2(n5577), .ZN(n5578) );
  NAND2_X1 U7044 ( .A1(n8830), .A2(n8761), .ZN(n6803) );
  NAND2_X1 U7045 ( .A1(n8771), .A2(n8781), .ZN(n5583) );
  INV_X1 U7046 ( .A(n8761), .ZN(n8503) );
  NAND2_X1 U7047 ( .A1(n8830), .A2(n8503), .ZN(n5582) );
  XNOR2_X1 U7048 ( .A(n5585), .B(n5584), .ZN(n7407) );
  NAND2_X1 U7049 ( .A1(n7407), .A2(n6875), .ZN(n5593) );
  OR2_X1 U7050 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  AND2_X1 U7051 ( .A1(n5589), .A2(n5588), .ZN(n8617) );
  AOI22_X1 U7052 ( .A1(n5591), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5590), .B2(
        n8617), .ZN(n5592) );
  NAND2_X1 U7053 ( .A1(n5594), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7054 ( .A1(n5596), .A2(n5595), .ZN(n8763) );
  NAND2_X1 U7055 ( .A1(n5719), .A2(n8763), .ZN(n5600) );
  INV_X1 U7056 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8765) );
  OR2_X1 U7057 ( .A1(n5339), .A2(n8765), .ZN(n5599) );
  INV_X1 U7058 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8898) );
  OR2_X1 U7059 ( .A1(n5343), .A2(n8898), .ZN(n5598) );
  INV_X1 U7060 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8827) );
  OR2_X1 U7061 ( .A1(n6881), .A2(n8827), .ZN(n5597) );
  NAND4_X1 U7062 ( .A1(n5600), .A2(n5599), .A3(n5598), .A4(n5597), .ZN(n8772)
         );
  AND2_X1 U7063 ( .A1(n8767), .A2(n8772), .ZN(n5602) );
  OR2_X1 U7064 ( .A1(n8767), .A2(n8772), .ZN(n5601) );
  NAND2_X1 U7065 ( .A1(n8892), .A2(n8759), .ZN(n8697) );
  NAND2_X1 U7066 ( .A1(n8444), .A2(n8745), .ZN(n8720) );
  NAND2_X1 U7067 ( .A1(n8699), .A2(n8720), .ZN(n8731) );
  XNOR2_X1 U7068 ( .A(n5603), .B(SI_21_), .ZN(n5604) );
  XNOR2_X1 U7069 ( .A(n5605), .B(n5604), .ZN(n7775) );
  NAND2_X1 U7070 ( .A1(n7775), .A2(n6875), .ZN(n5607) );
  OR2_X1 U7071 ( .A1(n6873), .A2(n7776), .ZN(n5606) );
  OR2_X1 U7072 ( .A1(n5608), .A2(n10441), .ZN(n5609) );
  NAND2_X1 U7073 ( .A1(n5617), .A2(n5609), .ZN(n8718) );
  NAND2_X1 U7074 ( .A1(n8718), .A2(n5719), .ZN(n5612) );
  AOI22_X1 U7075 ( .A1(n5775), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5776), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7076 ( .A1(n6876), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7077 ( .A1(n8719), .A2(n8708), .ZN(n6815) );
  NAND2_X1 U7078 ( .A1(n8701), .A2(n6815), .ZN(n6895) );
  XNOR2_X1 U7079 ( .A(n5614), .B(n5613), .ZN(n7849) );
  NAND2_X1 U7080 ( .A1(n7849), .A2(n6875), .ZN(n5616) );
  OR2_X1 U7081 ( .A1(n6873), .A2(n7852), .ZN(n5615) );
  NAND2_X1 U7082 ( .A1(n5617), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7083 ( .A1(n5619), .A2(n5618), .ZN(n8709) );
  NAND2_X1 U7084 ( .A1(n8709), .A2(n5719), .ZN(n5624) );
  INV_X1 U7085 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U7086 ( .A1(n5775), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7087 ( .A1(n5776), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5620) );
  OAI211_X1 U7088 ( .C1(n8877), .C2(n5343), .A(n5621), .B(n5620), .ZN(n5622)
         );
  INV_X1 U7089 ( .A(n5622), .ZN(n5623) );
  NAND2_X1 U7090 ( .A1(n5643), .A2(n5641), .ZN(n5628) );
  INV_X1 U7091 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7931) );
  INV_X1 U7092 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10418) );
  MUX2_X1 U7093 ( .A(n7931), .B(n10418), .S(n6965), .Z(n5625) );
  INV_X1 U7094 ( .A(SI_24_), .ZN(n10553) );
  NAND2_X1 U7095 ( .A1(n5625), .A2(n10553), .ZN(n5640) );
  INV_X1 U7096 ( .A(n5625), .ZN(n5626) );
  NAND2_X1 U7097 ( .A1(n5626), .A2(SI_24_), .ZN(n5644) );
  AND2_X1 U7098 ( .A1(n5640), .A2(n5644), .ZN(n5627) );
  NAND2_X1 U7099 ( .A1(n7930), .A2(n6875), .ZN(n5630) );
  OR2_X1 U7100 ( .A1(n6873), .A2(n7931), .ZN(n5629) );
  INV_X1 U7101 ( .A(n5651), .ZN(n5633) );
  NAND2_X1 U7102 ( .A1(n5631), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7103 ( .A1(n5633), .A2(n5632), .ZN(n8682) );
  NAND2_X1 U7104 ( .A1(n8682), .A2(n5719), .ZN(n5638) );
  INV_X1 U7105 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U7106 ( .A1(n5775), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7107 ( .A1(n5776), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5634) );
  OAI211_X1 U7108 ( .C1(n8865), .C2(n5343), .A(n5635), .B(n5634), .ZN(n5636)
         );
  INV_X1 U7109 ( .A(n5636), .ZN(n5637) );
  AND2_X1 U7110 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  INV_X1 U7111 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7962) );
  INV_X1 U7112 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10584) );
  MUX2_X1 U7113 ( .A(n7962), .B(n10584), .S(n4637), .Z(n5646) );
  INV_X1 U7114 ( .A(SI_25_), .ZN(n5645) );
  NAND2_X1 U7115 ( .A1(n5646), .A2(n5645), .ZN(n5676) );
  INV_X1 U7116 ( .A(n5646), .ZN(n5647) );
  NAND2_X1 U7117 ( .A1(n5647), .A2(SI_25_), .ZN(n5648) );
  AND2_X1 U7118 ( .A1(n5676), .A2(n5648), .ZN(n5673) );
  NAND2_X1 U7119 ( .A1(n7961), .A2(n6875), .ZN(n5650) );
  OR2_X1 U7120 ( .A1(n6873), .A2(n7962), .ZN(n5649) );
  INV_X1 U7121 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8409) );
  OR2_X1 U7122 ( .A1(n5651), .A2(n8409), .ZN(n5652) );
  NAND2_X1 U7123 ( .A1(n5663), .A2(n5652), .ZN(n8666) );
  INV_X1 U7124 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8859) );
  NAND2_X1 U7125 ( .A1(n5775), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7126 ( .A1(n5776), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5653) );
  OAI211_X1 U7127 ( .C1(n8859), .C2(n5343), .A(n5654), .B(n5653), .ZN(n5655)
         );
  NAND2_X1 U7128 ( .A1(n8860), .A2(n8653), .ZN(n6833) );
  INV_X1 U7129 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8039) );
  INV_X1 U7130 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10424) );
  MUX2_X1 U7131 ( .A(n8039), .B(n10424), .S(n6965), .Z(n5657) );
  INV_X1 U7132 ( .A(SI_26_), .ZN(n10421) );
  NAND2_X1 U7133 ( .A1(n5657), .A2(n10421), .ZN(n5678) );
  INV_X1 U7134 ( .A(n5657), .ZN(n5658) );
  NAND2_X1 U7135 ( .A1(n5658), .A2(SI_26_), .ZN(n5659) );
  NAND2_X1 U7136 ( .A1(n5678), .A2(n5659), .ZN(n5677) );
  INV_X1 U7137 ( .A(n5677), .ZN(n5672) );
  OR2_X1 U7138 ( .A1(n6873), .A2(n8039), .ZN(n5661) );
  NAND2_X1 U7139 ( .A1(n5663), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7140 ( .A1(n5687), .A2(n5664), .ZN(n8657) );
  NAND2_X1 U7141 ( .A1(n8657), .A2(n5719), .ZN(n5669) );
  INV_X1 U7142 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U7143 ( .A1(n5775), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7144 ( .A1(n5776), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5665) );
  OAI211_X1 U7145 ( .C1(n8854), .C2(n5343), .A(n5666), .B(n5665), .ZN(n5667)
         );
  INV_X1 U7146 ( .A(n5667), .ZN(n5668) );
  NAND2_X1 U7147 ( .A1(n8856), .A2(n8664), .ZN(n5671) );
  AND2_X1 U7148 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  OR2_X1 U7149 ( .A1(n5677), .A2(n5676), .ZN(n5679) );
  AND2_X1 U7150 ( .A1(n5679), .A2(n5678), .ZN(n5680) );
  INV_X1 U7151 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8320) );
  INV_X1 U7152 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10617) );
  MUX2_X1 U7153 ( .A(n8320), .B(n10617), .S(n6965), .Z(n5682) );
  INV_X1 U7154 ( .A(SI_27_), .ZN(n10431) );
  NAND2_X1 U7155 ( .A1(n5682), .A2(n10431), .ZN(n5698) );
  INV_X1 U7156 ( .A(n5682), .ZN(n5683) );
  NAND2_X1 U7157 ( .A1(n5683), .A2(SI_27_), .ZN(n5684) );
  AND2_X1 U7158 ( .A1(n5698), .A2(n5684), .ZN(n5696) );
  XNOR2_X1 U7159 ( .A(n5697), .B(n5696), .ZN(n8220) );
  OR2_X1 U7160 ( .A1(n6873), .A2(n8320), .ZN(n5685) );
  INV_X1 U7161 ( .A(n5704), .ZN(n5689) );
  NAND2_X1 U7162 ( .A1(n5687), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7163 ( .A1(n8648), .A2(n5719), .ZN(n5694) );
  INV_X1 U7164 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U7165 ( .A1(n5776), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7166 ( .A1(n5775), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5690) );
  OAI211_X1 U7167 ( .C1(n5343), .C2(n8848), .A(n5691), .B(n5690), .ZN(n5692)
         );
  INV_X1 U7168 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U7169 ( .A1(n8849), .A2(n8633), .ZN(n5695) );
  INV_X2 U7170 ( .A(n8633), .ZN(n8654) );
  INV_X1 U7171 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8102) );
  INV_X1 U7172 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10569) );
  MUX2_X1 U7173 ( .A(n8102), .B(n10569), .S(n4637), .Z(n5699) );
  INV_X1 U7174 ( .A(SI_28_), .ZN(n10420) );
  NAND2_X1 U7175 ( .A1(n5699), .A2(n10420), .ZN(n5715) );
  INV_X1 U7176 ( .A(n5699), .ZN(n5700) );
  NAND2_X1 U7177 ( .A1(n5700), .A2(SI_28_), .ZN(n5701) );
  AND2_X1 U7178 ( .A1(n5715), .A2(n5701), .ZN(n5713) );
  NAND2_X1 U7179 ( .A1(n8101), .A2(n6875), .ZN(n5703) );
  OR2_X1 U7180 ( .A1(n6873), .A2(n8102), .ZN(n5702) );
  INV_X1 U7181 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8335) );
  NOR2_X1 U7182 ( .A1(n5704), .A2(n8335), .ZN(n5705) );
  NAND2_X1 U7183 ( .A1(n8639), .A2(n5719), .ZN(n5710) );
  INV_X1 U7184 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U7185 ( .A1(n5776), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U7186 ( .A1(n5775), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5706) );
  OAI211_X1 U7187 ( .C1(n8842), .C2(n5343), .A(n5707), .B(n5706), .ZN(n5708)
         );
  INV_X1 U7188 ( .A(n5708), .ZN(n5709) );
  NAND2_X1 U7189 ( .A1(n5711), .A2(n5766), .ZN(n5712) );
  MUX2_X1 U7190 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6965), .Z(n6847) );
  INV_X1 U7191 ( .A(SI_29_), .ZN(n5717) );
  INV_X1 U7192 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8317) );
  OR2_X1 U7193 ( .A1(n6873), .A2(n8317), .ZN(n5718) );
  NAND2_X1 U7194 ( .A1(n8620), .A2(n5719), .ZN(n6884) );
  INV_X1 U7195 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U7196 ( .A1(n5776), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7197 ( .A1(n5775), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5720) );
  OAI211_X1 U7198 ( .C1(n5722), .C2(n5343), .A(n5721), .B(n5720), .ZN(n5723)
         );
  INV_X1 U7199 ( .A(n5723), .ZN(n5724) );
  NAND2_X1 U7200 ( .A1(n5828), .A2(n8499), .ZN(n6854) );
  XNOR2_X1 U7201 ( .A(n5725), .B(n6916), .ZN(n5785) );
  NOR2_X1 U7202 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5726) );
  INV_X1 U7203 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7204 ( .A1(n5730), .A2(n5728), .ZN(n5733) );
  NAND2_X1 U7205 ( .A1(n5733), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5729) );
  INV_X1 U7206 ( .A(n5730), .ZN(n5731) );
  NAND2_X1 U7207 ( .A1(n5731), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5732) );
  INV_X1 U7208 ( .A(n7700), .ZN(n6946) );
  NAND2_X1 U7209 ( .A1(n7175), .A2(n6946), .ZN(n5738) );
  INV_X1 U7210 ( .A(n5735), .ZN(n5736) );
  NAND2_X1 U7211 ( .A1(n5736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5737) );
  XNOR2_X1 U7212 ( .A(n5737), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6945) );
  NAND2_X1 U7213 ( .A1(n7346), .A2(n6945), .ZN(n5820) );
  NAND2_X1 U7214 ( .A1(n5738), .A2(n5820), .ZN(n10123) );
  NAND2_X1 U7215 ( .A1(n7500), .A2(n7422), .ZN(n6747) );
  NAND2_X1 U7216 ( .A1(n7620), .A2(n8513), .ZN(n6741) );
  NAND2_X1 U7217 ( .A1(n7331), .A2(n7332), .ZN(n7480) );
  NAND2_X1 U7218 ( .A1(n7480), .A2(n6747), .ZN(n5742) );
  NAND2_X1 U7219 ( .A1(n5741), .A2(n5740), .ZN(n7485) );
  NAND2_X1 U7220 ( .A1(n5742), .A2(n7485), .ZN(n7478) );
  NAND2_X1 U7221 ( .A1(n7554), .A2(n7490), .ZN(n6742) );
  NAND2_X1 U7222 ( .A1(n7555), .A2(n10119), .ZN(n10125) );
  NAND2_X1 U7223 ( .A1(n10157), .A2(n8512), .ZN(n6751) );
  NOR2_X1 U7224 ( .A1(n7555), .A2(n10119), .ZN(n10126) );
  NAND2_X1 U7225 ( .A1(n6749), .A2(n10126), .ZN(n5743) );
  INV_X1 U7226 ( .A(n8512), .ZN(n7805) );
  NAND2_X1 U7227 ( .A1(n7805), .A2(n10131), .ZN(n6753) );
  AND2_X1 U7228 ( .A1(n5743), .A2(n6753), .ZN(n6744) );
  NAND2_X1 U7229 ( .A1(n7830), .A2(n7823), .ZN(n6761) );
  INV_X1 U7230 ( .A(n7823), .ZN(n10161) );
  NAND2_X1 U7231 ( .A1(n10161), .A2(n10121), .ZN(n7856) );
  NAND2_X1 U7232 ( .A1(n6761), .A2(n7856), .ZN(n7814) );
  AND2_X1 U7233 ( .A1(n6755), .A2(n7856), .ZN(n6760) );
  NAND2_X1 U7234 ( .A1(n7811), .A2(n6760), .ZN(n5744) );
  NAND2_X1 U7235 ( .A1(n5744), .A2(n6762), .ZN(n7920) );
  NAND2_X1 U7236 ( .A1(n10176), .A2(n8024), .ZN(n8048) );
  NAND2_X1 U7237 ( .A1(n5746), .A2(n8077), .ZN(n8051) );
  XNOR2_X1 U7238 ( .A(n10194), .B(n8232), .ZN(n8124) );
  OR2_X1 U7239 ( .A1(n10194), .A2(n8232), .ZN(n5748) );
  INV_X1 U7240 ( .A(n8506), .ZN(n8226) );
  INV_X1 U7241 ( .A(n8237), .ZN(n8194) );
  OR2_X1 U7242 ( .A1(n8240), .A2(n5749), .ZN(n6788) );
  NAND2_X1 U7243 ( .A1(n8148), .A2(n6788), .ZN(n5750) );
  NAND2_X1 U7244 ( .A1(n8240), .A2(n5749), .ZN(n6787) );
  NAND2_X1 U7245 ( .A1(n5750), .A2(n6787), .ZN(n8142) );
  INV_X1 U7246 ( .A(n8504), .ZN(n8419) );
  AND2_X1 U7247 ( .A1(n8244), .A2(n8419), .ZN(n6790) );
  OR2_X1 U7248 ( .A1(n8244), .A2(n8419), .ZN(n6791) );
  INV_X1 U7249 ( .A(n8782), .ZN(n5753) );
  INV_X1 U7250 ( .A(n8781), .ZN(n5752) );
  AOI21_X1 U7251 ( .B1(n5753), .B2(n5752), .A(n5751), .ZN(n8754) );
  INV_X1 U7252 ( .A(n8772), .ZN(n8744) );
  NAND2_X1 U7253 ( .A1(n8767), .A2(n8744), .ZN(n6804) );
  NAND2_X1 U7254 ( .A1(n8754), .A2(n8755), .ZN(n8753) );
  INV_X1 U7255 ( .A(n6801), .ZN(n5754) );
  AND2_X1 U7256 ( .A1(n6815), .A2(n8720), .ZN(n8700) );
  AND2_X1 U7257 ( .A1(n8700), .A2(n6818), .ZN(n5756) );
  INV_X1 U7258 ( .A(n5760), .ZN(n6819) );
  NAND2_X1 U7259 ( .A1(n8872), .A2(n8707), .ZN(n6823) );
  AND2_X1 U7260 ( .A1(n8685), .A2(n6823), .ZN(n5763) );
  INV_X1 U7261 ( .A(n6823), .ZN(n6893) );
  AND2_X1 U7262 ( .A1(n8805), .A2(n8677), .ZN(n6894) );
  INV_X1 U7263 ( .A(n6894), .ZN(n6827) );
  NAND2_X1 U7264 ( .A1(n8668), .A2(n6833), .ZN(n5764) );
  XNOR2_X2 U7265 ( .A(n6836), .B(n8645), .ZN(n8656) );
  OR2_X2 U7266 ( .A1(n8849), .A2(n8654), .ZN(n6842) );
  NAND2_X1 U7267 ( .A1(n5765), .A2(n6842), .ZN(n8629) );
  AND2_X1 U7268 ( .A1(n7175), .A2(n7700), .ZN(n7347) );
  AND2_X1 U7269 ( .A1(n7547), .A2(n6945), .ZN(n5768) );
  NAND2_X1 U7270 ( .A1(n7347), .A2(n5768), .ZN(n7223) );
  INV_X1 U7271 ( .A(n6945), .ZN(n7850) );
  NAND2_X1 U7272 ( .A1(n4809), .A2(n7850), .ZN(n10183) );
  INV_X1 U7273 ( .A(n5768), .ZN(n5769) );
  NAND2_X1 U7274 ( .A1(n7216), .A2(n5769), .ZN(n5770) );
  AND2_X1 U7275 ( .A1(n10183), .A2(n5770), .ZN(n5771) );
  NAND2_X1 U7276 ( .A1(n7223), .A2(n5771), .ZN(n7817) );
  INV_X1 U7277 ( .A(n5772), .ZN(n6672) );
  NAND2_X1 U7278 ( .A1(n6672), .A2(n6925), .ZN(n6718) );
  NAND2_X1 U7279 ( .A1(n6678), .A2(n6718), .ZN(n7224) );
  INV_X1 U7280 ( .A(n7224), .ZN(n5774) );
  NAND2_X2 U7281 ( .A1(n7175), .A2(n6945), .ZN(n6948) );
  INV_X2 U7282 ( .A(n6948), .ZN(n6952) );
  INV_X1 U7283 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7284 ( .A1(n5775), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7285 ( .A1(n5776), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5777) );
  OAI211_X1 U7286 ( .C1(n5779), .C2(n5343), .A(n5778), .B(n5777), .ZN(n5780)
         );
  INV_X1 U7287 ( .A(n5780), .ZN(n5781) );
  NAND2_X1 U7288 ( .A1(n6884), .A2(n5781), .ZN(n8498) );
  NAND2_X1 U7289 ( .A1(n7224), .A2(n6952), .ZN(n8760) );
  AND2_X1 U7290 ( .A1(n6678), .A2(P2_B_REG_SCAN_IN), .ZN(n5782) );
  NOR2_X1 U7291 ( .A1(n8760), .A2(n5782), .ZN(n8621) );
  AOI22_X1 U7292 ( .A1(n8646), .A2(n10118), .B1(n8498), .B2(n8621), .ZN(n5783)
         );
  OAI21_X1 U7293 ( .B1(n8347), .B2(n7817), .A(n5783), .ZN(n5784) );
  NAND2_X1 U7294 ( .A1(n7700), .A2(n7346), .ZN(n5823) );
  NOR2_X1 U7295 ( .A1(n5823), .A2(n6945), .ZN(n10181) );
  INV_X1 U7296 ( .A(n10181), .ZN(n10162) );
  NAND2_X1 U7297 ( .A1(n8350), .A2(n5787), .ZN(n6955) );
  NAND2_X1 U7298 ( .A1(n5788), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7299 ( .A1(n5817), .A2(n5818), .ZN(n5789) );
  NAND2_X1 U7300 ( .A1(n5789), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7301 ( .A1(n5793), .A2(n5792), .ZN(n5795) );
  NAND2_X1 U7302 ( .A1(n5795), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5791) );
  OR2_X1 U7303 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  XNOR2_X1 U7304 ( .A(n7932), .B(P2_B_REG_SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7305 ( .A1(n7963), .A2(n5796), .ZN(n5800) );
  INV_X1 U7306 ( .A(n5797), .ZN(n5798) );
  NAND2_X1 U7307 ( .A1(n5798), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5799) );
  XNOR2_X1 U7308 ( .A(n5799), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5801) );
  OR2_X1 U7309 ( .A1(n5803), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5802) );
  INV_X1 U7310 ( .A(n5801), .ZN(n8040) );
  NAND2_X1 U7311 ( .A1(n7963), .A2(n8040), .ZN(n6995) );
  AND2_X1 U7312 ( .A1(n5802), .A2(n6995), .ZN(n6949) );
  NAND2_X1 U7313 ( .A1(n7932), .A2(n8040), .ZN(n6992) );
  INV_X1 U7314 ( .A(n7215), .ZN(n5824) );
  NOR2_X1 U7315 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5807) );
  NOR4_X1 U7316 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5806) );
  NOR4_X1 U7317 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5805) );
  NOR4_X1 U7318 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5804) );
  NAND4_X1 U7319 ( .A1(n5807), .A2(n5806), .A3(n5805), .A4(n5804), .ZN(n5813)
         );
  NOR4_X1 U7320 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5811) );
  NOR4_X1 U7321 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5810) );
  NOR4_X1 U7322 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5809) );
  NOR4_X1 U7323 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5808) );
  NAND4_X1 U7324 ( .A1(n5811), .A2(n5810), .A3(n5809), .A4(n5808), .ZN(n5812)
         );
  NOR2_X1 U7325 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  OR2_X1 U7326 ( .A1(n5803), .A2(n5814), .ZN(n7151) );
  INV_X1 U7327 ( .A(n7963), .ZN(n5816) );
  NOR2_X1 U7328 ( .A1(n7932), .A2(n8040), .ZN(n5815) );
  NAND2_X1 U7329 ( .A1(n5816), .A2(n5815), .ZN(n7176) );
  XNOR2_X1 U7330 ( .A(n5817), .B(n5818), .ZN(n6673) );
  AND2_X1 U7331 ( .A1(n7176), .A2(n6997), .ZN(n5819) );
  NAND2_X1 U7332 ( .A1(n7151), .A2(n5819), .ZN(n6953) );
  NOR2_X1 U7333 ( .A1(n7303), .A2(n6953), .ZN(n7226) );
  NOR2_X1 U7334 ( .A1(n7175), .A2(n7700), .ZN(n7213) );
  INV_X1 U7335 ( .A(n5820), .ZN(n5821) );
  NAND2_X1 U7336 ( .A1(n7213), .A2(n5821), .ZN(n7167) );
  AND2_X1 U7337 ( .A1(n6948), .A2(n10183), .ZN(n5822) );
  NAND2_X1 U7338 ( .A1(n7167), .A2(n5822), .ZN(n7169) );
  NAND2_X1 U7339 ( .A1(n10195), .A2(n5823), .ZN(n8679) );
  NAND2_X1 U7340 ( .A1(n7169), .A2(n8679), .ZN(n7155) );
  NAND2_X1 U7341 ( .A1(n7226), .A2(n7155), .ZN(n5827) );
  NAND2_X1 U7342 ( .A1(n5824), .A2(n6949), .ZN(n7157) );
  NOR2_X1 U7343 ( .A1(n7157), .A2(n6953), .ZN(n7173) );
  NAND2_X1 U7344 ( .A1(n7167), .A2(n7223), .ZN(n5825) );
  NAND2_X1 U7345 ( .A1(n7173), .A2(n5825), .ZN(n5826) );
  INV_X2 U7346 ( .A(n10198), .ZN(n10196) );
  NAND2_X1 U7347 ( .A1(n6955), .A2(n10196), .ZN(n5831) );
  INV_X1 U7348 ( .A(n5828), .ZN(n6956) );
  OR2_X1 U7349 ( .A1(n10198), .A2(n10183), .ZN(n8900) );
  NAND2_X1 U7350 ( .A1(n5831), .A2(n5830), .ZN(P2_U3456) );
  NAND2_X1 U7351 ( .A1(n6052), .A2(n5865), .ZN(n6071) );
  INV_X1 U7352 ( .A(n6071), .ZN(n5835) );
  NAND2_X1 U7353 ( .A1(n5835), .A2(n5834), .ZN(n6110) );
  INV_X2 U7354 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6168) );
  INV_X1 U7355 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7356 ( .A1(n6168), .A2(n5859), .ZN(n5836) );
  NAND3_X1 U7357 ( .A1(n6189), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7358 ( .A1(n5837), .A2(n6206), .ZN(n6246) );
  INV_X2 U7359 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7360 ( .A1(n5849), .A2(n6248), .ZN(n6267) );
  INV_X1 U7361 ( .A(n6267), .ZN(n5838) );
  INV_X2 U7362 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7363 ( .A1(n5861), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U7364 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_19__SCAN_IN), .ZN(
        n5839) );
  OAI21_X1 U7365 ( .B1(n6267), .B2(n5840), .A(n5839), .ZN(n5841) );
  AOI21_X1 U7366 ( .B1(n5843), .B2(n5164), .A(n5842), .ZN(n5844) );
  INV_X1 U7367 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6089) );
  AND4_X1 U7368 ( .A1(n6248), .A2(n5859), .A3(n6089), .A4(n5858), .ZN(n5848)
         );
  INV_X1 U7369 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5862) );
  INV_X1 U7370 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5870) );
  AND4_X1 U7371 ( .A1(n5862), .A2(n6168), .A3(n5870), .A4(n5861), .ZN(n5847)
         );
  NOR2_X1 U7372 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5846) );
  AND4_X1 U7373 ( .A1(n5849), .A2(n5848), .A3(n5847), .A4(n5846), .ZN(n5850)
         );
  NAND2_X1 U7374 ( .A1(n5850), .A2(n6052), .ZN(n5852) );
  NAND2_X1 U7375 ( .A1(n5852), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5851) );
  XNOR2_X1 U7376 ( .A(n5851), .B(n10606), .ZN(n9219) );
  NAND2_X1 U7377 ( .A1(n6286), .A2(n9219), .ZN(n6465) );
  INV_X1 U7378 ( .A(n5852), .ZN(n5853) );
  NAND2_X1 U7379 ( .A1(n5853), .A2(n10606), .ZN(n5854) );
  NAND2_X1 U7380 ( .A1(n9249), .A2(n9219), .ZN(n5914) );
  NAND2_X1 U7381 ( .A1(n6465), .A2(n5914), .ZN(n5857) );
  NAND2_X1 U7382 ( .A1(n5855), .A2(n5868), .ZN(n5856) );
  NAND2_X1 U7383 ( .A1(n5856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6445) );
  XNOR2_X1 U7384 ( .A(n6445), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9335) );
  NAND2_X1 U7385 ( .A1(n5857), .A2(n6542), .ZN(n5884) );
  NAND4_X1 U7386 ( .A1(n5860), .A2(n5859), .A3(n6089), .A4(n5858), .ZN(n5864)
         );
  NAND4_X1 U7387 ( .A1(n6248), .A2(n6168), .A3(n5862), .A4(n5861), .ZN(n5863)
         );
  NOR2_X1 U7388 ( .A1(n5864), .A2(n5863), .ZN(n5876) );
  INV_X1 U7389 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5866) );
  NAND4_X1 U7390 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(n5869)
         );
  NOR2_X1 U7391 ( .A1(n6246), .A2(n5869), .ZN(n5875) );
  NOR2_X1 U7392 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5871) );
  INV_X1 U7393 ( .A(n5951), .ZN(n5873) );
  NAND4_X1 U7394 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n5886)
         );
  INV_X1 U7396 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7397 ( .A1(n5880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5882) );
  INV_X1 U7398 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U7399 ( .A(n5882), .B(n5881), .ZN(n7934) );
  NOR2_X1 U7400 ( .A1(n7982), .A2(n7934), .ZN(n5883) );
  NAND2_X1 U7401 ( .A1(n5884), .A2(n7018), .ZN(n5918) );
  INV_X1 U7402 ( .A(n5886), .ZN(n5889) );
  NOR2_X1 U7403 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5887) );
  NAND2_X1 U7404 ( .A1(n5889), .A2(n5888), .ZN(n5899) );
  NAND2_X1 U7405 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5890) );
  NAND2_X1 U7406 ( .A1(n5892), .A2(n5890), .ZN(n5891) );
  INV_X1 U7407 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7408 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5894) );
  INV_X1 U7409 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5893) );
  INV_X1 U7410 ( .A(n5895), .ZN(n5896) );
  OR2_X1 U7411 ( .A1(n5948), .A2(n6982), .ZN(n5898) );
  INV_X1 U7412 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6966) );
  OR2_X1 U7413 ( .A1(n6190), .A2(n6966), .ZN(n5897) );
  NAND2_X1 U7414 ( .A1(n5970), .A2(n5919), .ZN(n5916) );
  INV_X1 U7415 ( .A(n5899), .ZN(n5901) );
  INV_X1 U7416 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7417 ( .A1(n5901), .A2(n5900), .ZN(n5906) );
  INV_X1 U7418 ( .A(n5906), .ZN(n5904) );
  INV_X1 U7419 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7420 ( .A1(n5904), .A2(n5155), .ZN(n9906) );
  XNOR2_X2 U7421 ( .A(n5905), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5909) );
  OAI21_X2 U7422 ( .B1(n5906), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7423 ( .A1(n6478), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7424 ( .A1(n5991), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5912) );
  INV_X1 U7425 ( .A(n5908), .ZN(n8315) );
  NAND2_X1 U7426 ( .A1(n4516), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5911) );
  INV_X1 U7427 ( .A(n5914), .ZN(n7517) );
  AND2_X4 U7428 ( .A1(n7517), .A2(n7018), .ZN(n6440) );
  NAND2_X1 U7429 ( .A1(n6493), .A2(n6440), .ZN(n5915) );
  INV_X1 U7430 ( .A(n5924), .ZN(n5921) );
  NAND2_X1 U7431 ( .A1(n5919), .A2(n6440), .ZN(n5920) );
  NAND2_X1 U7432 ( .A1(n5921), .A2(n5922), .ZN(n5925) );
  INV_X1 U7433 ( .A(n5922), .ZN(n5923) );
  NAND2_X1 U7434 ( .A1(n5924), .A2(n5923), .ZN(n5947) );
  NAND2_X1 U7435 ( .A1(n5925), .A2(n5947), .ZN(n7107) );
  NAND2_X1 U7436 ( .A1(n5991), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7437 ( .A1(n6478), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7438 ( .A1(n5926), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7439 ( .A1(n9998), .A2(n6440), .ZN(n5936) );
  INV_X1 U7440 ( .A(SI_0_), .ZN(n5932) );
  INV_X1 U7441 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5931) );
  OAI21_X1 U7442 ( .B1(n5176), .B2(n5932), .A(n5931), .ZN(n5934) );
  AND2_X1 U7443 ( .A1(n5934), .A2(n5933), .ZN(n9912) );
  NAND2_X1 U7444 ( .A1(n5970), .A2(n9748), .ZN(n5935) );
  NAND2_X1 U7445 ( .A1(n5936), .A2(n5935), .ZN(n5944) );
  INV_X1 U7446 ( .A(n5944), .ZN(n5938) );
  INV_X1 U7447 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7448 ( .A1(n5938), .A2(n5167), .ZN(n7104) );
  INV_X1 U7449 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5939) );
  NOR2_X1 U7450 ( .A1(n7018), .A2(n5939), .ZN(n5940) );
  NOR2_X1 U7451 ( .A1(n5941), .A2(n5940), .ZN(n5942) );
  NAND2_X1 U7452 ( .A1(n5159), .A2(n5942), .ZN(n7103) );
  NAND2_X1 U7453 ( .A1(n7104), .A2(n7103), .ZN(n5946) );
  NAND2_X1 U7454 ( .A1(n5946), .A2(n5945), .ZN(n7108) );
  INV_X1 U7455 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6967) );
  OR2_X1 U7456 ( .A1(n6190), .A2(n6967), .ZN(n5954) );
  NOR2_X1 U7457 ( .A1(n5895), .A2(n6130), .ZN(n5949) );
  MUX2_X1 U7458 ( .A(n6130), .B(n5949), .S(P1_IR_REG_2__SCAN_IN), .Z(n5950) );
  INV_X1 U7459 ( .A(n5950), .ZN(n5952) );
  NAND2_X1 U7460 ( .A1(n5952), .A2(n5951), .ZN(n7029) );
  OAI211_X1 U7461 ( .C1(n6535), .C2(n8221), .A(n5954), .B(n5953), .ZN(n6496)
         );
  NAND2_X1 U7462 ( .A1(n5970), .A2(n6496), .ZN(n5960) );
  NAND2_X1 U7463 ( .A1(n6478), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7464 ( .A1(n5991), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7465 ( .A1(n4516), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7466 ( .A1(n6034), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5955) );
  NAND4_X4 U7467 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n9997)
         );
  NAND2_X1 U7468 ( .A1(n9997), .A2(n6440), .ZN(n5959) );
  NAND2_X1 U7469 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  XNOR2_X1 U7470 ( .A(n5961), .B(n6438), .ZN(n5964) );
  INV_X1 U7471 ( .A(n9997), .ZN(n7646) );
  NAND2_X1 U7472 ( .A1(n6496), .A2(n6440), .ZN(n5962) );
  AND2_X1 U7473 ( .A1(n5963), .A2(n5962), .ZN(n5965) );
  NAND2_X1 U7474 ( .A1(n5964), .A2(n5965), .ZN(n5969) );
  INV_X1 U7475 ( .A(n5964), .ZN(n5967) );
  INV_X1 U7476 ( .A(n5965), .ZN(n5966) );
  NAND2_X1 U7477 ( .A1(n5967), .A2(n5966), .ZN(n5968) );
  AND2_X1 U7478 ( .A1(n5969), .A2(n5968), .ZN(n7124) );
  NAND2_X1 U7479 ( .A1(n7123), .A2(n7124), .ZN(n7122) );
  NAND2_X1 U7480 ( .A1(n7122), .A2(n5969), .ZN(n7183) );
  NAND2_X1 U7481 ( .A1(n5951), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5971) );
  XNOR2_X1 U7482 ( .A(n5971), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7030) );
  AOI22_X1 U7483 ( .A1(n6172), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n4526), .B2(
        n7030), .ZN(n5973) );
  OR2_X1 U7484 ( .A1(n6968), .A2(n6535), .ZN(n5972) );
  NAND2_X1 U7485 ( .A1(n5973), .A2(n5972), .ZN(n7628) );
  NAND2_X1 U7486 ( .A1(n5987), .A2(n7628), .ZN(n5979) );
  NAND2_X1 U7487 ( .A1(n5991), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5977) );
  INV_X1 U7488 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U7489 ( .A1(n6478), .A2(n7629), .ZN(n5976) );
  NAND2_X1 U7490 ( .A1(n6034), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7491 ( .A1(n4516), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5974) );
  NAND4_X1 U7492 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n9355)
         );
  NAND2_X1 U7493 ( .A1(n9355), .A2(n6440), .ZN(n5978) );
  NAND2_X1 U7494 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  XNOR2_X1 U7495 ( .A(n5980), .B(n6438), .ZN(n5985) );
  NAND2_X1 U7496 ( .A1(n7628), .A2(n6440), .ZN(n5981) );
  NAND2_X1 U7497 ( .A1(n5982), .A2(n5981), .ZN(n5983) );
  XNOR2_X1 U7498 ( .A(n5985), .B(n5983), .ZN(n7184) );
  NAND2_X1 U7499 ( .A1(n7183), .A2(n7184), .ZN(n7182) );
  INV_X1 U7500 ( .A(n5983), .ZN(n5984) );
  NAND2_X1 U7501 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7502 ( .A1(n7182), .A2(n5986), .ZN(n7255) );
  INV_X1 U7503 ( .A(n7255), .ZN(n6003) );
  OR2_X1 U7504 ( .A1(n6970), .A2(n6535), .ZN(n5990) );
  OR2_X1 U7505 ( .A1(n5951), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7506 ( .A1(n5988), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6008) );
  XNOR2_X1 U7507 ( .A(n6008), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9391) );
  AOI22_X1 U7508 ( .A1(n6172), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n4526), .B2(
        n9391), .ZN(n5989) );
  NAND2_X1 U7509 ( .A1(n5990), .A2(n5989), .ZN(n7583) );
  NAND2_X1 U7510 ( .A1(n5987), .A2(n7583), .ZN(n5998) );
  NAND2_X1 U7511 ( .A1(n6074), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5996) );
  INV_X1 U7512 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7259) );
  NAND2_X1 U7513 ( .A1(n7629), .A2(n7259), .ZN(n5992) );
  INV_X1 U7514 ( .A(n6013), .ZN(n6014) );
  AND2_X1 U7515 ( .A1(n5992), .A2(n6014), .ZN(n7584) );
  NAND2_X1 U7516 ( .A1(n6413), .A2(n7584), .ZN(n5995) );
  NAND2_X1 U7517 ( .A1(n6034), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7518 ( .A1(n5926), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7519 ( .A1(n9354), .A2(n6422), .ZN(n5997) );
  NAND2_X1 U7520 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  XNOR2_X1 U7521 ( .A(n5999), .B(n6387), .ZN(n6005) );
  INV_X1 U7522 ( .A(n9354), .ZN(n7384) );
  OR2_X1 U7523 ( .A1(n7384), .A2(n6400), .ZN(n6001) );
  NAND2_X1 U7524 ( .A1(n7583), .A2(n6440), .ZN(n6000) );
  NAND2_X1 U7525 ( .A1(n6001), .A2(n6000), .ZN(n6004) );
  XNOR2_X1 U7526 ( .A(n6005), .B(n6004), .ZN(n7256) );
  INV_X1 U7527 ( .A(n7256), .ZN(n6002) );
  NAND2_X1 U7528 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  OR2_X1 U7529 ( .A1(n6977), .A2(n6535), .ZN(n6012) );
  NAND2_X1 U7530 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  NAND2_X1 U7531 ( .A1(n6009), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7532 ( .A(n6010), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9408) );
  AOI22_X1 U7533 ( .A1(n6172), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n4526), .B2(
        n9408), .ZN(n6011) );
  NAND2_X1 U7534 ( .A1(n6012), .A2(n6011), .ZN(n10031) );
  NAND2_X1 U7535 ( .A1(n5987), .A2(n10031), .ZN(n6021) );
  NAND2_X1 U7536 ( .A1(n6074), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7537 ( .A1(n6013), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6032) );
  INV_X1 U7538 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7383) );
  NAND2_X1 U7539 ( .A1(n6014), .A2(n7383), .ZN(n6015) );
  AND2_X1 U7540 ( .A1(n6032), .A2(n6015), .ZN(n7606) );
  NAND2_X1 U7541 ( .A1(n6478), .A2(n7606), .ZN(n6018) );
  NAND2_X1 U7542 ( .A1(n6034), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7543 ( .A1(n5926), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6016) );
  NAND4_X1 U7544 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n9353)
         );
  NAND2_X1 U7545 ( .A1(n9353), .A2(n6440), .ZN(n6020) );
  NAND2_X1 U7546 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  XNOR2_X1 U7547 ( .A(n6022), .B(n6438), .ZN(n7380) );
  NAND2_X1 U7548 ( .A1(n10031), .A2(n6440), .ZN(n6024) );
  INV_X1 U7549 ( .A(n9353), .ZN(n7580) );
  OR2_X1 U7550 ( .A1(n7580), .A2(n6400), .ZN(n6023) );
  AND2_X1 U7551 ( .A1(n6024), .A2(n6023), .ZN(n6047) );
  NAND2_X1 U7552 ( .A1(n7380), .A2(n6047), .ZN(n6025) );
  NOR2_X1 U7553 ( .A1(n6026), .A2(n6130), .ZN(n6027) );
  MUX2_X1 U7554 ( .A(n6130), .B(n6027), .S(P1_IR_REG_6__SCAN_IN), .Z(n6028) );
  OR2_X1 U7555 ( .A1(n6028), .A2(n6052), .ZN(n7048) );
  INV_X1 U7556 ( .A(n7048), .ZN(n7043) );
  AOI22_X1 U7557 ( .A1(n6172), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n4526), .B2(
        n7043), .ZN(n6029) );
  NAND2_X1 U7558 ( .A1(n6030), .A2(n6029), .ZN(n10041) );
  NAND2_X1 U7559 ( .A1(n10041), .A2(n5987), .ZN(n6040) );
  NAND2_X1 U7560 ( .A1(n6074), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6038) );
  INV_X1 U7561 ( .A(n6056), .ZN(n6057) );
  NAND2_X1 U7562 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  AND2_X1 U7563 ( .A1(n6057), .A2(n6033), .ZN(n7658) );
  NAND2_X1 U7564 ( .A1(n6413), .A2(n7658), .ZN(n6037) );
  NAND2_X1 U7565 ( .A1(n6034), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7566 ( .A1(n5926), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7567 ( .A1(n10029), .A2(n6440), .ZN(n6039) );
  NAND2_X1 U7568 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  XNOR2_X1 U7569 ( .A(n6041), .B(n6438), .ZN(n6045) );
  NOR2_X1 U7570 ( .A1(n6400), .A2(n9971), .ZN(n6043) );
  AOI21_X1 U7571 ( .B1(n10041), .B2(n6422), .A(n6043), .ZN(n6044) );
  NAND2_X1 U7572 ( .A1(n6045), .A2(n6044), .ZN(n6051) );
  OR2_X1 U7573 ( .A1(n6045), .A2(n6044), .ZN(n6046) );
  NAND2_X1 U7574 ( .A1(n6051), .A2(n6046), .ZN(n7449) );
  INV_X1 U7575 ( .A(n7380), .ZN(n6048) );
  INV_X1 U7576 ( .A(n6047), .ZN(n7382) );
  AND2_X1 U7577 ( .A1(n6048), .A2(n7382), .ZN(n6049) );
  NOR2_X1 U7578 ( .A1(n7449), .A2(n6049), .ZN(n6050) );
  NAND2_X1 U7579 ( .A1(n7454), .A2(n6051), .ZN(n7354) );
  OR2_X1 U7580 ( .A1(n6985), .A2(n6535), .ZN(n6055) );
  OR2_X1 U7581 ( .A1(n6052), .A2(n6130), .ZN(n6053) );
  XNOR2_X1 U7582 ( .A(n6053), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7077) );
  AOI22_X1 U7583 ( .A1(n6172), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4526), .B2(
        n7077), .ZN(n6054) );
  NAND2_X1 U7584 ( .A1(n6055), .A2(n6054), .ZN(n9980) );
  NAND2_X1 U7585 ( .A1(n9980), .A2(n5987), .ZN(n6064) );
  NAND2_X1 U7586 ( .A1(n6074), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7587 ( .A1(n6056), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6076) );
  INV_X1 U7588 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U7589 ( .A1(n6057), .A2(n7055), .ZN(n6058) );
  AND2_X1 U7590 ( .A1(n6076), .A2(n6058), .ZN(n9978) );
  NAND2_X1 U7591 ( .A1(n6413), .A2(n9978), .ZN(n6061) );
  NAND2_X1 U7592 ( .A1(n6034), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7593 ( .A1(n5926), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6059) );
  NAND4_X1 U7594 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n9352)
         );
  NAND2_X1 U7595 ( .A1(n9352), .A2(n6422), .ZN(n6063) );
  NAND2_X1 U7596 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  XNOR2_X1 U7597 ( .A(n6065), .B(n6387), .ZN(n6067) );
  NOR2_X1 U7598 ( .A1(n6400), .A2(n7594), .ZN(n6066) );
  AOI21_X1 U7599 ( .B1(n9980), .B2(n6422), .A(n6066), .ZN(n6068) );
  XNOR2_X1 U7600 ( .A(n6067), .B(n6068), .ZN(n7355) );
  NAND2_X1 U7601 ( .A1(n7354), .A2(n7355), .ZN(n7353) );
  INV_X1 U7602 ( .A(n6067), .ZN(n6069) );
  NAND2_X1 U7603 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  INV_X2 U7604 ( .A(n6535), .ZN(n9058) );
  NAND2_X1 U7605 ( .A1(n6071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6090) );
  XNOR2_X1 U7606 ( .A(n6090), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7202) );
  AOI22_X1 U7607 ( .A1(n6172), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4526), .B2(
        n7202), .ZN(n6072) );
  NAND2_X1 U7608 ( .A1(n9131), .A2(n5987), .ZN(n6083) );
  NAND2_X1 U7609 ( .A1(n6074), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6081) );
  INV_X1 U7610 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7611 ( .A1(n6076), .A2(n6075), .ZN(n6077) );
  AND2_X1 U7612 ( .A1(n6095), .A2(n6077), .ZN(n7703) );
  NAND2_X1 U7613 ( .A1(n6478), .A2(n7703), .ZN(n6080) );
  NAND2_X1 U7614 ( .A1(n6034), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7615 ( .A1(n5926), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6078) );
  NAND4_X1 U7616 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n9351)
         );
  NAND2_X1 U7617 ( .A1(n9351), .A2(n6440), .ZN(n6082) );
  NAND2_X1 U7618 ( .A1(n6083), .A2(n6082), .ZN(n6084) );
  XNOR2_X1 U7619 ( .A(n6084), .B(n6387), .ZN(n6086) );
  INV_X1 U7620 ( .A(n9351), .ZN(n9969) );
  NOR2_X1 U7621 ( .A1(n6400), .A2(n9969), .ZN(n6085) );
  AOI21_X1 U7622 ( .B1(n9131), .B2(n6422), .A(n6085), .ZN(n7592) );
  NAND2_X1 U7623 ( .A1(n7591), .A2(n7592), .ZN(n7590) );
  INV_X1 U7624 ( .A(n6086), .ZN(n6087) );
  NAND2_X1 U7625 ( .A1(n6088), .A2(n6087), .ZN(n7710) );
  NAND2_X1 U7626 ( .A1(n7061), .A2(n9058), .ZN(n6094) );
  NAND2_X1 U7627 ( .A1(n6090), .A2(n6089), .ZN(n6091) );
  NAND2_X1 U7628 ( .A1(n6091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6092) );
  XNOR2_X1 U7629 ( .A(n6092), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9422) );
  AOI22_X1 U7630 ( .A1(n6172), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4526), .B2(
        n9422), .ZN(n6093) );
  NAND2_X1 U7631 ( .A1(n7442), .A2(n5987), .ZN(n6102) );
  NAND2_X1 U7632 ( .A1(n5991), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6100) );
  INV_X1 U7633 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7714) );
  INV_X1 U7634 ( .A(n6115), .ZN(n6117) );
  NAND2_X1 U7635 ( .A1(n6095), .A2(n7714), .ZN(n6096) );
  AND2_X1 U7636 ( .A1(n6117), .A2(n6096), .ZN(n7750) );
  NAND2_X1 U7637 ( .A1(n6478), .A2(n7750), .ZN(n6099) );
  NAND2_X1 U7638 ( .A1(n6034), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7639 ( .A1(n5926), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6097) );
  NAND4_X1 U7640 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(n9350)
         );
  NAND2_X1 U7641 ( .A1(n9350), .A2(n6422), .ZN(n6101) );
  NAND2_X1 U7642 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  XNOR2_X1 U7643 ( .A(n6103), .B(n6387), .ZN(n6106) );
  INV_X1 U7644 ( .A(n9350), .ZN(n7866) );
  NOR2_X1 U7645 ( .A1(n6400), .A2(n7866), .ZN(n6104) );
  AOI21_X1 U7646 ( .B1(n7442), .B2(n6422), .A(n6104), .ZN(n6107) );
  XNOR2_X1 U7647 ( .A(n6106), .B(n6107), .ZN(n7712) );
  NAND2_X1 U7648 ( .A1(n7590), .A2(n6105), .ZN(n7711) );
  INV_X1 U7649 ( .A(n6106), .ZN(n6108) );
  OR2_X1 U7650 ( .A1(n6108), .A2(n6107), .ZN(n6109) );
  NAND2_X1 U7651 ( .A1(n7065), .A2(n9058), .ZN(n6113) );
  NAND2_X1 U7652 ( .A1(n6110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6111) );
  XNOR2_X1 U7653 ( .A(n6111), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7322) );
  AOI22_X1 U7654 ( .A1(n6172), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4526), .B2(
        n7322), .ZN(n6112) );
  NAND2_X1 U7655 ( .A1(n7870), .A2(n5987), .ZN(n6124) );
  NAND2_X1 U7656 ( .A1(n5991), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6122) );
  INV_X1 U7657 ( .A(n6135), .ZN(n6136) );
  INV_X1 U7658 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7659 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  AND2_X1 U7660 ( .A1(n6136), .A2(n6118), .ZN(n7869) );
  NAND2_X1 U7661 ( .A1(n6413), .A2(n7869), .ZN(n6121) );
  NAND2_X1 U7662 ( .A1(n6034), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7663 ( .A1(n5926), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6119) );
  NAND4_X1 U7664 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n9349)
         );
  NAND2_X1 U7665 ( .A1(n9349), .A2(n6422), .ZN(n6123) );
  NAND2_X1 U7666 ( .A1(n6124), .A2(n6123), .ZN(n6125) );
  XNOR2_X1 U7667 ( .A(n6125), .B(n6387), .ZN(n6126) );
  NAND2_X1 U7668 ( .A1(n7870), .A2(n6422), .ZN(n6129) );
  INV_X1 U7669 ( .A(n9349), .ZN(n7886) );
  OR2_X1 U7670 ( .A1(n7886), .A2(n6400), .ZN(n6128) );
  NAND2_X1 U7671 ( .A1(n6129), .A2(n6128), .ZN(n7865) );
  NAND2_X1 U7672 ( .A1(n7070), .A2(n9058), .ZN(n6134) );
  OR2_X1 U7673 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  XNOR2_X1 U7674 ( .A(n6132), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9436) );
  AOI22_X1 U7675 ( .A1(n6172), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9436), .B2(
        n4526), .ZN(n6133) );
  NAND2_X1 U7676 ( .A1(n7543), .A2(n5987), .ZN(n6143) );
  NAND2_X1 U7677 ( .A1(n5991), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7678 ( .A1(n6135), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6153) );
  INV_X1 U7679 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U7680 ( .A1(n6136), .A2(n7885), .ZN(n6137) );
  AND2_X1 U7681 ( .A1(n6153), .A2(n6137), .ZN(n7888) );
  NAND2_X1 U7682 ( .A1(n6478), .A2(n7888), .ZN(n6140) );
  NAND2_X1 U7683 ( .A1(n6034), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7684 ( .A1(n5926), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6138) );
  NAND4_X1 U7685 ( .A1(n6141), .A2(n6140), .A3(n6139), .A4(n6138), .ZN(n9348)
         );
  NAND2_X1 U7686 ( .A1(n9348), .A2(n6422), .ZN(n6142) );
  NAND2_X1 U7687 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  XNOR2_X1 U7688 ( .A(n6144), .B(n6438), .ZN(n6147) );
  INV_X1 U7689 ( .A(n9348), .ZN(n7942) );
  NOR2_X1 U7690 ( .A1(n6400), .A2(n7942), .ZN(n6145) );
  AOI21_X1 U7691 ( .B1(n7543), .B2(n6422), .A(n6145), .ZN(n6146) );
  NAND2_X1 U7692 ( .A1(n6147), .A2(n6146), .ZN(n7935) );
  OR2_X1 U7693 ( .A1(n6147), .A2(n6146), .ZN(n6148) );
  AND2_X1 U7694 ( .A1(n7935), .A2(n6148), .ZN(n7881) );
  NAND2_X1 U7695 ( .A1(n7883), .A2(n7935), .ZN(n6166) );
  NAND2_X1 U7696 ( .A1(n7094), .A2(n9058), .ZN(n6151) );
  NAND2_X1 U7697 ( .A1(n6149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6169) );
  XNOR2_X1 U7698 ( .A(n6169), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9448) );
  AOI22_X1 U7699 ( .A1(n9448), .A2(n4526), .B1(n6172), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7700 ( .A1(n7791), .A2(n5987), .ZN(n6160) );
  NAND2_X1 U7701 ( .A1(n5991), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6158) );
  INV_X1 U7702 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7703 ( .A1(n6153), .A2(n6152), .ZN(n6154) );
  AND2_X1 U7704 ( .A1(n6175), .A2(n6154), .ZN(n7945) );
  NAND2_X1 U7705 ( .A1(n6478), .A2(n7945), .ZN(n6157) );
  NAND2_X1 U7706 ( .A1(n5926), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7707 ( .A1(n6034), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6155) );
  NAND4_X1 U7708 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n9347)
         );
  NAND2_X1 U7709 ( .A1(n9347), .A2(n6422), .ZN(n6159) );
  NAND2_X1 U7710 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  XNOR2_X1 U7711 ( .A(n6161), .B(n6438), .ZN(n6164) );
  INV_X1 U7712 ( .A(n9347), .ZN(n8003) );
  NOR2_X1 U7713 ( .A1(n6400), .A2(n8003), .ZN(n6162) );
  AOI21_X1 U7714 ( .B1(n7791), .B2(n6422), .A(n6162), .ZN(n6163) );
  NAND2_X1 U7715 ( .A1(n6164), .A2(n6163), .ZN(n6167) );
  OR2_X1 U7716 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  AND2_X1 U7717 ( .A1(n6167), .A2(n6165), .ZN(n7936) );
  NAND2_X1 U7718 ( .A1(n6166), .A2(n7936), .ZN(n7939) );
  NAND2_X1 U7719 ( .A1(n7939), .A2(n6167), .ZN(n7999) );
  NAND2_X1 U7720 ( .A1(n7101), .A2(n9058), .ZN(n6174) );
  NAND2_X1 U7721 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U7722 ( .A1(n6170), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6171) );
  XNOR2_X1 U7723 ( .A(n6171), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9462) );
  AOI22_X1 U7724 ( .A1(n9462), .A2(n4526), .B1(n6172), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7725 ( .A1(n7997), .A2(n5987), .ZN(n6182) );
  NAND2_X1 U7726 ( .A1(n5991), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6180) );
  INV_X1 U7727 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U7728 ( .A1(n6175), .A2(n8002), .ZN(n6176) );
  AND2_X1 U7729 ( .A1(n6195), .A2(n6176), .ZN(n8005) );
  NAND2_X1 U7730 ( .A1(n6413), .A2(n8005), .ZN(n6179) );
  NAND2_X1 U7731 ( .A1(n4527), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7732 ( .A1(n6034), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6177) );
  NAND4_X1 U7733 ( .A1(n6180), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(n10062)
         );
  NAND2_X1 U7734 ( .A1(n10062), .A2(n6422), .ZN(n6181) );
  NAND2_X1 U7735 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  XNOR2_X1 U7736 ( .A(n6183), .B(n6387), .ZN(n6185) );
  INV_X1 U7737 ( .A(n10062), .ZN(n8914) );
  NOR2_X1 U7738 ( .A1(n6400), .A2(n8914), .ZN(n6184) );
  AOI21_X1 U7739 ( .B1(n7997), .B2(n6422), .A(n6184), .ZN(n6186) );
  XNOR2_X1 U7740 ( .A(n6185), .B(n6186), .ZN(n8000) );
  INV_X1 U7741 ( .A(n6185), .ZN(n6187) );
  NAND2_X1 U7742 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  NAND2_X1 U7743 ( .A1(n7147), .A2(n9058), .ZN(n6193) );
  NAND2_X1 U7744 ( .A1(n6189), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6269) );
  XNOR2_X1 U7745 ( .A(n6269), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9480) );
  INV_X1 U7746 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10615) );
  NOR2_X1 U7747 ( .A1(n9060), .A2(n10615), .ZN(n6191) );
  AOI21_X1 U7748 ( .B1(n9480), .B2(n4526), .A(n6191), .ZN(n6192) );
  NAND2_X1 U7749 ( .A1(n9111), .A2(n5987), .ZN(n6200) );
  INV_X1 U7750 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6194) );
  INV_X1 U7751 ( .A(n6211), .ZN(n6213) );
  NAND2_X1 U7752 ( .A1(n6195), .A2(n6194), .ZN(n6196) );
  NAND2_X1 U7753 ( .A1(n6213), .A2(n6196), .ZN(n7780) );
  AOI22_X1 U7754 ( .A1(n5991), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n6034), .B2(
        P1_REG0_REG_14__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7755 ( .A1(n4527), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6197) );
  OAI211_X1 U7756 ( .C1(n7780), .C2(n6239), .A(n6198), .B(n6197), .ZN(n9346)
         );
  NAND2_X1 U7757 ( .A1(n9346), .A2(n6440), .ZN(n6199) );
  NAND2_X1 U7758 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  XNOR2_X1 U7759 ( .A(n6201), .B(n6438), .ZN(n6204) );
  INV_X1 U7760 ( .A(n9346), .ZN(n9110) );
  NOR2_X1 U7761 ( .A1(n6400), .A2(n9110), .ZN(n6203) );
  AOI21_X1 U7762 ( .B1(n9111), .B2(n6422), .A(n6203), .ZN(n8912) );
  NAND2_X1 U7763 ( .A1(n8911), .A2(n8912), .ZN(n6227) );
  NAND2_X1 U7764 ( .A1(n6205), .A2(n6204), .ZN(n8910) );
  NAND2_X1 U7765 ( .A1(n6227), .A2(n8910), .ZN(n6222) );
  NAND2_X1 U7766 ( .A1(n7210), .A2(n9058), .ZN(n6210) );
  NAND2_X1 U7767 ( .A1(n6269), .A2(n6206), .ZN(n6207) );
  NAND2_X1 U7768 ( .A1(n6207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6228) );
  XNOR2_X1 U7769 ( .A(n6228), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9488) );
  INV_X1 U7770 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10394) );
  NOR2_X1 U7771 ( .A1(n9060), .A2(n10394), .ZN(n6208) );
  AOI21_X1 U7772 ( .B1(n9488), .B2(n4526), .A(n6208), .ZN(n6209) );
  NAND2_X1 U7773 ( .A1(n9927), .A2(n5987), .ZN(n6220) );
  INV_X1 U7774 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7775 ( .A1(n6211), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6235) );
  INV_X1 U7776 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7777 ( .A1(n6213), .A2(n6212), .ZN(n6214) );
  NAND2_X1 U7778 ( .A1(n6235), .A2(n6214), .ZN(n9040) );
  OR2_X1 U7779 ( .A1(n9040), .A2(n6239), .ZN(n6216) );
  AOI22_X1 U7780 ( .A1(n5991), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n6034), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n6215) );
  OAI211_X1 U7781 ( .C1(n6218), .C2(n6217), .A(n6216), .B(n6215), .ZN(n10065)
         );
  NAND2_X1 U7782 ( .A1(n10065), .A2(n6440), .ZN(n6219) );
  NAND2_X1 U7783 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  XNOR2_X1 U7784 ( .A(n6221), .B(n6438), .ZN(n6225) );
  NAND2_X1 U7785 ( .A1(n9927), .A2(n6440), .ZN(n6224) );
  NAND2_X1 U7786 ( .A1(n6042), .A2(n10065), .ZN(n6223) );
  NAND2_X1 U7787 ( .A1(n6224), .A2(n6223), .ZN(n9043) );
  INV_X1 U7788 ( .A(n6225), .ZN(n6226) );
  NAND2_X1 U7789 ( .A1(n7263), .A2(n9058), .ZN(n6233) );
  NAND2_X1 U7790 ( .A1(n6228), .A2(n10664), .ZN(n6229) );
  NAND2_X1 U7791 ( .A1(n6229), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6230) );
  XNOR2_X1 U7792 ( .A(n6230), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9515) );
  NOR2_X1 U7793 ( .A1(n9060), .A2(n10374), .ZN(n6231) );
  AOI21_X1 U7794 ( .B1(n9515), .B2(n4526), .A(n6231), .ZN(n6232) );
  NAND2_X1 U7795 ( .A1(n8964), .A2(n5987), .ZN(n6241) );
  INV_X1 U7796 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7797 ( .A1(n6235), .A2(n6234), .ZN(n6236) );
  NAND2_X1 U7798 ( .A1(n8971), .A2(n6236), .ZN(n8962) );
  AOI22_X1 U7799 ( .A1(n5991), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n4527), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7800 ( .A1(n6034), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6237) );
  OAI211_X1 U7801 ( .C1(n8962), .C2(n6239), .A(n6238), .B(n6237), .ZN(n9345)
         );
  NAND2_X1 U7802 ( .A1(n9345), .A2(n6440), .ZN(n6240) );
  NAND2_X1 U7803 ( .A1(n6241), .A2(n6240), .ZN(n6242) );
  XNOR2_X1 U7804 ( .A(n6242), .B(n6438), .ZN(n6245) );
  AND2_X1 U7805 ( .A1(n9345), .A2(n6042), .ZN(n6243) );
  AOI21_X1 U7806 ( .B1(n8964), .B2(n6422), .A(n6243), .ZN(n6244) );
  NOR2_X1 U7807 ( .A1(n6245), .A2(n6244), .ZN(n8958) );
  NAND2_X1 U7808 ( .A1(n6245), .A2(n6244), .ZN(n8957) );
  NAND2_X1 U7809 ( .A1(n7294), .A2(n9058), .ZN(n6252) );
  NAND2_X1 U7810 ( .A1(n6246), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7811 ( .A1(n6269), .A2(n6247), .ZN(n6249) );
  XNOR2_X1 U7812 ( .A(n6249), .B(n6248), .ZN(n9532) );
  NOR2_X1 U7813 ( .A1(n9060), .A2(n10366), .ZN(n6250) );
  AOI21_X1 U7814 ( .B1(n9532), .B2(n4526), .A(n6250), .ZN(n6251) );
  NAND2_X1 U7815 ( .A1(n8977), .A2(n5987), .ZN(n6260) );
  XNOR2_X1 U7816 ( .A(n8971), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U7817 ( .A1(n7991), .A2(n6478), .ZN(n6258) );
  INV_X1 U7818 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7819 ( .A1(n6034), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7820 ( .A1(n4527), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6253) );
  OAI211_X1 U7821 ( .C1(n6114), .C2(n6255), .A(n6254), .B(n6253), .ZN(n6256)
         );
  INV_X1 U7822 ( .A(n6256), .ZN(n6257) );
  NAND2_X1 U7823 ( .A1(n6258), .A2(n6257), .ZN(n9918) );
  NAND2_X1 U7824 ( .A1(n9918), .A2(n6440), .ZN(n6259) );
  NAND2_X1 U7825 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  XNOR2_X1 U7826 ( .A(n6261), .B(n6438), .ZN(n8968) );
  AND2_X1 U7827 ( .A1(n9918), .A2(n6042), .ZN(n6262) );
  AOI21_X1 U7828 ( .B1(n8977), .B2(n6422), .A(n6262), .ZN(n8967) );
  INV_X1 U7829 ( .A(n8968), .ZN(n6264) );
  INV_X1 U7830 ( .A(n8967), .ZN(n6263) );
  NAND2_X1 U7831 ( .A1(n7407), .A2(n9058), .ZN(n6274) );
  NAND2_X1 U7832 ( .A1(n6267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7833 ( .A1(n6269), .A2(n6268), .ZN(n6270) );
  XNOR2_X1 U7834 ( .A(n6270), .B(n5861), .ZN(n9546) );
  INV_X1 U7835 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10379) );
  NOR2_X1 U7836 ( .A1(n9060), .A2(n10379), .ZN(n6271) );
  AOI21_X1 U7837 ( .B1(n9546), .B2(n4526), .A(n6271), .ZN(n6273) );
  INV_X1 U7838 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6275) );
  OR2_X1 U7839 ( .A1(n6276), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7840 ( .A1(n6276), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6291) );
  AND2_X1 U7841 ( .A1(n6277), .A2(n6291), .ZN(n9733) );
  NAND2_X1 U7842 ( .A1(n9733), .A2(n6478), .ZN(n6282) );
  INV_X1 U7843 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U7844 ( .A1(n6034), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7845 ( .A1(n4527), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6278) );
  OAI211_X1 U7846 ( .C1(n6114), .C2(n9853), .A(n6279), .B(n6278), .ZN(n6280)
         );
  INV_X1 U7847 ( .A(n6280), .ZN(n6281) );
  NAND2_X1 U7848 ( .A1(n6282), .A2(n6281), .ZN(n9711) );
  AOI22_X1 U7849 ( .A1(n9744), .A2(n6422), .B1(n6042), .B2(n9711), .ZN(n6284)
         );
  INV_X1 U7850 ( .A(n6284), .ZN(n9012) );
  AOI22_X1 U7851 ( .A1(n9744), .A2(n5987), .B1(n6440), .B2(n9711), .ZN(n6283)
         );
  XNOR2_X1 U7852 ( .A(n6283), .B(n6387), .ZN(n9013) );
  NAND2_X1 U7853 ( .A1(n7546), .A2(n9058), .ZN(n6289) );
  INV_X1 U7854 ( .A(n6287), .ZN(n6288) );
  NAND2_X1 U7855 ( .A1(n5991), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6297) );
  INV_X1 U7856 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7857 ( .A1(n6290), .A2(n6291), .ZN(n6293) );
  INV_X1 U7858 ( .A(n6291), .ZN(n6292) );
  AND2_X1 U7859 ( .A1(n6293), .A2(n6318), .ZN(n9716) );
  NAND2_X1 U7860 ( .A1(n6413), .A2(n9716), .ZN(n6296) );
  NAND2_X1 U7861 ( .A1(n4514), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7862 ( .A1(n4527), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6294) );
  NAND4_X1 U7863 ( .A1(n6297), .A2(n6296), .A3(n6295), .A4(n6294), .ZN(n9846)
         );
  AOI22_X1 U7864 ( .A1(n9843), .A2(n6422), .B1(n6042), .B2(n9846), .ZN(n6303)
         );
  NAND2_X1 U7865 ( .A1(n9843), .A2(n5987), .ZN(n6299) );
  NAND2_X1 U7866 ( .A1(n9846), .A2(n6440), .ZN(n6298) );
  NAND2_X1 U7867 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  XNOR2_X1 U7868 ( .A(n6300), .B(n6387), .ZN(n6301) );
  XOR2_X1 U7869 ( .A(n6303), .B(n6301), .Z(n8931) );
  INV_X1 U7870 ( .A(n6301), .ZN(n6302) );
  NAND2_X1 U7871 ( .A1(n7600), .A2(n9058), .ZN(n6306) );
  INV_X1 U7872 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6304) );
  OR2_X1 U7873 ( .A1(n9060), .A2(n6304), .ZN(n6305) );
  NAND2_X1 U7874 ( .A1(n5991), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6310) );
  XNOR2_X1 U7875 ( .A(n6318), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U7876 ( .A1(n6413), .A2(n9699), .ZN(n6309) );
  NAND2_X1 U7877 ( .A1(n6034), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U7878 ( .A1(n4527), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6307) );
  NAND4_X1 U7879 ( .A1(n6310), .A2(n6309), .A3(n6308), .A4(n6307), .ZN(n9828)
         );
  AOI22_X1 U7880 ( .A1(n9698), .A2(n5987), .B1(n6440), .B2(n9828), .ZN(n6311)
         );
  XNOR2_X1 U7881 ( .A(n6311), .B(n6387), .ZN(n6313) );
  AOI22_X1 U7882 ( .A1(n9698), .A2(n6422), .B1(n6042), .B2(n9828), .ZN(n6312)
         );
  NAND2_X1 U7883 ( .A1(n6313), .A2(n6312), .ZN(n8988) );
  NOR2_X1 U7884 ( .A1(n6313), .A2(n6312), .ZN(n8989) );
  NAND2_X1 U7885 ( .A1(n7775), .A2(n9058), .ZN(n6315) );
  OR2_X1 U7886 ( .A1(n9060), .A2(n7789), .ZN(n6314) );
  NAND2_X1 U7887 ( .A1(n9688), .A2(n5987), .ZN(n6325) );
  NAND2_X1 U7888 ( .A1(n5991), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6323) );
  INV_X1 U7889 ( .A(n6318), .ZN(n6316) );
  AOI21_X1 U7890 ( .B1(n6316), .B2(P1_REG3_REG_20__SCAN_IN), .A(
        P1_REG3_REG_21__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7891 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n6317) );
  OR2_X1 U7892 ( .A1(n6319), .A2(n6333), .ZN(n8943) );
  INV_X1 U7893 ( .A(n8943), .ZN(n9679) );
  NAND2_X1 U7894 ( .A1(n6413), .A2(n9679), .ZN(n6322) );
  NAND2_X1 U7895 ( .A1(n4514), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U7896 ( .A1(n4527), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6320) );
  NAND4_X1 U7897 ( .A1(n6323), .A2(n6322), .A3(n6321), .A4(n6320), .ZN(n9817)
         );
  NAND2_X1 U7898 ( .A1(n9817), .A2(n6440), .ZN(n6324) );
  NAND2_X1 U7899 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  XNOR2_X1 U7900 ( .A(n6326), .B(n6387), .ZN(n8939) );
  NAND2_X1 U7901 ( .A1(n9688), .A2(n6440), .ZN(n6328) );
  INV_X1 U7902 ( .A(n9817), .ZN(n9184) );
  OR2_X1 U7903 ( .A1(n9184), .A2(n6400), .ZN(n6327) );
  NAND2_X1 U7904 ( .A1(n6328), .A2(n6327), .ZN(n8938) );
  INV_X1 U7905 ( .A(n8939), .ZN(n6330) );
  INV_X1 U7906 ( .A(n8938), .ZN(n6329) );
  NAND2_X1 U7907 ( .A1(n7849), .A2(n9058), .ZN(n6332) );
  OR2_X1 U7908 ( .A1(n9060), .A2(n10642), .ZN(n6331) );
  NAND2_X1 U7909 ( .A1(n9670), .A2(n5987), .ZN(n6340) );
  NAND2_X1 U7910 ( .A1(n5991), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6338) );
  NOR2_X1 U7911 ( .A1(n6333), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6334) );
  OR2_X1 U7912 ( .A1(n6347), .A2(n6334), .ZN(n9007) );
  INV_X1 U7913 ( .A(n9007), .ZN(n9663) );
  NAND2_X1 U7914 ( .A1(n6478), .A2(n9663), .ZN(n6337) );
  NAND2_X1 U7915 ( .A1(n6034), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7916 ( .A1(n4527), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6335) );
  NAND4_X1 U7917 ( .A1(n6338), .A2(n6337), .A3(n6336), .A4(n6335), .ZN(n9827)
         );
  NAND2_X1 U7918 ( .A1(n9827), .A2(n6440), .ZN(n6339) );
  NAND2_X1 U7919 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  XNOR2_X1 U7920 ( .A(n6341), .B(n6387), .ZN(n8998) );
  NAND2_X1 U7921 ( .A1(n9670), .A2(n6440), .ZN(n6343) );
  INV_X1 U7922 ( .A(n9827), .ZN(n9682) );
  OR2_X1 U7923 ( .A1(n9682), .A2(n6400), .ZN(n6342) );
  NAND2_X1 U7924 ( .A1(n6343), .A2(n6342), .ZN(n9003) );
  NAND2_X1 U7925 ( .A1(n7877), .A2(n9058), .ZN(n6346) );
  OR2_X1 U7926 ( .A1(n9060), .A2(n6344), .ZN(n6345) );
  NAND2_X1 U7927 ( .A1(n9656), .A2(n5987), .ZN(n6354) );
  NAND2_X1 U7928 ( .A1(n6074), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6352) );
  OR2_X1 U7929 ( .A1(n6347), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U7930 ( .A1(n6347), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6362) );
  AND2_X1 U7931 ( .A1(n6348), .A2(n6362), .ZN(n9648) );
  NAND2_X1 U7932 ( .A1(n6478), .A2(n9648), .ZN(n6351) );
  NAND2_X1 U7933 ( .A1(n4514), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7934 ( .A1(n4527), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6349) );
  NAND4_X1 U7935 ( .A1(n6352), .A2(n6351), .A3(n6350), .A4(n6349), .ZN(n9816)
         );
  NAND2_X1 U7936 ( .A1(n9816), .A2(n6440), .ZN(n6353) );
  NAND2_X1 U7937 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  XNOR2_X1 U7938 ( .A(n6355), .B(n6438), .ZN(n6358) );
  INV_X1 U7939 ( .A(n9816), .ZN(n9666) );
  NOR2_X1 U7940 ( .A1(n6400), .A2(n9666), .ZN(n6356) );
  AOI21_X1 U7941 ( .B1(n9656), .B2(n6422), .A(n6356), .ZN(n6357) );
  NAND2_X1 U7942 ( .A1(n6358), .A2(n6357), .ZN(n8982) );
  OR2_X1 U7943 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NAND2_X1 U7944 ( .A1(n7930), .A2(n9058), .ZN(n6361) );
  OR2_X1 U7945 ( .A1(n9060), .A2(n10418), .ZN(n6360) );
  NAND2_X1 U7946 ( .A1(n9636), .A2(n5987), .ZN(n6369) );
  NAND2_X1 U7947 ( .A1(n5991), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6367) );
  INV_X1 U7948 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6363) );
  AOI21_X1 U7949 ( .B1(n6363), .B2(n6362), .A(n6379), .ZN(n9637) );
  NAND2_X1 U7950 ( .A1(n6413), .A2(n9637), .ZN(n6366) );
  NAND2_X1 U7951 ( .A1(n4514), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U7952 ( .A1(n4527), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6364) );
  NAND4_X1 U7953 ( .A1(n6367), .A2(n6366), .A3(n6365), .A4(n6364), .ZN(n9806)
         );
  NAND2_X1 U7954 ( .A1(n9806), .A2(n6440), .ZN(n6368) );
  NAND2_X1 U7955 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  XNOR2_X1 U7956 ( .A(n6370), .B(n6438), .ZN(n6373) );
  INV_X1 U7957 ( .A(n9806), .ZN(n9651) );
  NOR2_X1 U7958 ( .A1(n6400), .A2(n9651), .ZN(n6371) );
  AOI21_X1 U7959 ( .B1(n9636), .B2(n6440), .A(n6371), .ZN(n6372) );
  NAND2_X1 U7960 ( .A1(n6373), .A2(n6372), .ZN(n6375) );
  OR2_X1 U7961 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  NAND2_X1 U7962 ( .A1(n6375), .A2(n6374), .ZN(n8981) );
  INV_X1 U7963 ( .A(n6375), .ZN(n6376) );
  NAND2_X1 U7964 ( .A1(n7961), .A2(n9058), .ZN(n6378) );
  OR2_X1 U7965 ( .A1(n9060), .A2(n10584), .ZN(n6377) );
  NAND2_X1 U7966 ( .A1(n6074), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6384) );
  INV_X1 U7967 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8951) );
  INV_X1 U7968 ( .A(n6379), .ZN(n6380) );
  NAND2_X1 U7969 ( .A1(n6379), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6392) );
  INV_X1 U7970 ( .A(n6392), .ZN(n6391) );
  AOI21_X1 U7971 ( .B1(n8951), .B2(n6380), .A(n6391), .ZN(n9624) );
  NAND2_X1 U7972 ( .A1(n6413), .A2(n9624), .ZN(n6383) );
  NAND2_X1 U7973 ( .A1(n6034), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U7974 ( .A1(n4527), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6381) );
  NAND4_X1 U7975 ( .A1(n6384), .A2(n6383), .A3(n6382), .A4(n6381), .ZN(n9784)
         );
  AOI22_X1 U7976 ( .A1(n9878), .A2(n6422), .B1(n6042), .B2(n9784), .ZN(n6402)
         );
  NAND2_X1 U7977 ( .A1(n9878), .A2(n5987), .ZN(n6386) );
  NAND2_X1 U7978 ( .A1(n9784), .A2(n6440), .ZN(n6385) );
  NAND2_X1 U7979 ( .A1(n6386), .A2(n6385), .ZN(n6388) );
  XNOR2_X1 U7980 ( .A(n6388), .B(n6387), .ZN(n6404) );
  XOR2_X1 U7981 ( .A(n6402), .B(n6404), .Z(n8949) );
  NAND2_X1 U7982 ( .A1(n8038), .A2(n9058), .ZN(n6390) );
  OR2_X1 U7983 ( .A1(n9060), .A2(n10424), .ZN(n6389) );
  NAND2_X1 U7984 ( .A1(n9613), .A2(n5987), .ZN(n6398) );
  NAND2_X1 U7985 ( .A1(n6074), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6396) );
  INV_X1 U7986 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U7987 ( .A1(n6391), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6412) );
  INV_X1 U7988 ( .A(n6412), .ZN(n6427) );
  AOI21_X1 U7989 ( .B1(n9027), .B2(n6392), .A(n6427), .ZN(n9605) );
  NAND2_X1 U7990 ( .A1(n6478), .A2(n9605), .ZN(n6395) );
  NAND2_X1 U7991 ( .A1(n4514), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U7992 ( .A1(n4527), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6393) );
  NAND4_X1 U7993 ( .A1(n6396), .A2(n6395), .A3(n6394), .A4(n6393), .ZN(n9775)
         );
  NAND2_X1 U7994 ( .A1(n9775), .A2(n6440), .ZN(n6397) );
  NAND2_X1 U7995 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  XNOR2_X1 U7996 ( .A(n6399), .B(n6438), .ZN(n6406) );
  NOR2_X1 U7997 ( .A1(n6400), .A2(n9195), .ZN(n6401) );
  AOI21_X1 U7998 ( .B1(n9613), .B2(n6440), .A(n6401), .ZN(n6407) );
  XNOR2_X1 U7999 ( .A(n6406), .B(n6407), .ZN(n9021) );
  INV_X1 U8000 ( .A(n6402), .ZN(n6403) );
  INV_X1 U8001 ( .A(n6406), .ZN(n6409) );
  INV_X1 U8002 ( .A(n6407), .ZN(n6408) );
  NAND2_X1 U8003 ( .A1(n8220), .A2(n9058), .ZN(n6411) );
  OR2_X1 U8004 ( .A1(n9060), .A2(n10617), .ZN(n6410) );
  NAND2_X1 U8005 ( .A1(n9871), .A2(n5987), .ZN(n6419) );
  NAND2_X1 U8006 ( .A1(n6074), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6417) );
  XNOR2_X1 U8007 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n6412), .ZN(n9594) );
  NAND2_X1 U8008 ( .A1(n6413), .A2(n9594), .ZN(n6416) );
  NAND2_X1 U8009 ( .A1(n6034), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8010 ( .A1(n4527), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6414) );
  NAND4_X1 U8011 ( .A1(n6417), .A2(n6416), .A3(n6415), .A4(n6414), .ZN(n9783)
         );
  NAND2_X1 U8012 ( .A1(n9783), .A2(n6440), .ZN(n6418) );
  NAND2_X1 U8013 ( .A1(n6419), .A2(n6418), .ZN(n6420) );
  XNOR2_X1 U8014 ( .A(n6420), .B(n6438), .ZN(n6424) );
  NOR2_X1 U8015 ( .A1(n6400), .A2(n9608), .ZN(n6421) );
  AOI21_X1 U8016 ( .B1(n9871), .B2(n6422), .A(n6421), .ZN(n6423) );
  NAND2_X1 U8017 ( .A1(n6424), .A2(n6423), .ZN(n6485) );
  OAI21_X1 U8018 ( .B1(n6424), .B2(n6423), .A(n6485), .ZN(n6932) );
  NAND2_X1 U8019 ( .A1(n8101), .A2(n9058), .ZN(n6426) );
  OR2_X1 U8020 ( .A1(n9060), .A2(n10569), .ZN(n6425) );
  NAND2_X1 U8021 ( .A1(n9867), .A2(n5987), .ZN(n6437) );
  NAND2_X1 U8022 ( .A1(n5991), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6435) );
  AND2_X1 U8023 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n6427), .ZN(n6428) );
  NAND2_X1 U8024 ( .A1(n6428), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6477) );
  INV_X1 U8025 ( .A(n6428), .ZN(n6430) );
  INV_X1 U8026 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U8027 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  NAND2_X1 U8028 ( .A1(n6478), .A2(n9582), .ZN(n6434) );
  NAND2_X1 U8029 ( .A1(n4514), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U8030 ( .A1(n4527), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6432) );
  INV_X1 U8031 ( .A(n9597), .ZN(n9776) );
  NAND2_X1 U8032 ( .A1(n9776), .A2(n6440), .ZN(n6436) );
  NAND2_X1 U8033 ( .A1(n6437), .A2(n6436), .ZN(n6439) );
  XNOR2_X1 U8034 ( .A(n6439), .B(n6438), .ZN(n6443) );
  NAND2_X1 U8035 ( .A1(n9867), .A2(n6440), .ZN(n6441) );
  OAI21_X1 U8036 ( .B1(n9597), .B2(n5918), .A(n6441), .ZN(n6442) );
  XNOR2_X1 U8037 ( .A(n6443), .B(n6442), .ZN(n6468) );
  INV_X1 U8038 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8039 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  NAND2_X1 U8040 ( .A1(n6446), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6448) );
  INV_X1 U8041 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6447) );
  XNOR2_X1 U8042 ( .A(n6448), .B(n6447), .ZN(n7020) );
  AND2_X1 U8043 ( .A1(n7018), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6987) );
  NAND2_X1 U8044 ( .A1(n7982), .A2(P1_B_REG_SCAN_IN), .ZN(n6449) );
  INV_X1 U8045 ( .A(n7934), .ZN(n6452) );
  MUX2_X1 U8046 ( .A(n6449), .B(P1_B_REG_SCAN_IN), .S(n6452), .Z(n6451) );
  NAND2_X1 U8047 ( .A1(n6451), .A2(n6450), .ZN(n6973) );
  INV_X1 U8048 ( .A(n6973), .ZN(n6571) );
  INV_X1 U8049 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10601) );
  NOR2_X1 U8050 ( .A1(n6450), .A2(n6452), .ZN(n6453) );
  AOI21_X1 U8051 ( .B1(n6571), .B2(n10601), .A(n6453), .ZN(n7507) );
  NAND2_X1 U8052 ( .A1(n9995), .A2(n7507), .ZN(n9994) );
  NOR4_X1 U8053 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6457) );
  NOR4_X1 U8054 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6456) );
  NOR4_X1 U8055 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6455) );
  NOR4_X1 U8056 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6454) );
  AND4_X1 U8057 ( .A1(n6457), .A2(n6456), .A3(n6455), .A4(n6454), .ZN(n6463)
         );
  NOR2_X1 U8058 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6461) );
  NOR4_X1 U8059 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6460) );
  NOR4_X1 U8060 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6459) );
  NOR4_X1 U8061 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6458) );
  AND4_X1 U8062 ( .A1(n6461), .A2(n6460), .A3(n6459), .A4(n6458), .ZN(n6462)
         );
  NAND2_X1 U8063 ( .A1(n6463), .A2(n6462), .ZN(n6570) );
  INV_X1 U8064 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10611) );
  NOR2_X1 U8065 ( .A1(n6570), .A2(n10611), .ZN(n6464) );
  INV_X1 U8066 ( .A(n6450), .ZN(n8057) );
  NAND2_X1 U8067 ( .A1(n8057), .A2(n7982), .ZN(n6974) );
  OAI21_X1 U8068 ( .B1(n6973), .B2(n6464), .A(n6974), .ZN(n7506) );
  OR2_X1 U8069 ( .A1(n9994), .A2(n7506), .ZN(n6476) );
  INV_X1 U8070 ( .A(n9335), .ZN(n9299) );
  INV_X1 U8071 ( .A(n9249), .ZN(n9066) );
  AND2_X1 U8072 ( .A1(n9299), .A2(n9066), .ZN(n6566) );
  NAND2_X1 U8073 ( .A1(n6465), .A2(n6566), .ZN(n10068) );
  NAND2_X1 U8074 ( .A1(n9335), .A2(n9249), .ZN(n6540) );
  NAND2_X1 U8075 ( .A1(n10068), .A2(n6540), .ZN(n6466) );
  INV_X1 U8076 ( .A(n6468), .ZN(n6486) );
  INV_X1 U8077 ( .A(n9219), .ZN(n9306) );
  NOR2_X1 U8078 ( .A1(n9215), .A2(n9306), .ZN(n10054) );
  NAND2_X1 U8079 ( .A1(n10054), .A2(n9066), .ZN(n6573) );
  INV_X1 U8080 ( .A(n9995), .ZN(n6469) );
  INV_X1 U8081 ( .A(n6566), .ZN(n7090) );
  OR2_X1 U8082 ( .A1(n7090), .A2(n9219), .ZN(n7511) );
  OR2_X1 U8083 ( .A1(n6476), .A2(n7511), .ZN(n6470) );
  INV_X1 U8084 ( .A(n6465), .ZN(n9301) );
  INV_X1 U8085 ( .A(n6540), .ZN(n9323) );
  INV_X1 U8086 ( .A(n9378), .ZN(n9382) );
  AND2_X2 U8087 ( .A1(n9323), .A2(n9382), .ZN(n10063) );
  NAND2_X1 U8088 ( .A1(n9301), .A2(n10063), .ZN(n6472) );
  OR2_X2 U8089 ( .A1(n6476), .A2(n6472), .ZN(n9029) );
  AND2_X1 U8090 ( .A1(n9306), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7601) );
  INV_X1 U8091 ( .A(n7507), .ZN(n6575) );
  OAI22_X1 U8092 ( .A1(n10068), .A2(n7601), .B1(n7506), .B2(n6575), .ZN(n6474)
         );
  NAND2_X1 U8093 ( .A1(n7020), .A2(n7018), .ZN(n6473) );
  AOI21_X1 U8094 ( .B1(n6465), .B2(n9323), .A(n6473), .ZN(n6569) );
  NAND2_X1 U8095 ( .A1(n6474), .A2(n6569), .ZN(n8972) );
  NAND2_X1 U8096 ( .A1(n8972), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9041) );
  AOI22_X1 U8097 ( .A1(n9033), .A2(n9582), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6484) );
  AND2_X1 U8098 ( .A1(n9323), .A2(n9378), .ZN(n10030) );
  INV_X1 U8099 ( .A(n10030), .ZN(n9968) );
  INV_X1 U8100 ( .A(n9968), .ZN(n10064) );
  NAND2_X1 U8101 ( .A1(n9301), .A2(n10064), .ZN(n6475) );
  INV_X1 U8102 ( .A(n9028), .ZN(n9037) );
  NAND2_X1 U8103 ( .A1(n6074), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6482) );
  INV_X1 U8104 ( .A(n6477), .ZN(n8306) );
  NAND2_X1 U8105 ( .A1(n6478), .A2(n8306), .ZN(n6481) );
  NAND2_X1 U8106 ( .A1(n4514), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8107 ( .A1(n4527), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6479) );
  NAND4_X1 U8108 ( .A1(n6482), .A2(n6481), .A3(n6480), .A4(n6479), .ZN(n9573)
         );
  NAND2_X1 U8109 ( .A1(n9037), .A2(n9573), .ZN(n6483) );
  OAI211_X1 U8110 ( .C1(n9608), .C2(n9029), .A(n6484), .B(n6483), .ZN(n6488)
         );
  NOR3_X1 U8111 ( .A1(n6486), .A2(n9046), .A3(n6485), .ZN(n6487) );
  AOI211_X1 U8112 ( .C1(n9867), .C2(n9051), .A(n6488), .B(n6487), .ZN(n6489)
         );
  INV_X1 U8113 ( .A(n6489), .ZN(n6490) );
  NAND2_X1 U8114 ( .A1(n6492), .A2(n6491), .ZN(P1_U3220) );
  NAND2_X1 U8115 ( .A1(n9998), .A2(n9748), .ZN(n7650) );
  NAND2_X1 U8116 ( .A1(n7649), .A2(n7650), .ZN(n6495) );
  NAND2_X1 U8117 ( .A1(n6495), .A2(n6494), .ZN(n7741) );
  NAND2_X1 U8118 ( .A1(n7646), .A2(n6496), .ZN(n6547) );
  NAND2_X1 U8119 ( .A1(n10012), .A2(n9997), .ZN(n7577) );
  NAND2_X1 U8120 ( .A1(n7741), .A2(n9064), .ZN(n6498) );
  NAND2_X1 U8121 ( .A1(n7646), .A2(n10012), .ZN(n6497) );
  NAND2_X1 U8122 ( .A1(n6498), .A2(n6497), .ZN(n7626) );
  INV_X1 U8123 ( .A(n7628), .ZN(n10019) );
  NAND2_X1 U8124 ( .A1(n10019), .A2(n9355), .ZN(n9113) );
  NAND2_X1 U8125 ( .A1(n7579), .A2(n7628), .ZN(n9255) );
  NAND2_X1 U8126 ( .A1(n9113), .A2(n9255), .ZN(n9068) );
  NAND2_X1 U8127 ( .A1(n7626), .A2(n9068), .ZN(n6500) );
  NAND2_X1 U8128 ( .A1(n10019), .A2(n7579), .ZN(n6499) );
  NAND2_X1 U8129 ( .A1(n6500), .A2(n6499), .ZN(n7581) );
  INV_X1 U8130 ( .A(n7583), .ZN(n10024) );
  NAND2_X1 U8131 ( .A1(n10024), .A2(n9354), .ZN(n9114) );
  NAND2_X1 U8132 ( .A1(n7583), .A2(n7384), .ZN(n9135) );
  NAND2_X1 U8133 ( .A1(n9114), .A2(n9135), .ZN(n9069) );
  NAND2_X1 U8134 ( .A1(n7581), .A2(n9069), .ZN(n6502) );
  NAND2_X1 U8135 ( .A1(n10024), .A2(n7384), .ZN(n6501) );
  NAND2_X1 U8136 ( .A1(n6502), .A2(n6501), .ZN(n7603) );
  NAND2_X1 U8137 ( .A1(n10031), .A2(n7580), .ZN(n9136) );
  NAND2_X1 U8138 ( .A1(n9258), .A2(n9136), .ZN(n7611) );
  OR2_X1 U8139 ( .A1(n10031), .A2(n9353), .ZN(n6503) );
  NAND2_X1 U8140 ( .A1(n10041), .A2(n9971), .ZN(n9261) );
  NAND2_X1 U8141 ( .A1(n9119), .A2(n9261), .ZN(n7654) );
  XNOR2_X1 U8142 ( .A(n9980), .B(n7594), .ZN(n9128) );
  NAND2_X1 U8143 ( .A1(n9972), .A2(n9128), .ZN(n6505) );
  OR2_X1 U8144 ( .A1(n9980), .A2(n9352), .ZN(n6504) );
  NOR2_X1 U8145 ( .A1(n9131), .A2(n9351), .ZN(n7391) );
  NAND2_X1 U8146 ( .A1(n9131), .A2(n9351), .ZN(n7389) );
  NAND2_X1 U8147 ( .A1(n7442), .A2(n7866), .ZN(n9148) );
  OR2_X1 U8148 ( .A1(n7442), .A2(n9350), .ZN(n6506) );
  OR2_X1 U8149 ( .A1(n7870), .A2(n7886), .ZN(n9263) );
  NAND2_X1 U8150 ( .A1(n7870), .A2(n7886), .ZN(n9153) );
  NAND2_X1 U8151 ( .A1(n9263), .A2(n9153), .ZN(n9079) );
  NAND2_X1 U8152 ( .A1(n7462), .A2(n9079), .ZN(n7461) );
  OR2_X1 U8153 ( .A1(n7870), .A2(n9349), .ZN(n6507) );
  NAND2_X1 U8154 ( .A1(n7461), .A2(n6507), .ZN(n7527) );
  OR2_X1 U8155 ( .A1(n7543), .A2(n7942), .ZN(n9154) );
  NAND2_X1 U8156 ( .A1(n7543), .A2(n7942), .ZN(n9155) );
  NAND2_X1 U8157 ( .A1(n9154), .A2(n9155), .ZN(n9063) );
  NAND2_X1 U8158 ( .A1(n7527), .A2(n9063), .ZN(n7526) );
  OR2_X1 U8159 ( .A1(n7543), .A2(n9348), .ZN(n6508) );
  NAND2_X1 U8160 ( .A1(n7526), .A2(n6508), .ZN(n7681) );
  OR2_X1 U8161 ( .A1(n7791), .A2(n8003), .ZN(n9156) );
  NAND2_X1 U8162 ( .A1(n7791), .A2(n8003), .ZN(n9269) );
  NAND2_X1 U8163 ( .A1(n9156), .A2(n9269), .ZN(n7680) );
  NAND2_X1 U8164 ( .A1(n7681), .A2(n7680), .ZN(n7679) );
  OR2_X1 U8165 ( .A1(n7791), .A2(n9347), .ZN(n6509) );
  OR2_X1 U8166 ( .A1(n7997), .A2(n8914), .ZN(n9274) );
  NAND2_X1 U8167 ( .A1(n7997), .A2(n8914), .ZN(n9270) );
  NAND2_X1 U8168 ( .A1(n9274), .A2(n9270), .ZN(n9083) );
  OR2_X1 U8169 ( .A1(n7997), .A2(n10062), .ZN(n6510) );
  NAND2_X1 U8170 ( .A1(n9111), .A2(n9346), .ZN(n6511) );
  NAND2_X1 U8171 ( .A1(n6512), .A2(n6511), .ZN(n7837) );
  INV_X1 U8172 ( .A(n7837), .ZN(n6513) );
  OR2_X1 U8173 ( .A1(n9927), .A2(n10065), .ZN(n6514) );
  INV_X1 U8174 ( .A(n9345), .ZN(n8973) );
  OR2_X1 U8175 ( .A1(n8964), .A2(n8973), .ZN(n9277) );
  NAND2_X1 U8176 ( .A1(n8964), .A2(n8973), .ZN(n9280) );
  NAND2_X1 U8177 ( .A1(n8964), .A2(n9345), .ZN(n6516) );
  OR2_X1 U8178 ( .A1(n8977), .A2(n9918), .ZN(n6517) );
  INV_X1 U8179 ( .A(n9730), .ZN(n6518) );
  OR2_X1 U8180 ( .A1(n9744), .A2(n9711), .ZN(n6519) );
  NAND2_X1 U8181 ( .A1(n6520), .A2(n6519), .ZN(n9705) );
  NOR2_X1 U8182 ( .A1(n9843), .A2(n9846), .ZN(n6521) );
  INV_X1 U8183 ( .A(n9846), .ZN(n9737) );
  INV_X1 U8184 ( .A(n9843), .ZN(n9720) );
  OR2_X1 U8185 ( .A1(n9698), .A2(n9828), .ZN(n6522) );
  NOR2_X1 U8186 ( .A1(n9688), .A2(n9817), .ZN(n6523) );
  INV_X1 U8187 ( .A(n9688), .ZN(n9896) );
  OR2_X1 U8188 ( .A1(n9670), .A2(n9827), .ZN(n6524) );
  NAND2_X1 U8189 ( .A1(n9670), .A2(n9827), .ZN(n6525) );
  INV_X1 U8190 ( .A(n9647), .ZN(n6526) );
  OR2_X1 U8191 ( .A1(n9656), .A2(n9816), .ZN(n6527) );
  NAND2_X1 U8192 ( .A1(n9636), .A2(n9806), .ZN(n6528) );
  NAND2_X1 U8193 ( .A1(n6529), .A2(n6528), .ZN(n9629) );
  AND2_X1 U8194 ( .A1(n9878), .A2(n9784), .ZN(n6530) );
  OAI22_X2 U8195 ( .A1(n9629), .A2(n6530), .B1(n9784), .B2(n9878), .ZN(n9615)
         );
  NOR2_X1 U8196 ( .A1(n9613), .A2(n9775), .ZN(n6531) );
  NAND2_X1 U8197 ( .A1(n9613), .A2(n9775), .ZN(n6532) );
  NAND2_X1 U8198 ( .A1(n9871), .A2(n9608), .ZN(n9205) );
  NAND2_X1 U8199 ( .A1(n9867), .A2(n9597), .ZN(n9206) );
  NAND2_X1 U8200 ( .A1(n9867), .A2(n9776), .ZN(n6534) );
  NAND2_X1 U8201 ( .A1(n9579), .A2(n6534), .ZN(n6539) );
  INV_X1 U8202 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8316) );
  OR2_X1 U8203 ( .A1(n9060), .A2(n8316), .ZN(n6536) );
  INV_X1 U8204 ( .A(n9573), .ZN(n6538) );
  OR2_X1 U8205 ( .A1(n8307), .A2(n6538), .ZN(n9291) );
  NAND2_X1 U8206 ( .A1(n8307), .A2(n6538), .ZN(n9316) );
  OR2_X1 U8207 ( .A1(n6465), .A2(n6540), .ZN(n6541) );
  NAND2_X1 U8208 ( .A1(n6541), .A2(n7090), .ZN(n9754) );
  INV_X1 U8209 ( .A(n9754), .ZN(n6544) );
  NAND2_X1 U8210 ( .A1(n6465), .A2(n6542), .ZN(n6543) );
  NAND2_X1 U8211 ( .A1(n6544), .A2(n6543), .ZN(n9996) );
  INV_X1 U8212 ( .A(n10054), .ZN(n10005) );
  NAND2_X1 U8213 ( .A1(n9996), .A2(n10005), .ZN(n10060) );
  NAND2_X1 U8214 ( .A1(n8312), .A2(n10060), .ZN(n6568) );
  INV_X1 U8215 ( .A(n9748), .ZN(n7091) );
  NOR2_X1 U8216 ( .A1(n7091), .A2(n9998), .ZN(n7638) );
  NAND2_X1 U8217 ( .A1(n7125), .A2(n5919), .ZN(n6545) );
  AND2_X1 U8218 ( .A1(n9113), .A2(n7577), .ZN(n9251) );
  AND2_X1 U8219 ( .A1(n9135), .A2(n9255), .ZN(n6548) );
  INV_X1 U8220 ( .A(n9114), .ZN(n9254) );
  INV_X1 U8221 ( .A(n9118), .ZN(n6549) );
  INV_X1 U8222 ( .A(n7611), .ZN(n9072) );
  NAND2_X1 U8223 ( .A1(n6549), .A2(n9072), .ZN(n7614) );
  NAND2_X1 U8224 ( .A1(n7614), .A2(n9258), .ZN(n7655) );
  NAND2_X1 U8225 ( .A1(n9131), .A2(n9969), .ZN(n9141) );
  NAND2_X1 U8226 ( .A1(n9980), .A2(n7594), .ZN(n9140) );
  NAND4_X1 U8227 ( .A1(n7655), .A2(n9074), .A3(n9148), .A4(n9261), .ZN(n6553)
         );
  OR2_X1 U8228 ( .A1(n9131), .A2(n9969), .ZN(n9122) );
  INV_X1 U8229 ( .A(n9074), .ZN(n6550) );
  NAND3_X1 U8230 ( .A1(n9151), .A2(n9122), .A3(n6550), .ZN(n6551) );
  NAND2_X1 U8231 ( .A1(n6551), .A2(n9148), .ZN(n9266) );
  OR2_X1 U8232 ( .A1(n9980), .A2(n7594), .ZN(n9124) );
  AND2_X1 U8233 ( .A1(n9122), .A2(n9124), .ZN(n9076) );
  AND3_X1 U8234 ( .A1(n9076), .A2(n9151), .A3(n9119), .ZN(n6552) );
  AND2_X1 U8235 ( .A1(n6553), .A2(n9264), .ZN(n7465) );
  INV_X1 U8236 ( .A(n9079), .ZN(n7464) );
  NAND2_X1 U8237 ( .A1(n7463), .A2(n9153), .ZN(n7523) );
  INV_X1 U8238 ( .A(n7680), .ZN(n9081) );
  INV_X1 U8239 ( .A(n9083), .ZN(n7761) );
  NAND2_X1 U8240 ( .A1(n7762), .A2(n7761), .ZN(n7760) );
  AND2_X1 U8241 ( .A1(n7760), .A2(n9274), .ZN(n7779) );
  XNOR2_X1 U8242 ( .A(n9111), .B(n9346), .ZN(n9161) );
  NAND2_X1 U8243 ( .A1(n7779), .A2(n9161), .ZN(n7778) );
  NAND2_X1 U8244 ( .A1(n9111), .A2(n9110), .ZN(n9163) );
  INV_X1 U8245 ( .A(n10065), .ZN(n8915) );
  OR2_X1 U8246 ( .A1(n9927), .A2(n8915), .ZN(n9276) );
  NAND2_X1 U8247 ( .A1(n9927), .A2(n8915), .ZN(n9164) );
  INV_X1 U8248 ( .A(n9918), .ZN(n9017) );
  OR2_X1 U8249 ( .A1(n8977), .A2(n9017), .ZN(n9724) );
  NAND2_X1 U8250 ( .A1(n8977), .A2(n9017), .ZN(n9171) );
  NAND2_X1 U8251 ( .A1(n9724), .A2(n9171), .ZN(n9087) );
  INV_X1 U8252 ( .A(n9280), .ZN(n6554) );
  NOR2_X1 U8253 ( .A1(n9087), .A2(n6554), .ZN(n6555) );
  INV_X1 U8254 ( .A(n9711), .ZN(n8933) );
  OR2_X1 U8255 ( .A1(n9744), .A2(n8933), .ZN(n9170) );
  NAND2_X1 U8256 ( .A1(n9744), .A2(n8933), .ZN(n9172) );
  NAND2_X1 U8257 ( .A1(n9170), .A2(n9172), .ZN(n9729) );
  INV_X1 U8258 ( .A(n9724), .ZN(n6556) );
  NOR2_X1 U8259 ( .A1(n9729), .A2(n6556), .ZN(n6557) );
  NAND2_X1 U8260 ( .A1(n9726), .A2(n9172), .ZN(n9706) );
  OR2_X1 U8261 ( .A1(n9843), .A2(n9737), .ZN(n9180) );
  NAND2_X1 U8262 ( .A1(n9843), .A2(n9737), .ZN(n9173) );
  NAND2_X1 U8263 ( .A1(n9180), .A2(n9173), .ZN(n9707) );
  OR2_X2 U8264 ( .A1(n9706), .A2(n9707), .ZN(n9708) );
  NAND2_X2 U8265 ( .A1(n9708), .A2(n9180), .ZN(n9692) );
  INV_X1 U8266 ( .A(n9828), .ZN(n8944) );
  OR2_X1 U8267 ( .A1(n9698), .A2(n8944), .ZN(n9185) );
  NAND2_X1 U8268 ( .A1(n9698), .A2(n8944), .ZN(n9183) );
  XNOR2_X1 U8269 ( .A(n9688), .B(n9817), .ZN(n9677) );
  NAND2_X1 U8270 ( .A1(n9688), .A2(n9184), .ZN(n9186) );
  XNOR2_X1 U8271 ( .A(n9670), .B(n9827), .ZN(n9661) );
  NAND2_X1 U8272 ( .A1(n9660), .A2(n9661), .ZN(n6558) );
  NAND2_X1 U8273 ( .A1(n9670), .A2(n9682), .ZN(n9103) );
  NAND2_X1 U8274 ( .A1(n6558), .A2(n9103), .ZN(n9645) );
  OR2_X1 U8275 ( .A1(n9656), .A2(n9666), .ZN(n9190) );
  NAND2_X1 U8276 ( .A1(n9656), .A2(n9666), .ZN(n9224) );
  OR2_X1 U8277 ( .A1(n9636), .A2(n9651), .ZN(n9227) );
  NAND2_X1 U8278 ( .A1(n9636), .A2(n9651), .ZN(n9233) );
  NAND2_X1 U8279 ( .A1(n9227), .A2(n9233), .ZN(n9640) );
  INV_X1 U8280 ( .A(n9784), .ZN(n9030) );
  NAND2_X1 U8281 ( .A1(n9878), .A2(n9030), .ZN(n9237) );
  NAND2_X1 U8282 ( .A1(n9619), .A2(n9628), .ZN(n9618) );
  NAND2_X1 U8283 ( .A1(n9618), .A2(n9245), .ZN(n9604) );
  XNOR2_X1 U8284 ( .A(n9613), .B(n9195), .ZN(n9614) );
  OR2_X2 U8285 ( .A1(n9604), .A2(n9614), .ZN(n9602) );
  NAND2_X1 U8286 ( .A1(n9613), .A2(n9195), .ZN(n9308) );
  NAND2_X1 U8287 ( .A1(n9602), .A2(n9308), .ZN(n9588) );
  XNOR2_X1 U8288 ( .A(n6559), .B(n9212), .ZN(n6565) );
  NAND2_X1 U8289 ( .A1(n9249), .A2(n9306), .ZN(n9334) );
  OAI21_X1 U8290 ( .B1(n9340), .B2(n9299), .A(n9334), .ZN(n9821) );
  INV_X1 U8291 ( .A(n9821), .ZN(n9849) );
  INV_X1 U8292 ( .A(n10063), .ZN(n9970) );
  INV_X1 U8293 ( .A(P1_B_REG_SCAN_IN), .ZN(n9298) );
  OR2_X1 U8294 ( .A1(n9300), .A2(n9298), .ZN(n6560) );
  NAND2_X1 U8295 ( .A1(n10030), .A2(n6560), .ZN(n9558) );
  NAND2_X1 U8296 ( .A1(n6074), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U8297 ( .A1(n4527), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U8298 ( .A1(n4514), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6561) );
  AND3_X1 U8299 ( .A1(n6563), .A2(n6562), .A3(n6561), .ZN(n9099) );
  OAI22_X1 U8300 ( .A1(n9597), .A2(n9970), .B1(n9558), .B2(n9099), .ZN(n6564)
         );
  INV_X1 U8301 ( .A(n9867), .ZN(n9581) );
  INV_X1 U8302 ( .A(n9878), .ZN(n9626) );
  INV_X1 U8303 ( .A(n9670), .ZN(n9892) );
  INV_X1 U8304 ( .A(n9744), .ZN(n9905) );
  INV_X1 U8305 ( .A(n9111), .ZN(n10069) );
  INV_X1 U8306 ( .A(n7543), .ZN(n7891) );
  INV_X1 U8307 ( .A(n9980), .ZN(n10049) );
  INV_X1 U8308 ( .A(n7870), .ZN(n7472) );
  OR2_X2 U8309 ( .A1(n8964), .A2(n7912), .ZN(n7988) );
  NOR2_X2 U8310 ( .A1(n9688), .A2(n9683), .ZN(n9684) );
  NOR2_X2 U8311 ( .A1(n9871), .A2(n9609), .ZN(n9593) );
  NAND2_X1 U8312 ( .A1(n6566), .A2(n9219), .ZN(n9715) );
  AOI21_X1 U8313 ( .B1(n8307), .B2(n9580), .A(n9715), .ZN(n6567) );
  NAND2_X1 U8314 ( .A1(n6567), .A2(n9563), .ZN(n8310) );
  AND2_X1 U8315 ( .A1(n6569), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7509) );
  NAND2_X1 U8316 ( .A1(n6571), .A2(n10611), .ZN(n6572) );
  AOI22_X1 U8317 ( .A1(n6572), .A2(n6974), .B1(n6571), .B2(n6570), .ZN(n6574)
         );
  NAND3_X1 U8318 ( .A1(n7509), .A2(n6574), .A3(n6573), .ZN(n6724) );
  INV_X2 U8319 ( .A(n10092), .ZN(n10094) );
  INV_X1 U8320 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6576) );
  NOR2_X1 U8321 ( .A1(n10094), .A2(n6576), .ZN(n6577) );
  NOR2_X1 U8322 ( .A1(n10092), .A2(n10068), .ZN(n9798) );
  NAND2_X1 U8323 ( .A1(n7176), .A2(n6948), .ZN(n6580) );
  NAND2_X1 U8324 ( .A1(n6580), .A2(n6673), .ZN(n6610) );
  NAND2_X1 U8325 ( .A1(n6610), .A2(n6678), .ZN(n6581) );
  NAND2_X1 U8326 ( .A1(n6581), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8327 ( .A(n6997), .ZN(n7174) );
  INV_X1 U8328 ( .A(n8582), .ZN(n7265) );
  INV_X1 U8329 ( .A(n8549), .ZN(n7148) );
  INV_X1 U8330 ( .A(n8119), .ZN(n7096) );
  NAND2_X1 U8331 ( .A1(n5345), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8332 ( .A1(n6583), .A2(n6584), .ZN(n8205) );
  INV_X1 U8333 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U8334 ( .A1(n10111), .A2(n10112), .ZN(n10110) );
  INV_X1 U8335 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6585) );
  XNOR2_X1 U8336 ( .A(n6690), .B(n6585), .ZN(n7236) );
  AOI21_X1 U8337 ( .B1(n7235), .B2(n7237), .A(n7236), .ZN(n7234) );
  NOR2_X1 U8338 ( .A1(n7234), .A2(n6586), .ZN(n6587) );
  NAND2_X1 U8339 ( .A1(n6979), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6590) );
  OR2_X1 U8340 ( .A1(n6979), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6589) );
  NAND2_X1 U8341 ( .A1(n6590), .A2(n6589), .ZN(n7365) );
  INV_X1 U8342 ( .A(n6590), .ZN(n6591) );
  INV_X1 U8343 ( .A(n7733), .ZN(n7007) );
  NAND2_X1 U8344 ( .A1(n7007), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8345 ( .A1(n7733), .A2(n6593), .ZN(n6594) );
  NAND2_X1 U8346 ( .A1(n6595), .A2(n6594), .ZN(n7727) );
  XNOR2_X1 U8347 ( .A(n6596), .B(n7905), .ZN(n7893) );
  MUX2_X1 U8348 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10208), .S(n7978), .Z(n7964) );
  NOR2_X1 U8349 ( .A1(n8020), .A2(n6598), .ZN(n6599) );
  NOR2_X1 U8350 ( .A1(n8011), .A2(n5486), .ZN(n8010) );
  MUX2_X1 U8351 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6624), .S(n8119), .Z(n8105)
         );
  NOR2_X1 U8352 ( .A1(n8532), .A2(n6600), .ZN(n6601) );
  XNOR2_X1 U8353 ( .A(n8549), .B(n8155), .ZN(n8536) );
  XNOR2_X1 U8354 ( .A(n8582), .B(n8171), .ZN(n8569) );
  NOR2_X1 U8355 ( .A1(n8597), .A2(n6605), .ZN(n6606) );
  INV_X1 U8356 ( .A(n8617), .ZN(n8607) );
  NAND2_X1 U8357 ( .A1(n8607), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6607) );
  OAI21_X1 U8358 ( .B1(n8607), .B2(P2_REG1_REG_18__SCAN_IN), .A(n6607), .ZN(
        n8601) );
  INV_X1 U8359 ( .A(n6607), .ZN(n6608) );
  XNOR2_X1 U8360 ( .A(n7547), .B(n8820), .ZN(n6669) );
  XNOR2_X1 U8361 ( .A(n6609), .B(n6669), .ZN(n6611) );
  NAND2_X1 U8362 ( .A1(n6610), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6719) );
  OR2_X1 U8363 ( .A1(n6719), .A2(n5772), .ZN(n7114) );
  OR2_X1 U8364 ( .A1(n7114), .A2(n6925), .ZN(n8618) );
  INV_X2 U8365 ( .A(n6925), .ZN(n6638) );
  INV_X2 U8366 ( .A(n6925), .ZN(n8321) );
  NOR2_X1 U8367 ( .A1(n8321), .A2(n8778), .ZN(n6612) );
  AOI21_X1 U8368 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n6638), .A(n6612), .ZN(
        n6666) );
  XOR2_X1 U8369 ( .A(n8597), .B(n6666), .Z(n8589) );
  MUX2_X1 U8370 ( .A(n8175), .B(n8171), .S(n6638), .Z(n6613) );
  NAND2_X1 U8371 ( .A1(n8582), .A2(n6613), .ZN(n6664) );
  XNOR2_X1 U8372 ( .A(n6613), .B(n7265), .ZN(n8572) );
  INV_X1 U8373 ( .A(n6708), .ZN(n8562) );
  OR2_X1 U8374 ( .A1(n6638), .A2(n6614), .ZN(n6616) );
  NAND2_X1 U8375 ( .A1(n8321), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U8376 ( .A1(n6616), .A2(n6615), .ZN(n6617) );
  OR2_X1 U8377 ( .A1(n8562), .A2(n6617), .ZN(n6663) );
  XNOR2_X1 U8378 ( .A(n6708), .B(n6617), .ZN(n8556) );
  OR2_X1 U8379 ( .A1(n6638), .A2(n6618), .ZN(n6620) );
  NAND2_X1 U8380 ( .A1(n8321), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U8381 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  OR2_X1 U8382 ( .A1(n7148), .A2(n6621), .ZN(n6662) );
  XNOR2_X1 U8383 ( .A(n6621), .B(n8549), .ZN(n8539) );
  MUX2_X1 U8384 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8321), .Z(n6623) );
  INV_X1 U8385 ( .A(n6623), .ZN(n6622) );
  NAND2_X1 U8386 ( .A1(n8532), .A2(n6622), .ZN(n6661) );
  XNOR2_X1 U8387 ( .A(n6623), .B(n8532), .ZN(n8526) );
  MUX2_X1 U8388 ( .A(n8129), .B(n6624), .S(n8321), .Z(n6625) );
  NAND2_X1 U8389 ( .A1(n8119), .A2(n6625), .ZN(n6660) );
  XNOR2_X1 U8390 ( .A(n6625), .B(n7096), .ZN(n8109) );
  MUX2_X1 U8391 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n6638), .Z(n6627) );
  INV_X1 U8392 ( .A(n6627), .ZN(n6626) );
  NAND2_X1 U8393 ( .A1(n8020), .A2(n6626), .ZN(n6659) );
  XNOR2_X1 U8394 ( .A(n6627), .B(n8020), .ZN(n8014) );
  MUX2_X1 U8395 ( .A(n7956), .B(n10208), .S(n8321), .Z(n6628) );
  NAND2_X1 U8396 ( .A1(n7978), .A2(n6628), .ZN(n6658) );
  XNOR2_X1 U8397 ( .A(n6628), .B(n7067), .ZN(n7968) );
  MUX2_X1 U8398 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6638), .Z(n6630) );
  INV_X1 U8399 ( .A(n6630), .ZN(n6629) );
  NAND2_X1 U8400 ( .A1(n7905), .A2(n6629), .ZN(n6657) );
  XNOR2_X1 U8401 ( .A(n6630), .B(n7905), .ZN(n7896) );
  MUX2_X1 U8402 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8321), .Z(n6655) );
  OR2_X1 U8403 ( .A1(n7007), .A2(n6655), .ZN(n6656) );
  INV_X1 U8404 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6631) );
  OR2_X1 U8405 ( .A1(n8321), .A2(n6631), .ZN(n6633) );
  NAND2_X1 U8406 ( .A1(n6638), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U8407 ( .A1(n6633), .A2(n6632), .ZN(n6652) );
  INV_X1 U8408 ( .A(n6652), .ZN(n6653) );
  INV_X1 U8409 ( .A(n6979), .ZN(n7376) );
  MUX2_X1 U8410 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6638), .Z(n6650) );
  INV_X1 U8411 ( .A(n6650), .ZN(n6651) );
  MUX2_X1 U8412 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8321), .Z(n6648) );
  INV_X1 U8413 ( .A(n6648), .ZN(n6649) );
  MUX2_X1 U8414 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6638), .Z(n6646) );
  INV_X1 U8415 ( .A(n6646), .ZN(n6647) );
  MUX2_X1 U8416 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6638), .Z(n6643) );
  INV_X1 U8417 ( .A(n6643), .ZN(n6644) );
  OR2_X1 U8418 ( .A1(n8321), .A2(n6634), .ZN(n6636) );
  NAND2_X1 U8419 ( .A1(n6638), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U8420 ( .A1(n6636), .A2(n6635), .ZN(n6641) );
  OR2_X1 U8421 ( .A1(n6638), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U8422 ( .A1(n8321), .A2(n6582), .ZN(n6639) );
  NAND2_X1 U8423 ( .A1(n6640), .A2(n6639), .ZN(n7115) );
  NAND2_X1 U8424 ( .A1(n8213), .A2(n8212), .ZN(n8211) );
  NAND2_X1 U8425 ( .A1(n6641), .A2(n6685), .ZN(n6642) );
  NAND2_X1 U8426 ( .A1(n8211), .A2(n6642), .ZN(n10098) );
  XNOR2_X1 U8427 ( .A(n6643), .B(n6645), .ZN(n10097) );
  NAND2_X1 U8428 ( .A1(n10098), .A2(n10097), .ZN(n10096) );
  OAI21_X1 U8429 ( .B1(n6645), .B2(n6644), .A(n10096), .ZN(n7133) );
  XNOR2_X1 U8430 ( .A(n6646), .B(n6963), .ZN(n7134) );
  NOR2_X1 U8431 ( .A1(n7133), .A2(n7134), .ZN(n7132) );
  AOI21_X1 U8432 ( .B1(n4833), .B2(n6647), .A(n7132), .ZN(n7233) );
  XNOR2_X1 U8433 ( .A(n6648), .B(n6690), .ZN(n7232) );
  NAND2_X1 U8434 ( .A1(n7233), .A2(n7232), .ZN(n7231) );
  OAI21_X1 U8435 ( .B1(n6690), .B2(n6649), .A(n7231), .ZN(n7282) );
  XNOR2_X1 U8436 ( .A(n6650), .B(n6971), .ZN(n7281) );
  NAND2_X1 U8437 ( .A1(n7282), .A2(n7281), .ZN(n7280) );
  OAI21_X1 U8438 ( .B1(n6971), .B2(n6651), .A(n7280), .ZN(n7362) );
  XNOR2_X1 U8439 ( .A(n6652), .B(n6979), .ZN(n7363) );
  NOR2_X1 U8440 ( .A1(n7362), .A2(n7363), .ZN(n7361) );
  AOI21_X1 U8441 ( .B1(n6653), .B2(n7376), .A(n7361), .ZN(n7561) );
  MUX2_X1 U8442 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8321), .Z(n6654) );
  XNOR2_X1 U8443 ( .A(n6654), .B(n6983), .ZN(n7560) );
  OAI22_X1 U8444 ( .A1(n7561), .A2(n7560), .B1(n6654), .B2(n6983), .ZN(n7723)
         );
  XNOR2_X1 U8445 ( .A(n6655), .B(n7733), .ZN(n7724) );
  NAND2_X1 U8446 ( .A1(n7723), .A2(n7724), .ZN(n7722) );
  NAND2_X1 U8447 ( .A1(n6656), .A2(n7722), .ZN(n7895) );
  NAND2_X1 U8448 ( .A1(n7896), .A2(n7895), .ZN(n7894) );
  NAND2_X1 U8449 ( .A1(n6657), .A2(n7894), .ZN(n7967) );
  NAND2_X1 U8450 ( .A1(n7968), .A2(n7967), .ZN(n7966) );
  NAND2_X1 U8451 ( .A1(n6658), .A2(n7966), .ZN(n8013) );
  NAND2_X1 U8452 ( .A1(n8014), .A2(n8013), .ZN(n8012) );
  NAND2_X1 U8453 ( .A1(n6659), .A2(n8012), .ZN(n8108) );
  NAND2_X1 U8454 ( .A1(n8109), .A2(n8108), .ZN(n8107) );
  NAND2_X1 U8455 ( .A1(n6660), .A2(n8107), .ZN(n8525) );
  NAND2_X1 U8456 ( .A1(n8526), .A2(n8525), .ZN(n8524) );
  NAND2_X1 U8457 ( .A1(n6661), .A2(n8524), .ZN(n8538) );
  NAND2_X1 U8458 ( .A1(n8539), .A2(n8538), .ZN(n8537) );
  NAND2_X1 U8459 ( .A1(n6662), .A2(n8537), .ZN(n8555) );
  NAND2_X1 U8460 ( .A1(n8556), .A2(n8555), .ZN(n8554) );
  NAND2_X1 U8461 ( .A1(n6663), .A2(n8554), .ZN(n8571) );
  NAND2_X1 U8462 ( .A1(n8572), .A2(n8571), .ZN(n8570) );
  NAND2_X1 U8463 ( .A1(n6664), .A2(n8570), .ZN(n8588) );
  NAND2_X1 U8464 ( .A1(n8589), .A2(n8588), .ZN(n8587) );
  INV_X1 U8465 ( .A(n8587), .ZN(n6665) );
  AOI21_X1 U8466 ( .B1(n6666), .B2(n8597), .A(n6665), .ZN(n6668) );
  MUX2_X1 U8467 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8321), .Z(n6667) );
  NOR2_X1 U8468 ( .A1(n6668), .A2(n6667), .ZN(n8603) );
  NAND2_X1 U8469 ( .A1(n6668), .A2(n6667), .ZN(n8604) );
  OAI21_X1 U8470 ( .B1(n8603), .B2(n8617), .A(n8604), .ZN(n6671) );
  MUX2_X1 U8471 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8749), .S(n7547), .Z(n6715)
         );
  MUX2_X1 U8472 ( .A(n6669), .B(n6715), .S(n6925), .Z(n6670) );
  XNOR2_X1 U8473 ( .A(n6671), .B(n6670), .ZN(n6676) );
  OR2_X1 U8474 ( .A1(n8606), .A2(n6672), .ZN(n7378) );
  NAND2_X1 U8475 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8385) );
  INV_X1 U8476 ( .A(n6673), .ZN(n7152) );
  NOR2_X1 U8477 ( .A1(n7176), .A2(n7152), .ZN(n6674) );
  OR2_X1 U8478 ( .A1(P2_U3150), .A2(n6674), .ZN(n8611) );
  INV_X1 U8479 ( .A(n8611), .ZN(n10105) );
  NAND2_X1 U8480 ( .A1(n10105), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n6675) );
  OAI211_X1 U8481 ( .C1(n6676), .C2(n7378), .A(n8385), .B(n6675), .ZN(n6682)
         );
  INV_X1 U8482 ( .A(n6719), .ZN(n6677) );
  MUX2_X1 U8483 ( .A(P2_U3893), .B(n6677), .S(n5772), .Z(n6679) );
  AND2_X1 U8484 ( .A1(n6679), .A2(n6678), .ZN(n8596) );
  NOR2_X1 U8485 ( .A1(n6680), .A2(n7547), .ZN(n6681) );
  NOR2_X1 U8486 ( .A1(n6682), .A2(n6681), .ZN(n6722) );
  NAND2_X1 U8487 ( .A1(n5345), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U8488 ( .A1(n4837), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6687) );
  NOR2_X1 U8489 ( .A1(n5355), .A2(n7136), .ZN(n7135) );
  INV_X1 U8490 ( .A(n7135), .ZN(n7243) );
  XNOR2_X1 U8491 ( .A(n6690), .B(n7488), .ZN(n7242) );
  AOI21_X1 U8492 ( .B1(n7243), .B2(n7241), .A(n7242), .ZN(n7245) );
  NOR2_X1 U8493 ( .A1(n7245), .A2(n6691), .ZN(n6692) );
  NAND2_X1 U8494 ( .A1(n6979), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6696) );
  OR2_X1 U8495 ( .A1(n6979), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U8496 ( .A1(n6696), .A2(n6695), .ZN(n7368) );
  INV_X1 U8497 ( .A(n6696), .ZN(n6697) );
  NOR2_X1 U8498 ( .A1(n7570), .A2(n6698), .ZN(n6699) );
  XNOR2_X1 U8499 ( .A(n6698), .B(n7570), .ZN(n7566) );
  NAND2_X1 U8500 ( .A1(n7007), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6702) );
  INV_X1 U8501 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6700) );
  NAND2_X1 U8502 ( .A1(n7733), .A2(n6700), .ZN(n6701) );
  NAND2_X1 U8503 ( .A1(n6702), .A2(n6701), .ZN(n7720) );
  NOR2_X1 U8504 ( .A1(n7905), .A2(n6703), .ZN(n6704) );
  NOR2_X1 U8505 ( .A1(n5446), .A2(n7901), .ZN(n7900) );
  NOR2_X1 U8506 ( .A1(n6704), .A2(n7900), .ZN(n7974) );
  AOI22_X1 U8507 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7978), .B1(n7067), .B2(
        n7956), .ZN(n7973) );
  NOR2_X1 U8508 ( .A1(n7974), .A2(n7973), .ZN(n7972) );
  NOR2_X1 U8509 ( .A1(n8020), .A2(n6705), .ZN(n6706) );
  AOI22_X1 U8510 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8119), .B1(n7096), .B2(
        n8129), .ZN(n8115) );
  AOI22_X1 U8511 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8549), .B1(n7148), .B2(
        n6618), .ZN(n8544) );
  NOR2_X1 U8512 ( .A1(n6708), .A2(n6709), .ZN(n6710) );
  AOI22_X1 U8513 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8582), .B1(n7265), .B2(
        n8175), .ZN(n8577) );
  NOR2_X1 U8514 ( .A1(n8597), .A2(n6711), .ZN(n6712) );
  NAND2_X1 U8515 ( .A1(n8607), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6713) );
  OAI21_X1 U8516 ( .B1(n8607), .B2(P2_REG2_REG_18__SCAN_IN), .A(n6713), .ZN(
        n8613) );
  INV_X1 U8517 ( .A(n6713), .ZN(n6714) );
  INV_X1 U8518 ( .A(n6715), .ZN(n6716) );
  XNOR2_X1 U8519 ( .A(n6717), .B(n6716), .ZN(n6721) );
  NAND3_X1 U8520 ( .A1(n6723), .A2(n6722), .A3(n5158), .ZN(P2_U3201) );
  INV_X2 U8521 ( .A(n10076), .ZN(n10078) );
  INV_X1 U8522 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6726) );
  NOR2_X1 U8523 ( .A1(n10076), .A2(n10068), .ZN(n9879) );
  MUX2_X1 U8524 ( .A(n8646), .B(n8843), .S(n6948), .Z(n6859) );
  XNOR2_X1 U8525 ( .A(n6728), .B(n6952), .ZN(n6798) );
  INV_X1 U8526 ( .A(n7308), .ZN(n7191) );
  NAND2_X1 U8527 ( .A1(n6896), .A2(n7175), .ZN(n6729) );
  NAND2_X1 U8528 ( .A1(n6729), .A2(n6948), .ZN(n6731) );
  NAND3_X1 U8529 ( .A1(n6896), .A2(n6732), .A3(n6945), .ZN(n6730) );
  NAND2_X1 U8530 ( .A1(n6741), .A2(n6733), .ZN(n6736) );
  NAND2_X1 U8531 ( .A1(n6747), .A2(n6734), .ZN(n6735) );
  MUX2_X1 U8532 ( .A(n6736), .B(n6735), .S(n6948), .Z(n6737) );
  INV_X1 U8533 ( .A(n6737), .ZN(n6738) );
  NAND2_X1 U8534 ( .A1(n6739), .A2(n6738), .ZN(n6740) );
  NAND2_X1 U8535 ( .A1(n6740), .A2(n7485), .ZN(n6750) );
  INV_X1 U8536 ( .A(n6741), .ZN(n6743) );
  OAI21_X1 U8537 ( .B1(n6750), .B2(n6743), .A(n6742), .ZN(n6746) );
  INV_X1 U8538 ( .A(n6744), .ZN(n6745) );
  INV_X1 U8539 ( .A(n6747), .ZN(n7477) );
  NAND2_X1 U8540 ( .A1(n7666), .A2(n10147), .ZN(n6748) );
  OAI211_X1 U8541 ( .C1(n6750), .C2(n7477), .A(n6749), .B(n6748), .ZN(n6754)
         );
  NAND2_X1 U8542 ( .A1(n10126), .A2(n6751), .ZN(n6752) );
  NAND2_X1 U8543 ( .A1(n6759), .A2(n6755), .ZN(n6757) );
  NAND2_X1 U8544 ( .A1(n6763), .A2(n6762), .ZN(n6756) );
  MUX2_X1 U8545 ( .A(n6757), .B(n6756), .S(n6948), .Z(n6765) );
  NOR2_X1 U8546 ( .A1(n6765), .A2(n7814), .ZN(n6758) );
  OAI211_X1 U8547 ( .C1(n6765), .C2(n6760), .A(n8073), .B(n6759), .ZN(n6767)
         );
  AND2_X1 U8548 ( .A1(n6762), .A2(n6761), .ZN(n6764) );
  OAI211_X1 U8549 ( .C1(n6765), .C2(n6764), .A(n6763), .B(n8048), .ZN(n6766)
         );
  MUX2_X1 U8550 ( .A(n6767), .B(n6766), .S(n6952), .Z(n6768) );
  INV_X1 U8551 ( .A(n6768), .ZN(n6769) );
  NAND3_X1 U8552 ( .A1(n6771), .A2(n8048), .A3(n6774), .ZN(n6770) );
  NAND2_X1 U8553 ( .A1(n6770), .A2(n6772), .ZN(n6777) );
  NAND2_X1 U8554 ( .A1(n6771), .A2(n8073), .ZN(n6775) );
  INV_X1 U8555 ( .A(n6772), .ZN(n6773) );
  AOI21_X1 U8556 ( .B1(n6775), .B2(n6774), .A(n6773), .ZN(n6776) );
  MUX2_X1 U8557 ( .A(n6777), .B(n6776), .S(n6952), .Z(n6782) );
  AND2_X1 U8558 ( .A1(n10194), .A2(n6948), .ZN(n6779) );
  NOR2_X1 U8559 ( .A1(n10194), .A2(n6948), .ZN(n6778) );
  MUX2_X1 U8560 ( .A(n6779), .B(n6778), .S(n8507), .Z(n6780) );
  INV_X1 U8561 ( .A(n6780), .ZN(n6781) );
  OAI21_X1 U8562 ( .B1(n6782), .B2(n8124), .A(n6781), .ZN(n6784) );
  MUX2_X1 U8563 ( .A(n8194), .B(n8226), .S(n6948), .Z(n6786) );
  NAND2_X1 U8564 ( .A1(n6788), .A2(n6787), .ZN(n8149) );
  MUX2_X1 U8565 ( .A(n6788), .B(n6787), .S(n6948), .Z(n6789) );
  INV_X1 U8566 ( .A(n6790), .ZN(n6794) );
  AND2_X1 U8567 ( .A1(n6794), .A2(n6791), .ZN(n8141) );
  INV_X1 U8568 ( .A(n6907), .ZN(n8165) );
  NAND3_X1 U8569 ( .A1(n6795), .A2(n8165), .A3(n6791), .ZN(n6797) );
  INV_X1 U8570 ( .A(n6792), .ZN(n6793) );
  AOI211_X1 U8571 ( .C1(n6795), .C2(n6794), .A(n6952), .B(n6793), .ZN(n6796)
         );
  AOI211_X1 U8572 ( .C1(n6798), .C2(n6797), .A(n8781), .B(n6796), .ZN(n6807)
         );
  NAND2_X1 U8573 ( .A1(n6805), .A2(n6799), .ZN(n6800) );
  OAI211_X1 U8574 ( .C1(n6807), .C2(n6800), .A(n6804), .B(n8697), .ZN(n6802)
         );
  NAND3_X1 U8575 ( .A1(n6802), .A2(n8699), .A3(n6801), .ZN(n6810) );
  NAND2_X1 U8576 ( .A1(n6804), .A2(n6803), .ZN(n6806) );
  OAI211_X1 U8577 ( .C1(n6807), .C2(n6806), .A(n8739), .B(n6805), .ZN(n6808)
         );
  NAND2_X1 U8578 ( .A1(n6808), .A2(n8697), .ZN(n6809) );
  MUX2_X1 U8579 ( .A(n6810), .B(n6809), .S(n6952), .Z(n6814) );
  INV_X1 U8580 ( .A(n8720), .ZN(n6813) );
  AND2_X1 U8581 ( .A1(n8699), .A2(n8701), .ZN(n6811) );
  MUX2_X1 U8582 ( .A(n6811), .B(n8700), .S(n6948), .Z(n6812) );
  OAI21_X1 U8583 ( .B1(n6814), .B2(n6813), .A(n6812), .ZN(n6817) );
  MUX2_X1 U8584 ( .A(n8701), .B(n6815), .S(n6952), .Z(n6816) );
  NAND3_X1 U8585 ( .A1(n6817), .A2(n8705), .A3(n6816), .ZN(n6832) );
  INV_X1 U8586 ( .A(n6826), .ZN(n6822) );
  NAND2_X1 U8587 ( .A1(n6823), .A2(n6818), .ZN(n6820) );
  MUX2_X1 U8588 ( .A(n6820), .B(n6819), .S(n6952), .Z(n6821) );
  NOR3_X1 U8589 ( .A1(n8674), .A2(n6894), .A3(n6821), .ZN(n6831) );
  INV_X1 U8590 ( .A(n6825), .ZN(n6824) );
  AOI21_X1 U8591 ( .B1(n6824), .B2(n6823), .A(n6822), .ZN(n6829) );
  AOI21_X1 U8592 ( .B1(n6827), .B2(n6826), .A(n6825), .ZN(n6828) );
  MUX2_X1 U8593 ( .A(n6829), .B(n6828), .S(n6948), .Z(n6830) );
  AOI211_X1 U8594 ( .C1(n6832), .C2(n6831), .A(n6830), .B(n8667), .ZN(n6841)
         );
  MUX2_X1 U8595 ( .A(n6834), .B(n6833), .S(n6948), .Z(n6835) );
  NAND2_X1 U8596 ( .A1(n6835), .A2(n8656), .ZN(n6840) );
  NAND2_X1 U8597 ( .A1(n6836), .A2(n8664), .ZN(n6837) );
  MUX2_X1 U8598 ( .A(n6838), .B(n6837), .S(n6952), .Z(n6839) );
  INV_X1 U8599 ( .A(n6842), .ZN(n6844) );
  NOR2_X1 U8600 ( .A1(n8360), .A2(n8633), .ZN(n6843) );
  MUX2_X1 U8601 ( .A(n6844), .B(n6843), .S(n6952), .Z(n6845) );
  MUX2_X1 U8602 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n5176), .Z(n6865) );
  XNOR2_X1 U8603 ( .A(n6865), .B(SI_30_), .ZN(n6866) );
  NAND2_X1 U8604 ( .A1(n9059), .A2(n6875), .ZN(n6853) );
  INV_X1 U8605 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6851) );
  OR2_X1 U8606 ( .A1(n6873), .A2(n6851), .ZN(n6852) );
  INV_X1 U8607 ( .A(n8498), .ZN(n6855) );
  NAND2_X1 U8608 ( .A1(n8838), .A2(n6855), .ZN(n6917) );
  AND2_X1 U8609 ( .A1(n6917), .A2(n6854), .ZN(n6887) );
  OAI21_X1 U8610 ( .B1(n6856), .B2(n8646), .A(n6887), .ZN(n6858) );
  MUX2_X1 U8611 ( .A(n6858), .B(n6857), .S(n6952), .Z(n6862) );
  AND2_X1 U8612 ( .A1(n6860), .A2(n6859), .ZN(n6861) );
  INV_X1 U8613 ( .A(n6918), .ZN(n6863) );
  AOI21_X1 U8614 ( .B1(n6952), .B2(n6917), .A(n6863), .ZN(n6864) );
  MUX2_X1 U8615 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5176), .Z(n6869) );
  INV_X1 U8616 ( .A(SI_31_), .ZN(n6868) );
  XNOR2_X1 U8617 ( .A(n6869), .B(n6868), .ZN(n6870) );
  INV_X1 U8618 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6872) );
  NOR2_X1 U8619 ( .A1(n6873), .A2(n6872), .ZN(n6874) );
  INV_X1 U8620 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U8621 ( .A1(n6876), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6879) );
  INV_X1 U8622 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6877) );
  OR2_X1 U8623 ( .A1(n5339), .A2(n6877), .ZN(n6878) );
  OAI211_X1 U8624 ( .C1(n6881), .C2(n6880), .A(n6879), .B(n6878), .ZN(n6882)
         );
  INV_X1 U8625 ( .A(n6882), .ZN(n6883) );
  NAND2_X1 U8626 ( .A1(n6884), .A2(n6883), .ZN(n8622) );
  AND2_X1 U8627 ( .A1(n8625), .A2(n8622), .ZN(n6889) );
  INV_X1 U8628 ( .A(n8622), .ZN(n6885) );
  INV_X1 U8629 ( .A(n8838), .ZN(n8628) );
  INV_X1 U8630 ( .A(n6889), .ZN(n6920) );
  OAI211_X1 U8631 ( .C1(n8628), .C2(n8834), .A(n6890), .B(n6920), .ZN(n6892)
         );
  NAND2_X1 U8632 ( .A1(n6892), .A2(n6891), .ZN(n6924) );
  NOR2_X1 U8633 ( .A1(n6894), .A2(n6893), .ZN(n8689) );
  INV_X1 U8634 ( .A(n6895), .ZN(n8722) );
  INV_X1 U8635 ( .A(n8141), .ZN(n8135) );
  AND2_X1 U8636 ( .A1(n7341), .A2(n6896), .ZN(n7299) );
  AND2_X1 U8637 ( .A1(n7332), .A2(n7299), .ZN(n6900) );
  NOR2_X1 U8638 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  XNOR2_X1 U8639 ( .A(n7693), .B(n7555), .ZN(n7664) );
  NAND4_X1 U8640 ( .A1(n6900), .A2(n6899), .A3(n7485), .A4(n7664), .ZN(n6901)
         );
  XNOR2_X1 U8641 ( .A(n10157), .B(n8512), .ZN(n10128) );
  NOR4_X1 U8642 ( .A1(n6901), .A2(n10128), .A3(n7857), .A4(n7814), .ZN(n6903)
         );
  NAND4_X1 U8643 ( .A1(n8077), .A2(n6903), .A3(n7951), .A4(n5745), .ZN(n6904)
         );
  NOR2_X1 U8644 ( .A1(n8124), .A2(n6904), .ZN(n6905) );
  XNOR2_X1 U8645 ( .A(n8237), .B(n8506), .ZN(n8184) );
  NAND3_X1 U8646 ( .A1(n4803), .A2(n6905), .A3(n8184), .ZN(n6906) );
  OR3_X1 U8647 ( .A1(n6907), .A2(n8135), .A3(n6906), .ZN(n6908) );
  NOR2_X1 U8648 ( .A1(n8781), .A2(n6908), .ZN(n6909) );
  NAND3_X1 U8649 ( .A1(n8739), .A2(n8755), .A3(n6909), .ZN(n6910) );
  NOR2_X1 U8650 ( .A1(n8731), .A2(n6910), .ZN(n6911) );
  NAND4_X1 U8651 ( .A1(n8689), .A2(n8705), .A3(n8722), .A4(n6911), .ZN(n6912)
         );
  OR2_X1 U8652 ( .A1(n8674), .A2(n6912), .ZN(n6913) );
  NOR2_X1 U8653 ( .A1(n6913), .A2(n8667), .ZN(n6914) );
  NAND4_X1 U8654 ( .A1(n8630), .A2(n6914), .A3(n8644), .A4(n8656), .ZN(n6915)
         );
  NOR2_X1 U8655 ( .A1(n6916), .A2(n6915), .ZN(n6919) );
  NAND4_X1 U8656 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n6921)
         );
  OAI21_X1 U8657 ( .B1(n6921), .B2(n7175), .A(n6946), .ZN(n6922) );
  INV_X1 U8658 ( .A(n6922), .ZN(n6923) );
  NAND2_X1 U8659 ( .A1(n7152), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7878) );
  INV_X1 U8660 ( .A(n7223), .ZN(n7298) );
  NAND3_X1 U8661 ( .A1(n7298), .A2(n6997), .A3(n7176), .ZN(n7162) );
  NOR3_X1 U8662 ( .A1(n7162), .A2(n6925), .A3(n5772), .ZN(n6927) );
  OAI21_X1 U8663 ( .B1(n7878), .B2(n6945), .A(P2_B_REG_SCAN_IN), .ZN(n6926) );
  OR2_X1 U8664 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  OAI21_X1 U8665 ( .B1(n6929), .B2(n7878), .A(n6928), .ZN(P2_U3296) );
  INV_X1 U8666 ( .A(n6930), .ZN(n9026) );
  INV_X1 U8667 ( .A(n6931), .ZN(n6934) );
  INV_X1 U8668 ( .A(n6932), .ZN(n6933) );
  AOI21_X1 U8669 ( .B1(n9026), .B2(n6934), .A(n6933), .ZN(n6936) );
  OAI21_X1 U8670 ( .B1(n6936), .B2(n6935), .A(n9025), .ZN(n6944) );
  INV_X1 U8671 ( .A(n9871), .ZN(n6941) );
  OAI22_X1 U8672 ( .A1(n9195), .A2(n9029), .B1(n9028), .B2(n9597), .ZN(n6939)
         );
  INV_X1 U8673 ( .A(n9594), .ZN(n6937) );
  NOR2_X1 U8674 ( .A1(n9041), .A2(n6937), .ZN(n6938) );
  AOI211_X1 U8675 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n6939), 
        .B(n6938), .ZN(n6940) );
  OAI21_X1 U8676 ( .B1(n6941), .B2(n9036), .A(n6940), .ZN(n6942) );
  NAND2_X1 U8677 ( .A1(n6944), .A2(n6943), .ZN(P1_U3214) );
  NAND3_X1 U8678 ( .A1(n6946), .A2(n6945), .A3(n7547), .ZN(n6947) );
  NAND2_X1 U8679 ( .A1(n6948), .A2(n6947), .ZN(n6951) );
  NAND2_X1 U8680 ( .A1(n6949), .A2(n6951), .ZN(n6950) );
  OAI21_X1 U8681 ( .B1(n7215), .B2(n6951), .A(n6950), .ZN(n7304) );
  AND2_X1 U8682 ( .A1(n6952), .A2(n7216), .ZN(n7154) );
  NOR2_X1 U8683 ( .A1(n6953), .A2(n7154), .ZN(n7302) );
  NAND2_X1 U8684 ( .A1(n10181), .A2(n4809), .ZN(n6954) );
  AND4_X2 U8685 ( .A1(n7304), .A2(n7302), .A3(n7157), .A4(n6954), .ZN(n10213)
         );
  NAND2_X1 U8686 ( .A1(n6955), .A2(n10213), .ZN(n6961) );
  NAND2_X1 U8687 ( .A1(n10213), .A2(n10195), .ZN(n8829) );
  INV_X1 U8688 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6957) );
  NOR2_X1 U8689 ( .A1(n10213), .A2(n6957), .ZN(n6958) );
  NAND2_X1 U8690 ( .A1(n6961), .A2(n6960), .ZN(P2_U3488) );
  NOR2_X1 U8691 ( .A1(n7018), .A2(P1_U3086), .ZN(n6962) );
  AND2_X1 U8692 ( .A1(n4637), .A2(P2_U3151), .ZN(n7295) );
  NAND2_X1 U8693 ( .A1(n5176), .A2(P2_U3151), .ZN(n8908) );
  OAI222_X1 U8694 ( .A1(n4517), .A2(n5020), .B1(n8908), .B2(n6968), .C1(
        P2_U3151), .C2(n6963), .ZN(P2_U3292) );
  OAI222_X1 U8695 ( .A1(n4517), .A2(n6964), .B1(n8908), .B2(n6970), .C1(
        P2_U3151), .C2(n7254), .ZN(P2_U3291) );
  NAND2_X1 U8696 ( .A1(n5176), .A2(P1_U3086), .ZN(n8343) );
  AND2_X1 U8697 ( .A1(n6965), .A2(P1_U3086), .ZN(n7874) );
  INV_X2 U8698 ( .A(n7874), .ZN(n9910) );
  OAI222_X1 U8699 ( .A1(n8343), .A2(n6966), .B1(n9910), .B2(n6982), .C1(
        P1_U3086), .C2(n7028), .ZN(P1_U3354) );
  OAI222_X1 U8700 ( .A1(n8343), .A2(n6967), .B1(n9910), .B2(n8221), .C1(
        P1_U3086), .C2(n7029), .ZN(P1_U3353) );
  INV_X1 U8701 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6969) );
  INV_X1 U8702 ( .A(n7030), .ZN(n9365) );
  OAI222_X1 U8703 ( .A1(n8343), .A2(n6969), .B1(n9910), .B2(n6968), .C1(
        P1_U3086), .C2(n9365), .ZN(P1_U3352) );
  INV_X1 U8704 ( .A(n9391), .ZN(n9385) );
  INV_X1 U8705 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7098) );
  OAI222_X1 U8706 ( .A1(P1_U3086), .A2(n9385), .B1(n9910), .B2(n6970), .C1(
        n8343), .C2(n7098), .ZN(P1_U3351) );
  INV_X1 U8707 ( .A(n6971), .ZN(n7293) );
  OAI222_X1 U8708 ( .A1(n4517), .A2(n6972), .B1(n8908), .B2(n6977), .C1(
        P2_U3151), .C2(n7293), .ZN(P2_U3290) );
  AND2_X1 U8709 ( .A1(n9995), .A2(n6973), .ZN(n9993) );
  NAND2_X1 U8710 ( .A1(n9993), .A2(n6974), .ZN(n6975) );
  OAI21_X1 U8711 ( .B1(n9993), .B2(n10611), .A(n6975), .ZN(P1_U3440) );
  INV_X1 U8712 ( .A(n8343), .ZN(n9908) );
  AOI22_X1 U8713 ( .A1(n9408), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9908), .ZN(n6976) );
  OAI21_X1 U8714 ( .B1(n6977), .B2(n9910), .A(n6976), .ZN(P1_U3350) );
  INV_X1 U8715 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6978) );
  OAI222_X1 U8716 ( .A1(n8343), .A2(n6978), .B1(n9910), .B2(n6980), .C1(
        P1_U3086), .C2(n7048), .ZN(P1_U3349) );
  OAI222_X1 U8717 ( .A1(n4517), .A2(n6981), .B1(n8908), .B2(n6980), .C1(
        P2_U3151), .C2(n6979), .ZN(P2_U3289) );
  INV_X1 U8718 ( .A(n8908), .ZN(n7876) );
  INV_X1 U8719 ( .A(n7876), .ZN(n8323) );
  INV_X1 U8720 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7006) );
  OAI222_X1 U8721 ( .A1(n6685), .A2(P2_U3151), .B1(n8323), .B2(n6982), .C1(
        n4517), .C2(n7006), .ZN(P2_U3294) );
  OAI222_X1 U8722 ( .A1(n4517), .A2(n6984), .B1(n8908), .B2(n6985), .C1(
        P2_U3151), .C2(n6983), .ZN(P2_U3288) );
  INV_X1 U8723 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10407) );
  INV_X1 U8724 ( .A(n7077), .ZN(n7058) );
  OAI222_X1 U8725 ( .A1(n8343), .A2(n10407), .B1(n9910), .B2(n6985), .C1(
        P1_U3086), .C2(n7058), .ZN(P1_U3348) );
  NAND2_X1 U8726 ( .A1(n9323), .A2(n7020), .ZN(n6986) );
  OR2_X1 U8727 ( .A1(n7020), .A2(P1_U3086), .ZN(n9336) );
  INV_X1 U8728 ( .A(n6987), .ZN(n6988) );
  NAND2_X1 U8729 ( .A1(n9336), .A2(n6988), .ZN(n6989) );
  AND2_X1 U8730 ( .A1(n7022), .A2(n6989), .ZN(n9946) );
  NOR2_X1 U8731 ( .A1(n9946), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8732 ( .A(n6990), .ZN(n7008) );
  AOI22_X1 U8733 ( .A1(n7202), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9908), .ZN(n6991) );
  OAI21_X1 U8734 ( .B1(n7008), .B2(n9910), .A(n6991), .ZN(P1_U3347) );
  NAND2_X1 U8735 ( .A1(n5803), .A2(n6997), .ZN(n7010) );
  INV_X1 U8736 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6994) );
  INV_X1 U8737 ( .A(n6992), .ZN(n6993) );
  AOI22_X1 U8738 ( .A1(n7010), .A2(n6994), .B1(n6997), .B2(n6993), .ZN(
        P2_U3376) );
  INV_X1 U8739 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6998) );
  INV_X1 U8740 ( .A(n6995), .ZN(n6996) );
  AOI22_X1 U8741 ( .A1(n7010), .A2(n6998), .B1(n6997), .B2(n6996), .ZN(
        P2_U3377) );
  NAND2_X1 U8742 ( .A1(n6074), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U8743 ( .A1(n4527), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U8744 ( .A1(n4514), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6999) );
  NAND3_X1 U8745 ( .A1(n7001), .A2(n7000), .A3(n6999), .ZN(n9057) );
  NAND2_X1 U8746 ( .A1(n9057), .A2(P1_U3973), .ZN(n7002) );
  OAI21_X1 U8747 ( .B1(P1_U3973), .B2(n6872), .A(n7002), .ZN(P1_U3585) );
  INV_X1 U8748 ( .A(n9099), .ZN(n7003) );
  NAND2_X1 U8749 ( .A1(n7003), .A2(P1_U3973), .ZN(n7004) );
  OAI21_X1 U8750 ( .B1(n6851), .B2(P1_U3973), .A(n7004), .ZN(P1_U3584) );
  NAND2_X1 U8751 ( .A1(n9750), .A2(P1_U3973), .ZN(n7005) );
  OAI21_X1 U8752 ( .B1(P1_U3973), .B2(n7006), .A(n7005), .ZN(P1_U3555) );
  OAI222_X1 U8753 ( .A1(n4517), .A2(n7009), .B1(n8323), .B2(n7008), .C1(
        P2_U3151), .C2(n7007), .ZN(P2_U3287) );
  AND2_X1 U8754 ( .A1(n7010), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8755 ( .A1(n7010), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8756 ( .A1(n7010), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8757 ( .A1(n7010), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8758 ( .A1(n7010), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8759 ( .A1(n7010), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8760 ( .A1(n7010), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8761 ( .A1(n7010), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8762 ( .A1(n7010), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8763 ( .A1(n7010), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8764 ( .A1(n7010), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8765 ( .A1(n7010), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8766 ( .A1(n7010), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8767 ( .A1(n7010), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8768 ( .A1(n7010), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8769 ( .A1(n7010), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8770 ( .A1(n7010), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8771 ( .A1(n7010), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8772 ( .A1(n7010), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8773 ( .A1(n7010), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8774 ( .A1(n7010), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8775 ( .A1(n7010), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8776 ( .A1(n7010), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8777 ( .A1(n7010), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8778 ( .A1(n7010), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8779 ( .A1(n7010), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8780 ( .A1(n7010), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8781 ( .A1(n7010), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8782 ( .A1(n7010), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8783 ( .A1(n7010), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8784 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7014) );
  INV_X1 U8785 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7013) );
  INV_X1 U8786 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7012) );
  MUX2_X1 U8787 ( .A(n7012), .B(P1_REG2_REG_2__SCAN_IN), .S(n7029), .Z(n9947)
         );
  INV_X1 U8788 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7641) );
  AND2_X1 U8789 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9380) );
  NAND2_X1 U8790 ( .A1(n9356), .A2(n9380), .ZN(n9948) );
  INV_X1 U8791 ( .A(n7028), .ZN(n9360) );
  NAND2_X1 U8792 ( .A1(n9360), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U8793 ( .A1(n9948), .A2(n9949), .ZN(n7011) );
  NAND2_X1 U8794 ( .A1(n9947), .A2(n7011), .ZN(n9951) );
  OAI21_X1 U8795 ( .B1(n7029), .B2(n7012), .A(n9951), .ZN(n9369) );
  XOR2_X1 U8796 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7030), .Z(n9370) );
  NAND2_X1 U8797 ( .A1(n9369), .A2(n9370), .ZN(n9368) );
  OAI21_X1 U8798 ( .B1(n7013), .B2(n9365), .A(n9368), .ZN(n9389) );
  XOR2_X1 U8799 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9391), .Z(n9390) );
  NAND2_X1 U8800 ( .A1(n9389), .A2(n9390), .ZN(n9388) );
  OAI21_X1 U8801 ( .B1(n9385), .B2(n7014), .A(n9388), .ZN(n9400) );
  INV_X1 U8802 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7015) );
  MUX2_X1 U8803 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7015), .S(n9408), .Z(n9401)
         );
  INV_X1 U8804 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7016) );
  MUX2_X1 U8805 ( .A(n7016), .B(P1_REG2_REG_6__SCAN_IN), .S(n7048), .Z(n7017)
         );
  INV_X1 U8806 ( .A(n7017), .ZN(n7024) );
  INV_X1 U8807 ( .A(n7018), .ZN(n7019) );
  AND2_X1 U8808 ( .A1(n7020), .A2(n7019), .ZN(n7021) );
  OR3_X1 U8809 ( .A1(n7022), .A2(n7021), .A3(P1_U3086), .ZN(n9944) );
  INV_X1 U8810 ( .A(n9944), .ZN(n7026) );
  NOR2_X1 U8811 ( .A1(n9378), .A2(n9300), .ZN(n7023) );
  NAND2_X1 U8812 ( .A1(n7026), .A2(n7023), .ZN(n9962) );
  AOI211_X1 U8813 ( .C1(n7025), .C2(n7024), .A(n9962), .B(n7042), .ZN(n7041)
         );
  NOR2_X1 U8814 ( .A1(n9944), .A2(n9382), .ZN(n9958) );
  INV_X1 U8815 ( .A(n9958), .ZN(n9457) );
  NAND2_X1 U8816 ( .A1(n7026), .A2(n9300), .ZN(n9957) );
  INV_X1 U8817 ( .A(n9957), .ZN(n9551) );
  INV_X1 U8818 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7027) );
  MUX2_X1 U8819 ( .A(n7027), .B(P1_REG1_REG_2__SCAN_IN), .S(n7029), .Z(n9955)
         );
  INV_X1 U8820 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10079) );
  MUX2_X1 U8821 ( .A(n10079), .B(P1_REG1_REG_1__SCAN_IN), .S(n7028), .Z(n9358)
         );
  AND2_X1 U8822 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9359) );
  NAND2_X1 U8823 ( .A1(n9358), .A2(n9359), .ZN(n9357) );
  OAI21_X1 U8824 ( .B1(n10079), .B2(n7028), .A(n9357), .ZN(n9954) );
  NAND2_X1 U8825 ( .A1(n9955), .A2(n9954), .ZN(n9953) );
  NAND2_X1 U8826 ( .A1(n4647), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9372) );
  INV_X1 U8827 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10082) );
  MUX2_X1 U8828 ( .A(n10082), .B(P1_REG1_REG_3__SCAN_IN), .S(n7030), .Z(n9371)
         );
  AOI21_X1 U8829 ( .B1(n9953), .B2(n9372), .A(n9371), .ZN(n9396) );
  NOR2_X1 U8830 ( .A1(n9365), .A2(n10082), .ZN(n9392) );
  INV_X1 U8831 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7031) );
  MUX2_X1 U8832 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7031), .S(n9391), .Z(n7032)
         );
  OAI21_X1 U8833 ( .B1(n9396), .B2(n9392), .A(n7032), .ZN(n9404) );
  NAND2_X1 U8834 ( .A1(n9391), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9403) );
  INV_X1 U8835 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10085) );
  MUX2_X1 U8836 ( .A(n10085), .B(P1_REG1_REG_5__SCAN_IN), .S(n9408), .Z(n9402)
         );
  AOI21_X1 U8837 ( .B1(n9404), .B2(n9403), .A(n9402), .ZN(n7033) );
  INV_X1 U8838 ( .A(n7033), .ZN(n9406) );
  NAND2_X1 U8839 ( .A1(n9408), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7035) );
  INV_X1 U8840 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10087) );
  MUX2_X1 U8841 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10087), .S(n7048), .Z(n7034)
         );
  AOI21_X1 U8842 ( .B1(n9406), .B2(n7035), .A(n7034), .ZN(n7054) );
  INV_X1 U8843 ( .A(n7054), .ZN(n7037) );
  NAND3_X1 U8844 ( .A1(n9406), .A2(n7035), .A3(n7034), .ZN(n7036) );
  NAND3_X1 U8845 ( .A1(n9551), .A2(n7037), .A3(n7036), .ZN(n7039) );
  AND2_X1 U8846 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7458) );
  AOI21_X1 U8847 ( .B1(n9946), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7458), .ZN(
        n7038) );
  OAI211_X1 U8848 ( .C1(n9457), .C2(n7048), .A(n7039), .B(n7038), .ZN(n7040)
         );
  OR2_X1 U8849 ( .A1(n7041), .A2(n7040), .ZN(P1_U3249) );
  INV_X1 U8850 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7044) );
  MUX2_X1 U8851 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7044), .S(n7077), .Z(n7045)
         );
  INV_X1 U8852 ( .A(n7045), .ZN(n7046) );
  NOR2_X1 U8853 ( .A1(n7047), .A2(n7046), .ZN(n7072) );
  AOI211_X1 U8854 ( .C1(n7047), .C2(n7046), .A(n9962), .B(n7072), .ZN(n7060)
         );
  INV_X1 U8855 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10089) );
  MUX2_X1 U8856 ( .A(n10089), .B(P1_REG1_REG_7__SCAN_IN), .S(n7077), .Z(n7050)
         );
  NOR2_X1 U8857 ( .A1(n7048), .A2(n10087), .ZN(n7052) );
  INV_X1 U8858 ( .A(n7052), .ZN(n7049) );
  NAND2_X1 U8859 ( .A1(n7050), .A2(n7049), .ZN(n7053) );
  MUX2_X1 U8860 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10089), .S(n7077), .Z(n7051)
         );
  OAI21_X1 U8861 ( .B1(n7054), .B2(n7052), .A(n7051), .ZN(n7081) );
  OAI211_X1 U8862 ( .C1(n7054), .C2(n7053), .A(n7081), .B(n9551), .ZN(n7057)
         );
  NOR2_X1 U8863 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7055), .ZN(n7358) );
  AOI21_X1 U8864 ( .B1(n9946), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7358), .ZN(
        n7056) );
  OAI211_X1 U8865 ( .C1(n9457), .C2(n7058), .A(n7057), .B(n7056), .ZN(n7059)
         );
  OR2_X1 U8866 ( .A1(n7060), .A2(n7059), .ZN(P1_U3250) );
  INV_X1 U8867 ( .A(n7061), .ZN(n7064) );
  AOI22_X1 U8868 ( .A1(n7905), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n7295), .ZN(n7062) );
  OAI21_X1 U8869 ( .B1(n7064), .B2(n8908), .A(n7062), .ZN(P2_U3286) );
  AOI22_X1 U8870 ( .A1(n9422), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9908), .ZN(n7063) );
  OAI21_X1 U8871 ( .B1(n7064), .B2(n9910), .A(n7063), .ZN(P1_U3346) );
  INV_X1 U8872 ( .A(n7065), .ZN(n7068) );
  INV_X1 U8873 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7066) );
  OAI222_X1 U8874 ( .A1(n8323), .A2(n7068), .B1(n7067), .B2(P2_U3151), .C1(
        n7066), .C2(n4517), .ZN(P2_U3285) );
  CLKBUF_X1 U8875 ( .A(n8343), .Z(n8225) );
  INV_X1 U8876 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7069) );
  INV_X1 U8877 ( .A(n7322), .ZN(n7200) );
  OAI222_X1 U8878 ( .A1(n8225), .A2(n7069), .B1(n9910), .B2(n7068), .C1(n7200), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8879 ( .A(n7070), .ZN(n7088) );
  AOI22_X1 U8880 ( .A1(n8020), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n7295), .ZN(n7071) );
  OAI21_X1 U8881 ( .B1(n7088), .B2(n8908), .A(n7071), .ZN(P2_U3284) );
  INV_X1 U8882 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7073) );
  MUX2_X1 U8883 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7073), .S(n7202), .Z(n7074)
         );
  INV_X1 U8884 ( .A(n7074), .ZN(n7075) );
  AOI211_X1 U8885 ( .C1(n7076), .C2(n7075), .A(n9962), .B(n7201), .ZN(n7087)
         );
  NAND2_X1 U8886 ( .A1(n7077), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7080) );
  INV_X1 U8887 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7078) );
  MUX2_X1 U8888 ( .A(n7078), .B(P1_REG1_REG_8__SCAN_IN), .S(n7202), .Z(n7079)
         );
  AOI21_X1 U8889 ( .B1(n7081), .B2(n7080), .A(n7079), .ZN(n7197) );
  AND3_X1 U8890 ( .A1(n7081), .A2(n7080), .A3(n7079), .ZN(n7082) );
  NOR3_X1 U8891 ( .A1(n7197), .A2(n7082), .A3(n9957), .ZN(n7086) );
  INV_X1 U8892 ( .A(n7202), .ZN(n7084) );
  AND2_X1 U8893 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7596) );
  AOI21_X1 U8894 ( .B1(n9946), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7596), .ZN(
        n7083) );
  OAI21_X1 U8895 ( .B1(n9457), .B2(n7084), .A(n7083), .ZN(n7085) );
  OR3_X1 U8896 ( .A1(n7087), .A2(n7086), .A3(n7085), .ZN(P1_U3251) );
  INV_X1 U8897 ( .A(n9436), .ZN(n7316) );
  OAI222_X1 U8898 ( .A1(n8225), .A2(n10457), .B1(n9910), .B2(n7088), .C1(
        P1_U3086), .C2(n7316), .ZN(P1_U3344) );
  INV_X1 U8899 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7093) );
  AND2_X1 U8900 ( .A1(n9998), .A2(n7091), .ZN(n9247) );
  NOR2_X1 U8901 ( .A1(n7638), .A2(n9247), .ZN(n9755) );
  NOR2_X1 U8902 ( .A1(n10060), .A2(n9821), .ZN(n7089) );
  OAI222_X1 U8903 ( .A1(n7091), .A2(n7090), .B1(n9755), .B2(n7089), .C1(n9968), 
        .C2(n7125), .ZN(n9856) );
  NAND2_X1 U8904 ( .A1(n9856), .A2(n10078), .ZN(n7092) );
  OAI21_X1 U8905 ( .B1(n10078), .B2(n7093), .A(n7092), .ZN(P1_U3453) );
  INV_X1 U8906 ( .A(n7094), .ZN(n7099) );
  INV_X1 U8907 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7095) );
  OAI222_X1 U8908 ( .A1(n8323), .A2(n7099), .B1(n7096), .B2(P2_U3151), .C1(
        n7095), .C2(n4517), .ZN(P2_U3283) );
  NAND2_X1 U8909 ( .A1(n7666), .A2(P2_U3893), .ZN(n7097) );
  OAI21_X1 U8910 ( .B1(P2_U3893), .B2(n7098), .A(n7097), .ZN(P2_U3495) );
  INV_X1 U8911 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7100) );
  INV_X1 U8912 ( .A(n9448), .ZN(n9442) );
  OAI222_X1 U8913 ( .A1(n8225), .A2(n7100), .B1(n9910), .B2(n7099), .C1(n9442), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8914 ( .A(n7101), .ZN(n7121) );
  AOI22_X1 U8915 ( .A1(n8532), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n7295), .ZN(n7102) );
  OAI21_X1 U8916 ( .B1(n7121), .B2(n8908), .A(n7102), .ZN(P2_U3282) );
  XNOR2_X1 U8917 ( .A(n7104), .B(n7103), .ZN(n9381) );
  NOR2_X1 U8918 ( .A1(n8972), .A2(P1_U3086), .ZN(n7127) );
  INV_X1 U8919 ( .A(n7127), .ZN(n7109) );
  AOI22_X1 U8920 ( .A1(n7109), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9037), .B2(
        n9750), .ZN(n7106) );
  NAND2_X1 U8921 ( .A1(n9051), .A2(n9748), .ZN(n7105) );
  OAI211_X1 U8922 ( .C1(n9381), .C2(n9046), .A(n7106), .B(n7105), .ZN(P1_U3232) );
  AOI21_X1 U8923 ( .B1(n7108), .B2(n7107), .A(n4629), .ZN(n7112) );
  INV_X1 U8924 ( .A(n9029), .ZN(n9038) );
  AOI22_X1 U8925 ( .A1(n7109), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9038), .B2(
        n9998), .ZN(n7111) );
  AOI22_X1 U8926 ( .A1(n9051), .A2(n5919), .B1(n9037), .B2(n9997), .ZN(n7110)
         );
  OAI211_X1 U8927 ( .C1(n7112), .C2(n9046), .A(n7111), .B(n7110), .ZN(P1_U3222) );
  NAND2_X1 U8928 ( .A1(n9816), .A2(P1_U3973), .ZN(n7113) );
  OAI21_X1 U8929 ( .B1(n5275), .B2(P1_U3973), .A(n7113), .ZN(P1_U3577) );
  INV_X1 U8930 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7120) );
  NAND2_X1 U8931 ( .A1(n7114), .A2(n7378), .ZN(n7117) );
  AOI22_X1 U8932 ( .A1(n7117), .A2(n7116), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n7118) );
  OAI211_X1 U8933 ( .C1(n8611), .C2(n7120), .A(n7119), .B(n7118), .ZN(P2_U3182) );
  INV_X1 U8934 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10605) );
  INV_X1 U8935 ( .A(n9462), .ZN(n9468) );
  OAI222_X1 U8936 ( .A1(n8225), .A2(n10605), .B1(n9910), .B2(n7121), .C1(
        P1_U3086), .C2(n9468), .ZN(P1_U3342) );
  OAI21_X1 U8937 ( .B1(n7124), .B2(n7123), .A(n7122), .ZN(n7130) );
  INV_X1 U8938 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7126) );
  OAI22_X1 U8939 ( .A1(n7127), .A2(n7126), .B1(n7125), .B2(n9029), .ZN(n7129)
         );
  OAI22_X1 U8940 ( .A1(n9036), .A2(n10012), .B1(n7579), .B2(n9028), .ZN(n7128)
         );
  AOI211_X1 U8941 ( .C1(n7130), .C2(n9025), .A(n7129), .B(n7128), .ZN(n7131)
         );
  INV_X1 U8942 ( .A(n7131), .ZN(P1_U3237) );
  AOI21_X1 U8943 ( .B1(n7134), .B2(n7133), .A(n7132), .ZN(n7146) );
  AOI21_X1 U8944 ( .B1(n7136), .B2(n5355), .A(n7135), .ZN(n7138) );
  INV_X1 U8945 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10633) );
  NOR2_X1 U8946 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10633), .ZN(n7430) );
  INV_X1 U8947 ( .A(n7430), .ZN(n7137) );
  OAI21_X1 U8948 ( .B1(n10100), .B2(n7138), .A(n7137), .ZN(n7143) );
  AOI21_X1 U8949 ( .B1(n7140), .B2(n5354), .A(n7139), .ZN(n7141) );
  NOR2_X1 U8950 ( .A1(n8618), .A2(n7141), .ZN(n7142) );
  AOI211_X1 U8951 ( .C1(n10105), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n7143), .B(
        n7142), .ZN(n7145) );
  NAND2_X1 U8952 ( .A1(n8596), .A2(n4833), .ZN(n7144) );
  OAI211_X1 U8953 ( .C1(n7146), .C2(n7378), .A(n7145), .B(n7144), .ZN(P2_U3185) );
  INV_X1 U8954 ( .A(n7147), .ZN(n7149) );
  INV_X1 U8955 ( .A(n9480), .ZN(n9475) );
  OAI222_X1 U8956 ( .A1(n8225), .A2(n10615), .B1(n9910), .B2(n7149), .C1(
        P1_U3086), .C2(n9475), .ZN(P1_U3341) );
  INV_X1 U8957 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7150) );
  OAI222_X1 U8958 ( .A1(n4517), .A2(n7150), .B1(n8323), .B2(n7149), .C1(
        P2_U3151), .C2(n7148), .ZN(P2_U3281) );
  INV_X1 U8959 ( .A(n7151), .ZN(n7156) );
  NOR2_X1 U8960 ( .A1(n7303), .A2(n7156), .ZN(n7161) );
  INV_X1 U8961 ( .A(n7176), .ZN(n7153) );
  NOR3_X1 U8962 ( .A1(n7154), .A2(n7153), .A3(n7152), .ZN(n7159) );
  OAI21_X1 U8963 ( .B1(n7157), .B2(n7156), .A(n7155), .ZN(n7158) );
  OAI211_X1 U8964 ( .C1(n7161), .C2(n7167), .A(n7159), .B(n7158), .ZN(n7160)
         );
  NAND2_X1 U8965 ( .A1(n7160), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7166) );
  INV_X1 U8966 ( .A(n7161), .ZN(n7164) );
  INV_X1 U8967 ( .A(n7162), .ZN(n7163) );
  NAND2_X1 U8968 ( .A1(n7164), .A2(n7163), .ZN(n7165) );
  NOR2_X1 U8969 ( .A1(n8479), .A2(P2_U3151), .ZN(n7277) );
  INV_X1 U8970 ( .A(n7299), .ZN(n7189) );
  INV_X1 U8971 ( .A(n7167), .ZN(n7168) );
  NAND2_X1 U8972 ( .A1(n7226), .A2(n7168), .ZN(n7172) );
  INV_X1 U8973 ( .A(n7169), .ZN(n7170) );
  NAND2_X1 U8974 ( .A1(n7173), .A2(n7170), .ZN(n7171) );
  NAND2_X1 U8975 ( .A1(n7173), .A2(n10195), .ZN(n7178) );
  NOR2_X1 U8976 ( .A1(n7175), .A2(n7174), .ZN(n7177) );
  NAND2_X1 U8977 ( .A1(n7178), .A2(n8776), .ZN(n8378) );
  AND2_X1 U8978 ( .A1(n7224), .A2(n7298), .ZN(n7179) );
  NAND2_X1 U8979 ( .A1(n7226), .A2(n7179), .ZN(n8488) );
  OAI22_X1 U8980 ( .A1(n8496), .A2(n7191), .B1(n7271), .B2(n8488), .ZN(n7180)
         );
  AOI21_X1 U8981 ( .B1(n7189), .B2(n8472), .A(n7180), .ZN(n7181) );
  OAI21_X1 U8982 ( .B1(n7277), .B2(n10630), .A(n7181), .ZN(P2_U3172) );
  OAI21_X1 U8983 ( .B1(n7184), .B2(n7183), .A(n7182), .ZN(n7185) );
  NAND2_X1 U8984 ( .A1(n7185), .A2(n9025), .ZN(n7188) );
  NOR2_X1 U8985 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7629), .ZN(n9367) );
  OAI22_X1 U8986 ( .A1(n7384), .A2(n9028), .B1(n9029), .B2(n7646), .ZN(n7186)
         );
  AOI211_X1 U8987 ( .C1(n9033), .C2(n7629), .A(n9367), .B(n7186), .ZN(n7187)
         );
  OAI211_X1 U8988 ( .C1(n10019), .C2(n9036), .A(n7188), .B(n7187), .ZN(
        P1_U3218) );
  INV_X1 U8989 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U8990 ( .A1(n7817), .A2(n10162), .ZN(n10188) );
  OAI21_X1 U8991 ( .B1(n10123), .B2(n10188), .A(n7189), .ZN(n7190) );
  OR2_X1 U8992 ( .A1(n7271), .A2(n8760), .ZN(n7297) );
  OAI211_X1 U8993 ( .C1(n10183), .C2(n7191), .A(n7190), .B(n7297), .ZN(n7194)
         );
  NAND2_X1 U8994 ( .A1(n7194), .A2(n10196), .ZN(n7192) );
  OAI21_X1 U8995 ( .B1(n7193), .B2(n10196), .A(n7192), .ZN(P2_U3390) );
  NAND2_X1 U8996 ( .A1(n7194), .A2(n10213), .ZN(n7195) );
  OAI21_X1 U8997 ( .B1(n10213), .B2(n6582), .A(n7195), .ZN(P2_U3459) );
  INV_X1 U8998 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7196) );
  MUX2_X1 U8999 ( .A(n7196), .B(P1_REG1_REG_10__SCAN_IN), .S(n7322), .Z(n7312)
         );
  AOI21_X1 U9000 ( .B1(n7202), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7197), .ZN(
        n9419) );
  INV_X1 U9001 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7198) );
  MUX2_X1 U9002 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7198), .S(n9422), .Z(n9420)
         );
  NAND2_X1 U9003 ( .A1(n9419), .A2(n9420), .ZN(n9418) );
  OAI21_X1 U9004 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9422), .A(n9418), .ZN(
        n7313) );
  XOR2_X1 U9005 ( .A(n7312), .B(n7313), .Z(n7208) );
  AND2_X1 U9006 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7868) );
  AOI21_X1 U9007 ( .B1(n9946), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7868), .ZN(
        n7199) );
  OAI21_X1 U9008 ( .B1(n9457), .B2(n7200), .A(n7199), .ZN(n7207) );
  XOR2_X1 U9009 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9422), .Z(n9415) );
  OAI21_X1 U9010 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9422), .A(n9413), .ZN(
        n7205) );
  NAND2_X1 U9011 ( .A1(n7322), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7203) );
  OAI21_X1 U9012 ( .B1(n7322), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7203), .ZN(
        n7204) );
  NOR2_X1 U9013 ( .A1(n7205), .A2(n7204), .ZN(n7321) );
  AOI211_X1 U9014 ( .C1(n7205), .C2(n7204), .A(n9962), .B(n7321), .ZN(n7206)
         );
  AOI211_X1 U9015 ( .C1(n9551), .C2(n7208), .A(n7207), .B(n7206), .ZN(n7209)
         );
  INV_X1 U9016 ( .A(n7209), .ZN(P1_U3253) );
  INV_X1 U9017 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7211) );
  INV_X1 U9018 ( .A(n7210), .ZN(n7212) );
  OAI222_X1 U9019 ( .A1(n4517), .A2(n7211), .B1(n8323), .B2(n7212), .C1(
        P2_U3151), .C2(n8562), .ZN(P2_U3280) );
  INV_X1 U9020 ( .A(n9488), .ZN(n9494) );
  OAI222_X1 U9021 ( .A1(n8225), .A2(n10394), .B1(n9910), .B2(n7212), .C1(
        P1_U3086), .C2(n9494), .ZN(P1_U3340) );
  INV_X1 U9022 ( .A(n7213), .ZN(n7214) );
  INV_X1 U9023 ( .A(n7216), .ZN(n7217) );
  NOR2_X1 U9024 ( .A1(n7347), .A2(n7217), .ZN(n7218) );
  XNOR2_X1 U9025 ( .A(n7345), .B(n8281), .ZN(n7219) );
  OAI21_X1 U9026 ( .B1(n7308), .B2(n7421), .A(n7341), .ZN(n7220) );
  OAI21_X1 U9027 ( .B1(n7221), .B2(n7220), .A(n7267), .ZN(n7222) );
  NAND2_X1 U9028 ( .A1(n7222), .A2(n8472), .ZN(n7230) );
  NOR2_X1 U9029 ( .A1(n7224), .A2(n7223), .ZN(n7225) );
  NAND2_X1 U9030 ( .A1(n7226), .A2(n7225), .ZN(n8477) );
  OAI22_X1 U9031 ( .A1(n7227), .A2(n8477), .B1(n8488), .B2(n5351), .ZN(n7228)
         );
  AOI21_X1 U9032 ( .B1(n7345), .B2(n8378), .A(n7228), .ZN(n7229) );
  OAI211_X1 U9033 ( .C1(n7277), .C2(n8209), .A(n7230), .B(n7229), .ZN(P2_U3162) );
  OAI211_X1 U9034 ( .C1(n7233), .C2(n7232), .A(n7231), .B(n10095), .ZN(n7253)
         );
  INV_X1 U9035 ( .A(n7234), .ZN(n7239) );
  NAND3_X1 U9036 ( .A1(n7237), .A2(n7236), .A3(n7235), .ZN(n7238) );
  AOI21_X1 U9037 ( .B1(n7239), .B2(n7238), .A(n8618), .ZN(n7251) );
  INV_X1 U9038 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7240) );
  NOR2_X1 U9039 ( .A1(n8611), .A2(n7240), .ZN(n7250) );
  AND3_X1 U9040 ( .A1(n7243), .A2(n7242), .A3(n7241), .ZN(n7244) );
  NOR2_X1 U9041 ( .A1(n7245), .A2(n7244), .ZN(n7248) );
  INV_X1 U9042 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7246) );
  NOR2_X1 U9043 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7246), .ZN(n7502) );
  INV_X1 U9044 ( .A(n7502), .ZN(n7247) );
  OAI21_X1 U9045 ( .B1(n10100), .B2(n7248), .A(n7247), .ZN(n7249) );
  NOR3_X1 U9046 ( .A1(n7251), .A2(n7250), .A3(n7249), .ZN(n7252) );
  OAI211_X1 U9047 ( .C1(n6680), .C2(n7254), .A(n7253), .B(n7252), .ZN(P2_U3186) );
  AOI21_X1 U9048 ( .B1(n7255), .B2(n7256), .A(n9046), .ZN(n7258) );
  NAND2_X1 U9049 ( .A1(n7258), .A2(n7257), .ZN(n7262) );
  NOR2_X1 U9050 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7259), .ZN(n9387) );
  OAI22_X1 U9051 ( .A1(n7579), .A2(n9029), .B1(n9028), .B2(n7580), .ZN(n7260)
         );
  AOI211_X1 U9052 ( .C1(n9033), .C2(n7584), .A(n9387), .B(n7260), .ZN(n7261)
         );
  OAI211_X1 U9053 ( .C1(n10024), .C2(n9036), .A(n7262), .B(n7261), .ZN(
        P1_U3230) );
  INV_X1 U9054 ( .A(n7263), .ZN(n7278) );
  OAI222_X1 U9055 ( .A1(n8323), .A2(n7278), .B1(n7265), .B2(P2_U3151), .C1(
        n7264), .C2(n4517), .ZN(P2_U3279) );
  XNOR2_X1 U9056 ( .A(n7421), .B(n7273), .ZN(n7423) );
  XNOR2_X1 U9057 ( .A(n7423), .B(n8514), .ZN(n7269) );
  NAND2_X1 U9058 ( .A1(n7269), .A2(n7268), .ZN(n7424) );
  OAI21_X1 U9059 ( .B1(n7269), .B2(n7268), .A(n7424), .ZN(n7270) );
  NAND2_X1 U9060 ( .A1(n7270), .A2(n8472), .ZN(n7275) );
  OAI22_X1 U9061 ( .A1(n7271), .A2(n8477), .B1(n8488), .B2(n7500), .ZN(n7272)
         );
  AOI21_X1 U9062 ( .B1(n7273), .B2(n8378), .A(n7272), .ZN(n7274) );
  OAI211_X1 U9063 ( .C1(n7277), .C2(n7276), .A(n7275), .B(n7274), .ZN(P2_U3177) );
  INV_X1 U9064 ( .A(n9515), .ZN(n9509) );
  OAI222_X1 U9065 ( .A1(n8225), .A2(n10374), .B1(n9910), .B2(n7278), .C1(n9509), .C2(P1_U3086), .ZN(P1_U3339) );
  NAND2_X1 U9066 ( .A1(n8677), .A2(P2_U3893), .ZN(n7279) );
  OAI21_X1 U9067 ( .B1(P2_U3893), .B2(n6344), .A(n7279), .ZN(P2_U3514) );
  OAI211_X1 U9068 ( .C1(n7282), .C2(n7281), .A(n7280), .B(n10095), .ZN(n7292)
         );
  AOI21_X1 U9069 ( .B1(n7283), .B2(n7670), .A(n4630), .ZN(n7285) );
  NOR2_X1 U9070 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5385), .ZN(n7557) );
  INV_X1 U9071 ( .A(n7557), .ZN(n7284) );
  OAI21_X1 U9072 ( .B1(n7285), .B2(n10100), .A(n7284), .ZN(n7290) );
  AOI21_X1 U9073 ( .B1(n7287), .B2(n5383), .A(n7286), .ZN(n7288) );
  NOR2_X1 U9074 ( .A1(n8618), .A2(n7288), .ZN(n7289) );
  AOI211_X1 U9075 ( .C1(n10105), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7290), .B(
        n7289), .ZN(n7291) );
  OAI211_X1 U9076 ( .C1(n6680), .C2(n7293), .A(n7292), .B(n7291), .ZN(P2_U3187) );
  INV_X1 U9077 ( .A(n7294), .ZN(n7352) );
  AOI22_X1 U9078 ( .A1(n8597), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n7295), .ZN(n7296) );
  OAI21_X1 U9079 ( .B1(n7352), .B2(n8908), .A(n7296), .ZN(P2_U3278) );
  INV_X1 U9080 ( .A(n7297), .ZN(n7301) );
  NOR3_X1 U9081 ( .A1(n7299), .A2(n7298), .A3(n10195), .ZN(n7300) );
  AOI211_X1 U9082 ( .C1(n10133), .C2(P2_REG3_REG_0__SCAN_IN), .A(n7301), .B(
        n7300), .ZN(n7310) );
  AND2_X1 U9083 ( .A1(n7303), .A2(n7302), .ZN(n7306) );
  INV_X1 U9084 ( .A(n7304), .ZN(n7305) );
  NAND2_X1 U9085 ( .A1(n7306), .A2(n7305), .ZN(n7307) );
  NAND2_X2 U9086 ( .A1(n7307), .A2(n8776), .ZN(n8779) );
  INV_X2 U9087 ( .A(n8779), .ZN(n10136) );
  NOR2_X2 U9088 ( .A1(n7307), .A2(n8679), .ZN(n10130) );
  AOI22_X1 U9089 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n10136), .B1(n10130), .B2(
        n7308), .ZN(n7309) );
  OAI21_X1 U9090 ( .B1(n7310), .B2(n10136), .A(n7309), .ZN(P2_U3233) );
  INV_X1 U9091 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7311) );
  MUX2_X1 U9092 ( .A(n7311), .B(P1_REG1_REG_12__SCAN_IN), .S(n9448), .Z(n7319)
         );
  INV_X1 U9093 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7317) );
  NAND2_X1 U9094 ( .A1(n7322), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7315) );
  OR2_X1 U9095 ( .A1(n7313), .A2(n7312), .ZN(n7314) );
  NAND2_X1 U9096 ( .A1(n7315), .A2(n7314), .ZN(n9429) );
  MUX2_X1 U9097 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7317), .S(n9436), .Z(n9428)
         );
  NAND2_X1 U9098 ( .A1(n9429), .A2(n9428), .ZN(n9427) );
  OAI21_X1 U9099 ( .B1(n7317), .B2(n7316), .A(n9427), .ZN(n7318) );
  NOR2_X1 U9100 ( .A1(n7318), .A2(n7319), .ZN(n9441) );
  AOI21_X1 U9101 ( .B1(n7319), .B2(n7318), .A(n9441), .ZN(n7330) );
  INV_X1 U9102 ( .A(n9962), .ZN(n9528) );
  INV_X1 U9103 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7320) );
  XNOR2_X1 U9104 ( .A(n9436), .B(n7320), .ZN(n9434) );
  NOR2_X1 U9105 ( .A1(n9448), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7323) );
  AOI21_X1 U9106 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9448), .A(n7323), .ZN(
        n7324) );
  NAND2_X1 U9107 ( .A1(n7324), .A2(n7325), .ZN(n9447) );
  OAI21_X1 U9108 ( .B1(n7325), .B2(n7324), .A(n9447), .ZN(n7328) );
  AND2_X1 U9109 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7944) );
  AOI21_X1 U9110 ( .B1(n9946), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7944), .ZN(
        n7326) );
  OAI21_X1 U9111 ( .B1(n9457), .B2(n9442), .A(n7326), .ZN(n7327) );
  AOI21_X1 U9112 ( .B1(n9528), .B2(n7328), .A(n7327), .ZN(n7329) );
  OAI21_X1 U9113 ( .B1(n7330), .B2(n9957), .A(n7329), .ZN(P1_U3255) );
  OAI21_X1 U9114 ( .B1(n7331), .B2(n7332), .A(n7480), .ZN(n7624) );
  INV_X1 U9115 ( .A(n10123), .ZN(n8757) );
  XNOR2_X1 U9116 ( .A(n7333), .B(n7332), .ZN(n7334) );
  OAI222_X1 U9117 ( .A1(n8760), .A2(n7554), .B1(n8762), .B2(n5351), .C1(n8757), 
        .C2(n7334), .ZN(n7621) );
  AOI21_X1 U9118 ( .B1(n10188), .B2(n7624), .A(n7621), .ZN(n7339) );
  INV_X1 U9119 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7335) );
  OAI22_X1 U9120 ( .A1(n7620), .A2(n8900), .B1(n10196), .B2(n7335), .ZN(n7336)
         );
  INV_X1 U9121 ( .A(n7336), .ZN(n7337) );
  OAI21_X1 U9122 ( .B1(n7339), .B2(n10198), .A(n7337), .ZN(P2_U3399) );
  AOI22_X1 U9123 ( .A1(n6959), .A2(n7422), .B1(n10211), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7338) );
  OAI21_X1 U9124 ( .B1(n7339), .B2(n10211), .A(n7338), .ZN(P2_U3462) );
  XOR2_X1 U9125 ( .A(n7340), .B(n6897), .Z(n7344) );
  AOI22_X1 U9126 ( .A1(n8514), .A2(n10120), .B1(n10118), .B2(n8516), .ZN(n7343) );
  XNOR2_X1 U9127 ( .A(n6897), .B(n7341), .ZN(n10140) );
  INV_X1 U9128 ( .A(n7817), .ZN(n7953) );
  NAND2_X1 U9129 ( .A1(n10140), .A2(n7953), .ZN(n7342) );
  OAI211_X1 U9130 ( .C1(n7344), .C2(n8757), .A(n7343), .B(n7342), .ZN(n10138)
         );
  AOI22_X1 U9131 ( .A1(n10130), .A2(n7345), .B1(n10133), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7349) );
  AND2_X1 U9132 ( .A1(n7347), .A2(n7346), .ZN(n7482) );
  NAND2_X1 U9133 ( .A1(n8779), .A2(n7482), .ZN(n8346) );
  INV_X1 U9134 ( .A(n8346), .ZN(n7927) );
  NAND2_X1 U9135 ( .A1(n10140), .A2(n7927), .ZN(n7348) );
  OAI211_X1 U9136 ( .C1(n6634), .C2(n8779), .A(n7349), .B(n7348), .ZN(n7350)
         );
  AOI21_X1 U9137 ( .B1(n10138), .B2(n8779), .A(n7350), .ZN(n7351) );
  INV_X1 U9138 ( .A(n7351), .ZN(P2_U3232) );
  INV_X1 U9139 ( .A(n9532), .ZN(n9510) );
  OAI222_X1 U9140 ( .A1(n10366), .A2(n8343), .B1(P1_U3086), .B2(n9510), .C1(
        n9910), .C2(n7352), .ZN(P1_U3338) );
  OAI21_X1 U9141 ( .B1(n7355), .B2(n7354), .A(n7353), .ZN(n7356) );
  NAND2_X1 U9142 ( .A1(n7356), .A2(n9025), .ZN(n7360) );
  OAI22_X1 U9143 ( .A1(n9971), .A2(n9029), .B1(n9028), .B2(n9969), .ZN(n7357)
         );
  AOI211_X1 U9144 ( .C1(n9033), .C2(n9978), .A(n7358), .B(n7357), .ZN(n7359)
         );
  OAI211_X1 U9145 ( .C1(n10049), .C2(n9036), .A(n7360), .B(n7359), .ZN(
        P1_U3213) );
  AOI21_X1 U9146 ( .B1(n7363), .B2(n7362), .A(n7361), .ZN(n7379) );
  AOI21_X1 U9147 ( .B1(n7366), .B2(n7365), .A(n7364), .ZN(n7374) );
  AOI21_X1 U9148 ( .B1(n7369), .B2(n7368), .A(n7367), .ZN(n7371) );
  INV_X1 U9149 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7370) );
  OR2_X1 U9150 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7370), .ZN(n7694) );
  OAI21_X1 U9151 ( .B1(n10100), .B2(n7371), .A(n7694), .ZN(n7372) );
  AOI21_X1 U9152 ( .B1(n10105), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7372), .ZN(
        n7373) );
  OAI21_X1 U9153 ( .B1(n7374), .B2(n8618), .A(n7373), .ZN(n7375) );
  AOI21_X1 U9154 ( .B1(n7376), .B2(n8596), .A(n7375), .ZN(n7377) );
  OAI21_X1 U9155 ( .B1(n7379), .B2(n7378), .A(n7377), .ZN(P2_U3188) );
  NAND2_X1 U9156 ( .A1(n4625), .A2(n7380), .ZN(n7450) );
  OAI21_X1 U9157 ( .B1(n4625), .B2(n7380), .A(n7450), .ZN(n7381) );
  NOR2_X1 U9158 ( .A1(n7381), .A2(n7382), .ZN(n7453) );
  AOI21_X1 U9159 ( .B1(n7382), .B2(n7381), .A(n7453), .ZN(n7388) );
  NOR2_X1 U9160 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7383), .ZN(n9407) );
  OAI22_X1 U9161 ( .A1(n7384), .A2(n9029), .B1(n9028), .B2(n9971), .ZN(n7385)
         );
  AOI211_X1 U9162 ( .C1(n9033), .C2(n7606), .A(n9407), .B(n7385), .ZN(n7387)
         );
  NAND2_X1 U9163 ( .A1(n9051), .A2(n10031), .ZN(n7386) );
  OAI211_X1 U9164 ( .C1(n7388), .C2(n9046), .A(n7387), .B(n7386), .ZN(P1_U3227) );
  INV_X1 U9165 ( .A(n7389), .ZN(n7390) );
  OR2_X1 U9166 ( .A1(n7391), .A2(n7390), .ZN(n9129) );
  XNOR2_X1 U9167 ( .A(n7392), .B(n9129), .ZN(n7709) );
  INV_X1 U9168 ( .A(n7709), .ZN(n7401) );
  INV_X1 U9169 ( .A(n7436), .ZN(n7393) );
  AOI211_X1 U9170 ( .C1(n9131), .C2(n9984), .A(n9715), .B(n7393), .ZN(n7706)
         );
  INV_X1 U9171 ( .A(n9119), .ZN(n7394) );
  OAI21_X1 U9172 ( .B1(n7655), .B2(n7394), .A(n9261), .ZN(n9967) );
  INV_X1 U9173 ( .A(n9128), .ZN(n9973) );
  INV_X1 U9174 ( .A(n9140), .ZN(n7395) );
  AOI21_X1 U9175 ( .B1(n9967), .B2(n9973), .A(n7395), .ZN(n7434) );
  INV_X1 U9176 ( .A(n9129), .ZN(n7396) );
  XNOR2_X1 U9177 ( .A(n7434), .B(n7396), .ZN(n7397) );
  NAND2_X1 U9178 ( .A1(n7397), .A2(n10075), .ZN(n7399) );
  AOI22_X1 U9179 ( .A1(n10063), .A2(n9352), .B1(n9350), .B2(n10030), .ZN(n7398) );
  AND2_X1 U9180 ( .A1(n7399), .A2(n7398), .ZN(n7702) );
  INV_X1 U9181 ( .A(n7702), .ZN(n7400) );
  AOI211_X1 U9182 ( .C1(n7401), .C2(n10060), .A(n7706), .B(n7400), .ZN(n7406)
         );
  INV_X1 U9183 ( .A(n9879), .ZN(n9904) );
  INV_X1 U9184 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7402) );
  OAI22_X1 U9185 ( .A1(n9904), .A2(n4968), .B1(n10078), .B2(n7402), .ZN(n7403)
         );
  INV_X1 U9186 ( .A(n7403), .ZN(n7404) );
  OAI21_X1 U9187 ( .B1(n7406), .B2(n10076), .A(n7404), .ZN(P1_U3477) );
  AOI22_X1 U9188 ( .A1(n9798), .A2(n9131), .B1(n10092), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7405) );
  OAI21_X1 U9189 ( .B1(n7406), .B2(n10092), .A(n7405), .ZN(P1_U3530) );
  INV_X1 U9190 ( .A(n9546), .ZN(n7408) );
  INV_X1 U9191 ( .A(n7407), .ZN(n7447) );
  OAI222_X1 U9192 ( .A1(n8343), .A2(n10379), .B1(P1_U3086), .B2(n7408), .C1(
        n7447), .C2(n9910), .ZN(P1_U3337) );
  OAI21_X1 U9193 ( .B1(n7410), .B2(n7411), .A(n7409), .ZN(n7413) );
  INV_X1 U9194 ( .A(n7413), .ZN(n10143) );
  XNOR2_X1 U9195 ( .A(n7412), .B(n7411), .ZN(n7416) );
  NAND2_X1 U9196 ( .A1(n7413), .A2(n7953), .ZN(n7415) );
  AOI22_X1 U9197 ( .A1(n8515), .A2(n10118), .B1(n10120), .B2(n8513), .ZN(n7414) );
  OAI211_X1 U9198 ( .C1(n8757), .C2(n7416), .A(n7415), .B(n7414), .ZN(n10144)
         );
  OAI22_X1 U9199 ( .A1(n10142), .A2(n8679), .B1(n7276), .B2(n8776), .ZN(n7417)
         );
  NOR2_X1 U9200 ( .A1(n10144), .A2(n7417), .ZN(n7419) );
  MUX2_X1 U9201 ( .A(n7419), .B(n7418), .S(n10136), .Z(n7420) );
  OAI21_X1 U9202 ( .B1(n10143), .B2(n8346), .A(n7420), .ZN(P2_U3231) );
  XNOR2_X1 U9203 ( .A(n7421), .B(n7422), .ZN(n7493) );
  XNOR2_X1 U9204 ( .A(n7493), .B(n7500), .ZN(n7427) );
  INV_X1 U9205 ( .A(n7423), .ZN(n7425) );
  OAI21_X1 U9206 ( .B1(n7425), .B2(n8514), .A(n7424), .ZN(n7426) );
  AOI211_X1 U9207 ( .C1(n7427), .C2(n7426), .A(n8482), .B(n7494), .ZN(n7428)
         );
  INV_X1 U9208 ( .A(n7428), .ZN(n7432) );
  INV_X1 U9209 ( .A(n8488), .ZN(n8475) );
  OAI22_X1 U9210 ( .A1(n8496), .A2(n7620), .B1(n5351), .B2(n8477), .ZN(n7429)
         );
  AOI211_X1 U9211 ( .C1(n8475), .C2(n7666), .A(n7430), .B(n7429), .ZN(n7431)
         );
  OAI211_X1 U9212 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8490), .A(n7432), .B(
        n7431), .ZN(P2_U3158) );
  INV_X1 U9213 ( .A(n9122), .ZN(n7433) );
  AOI21_X1 U9214 ( .B1(n7434), .B2(n9141), .A(n7433), .ZN(n7435) );
  XNOR2_X1 U9215 ( .A(n7435), .B(n9077), .ZN(n7749) );
  AOI211_X1 U9216 ( .C1(n7442), .C2(n7436), .A(n9715), .B(n7468), .ZN(n7437)
         );
  AOI21_X1 U9217 ( .B1(n10030), .B2(n9349), .A(n7437), .ZN(n7754) );
  XNOR2_X1 U9218 ( .A(n7438), .B(n9077), .ZN(n7757) );
  NAND2_X1 U9219 ( .A1(n7757), .A2(n10060), .ZN(n7439) );
  OAI211_X1 U9220 ( .C1(n9969), .C2(n9970), .A(n7754), .B(n7439), .ZN(n7440)
         );
  AOI21_X1 U9221 ( .B1(n7749), .B2(n9821), .A(n7440), .ZN(n7446) );
  AOI22_X1 U9222 ( .A1(n7442), .A2(n9798), .B1(n10092), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7441) );
  OAI21_X1 U9223 ( .B1(n7446), .B2(n10092), .A(n7441), .ZN(P1_U3531) );
  INV_X1 U9224 ( .A(n7442), .ZN(n7753) );
  INV_X1 U9225 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7443) );
  OAI22_X1 U9226 ( .A1(n7753), .A2(n9904), .B1(n10078), .B2(n7443), .ZN(n7444)
         );
  INV_X1 U9227 ( .A(n7444), .ZN(n7445) );
  OAI21_X1 U9228 ( .B1(n7446), .B2(n10076), .A(n7445), .ZN(P1_U3480) );
  INV_X1 U9229 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7448) );
  OAI222_X1 U9230 ( .A1(n4517), .A2(n7448), .B1(n8607), .B2(P2_U3151), .C1(
        n8323), .C2(n7447), .ZN(P2_U3277) );
  INV_X1 U9231 ( .A(n10041), .ZN(n7660) );
  INV_X1 U9232 ( .A(n7449), .ZN(n7452) );
  INV_X1 U9233 ( .A(n7450), .ZN(n7451) );
  NOR3_X1 U9234 ( .A1(n7453), .A2(n7452), .A3(n7451), .ZN(n7456) );
  INV_X1 U9235 ( .A(n7454), .ZN(n7455) );
  OAI21_X1 U9236 ( .B1(n7456), .B2(n7455), .A(n9025), .ZN(n7460) );
  OAI22_X1 U9237 ( .A1(n7580), .A2(n9029), .B1(n9028), .B2(n7594), .ZN(n7457)
         );
  AOI211_X1 U9238 ( .C1(n9033), .C2(n7658), .A(n7458), .B(n7457), .ZN(n7459)
         );
  OAI211_X1 U9239 ( .C1(n7660), .C2(n9036), .A(n7460), .B(n7459), .ZN(P1_U3239) );
  OAI21_X1 U9240 ( .B1(n7462), .B2(n9079), .A(n7461), .ZN(n7519) );
  OAI21_X1 U9241 ( .B1(n7465), .B2(n7464), .A(n7463), .ZN(n7466) );
  INV_X1 U9242 ( .A(n7466), .ZN(n7522) );
  AOI22_X1 U9243 ( .A1(n10063), .A2(n9350), .B1(n9348), .B2(n10030), .ZN(n7469) );
  INV_X1 U9244 ( .A(n7530), .ZN(n7467) );
  INV_X1 U9245 ( .A(n9715), .ZN(n9983) );
  OAI211_X1 U9246 ( .C1(n7472), .C2(n7468), .A(n7467), .B(n9983), .ZN(n7514)
         );
  OAI211_X1 U9247 ( .C1(n7522), .C2(n9849), .A(n7469), .B(n7514), .ZN(n7470)
         );
  AOI21_X1 U9248 ( .B1(n10060), .B2(n7519), .A(n7470), .ZN(n7476) );
  INV_X1 U9249 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7471) );
  OAI22_X1 U9250 ( .A1(n7472), .A2(n9904), .B1(n10078), .B2(n7471), .ZN(n7473)
         );
  INV_X1 U9251 ( .A(n7473), .ZN(n7474) );
  OAI21_X1 U9252 ( .B1(n7476), .B2(n10076), .A(n7474), .ZN(P1_U3483) );
  AOI22_X1 U9253 ( .A1(n7870), .A2(n9798), .B1(n10092), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7475) );
  OAI21_X1 U9254 ( .B1(n7476), .B2(n10092), .A(n7475), .ZN(P1_U3532) );
  NOR2_X1 U9255 ( .A1(n7485), .A2(n7477), .ZN(n7481) );
  INV_X1 U9256 ( .A(n7478), .ZN(n7479) );
  AOI21_X1 U9257 ( .B1(n7481), .B2(n7480), .A(n7479), .ZN(n10148) );
  INV_X1 U9258 ( .A(n7482), .ZN(n7483) );
  NAND2_X1 U9259 ( .A1(n7483), .A2(n7817), .ZN(n7484) );
  NAND2_X1 U9260 ( .A1(n8779), .A2(n7484), .ZN(n8770) );
  XNOR2_X1 U9261 ( .A(n7486), .B(n7485), .ZN(n7487) );
  AOI222_X1 U9262 ( .A1(n10123), .A2(n7487), .B1(n10119), .B2(n10120), .C1(
        n8513), .C2(n10118), .ZN(n10146) );
  MUX2_X1 U9263 ( .A(n7488), .B(n10146), .S(n8779), .Z(n7492) );
  INV_X1 U9264 ( .A(n7505), .ZN(n7489) );
  AOI22_X1 U9265 ( .A1(n10130), .A2(n7490), .B1(n10133), .B2(n7489), .ZN(n7491) );
  OAI211_X1 U9266 ( .C1(n10148), .C2(n8770), .A(n7492), .B(n7491), .ZN(
        P2_U3229) );
  INV_X1 U9267 ( .A(n7493), .ZN(n7495) );
  AOI21_X1 U9268 ( .B1(n7495), .B2(n8513), .A(n7494), .ZN(n7498) );
  XNOR2_X1 U9269 ( .A(n10147), .B(n7421), .ZN(n7496) );
  NOR2_X1 U9270 ( .A1(n7496), .A2(n7666), .ZN(n7549) );
  AOI21_X1 U9271 ( .B1(n7496), .B2(n7666), .A(n7549), .ZN(n7497) );
  OAI21_X1 U9272 ( .B1(n7498), .B2(n7497), .A(n7552), .ZN(n7499) );
  NAND2_X1 U9273 ( .A1(n7499), .A2(n8472), .ZN(n7504) );
  OAI22_X1 U9274 ( .A1(n8496), .A2(n10147), .B1(n7500), .B2(n8477), .ZN(n7501)
         );
  AOI211_X1 U9275 ( .C1(n8475), .C2(n10119), .A(n7502), .B(n7501), .ZN(n7503)
         );
  OAI211_X1 U9276 ( .C1(n7505), .C2(n8490), .A(n7504), .B(n7503), .ZN(P2_U3170) );
  NOR2_X1 U9277 ( .A1(n7507), .A2(n7506), .ZN(n7508) );
  NAND2_X1 U9278 ( .A1(n7509), .A2(n7508), .ZN(n7510) );
  NAND2_X1 U9279 ( .A1(n9757), .A2(n9821), .ZN(n9747) );
  INV_X2 U9280 ( .A(n9757), .ZN(n9991) );
  NAND2_X1 U9281 ( .A1(n9757), .A2(n10064), .ZN(n9738) );
  NOR2_X1 U9282 ( .A1(n9991), .A2(n9970), .ZN(n9732) );
  NAND2_X1 U9283 ( .A1(n9732), .A2(n9350), .ZN(n7513) );
  INV_X2 U9284 ( .A(n9753), .ZN(n9977) );
  AOI22_X1 U9285 ( .A1(n9991), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9977), .B2(
        n7869), .ZN(n7512) );
  OAI211_X1 U9286 ( .C1(n9738), .C2(n7942), .A(n7513), .B(n7512), .ZN(n7516)
         );
  NAND2_X1 U9287 ( .A1(n9757), .A2(n9340), .ZN(n9741) );
  NOR2_X1 U9288 ( .A1(n7514), .A2(n9741), .ZN(n7515) );
  AOI211_X1 U9289 ( .C1(n4511), .C2(n7870), .A(n7516), .B(n7515), .ZN(n7521)
         );
  INV_X1 U9290 ( .A(n9340), .ZN(n9555) );
  NAND2_X1 U9291 ( .A1(n9555), .A2(n7517), .ZN(n9982) );
  AND2_X1 U9292 ( .A1(n9996), .A2(n9982), .ZN(n7518) );
  NAND2_X1 U9293 ( .A1(n7519), .A2(n9731), .ZN(n7520) );
  OAI211_X1 U9294 ( .C1(n7522), .C2(n9747), .A(n7521), .B(n7520), .ZN(P1_U3283) );
  AOI21_X1 U9295 ( .B1(n7523), .B2(n9063), .A(n9849), .ZN(n7525) );
  NAND2_X1 U9296 ( .A1(n7525), .A2(n7524), .ZN(n7537) );
  OAI21_X1 U9297 ( .B1(n7527), .B2(n9063), .A(n7526), .ZN(n7539) );
  NAND2_X1 U9298 ( .A1(n7539), .A2(n9731), .ZN(n7534) );
  NAND2_X1 U9299 ( .A1(n9732), .A2(n9349), .ZN(n7529) );
  AOI22_X1 U9300 ( .A1(n9734), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9977), .B2(
        n7888), .ZN(n7528) );
  OAI211_X1 U9301 ( .C1(n9738), .C2(n8003), .A(n7529), .B(n7528), .ZN(n7532)
         );
  OAI211_X1 U9302 ( .C1(n7891), .C2(n7530), .A(n9983), .B(n7682), .ZN(n7535)
         );
  NOR2_X1 U9303 ( .A1(n7535), .A2(n9741), .ZN(n7531) );
  AOI211_X1 U9304 ( .C1(n4511), .C2(n7543), .A(n7532), .B(n7531), .ZN(n7533)
         );
  OAI211_X1 U9305 ( .C1(n9991), .C2(n7537), .A(n7534), .B(n7533), .ZN(P1_U3282) );
  AOI22_X1 U9306 ( .A1(n10063), .A2(n9349), .B1(n9347), .B2(n10030), .ZN(n7536) );
  NAND3_X1 U9307 ( .A1(n7537), .A2(n7536), .A3(n7535), .ZN(n7538) );
  AOI21_X1 U9308 ( .B1(n7539), .B2(n10060), .A(n7538), .ZN(n7545) );
  INV_X1 U9309 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7540) );
  OAI22_X1 U9310 ( .A1(n7891), .A2(n9904), .B1(n10078), .B2(n7540), .ZN(n7541)
         );
  INV_X1 U9311 ( .A(n7541), .ZN(n7542) );
  OAI21_X1 U9312 ( .B1(n7545), .B2(n10076), .A(n7542), .ZN(P1_U3486) );
  AOI22_X1 U9313 ( .A1(n7543), .A2(n9798), .B1(n10092), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7544) );
  OAI21_X1 U9314 ( .B1(n7545), .B2(n10092), .A(n7544), .ZN(P1_U3533) );
  INV_X1 U9315 ( .A(n7546), .ZN(n8341) );
  OAI222_X1 U9316 ( .A1(n4517), .A2(n7548), .B1(n8323), .B2(n8341), .C1(n7547), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  INV_X1 U9317 ( .A(n7549), .ZN(n7550) );
  XNOR2_X1 U9318 ( .A(n7555), .B(n7421), .ZN(n7688) );
  XNOR2_X1 U9319 ( .A(n7688), .B(n10119), .ZN(n7551) );
  AND3_X1 U9320 ( .A1(n7552), .A2(n7551), .A3(n7550), .ZN(n7553) );
  OAI21_X1 U9321 ( .B1(n7689), .B2(n7553), .A(n8472), .ZN(n7559) );
  OAI22_X1 U9322 ( .A1(n8496), .A2(n7555), .B1(n7554), .B2(n8477), .ZN(n7556)
         );
  AOI211_X1 U9323 ( .C1(n8475), .C2(n8512), .A(n7557), .B(n7556), .ZN(n7558)
         );
  OAI211_X1 U9324 ( .C1(n7671), .C2(n8490), .A(n7559), .B(n7558), .ZN(P2_U3167) );
  XNOR2_X1 U9325 ( .A(n7561), .B(n7560), .ZN(n7575) );
  AOI21_X1 U9326 ( .B1(n5418), .B2(n7563), .A(n7562), .ZN(n7564) );
  NOR2_X1 U9327 ( .A1(n7564), .A2(n8618), .ZN(n7574) );
  AOI21_X1 U9328 ( .B1(n7820), .B2(n7566), .A(n7565), .ZN(n7572) );
  INV_X1 U9329 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7568) );
  INV_X1 U9330 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10443) );
  NOR2_X1 U9331 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10443), .ZN(n7804) );
  INV_X1 U9332 ( .A(n7804), .ZN(n7567) );
  OAI21_X1 U9333 ( .B1(n8611), .B2(n7568), .A(n7567), .ZN(n7569) );
  AOI21_X1 U9334 ( .B1(n7570), .B2(n8596), .A(n7569), .ZN(n7571) );
  OAI21_X1 U9335 ( .B1(n7572), .B2(n10100), .A(n7571), .ZN(n7573) );
  AOI211_X1 U9336 ( .C1(n7575), .C2(n10095), .A(n7574), .B(n7573), .ZN(n7576)
         );
  INV_X1 U9337 ( .A(n7576), .ZN(P2_U3189) );
  AND2_X1 U9338 ( .A1(n9253), .A2(n7577), .ZN(n9116) );
  INV_X1 U9339 ( .A(n9068), .ZN(n7633) );
  NAND2_X1 U9340 ( .A1(n9116), .A2(n7633), .ZN(n7632) );
  NAND2_X1 U9341 ( .A1(n7632), .A2(n9255), .ZN(n7610) );
  XNOR2_X1 U9342 ( .A(n7610), .B(n9069), .ZN(n7578) );
  OAI222_X1 U9343 ( .A1(n9968), .A2(n7580), .B1(n9970), .B2(n7579), .C1(n7578), 
        .C2(n9849), .ZN(n10025) );
  INV_X1 U9344 ( .A(n10025), .ZN(n7589) );
  XNOR2_X1 U9345 ( .A(n7581), .B(n9069), .ZN(n10027) );
  INV_X1 U9346 ( .A(n7627), .ZN(n7582) );
  OAI211_X1 U9347 ( .C1(n7582), .C2(n10024), .A(n9983), .B(n7604), .ZN(n10023)
         );
  NAND2_X1 U9348 ( .A1(n4511), .A2(n7583), .ZN(n7586) );
  AOI22_X1 U9349 ( .A1(n9991), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9977), .B2(
        n7584), .ZN(n7585) );
  OAI211_X1 U9350 ( .C1(n9741), .C2(n10023), .A(n7586), .B(n7585), .ZN(n7587)
         );
  AOI21_X1 U9351 ( .B1(n10027), .B2(n9731), .A(n7587), .ZN(n7588) );
  OAI21_X1 U9352 ( .B1(n7589), .B2(n9991), .A(n7588), .ZN(P1_U3289) );
  OAI21_X1 U9353 ( .B1(n7592), .B2(n7591), .A(n7590), .ZN(n7593) );
  NAND2_X1 U9354 ( .A1(n7593), .A2(n9025), .ZN(n7598) );
  OAI22_X1 U9355 ( .A1(n7594), .A2(n9029), .B1(n9028), .B2(n7866), .ZN(n7595)
         );
  AOI211_X1 U9356 ( .C1(n9033), .C2(n7703), .A(n7596), .B(n7595), .ZN(n7597)
         );
  OAI211_X1 U9357 ( .C1(n4968), .C2(n9036), .A(n7598), .B(n7597), .ZN(P1_U3221) );
  INV_X1 U9358 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10455) );
  NAND2_X1 U9359 ( .A1(n8622), .A2(P2_U3893), .ZN(n7599) );
  OAI21_X1 U9360 ( .B1(P2_U3893), .B2(n10455), .A(n7599), .ZN(P2_U3522) );
  INV_X1 U9361 ( .A(n7600), .ZN(n7701) );
  AOI21_X1 U9362 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(n9908), .A(n7601), .ZN(
        n7602) );
  OAI21_X1 U9363 ( .B1(n7701), .B2(n9910), .A(n7602), .ZN(P1_U3335) );
  XNOR2_X1 U9364 ( .A(n7603), .B(n7611), .ZN(n10036) );
  AOI21_X1 U9365 ( .B1(n7604), .B2(n10031), .A(n9715), .ZN(n7605) );
  NAND2_X1 U9366 ( .A1(n7605), .A2(n7657), .ZN(n10033) );
  INV_X1 U9367 ( .A(n9738), .ZN(n9751) );
  AOI22_X1 U9368 ( .A1(n9751), .A2(n10029), .B1(n9977), .B2(n7606), .ZN(n7608)
         );
  NAND2_X1 U9369 ( .A1(n4511), .A2(n10031), .ZN(n7607) );
  OAI211_X1 U9370 ( .C1(n10033), .C2(n9741), .A(n7608), .B(n7607), .ZN(n7618)
         );
  INV_X1 U9371 ( .A(n9135), .ZN(n7609) );
  OR2_X1 U9372 ( .A1(n7610), .A2(n7609), .ZN(n7612) );
  NAND3_X1 U9373 ( .A1(n7612), .A2(n9114), .A3(n7611), .ZN(n7613) );
  NAND3_X1 U9374 ( .A1(n7614), .A2(n10075), .A3(n7613), .ZN(n7616) );
  NAND2_X1 U9375 ( .A1(n9354), .A2(n10063), .ZN(n7615) );
  NAND2_X1 U9376 ( .A1(n7616), .A2(n7615), .ZN(n10035) );
  MUX2_X1 U9377 ( .A(n10035), .B(P1_REG2_REG_5__SCAN_IN), .S(n9734), .Z(n7617)
         );
  AOI211_X1 U9378 ( .C1(n9731), .C2(n10036), .A(n7618), .B(n7617), .ZN(n7619)
         );
  INV_X1 U9379 ( .A(n7619), .ZN(P1_U3288) );
  INV_X1 U9380 ( .A(n10130), .ZN(n8735) );
  OAI22_X1 U9381 ( .A1(n8735), .A2(n7620), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8776), .ZN(n7623) );
  MUX2_X1 U9382 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7621), .S(n8779), .Z(n7622)
         );
  AOI211_X1 U9383 ( .C1(n10132), .C2(n7624), .A(n7623), .B(n7622), .ZN(n7625)
         );
  INV_X1 U9384 ( .A(n7625), .ZN(P2_U3230) );
  XNOR2_X1 U9385 ( .A(n7626), .B(n9068), .ZN(n10021) );
  OAI211_X1 U9386 ( .C1(n7742), .C2(n10019), .A(n9983), .B(n7627), .ZN(n10017)
         );
  NAND2_X1 U9387 ( .A1(n4511), .A2(n7628), .ZN(n7631) );
  AOI22_X1 U9388 ( .A1(n9734), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9977), .B2(
        n7629), .ZN(n7630) );
  OAI211_X1 U9389 ( .C1(n9741), .C2(n10017), .A(n7631), .B(n7630), .ZN(n7636)
         );
  OAI21_X1 U9390 ( .B1(n9116), .B2(n7633), .A(n7632), .ZN(n7634) );
  AOI222_X1 U9391 ( .A1(n10075), .A2(n7634), .B1(n9997), .B2(n10063), .C1(
        n9354), .C2(n10064), .ZN(n10018) );
  NOR2_X1 U9392 ( .A1(n10018), .A2(n9991), .ZN(n7635) );
  AOI211_X1 U9393 ( .C1(n9731), .C2(n10021), .A(n7636), .B(n7635), .ZN(n7637)
         );
  INV_X1 U9394 ( .A(n7637), .ZN(P1_U3290) );
  INV_X1 U9395 ( .A(n7638), .ZN(n7639) );
  XNOR2_X1 U9396 ( .A(n7639), .B(n7649), .ZN(n7640) );
  NAND2_X1 U9397 ( .A1(n7640), .A2(n9821), .ZN(n10003) );
  NAND2_X1 U9398 ( .A1(n4511), .A2(n5919), .ZN(n7643) );
  AOI22_X1 U9399 ( .A1(n9734), .A2(P1_REG2_REG_1__SCAN_IN), .B1(n9977), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7642) );
  NAND2_X1 U9400 ( .A1(n7643), .A2(n7642), .ZN(n7648) );
  NAND2_X1 U9401 ( .A1(n5919), .A2(n9748), .ZN(n7644) );
  NAND2_X1 U9402 ( .A1(n9983), .A2(n7644), .ZN(n7645) );
  OR2_X1 U9403 ( .A1(n7645), .A2(n7744), .ZN(n9999) );
  OAI22_X1 U9404 ( .A1(n7646), .A2(n9738), .B1(n9741), .B2(n9999), .ZN(n7647)
         );
  AOI211_X1 U9405 ( .C1(n9732), .C2(n9998), .A(n7648), .B(n7647), .ZN(n7652)
         );
  XNOR2_X1 U9406 ( .A(n7650), .B(n7649), .ZN(n10008) );
  NAND2_X1 U9407 ( .A1(n9731), .A2(n10008), .ZN(n7651) );
  OAI211_X1 U9408 ( .C1(n9734), .C2(n10003), .A(n7652), .B(n7651), .ZN(
        P1_U3292) );
  INV_X1 U9409 ( .A(n7654), .ZN(n9073) );
  XNOR2_X1 U9410 ( .A(n7653), .B(n9073), .ZN(n10045) );
  INV_X1 U9411 ( .A(n9731), .ZN(n9723) );
  XNOR2_X1 U9412 ( .A(n7655), .B(n7654), .ZN(n7656) );
  AOI222_X1 U9413 ( .A1(n10075), .A2(n7656), .B1(n9352), .B2(n10064), .C1(
        n9353), .C2(n10063), .ZN(n10044) );
  MUX2_X1 U9414 ( .A(n7016), .B(n10044), .S(n9757), .Z(n7663) );
  AOI211_X1 U9415 ( .C1(n10041), .C2(n7657), .A(n9715), .B(n9985), .ZN(n10040)
         );
  INV_X1 U9416 ( .A(n9741), .ZN(n9987) );
  INV_X1 U9417 ( .A(n7658), .ZN(n7659) );
  OAI22_X1 U9418 ( .A1(n9719), .A2(n7660), .B1(n7659), .B2(n9753), .ZN(n7661)
         );
  AOI21_X1 U9419 ( .B1(n10040), .B2(n9987), .A(n7661), .ZN(n7662) );
  OAI211_X1 U9420 ( .C1(n10045), .C2(n9723), .A(n7663), .B(n7662), .ZN(
        P1_U3287) );
  XNOR2_X1 U9421 ( .A(n10127), .B(n7664), .ZN(n10152) );
  INV_X1 U9422 ( .A(n10152), .ZN(n7675) );
  XOR2_X1 U9423 ( .A(n7665), .B(n7664), .Z(n7668) );
  AOI22_X1 U9424 ( .A1(n7666), .A2(n10118), .B1(n10120), .B2(n8512), .ZN(n7667) );
  OAI21_X1 U9425 ( .B1(n7668), .B2(n8757), .A(n7667), .ZN(n7669) );
  AOI21_X1 U9426 ( .B1(n7953), .B2(n10152), .A(n7669), .ZN(n10154) );
  MUX2_X1 U9427 ( .A(n7670), .B(n10154), .S(n8779), .Z(n7674) );
  INV_X1 U9428 ( .A(n7671), .ZN(n7672) );
  AOI22_X1 U9429 ( .A1(n10130), .A2(n10151), .B1(n10133), .B2(n7672), .ZN(
        n7673) );
  OAI211_X1 U9430 ( .C1(n7675), .C2(n8346), .A(n7674), .B(n7673), .ZN(P2_U3228) );
  OAI21_X1 U9431 ( .B1(n9081), .B2(n7677), .A(n7676), .ZN(n7678) );
  AOI222_X1 U9432 ( .A1(n10075), .A2(n7678), .B1(n10062), .B2(n10064), .C1(
        n9348), .C2(n10063), .ZN(n7794) );
  OAI21_X1 U9433 ( .B1(n7681), .B2(n7680), .A(n7679), .ZN(n7790) );
  INV_X1 U9434 ( .A(n7791), .ZN(n7948) );
  NAND2_X1 U9435 ( .A1(n7682), .A2(n7791), .ZN(n7683) );
  AND2_X1 U9436 ( .A1(n7767), .A2(n7683), .ZN(n7792) );
  NOR2_X1 U9437 ( .A1(n9741), .A2(n9715), .ZN(n9749) );
  NAND2_X1 U9438 ( .A1(n7792), .A2(n9749), .ZN(n7685) );
  AOI22_X1 U9439 ( .A1(n9991), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9977), .B2(
        n7945), .ZN(n7684) );
  OAI211_X1 U9440 ( .C1(n7948), .C2(n9719), .A(n7685), .B(n7684), .ZN(n7686)
         );
  AOI21_X1 U9441 ( .B1(n7790), .B2(n9731), .A(n7686), .ZN(n7687) );
  OAI21_X1 U9442 ( .B1(n7794), .B2(n9991), .A(n7687), .ZN(P1_U3281) );
  INV_X1 U9443 ( .A(n7688), .ZN(n7690) );
  XNOR2_X1 U9444 ( .A(n7421), .B(n10131), .ZN(n7801) );
  XNOR2_X1 U9445 ( .A(n7801), .B(n8512), .ZN(n7691) );
  OAI211_X1 U9446 ( .C1(n7692), .C2(n7691), .A(n7800), .B(n8472), .ZN(n7698)
         );
  NOR2_X1 U9447 ( .A1(n8477), .A2(n7693), .ZN(n7696) );
  OAI21_X1 U9448 ( .B1(n8488), .B2(n7830), .A(n7694), .ZN(n7695) );
  AOI211_X1 U9449 ( .C1(n10131), .C2(n8378), .A(n7696), .B(n7695), .ZN(n7697)
         );
  OAI211_X1 U9450 ( .C1(n10124), .C2(n8490), .A(n7698), .B(n7697), .ZN(
        P2_U3179) );
  OAI222_X1 U9451 ( .A1(n8323), .A2(n7701), .B1(P2_U3151), .B2(n7700), .C1(
        n7699), .C2(n4517), .ZN(P2_U3275) );
  MUX2_X1 U9452 ( .A(n7073), .B(n7702), .S(n9757), .Z(n7708) );
  INV_X1 U9453 ( .A(n7703), .ZN(n7704) );
  OAI22_X1 U9454 ( .A1(n9719), .A2(n4968), .B1(n7704), .B2(n9753), .ZN(n7705)
         );
  AOI21_X1 U9455 ( .B1(n7706), .B2(n9987), .A(n7705), .ZN(n7707) );
  OAI211_X1 U9456 ( .C1(n9723), .C2(n7709), .A(n7708), .B(n7707), .ZN(P1_U3285) );
  AND2_X1 U9457 ( .A1(n7590), .A2(n7710), .ZN(n7713) );
  OAI211_X1 U9458 ( .C1(n7713), .C2(n7712), .A(n9025), .B(n7711), .ZN(n7717)
         );
  NOR2_X1 U9459 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7714), .ZN(n9417) );
  OAI22_X1 U9460 ( .A1(n9969), .A2(n9029), .B1(n9028), .B2(n7886), .ZN(n7715)
         );
  AOI211_X1 U9461 ( .C1(n9033), .C2(n7750), .A(n9417), .B(n7715), .ZN(n7716)
         );
  OAI211_X1 U9462 ( .C1(n7753), .C2(n9036), .A(n7717), .B(n7716), .ZN(P1_U3231) );
  INV_X1 U9463 ( .A(n7718), .ZN(n7719) );
  AOI21_X1 U9464 ( .B1(n7721), .B2(n7720), .A(n7719), .ZN(n7736) );
  OAI21_X1 U9465 ( .B1(n7724), .B2(n7723), .A(n7722), .ZN(n7725) );
  NAND2_X1 U9466 ( .A1(n7725), .A2(n10095), .ZN(n7735) );
  INV_X1 U9467 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10232) );
  NOR2_X1 U9468 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10566), .ZN(n7829) );
  INV_X1 U9469 ( .A(n7829), .ZN(n7726) );
  OAI21_X1 U9470 ( .B1(n8611), .B2(n10232), .A(n7726), .ZN(n7732) );
  NAND2_X1 U9471 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  AOI21_X1 U9472 ( .B1(n7730), .B2(n7729), .A(n8618), .ZN(n7731) );
  AOI211_X1 U9473 ( .C1(n8596), .C2(n7733), .A(n7732), .B(n7731), .ZN(n7734)
         );
  OAI211_X1 U9474 ( .C1(n7736), .C2(n10100), .A(n7735), .B(n7734), .ZN(
        P2_U3190) );
  XNOR2_X1 U9475 ( .A(n9064), .B(n7737), .ZN(n7738) );
  NAND2_X1 U9476 ( .A1(n7738), .A2(n9821), .ZN(n7740) );
  AOI22_X1 U9477 ( .A1(n10063), .A2(n9750), .B1(n9355), .B2(n10030), .ZN(n7739) );
  NAND2_X1 U9478 ( .A1(n7740), .A2(n7739), .ZN(n10013) );
  AOI21_X1 U9479 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n9977), .A(n10013), .ZN(
        n7748) );
  XNOR2_X1 U9480 ( .A(n7741), .B(n9064), .ZN(n10015) );
  INV_X1 U9481 ( .A(n7742), .ZN(n7743) );
  OAI211_X1 U9482 ( .C1(n10012), .C2(n7744), .A(n7743), .B(n9983), .ZN(n10011)
         );
  NOR2_X1 U9483 ( .A1(n9741), .A2(n10011), .ZN(n7746) );
  OAI22_X1 U9484 ( .A1(n9719), .A2(n10012), .B1(n7012), .B2(n9757), .ZN(n7745)
         );
  AOI211_X1 U9485 ( .C1(n9731), .C2(n10015), .A(n7746), .B(n7745), .ZN(n7747)
         );
  OAI21_X1 U9486 ( .B1(n9991), .B2(n7748), .A(n7747), .ZN(P1_U3291) );
  INV_X1 U9487 ( .A(n7749), .ZN(n7759) );
  AOI22_X1 U9488 ( .A1(n9734), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9977), .B2(
        n7750), .ZN(n7752) );
  NAND2_X1 U9489 ( .A1(n9732), .A2(n9351), .ZN(n7751) );
  OAI211_X1 U9490 ( .C1(n7753), .C2(n9719), .A(n7752), .B(n7751), .ZN(n7756)
         );
  NOR2_X1 U9491 ( .A1(n7754), .A2(n9741), .ZN(n7755) );
  AOI211_X1 U9492 ( .C1(n7757), .C2(n9731), .A(n7756), .B(n7755), .ZN(n7758)
         );
  OAI21_X1 U9493 ( .B1(n7759), .B2(n9747), .A(n7758), .ZN(P1_U3284) );
  OAI211_X1 U9494 ( .C1(n7762), .C2(n7761), .A(n7760), .B(n10075), .ZN(n7764)
         );
  AOI22_X1 U9495 ( .A1(n9346), .A2(n10064), .B1(n10063), .B2(n9347), .ZN(n7763) );
  NAND2_X1 U9496 ( .A1(n7764), .A2(n7763), .ZN(n10057) );
  INV_X1 U9497 ( .A(n10057), .ZN(n7774) );
  OAI21_X1 U9498 ( .B1(n7766), .B2(n9083), .A(n7765), .ZN(n10059) );
  NAND2_X1 U9499 ( .A1(n7997), .A2(n7767), .ZN(n7768) );
  NAND2_X1 U9500 ( .A1(n7768), .A2(n9983), .ZN(n7769) );
  OR2_X1 U9501 ( .A1(n4607), .A2(n7769), .ZN(n10056) );
  AOI22_X1 U9502 ( .A1(n9734), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9977), .B2(
        n8005), .ZN(n7771) );
  NAND2_X1 U9503 ( .A1(n7997), .A2(n4511), .ZN(n7770) );
  OAI211_X1 U9504 ( .C1(n10056), .C2(n9741), .A(n7771), .B(n7770), .ZN(n7772)
         );
  AOI21_X1 U9505 ( .B1(n10059), .B2(n9731), .A(n7772), .ZN(n7773) );
  OAI21_X1 U9506 ( .B1(n9734), .B2(n7774), .A(n7773), .ZN(P1_U3280) );
  INV_X1 U9507 ( .A(n7775), .ZN(n7788) );
  OAI222_X1 U9508 ( .A1(n8323), .A2(n7788), .B1(P2_U3151), .B2(n4809), .C1(
        n7776), .C2(n4517), .ZN(P2_U3274) );
  XNOR2_X1 U9509 ( .A(n7777), .B(n9161), .ZN(n10071) );
  OAI21_X1 U9510 ( .B1(n7779), .B2(n9161), .A(n7778), .ZN(n10074) );
  INV_X1 U9511 ( .A(n9747), .ZN(n7786) );
  OAI211_X1 U9512 ( .C1(n10069), .C2(n4607), .A(n9983), .B(n7841), .ZN(n10067)
         );
  NAND2_X1 U9513 ( .A1(n9732), .A2(n10062), .ZN(n7782) );
  INV_X1 U9514 ( .A(n7780), .ZN(n8917) );
  AOI22_X1 U9515 ( .A1(n9991), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9977), .B2(
        n8917), .ZN(n7781) );
  OAI211_X1 U9516 ( .C1(n9738), .C2(n8915), .A(n7782), .B(n7781), .ZN(n7783)
         );
  AOI21_X1 U9517 ( .B1(n9111), .B2(n4511), .A(n7783), .ZN(n7784) );
  OAI21_X1 U9518 ( .B1(n10067), .B2(n9741), .A(n7784), .ZN(n7785) );
  AOI21_X1 U9519 ( .B1(n10074), .B2(n7786), .A(n7785), .ZN(n7787) );
  OAI21_X1 U9520 ( .B1(n10071), .B2(n9723), .A(n7787), .ZN(P1_U3279) );
  OAI222_X1 U9521 ( .A1(n8343), .A2(n7789), .B1(n9910), .B2(n7788), .C1(n9066), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U9522 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7797) );
  INV_X1 U9523 ( .A(n10060), .ZN(n10070) );
  INV_X1 U9524 ( .A(n7790), .ZN(n7795) );
  INV_X1 U9525 ( .A(n10068), .ZN(n10042) );
  AOI22_X1 U9526 ( .A1(n7792), .A2(n9983), .B1(n10042), .B2(n7791), .ZN(n7793)
         );
  OAI211_X1 U9527 ( .C1(n10070), .C2(n7795), .A(n7794), .B(n7793), .ZN(n7798)
         );
  NAND2_X1 U9528 ( .A1(n7798), .A2(n10078), .ZN(n7796) );
  OAI21_X1 U9529 ( .B1(n10078), .B2(n7797), .A(n7796), .ZN(P1_U3489) );
  NAND2_X1 U9530 ( .A1(n7798), .A2(n10094), .ZN(n7799) );
  OAI21_X1 U9531 ( .B1(n10094), .B2(n7311), .A(n7799), .ZN(P1_U3534) );
  XNOR2_X1 U9532 ( .A(n7421), .B(n7823), .ZN(n7827) );
  XNOR2_X1 U9533 ( .A(n7827), .B(n7830), .ZN(n7803) );
  OAI21_X1 U9534 ( .B1(n7805), .B2(n7801), .A(n7800), .ZN(n7802) );
  AOI21_X1 U9535 ( .B1(n7803), .B2(n7802), .A(n7826), .ZN(n7810) );
  AOI21_X1 U9536 ( .B1(n8475), .B2(n8511), .A(n7804), .ZN(n7807) );
  OR2_X1 U9537 ( .A1(n8477), .A2(n7805), .ZN(n7806) );
  OAI211_X1 U9538 ( .C1(n8490), .C2(n7821), .A(n7807), .B(n7806), .ZN(n7808)
         );
  AOI21_X1 U9539 ( .B1(n7823), .B2(n8378), .A(n7808), .ZN(n7809) );
  OAI21_X1 U9540 ( .B1(n7810), .B2(n8482), .A(n7809), .ZN(P2_U3153) );
  NAND2_X1 U9541 ( .A1(n7812), .A2(n7814), .ZN(n7813) );
  NAND2_X1 U9542 ( .A1(n7811), .A2(n7813), .ZN(n10163) );
  XNOR2_X1 U9543 ( .A(n7815), .B(n7814), .ZN(n7819) );
  AOI22_X1 U9544 ( .A1(n10118), .A2(n8512), .B1(n8511), .B2(n10120), .ZN(n7816) );
  OAI21_X1 U9545 ( .B1(n10163), .B2(n7817), .A(n7816), .ZN(n7818) );
  AOI21_X1 U9546 ( .B1(n10123), .B2(n7819), .A(n7818), .ZN(n10160) );
  MUX2_X1 U9547 ( .A(n7820), .B(n10160), .S(n8779), .Z(n7825) );
  INV_X1 U9548 ( .A(n7821), .ZN(n7822) );
  AOI22_X1 U9549 ( .A1(n10130), .A2(n7823), .B1(n10133), .B2(n7822), .ZN(n7824) );
  OAI211_X1 U9550 ( .C1(n10163), .C2(n8346), .A(n7825), .B(n7824), .ZN(
        P2_U3226) );
  XNOR2_X1 U9551 ( .A(n10167), .B(n7421), .ZN(n8029) );
  XNOR2_X1 U9552 ( .A(n8029), .B(n8511), .ZN(n7828) );
  XNOR2_X1 U9553 ( .A(n8031), .B(n7828), .ZN(n7836) );
  AOI21_X1 U9554 ( .B1(n8475), .B2(n8510), .A(n7829), .ZN(n7832) );
  OR2_X1 U9555 ( .A1(n8477), .A2(n7830), .ZN(n7831) );
  OAI211_X1 U9556 ( .C1(n8490), .C2(n7833), .A(n7832), .B(n7831), .ZN(n7834)
         );
  AOI21_X1 U9557 ( .B1(n10167), .B2(n8378), .A(n7834), .ZN(n7835) );
  OAI21_X1 U9558 ( .B1(n7836), .B2(n8482), .A(n7835), .ZN(P2_U3161) );
  XNOR2_X1 U9559 ( .A(n7837), .B(n4552), .ZN(n9932) );
  INV_X1 U9560 ( .A(n9932), .ZN(n7848) );
  OAI211_X1 U9561 ( .C1(n5171), .C2(n4552), .A(n9821), .B(n7838), .ZN(n7840)
         );
  AOI22_X1 U9562 ( .A1(n9345), .A2(n10064), .B1(n10063), .B2(n9346), .ZN(n7839) );
  NAND2_X1 U9563 ( .A1(n7840), .A2(n7839), .ZN(n9930) );
  AOI21_X1 U9564 ( .B1(n7841), .B2(n9927), .A(n9715), .ZN(n7842) );
  NAND2_X1 U9565 ( .A1(n7842), .A2(n7912), .ZN(n9928) );
  INV_X1 U9566 ( .A(n9040), .ZN(n7843) );
  AOI22_X1 U9567 ( .A1(n9734), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9977), .B2(
        n7843), .ZN(n7845) );
  NAND2_X1 U9568 ( .A1(n9927), .A2(n4511), .ZN(n7844) );
  OAI211_X1 U9569 ( .C1(n9928), .C2(n9741), .A(n7845), .B(n7844), .ZN(n7846)
         );
  AOI21_X1 U9570 ( .B1(n9930), .B2(n9757), .A(n7846), .ZN(n7847) );
  OAI21_X1 U9571 ( .B1(n9723), .B2(n7848), .A(n7847), .ZN(P1_U3278) );
  INV_X1 U9572 ( .A(n7849), .ZN(n7851) );
  OAI222_X1 U9573 ( .A1(n8343), .A2(n10642), .B1(n9910), .B2(n7851), .C1(
        P1_U3086), .C2(n9299), .ZN(P1_U3333) );
  OAI222_X1 U9574 ( .A1(n4517), .A2(n7852), .B1(n8323), .B2(n7851), .C1(n7850), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI21_X1 U9575 ( .B1(n7854), .B2(n7857), .A(n7853), .ZN(n7855) );
  AOI222_X1 U9576 ( .A1(n10123), .A2(n7855), .B1(n10121), .B2(n10118), .C1(
        n8510), .C2(n10120), .ZN(n10170) );
  NAND2_X1 U9577 ( .A1(n7811), .A2(n7856), .ZN(n7858) );
  XNOR2_X1 U9578 ( .A(n7858), .B(n7857), .ZN(n10168) );
  AOI22_X1 U9579 ( .A1(n10136), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10133), .B2(
        n7859), .ZN(n7860) );
  OAI21_X1 U9580 ( .B1(n7861), .B2(n8735), .A(n7860), .ZN(n7862) );
  AOI21_X1 U9581 ( .B1(n10168), .B2(n10132), .A(n7862), .ZN(n7863) );
  OAI21_X1 U9582 ( .B1(n10170), .B2(n10136), .A(n7863), .ZN(P2_U3225) );
  AOI21_X1 U9583 ( .B1(n7865), .B2(n7864), .A(n4546), .ZN(n7873) );
  OAI22_X1 U9584 ( .A1(n7866), .A2(n9029), .B1(n9028), .B2(n7942), .ZN(n7867)
         );
  AOI211_X1 U9585 ( .C1(n9033), .C2(n7869), .A(n7868), .B(n7867), .ZN(n7872)
         );
  NAND2_X1 U9586 ( .A1(n7870), .A2(n9051), .ZN(n7871) );
  OAI211_X1 U9587 ( .C1(n7873), .C2(n9046), .A(n7872), .B(n7871), .ZN(P1_U3217) );
  NAND2_X1 U9588 ( .A1(n7877), .A2(n7874), .ZN(n7875) );
  OAI211_X1 U9589 ( .C1(n6344), .C2(n8343), .A(n7875), .B(n9336), .ZN(P1_U3332) );
  NAND2_X1 U9590 ( .A1(n7877), .A2(n7876), .ZN(n7879) );
  OAI211_X1 U9591 ( .C1(n5275), .C2(n4517), .A(n7879), .B(n7878), .ZN(P2_U3272) );
  INV_X1 U9592 ( .A(n7880), .ZN(n7882) );
  NOR3_X1 U9593 ( .A1(n4546), .A2(n7882), .A3(n7881), .ZN(n7884) );
  INV_X1 U9594 ( .A(n7883), .ZN(n7938) );
  OAI21_X1 U9595 ( .B1(n7884), .B2(n7938), .A(n9025), .ZN(n7890) );
  NOR2_X1 U9596 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7885), .ZN(n9430) );
  OAI22_X1 U9597 ( .A1(n7886), .A2(n9029), .B1(n9028), .B2(n8003), .ZN(n7887)
         );
  AOI211_X1 U9598 ( .C1(n9033), .C2(n7888), .A(n9430), .B(n7887), .ZN(n7889)
         );
  OAI211_X1 U9599 ( .C1(n7891), .C2(n9036), .A(n7890), .B(n7889), .ZN(P1_U3236) );
  AOI21_X1 U9600 ( .B1(n7893), .B2(n5445), .A(n7892), .ZN(n7907) );
  INV_X1 U9601 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10236) );
  OAI21_X1 U9602 ( .B1(n7896), .B2(n7895), .A(n7894), .ZN(n7897) );
  NAND2_X1 U9603 ( .A1(n7897), .A2(n10095), .ZN(n7899) );
  AND2_X1 U9604 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8023) );
  INV_X1 U9605 ( .A(n8023), .ZN(n7898) );
  OAI211_X1 U9606 ( .C1(n10236), .C2(n8611), .A(n7899), .B(n7898), .ZN(n7904)
         );
  AOI21_X1 U9607 ( .B1(n5446), .B2(n7901), .A(n7900), .ZN(n7902) );
  NOR2_X1 U9608 ( .A1(n7902), .A2(n10100), .ZN(n7903) );
  AOI211_X1 U9609 ( .C1(n8596), .C2(n7905), .A(n7904), .B(n7903), .ZN(n7906)
         );
  OAI21_X1 U9610 ( .B1(n7907), .B2(n8618), .A(n7906), .ZN(P2_U3191) );
  OAI21_X1 U9611 ( .B1(n7908), .B2(n9085), .A(n7984), .ZN(n9926) );
  INV_X1 U9612 ( .A(n9926), .ZN(n7919) );
  NAND2_X1 U9613 ( .A1(n9732), .A2(n10065), .ZN(n7911) );
  INV_X1 U9614 ( .A(n8962), .ZN(n7909) );
  AOI22_X1 U9615 ( .A1(n9991), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9977), .B2(
        n7909), .ZN(n7910) );
  OAI211_X1 U9616 ( .C1(n9738), .C2(n9017), .A(n7911), .B(n7910), .ZN(n7915)
         );
  INV_X1 U9617 ( .A(n8964), .ZN(n9921) );
  INV_X1 U9618 ( .A(n7912), .ZN(n7913) );
  OAI211_X1 U9619 ( .C1(n9921), .C2(n7913), .A(n9983), .B(n7988), .ZN(n9920)
         );
  NOR2_X1 U9620 ( .A1(n9920), .A2(n9741), .ZN(n7914) );
  AOI211_X1 U9621 ( .C1(n4511), .C2(n8964), .A(n7915), .B(n7914), .ZN(n7918)
         );
  NAND2_X1 U9622 ( .A1(n7916), .A2(n9085), .ZN(n9922) );
  NAND3_X1 U9623 ( .A1(n9923), .A2(n9922), .A3(n9731), .ZN(n7917) );
  OAI211_X1 U9624 ( .C1(n7919), .C2(n9747), .A(n7918), .B(n7917), .ZN(P1_U3277) );
  XNOR2_X1 U9625 ( .A(n7920), .B(n5745), .ZN(n10172) );
  OAI22_X1 U9626 ( .A1(n8024), .A2(n8760), .B1(n8028), .B2(n8762), .ZN(n7925)
         );
  NAND3_X1 U9627 ( .A1(n7853), .A2(n5745), .A3(n7922), .ZN(n7923) );
  AOI21_X1 U9628 ( .B1(n7921), .B2(n7923), .A(n8757), .ZN(n7924) );
  AOI211_X1 U9629 ( .C1(n7953), .C2(n10172), .A(n7925), .B(n7924), .ZN(n10174)
         );
  OAI22_X1 U9630 ( .A1(n8779), .A2(n5446), .B1(n8027), .B2(n8776), .ZN(n7926)
         );
  AOI21_X1 U9631 ( .B1(n10130), .B2(n10171), .A(n7926), .ZN(n7929) );
  NAND2_X1 U9632 ( .A1(n10172), .A2(n7927), .ZN(n7928) );
  OAI211_X1 U9633 ( .C1(n10174), .C2(n10136), .A(n7929), .B(n7928), .ZN(
        P2_U3224) );
  INV_X1 U9634 ( .A(n7930), .ZN(n7933) );
  OAI222_X1 U9635 ( .A1(n8323), .A2(n7933), .B1(P2_U3151), .B2(n7932), .C1(
        n7931), .C2(n4517), .ZN(P2_U3271) );
  OAI222_X1 U9636 ( .A1(n7934), .A2(P1_U3086), .B1(n9910), .B2(n7933), .C1(
        n10418), .C2(n8225), .ZN(P1_U3331) );
  INV_X1 U9637 ( .A(n7935), .ZN(n7937) );
  NOR3_X1 U9638 ( .A1(n7938), .A2(n7937), .A3(n7936), .ZN(n7941) );
  INV_X1 U9639 ( .A(n7939), .ZN(n7940) );
  OAI21_X1 U9640 ( .B1(n7941), .B2(n7940), .A(n9025), .ZN(n7947) );
  OAI22_X1 U9641 ( .A1(n7942), .A2(n9029), .B1(n9028), .B2(n8914), .ZN(n7943)
         );
  AOI211_X1 U9642 ( .C1(n9033), .C2(n7945), .A(n7944), .B(n7943), .ZN(n7946)
         );
  OAI211_X1 U9643 ( .C1(n7948), .C2(n9036), .A(n7947), .B(n7946), .ZN(P1_U3224) );
  OAI21_X1 U9644 ( .B1(n7949), .B2(n7951), .A(n8049), .ZN(n10180) );
  INV_X1 U9645 ( .A(n10180), .ZN(n7960) );
  XNOR2_X1 U9646 ( .A(n8041), .B(n7951), .ZN(n7955) );
  OAI22_X1 U9647 ( .A1(n8059), .A2(n8762), .B1(n8127), .B2(n8760), .ZN(n7952)
         );
  AOI21_X1 U9648 ( .B1(n10180), .B2(n7953), .A(n7952), .ZN(n7954) );
  OAI21_X1 U9649 ( .B1(n7955), .B2(n8757), .A(n7954), .ZN(n10178) );
  NAND2_X1 U9650 ( .A1(n10178), .A2(n8779), .ZN(n7959) );
  OAI22_X1 U9651 ( .A1(n8779), .A2(n7956), .B1(n8066), .B2(n8776), .ZN(n7957)
         );
  AOI21_X1 U9652 ( .B1(n10130), .B2(n10176), .A(n7957), .ZN(n7958) );
  OAI211_X1 U9653 ( .C1(n7960), .C2(n8346), .A(n7959), .B(n7958), .ZN(P2_U3223) );
  INV_X1 U9654 ( .A(n7961), .ZN(n7981) );
  OAI222_X1 U9655 ( .A1(n8908), .A2(n7981), .B1(P2_U3151), .B2(n7963), .C1(
        n7962), .C2(n4517), .ZN(P2_U3270) );
  AOI21_X1 U9656 ( .B1(n7965), .B2(n7964), .A(n4628), .ZN(n7980) );
  INV_X1 U9657 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10240) );
  OAI21_X1 U9658 ( .B1(n7968), .B2(n7967), .A(n7966), .ZN(n7969) );
  NAND2_X1 U9659 ( .A1(n7969), .A2(n10095), .ZN(n7971) );
  INV_X1 U9660 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10390) );
  NOR2_X1 U9661 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10390), .ZN(n8063) );
  INV_X1 U9662 ( .A(n8063), .ZN(n7970) );
  OAI211_X1 U9663 ( .C1(n10240), .C2(n8611), .A(n7971), .B(n7970), .ZN(n7977)
         );
  AOI21_X1 U9664 ( .B1(n7974), .B2(n7973), .A(n7972), .ZN(n7975) );
  NOR2_X1 U9665 ( .A1(n7975), .A2(n10100), .ZN(n7976) );
  AOI211_X1 U9666 ( .C1(n8596), .C2(n7978), .A(n7977), .B(n7976), .ZN(n7979)
         );
  OAI21_X1 U9667 ( .B1(n7980), .B2(n8618), .A(n7979), .ZN(P2_U3192) );
  OAI222_X1 U9668 ( .A1(n7982), .A2(P1_U3086), .B1(n9910), .B2(n7981), .C1(
        n10584), .C2(n8225), .ZN(P1_U3330) );
  INV_X1 U9669 ( .A(n9087), .ZN(n9166) );
  XNOR2_X1 U9670 ( .A(n7983), .B(n9166), .ZN(n9917) );
  INV_X1 U9671 ( .A(n9917), .ZN(n7996) );
  NAND2_X1 U9672 ( .A1(n9725), .A2(n9821), .ZN(n7987) );
  AOI21_X1 U9673 ( .B1(n7984), .B2(n9280), .A(n9166), .ZN(n7986) );
  AOI22_X1 U9674 ( .A1(n9711), .A2(n10064), .B1(n10063), .B2(n9345), .ZN(n7985) );
  OAI21_X1 U9675 ( .B1(n7987), .B2(n7986), .A(n7985), .ZN(n9915) );
  INV_X1 U9676 ( .A(n8977), .ZN(n9914) );
  INV_X1 U9677 ( .A(n7988), .ZN(n7990) );
  INV_X1 U9678 ( .A(n9740), .ZN(n7989) );
  OAI211_X1 U9679 ( .C1(n9914), .C2(n7990), .A(n7989), .B(n9983), .ZN(n9913)
         );
  AOI22_X1 U9680 ( .A1(n9734), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9977), .B2(
        n7991), .ZN(n7993) );
  NAND2_X1 U9681 ( .A1(n8977), .A2(n4511), .ZN(n7992) );
  OAI211_X1 U9682 ( .C1(n9913), .C2(n9741), .A(n7993), .B(n7992), .ZN(n7994)
         );
  AOI21_X1 U9683 ( .B1(n9915), .B2(n9757), .A(n7994), .ZN(n7995) );
  OAI21_X1 U9684 ( .B1(n9723), .B2(n7996), .A(n7995), .ZN(P1_U3276) );
  OAI21_X1 U9685 ( .B1(n8000), .B2(n7999), .A(n7998), .ZN(n8001) );
  NAND2_X1 U9686 ( .A1(n8001), .A2(n9025), .ZN(n8007) );
  NOR2_X1 U9687 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8002), .ZN(n9446) );
  OAI22_X1 U9688 ( .A1(n9110), .A2(n9028), .B1(n9029), .B2(n8003), .ZN(n8004)
         );
  AOI211_X1 U9689 ( .C1(n9033), .C2(n8005), .A(n9446), .B(n8004), .ZN(n8006)
         );
  OAI211_X1 U9690 ( .C1(n4974), .C2(n9036), .A(n8007), .B(n8006), .ZN(P1_U3234) );
  AOI21_X1 U9691 ( .B1(n5487), .B2(n8009), .A(n8008), .ZN(n8022) );
  AOI21_X1 U9692 ( .B1(n8011), .B2(n5486), .A(n8010), .ZN(n8018) );
  AND2_X1 U9693 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8093) );
  AOI21_X1 U9694 ( .B1(n10105), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8093), .ZN(
        n8017) );
  OAI21_X1 U9695 ( .B1(n8014), .B2(n8013), .A(n8012), .ZN(n8015) );
  NAND2_X1 U9696 ( .A1(n8015), .A2(n10095), .ZN(n8016) );
  OAI211_X1 U9697 ( .C1(n8018), .C2(n8618), .A(n8017), .B(n8016), .ZN(n8019)
         );
  AOI21_X1 U9698 ( .B1(n8020), .B2(n8596), .A(n8019), .ZN(n8021) );
  OAI21_X1 U9699 ( .B1(n8022), .B2(n10100), .A(n8021), .ZN(P2_U3193) );
  INV_X1 U9700 ( .A(n8477), .ZN(n8493) );
  AOI21_X1 U9701 ( .B1(n8493), .B2(n8511), .A(n8023), .ZN(n8026) );
  OR2_X1 U9702 ( .A1(n8488), .A2(n8024), .ZN(n8025) );
  OAI211_X1 U9703 ( .C1(n8490), .C2(n8027), .A(n8026), .B(n8025), .ZN(n8036)
         );
  XNOR2_X1 U9704 ( .A(n10171), .B(n7421), .ZN(n8058) );
  XNOR2_X1 U9705 ( .A(n8058), .B(n8059), .ZN(n8034) );
  NOR2_X1 U9706 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  INV_X1 U9707 ( .A(n8062), .ZN(n8032) );
  AOI211_X1 U9708 ( .C1(n8034), .C2(n8033), .A(n8482), .B(n8032), .ZN(n8035)
         );
  AOI211_X1 U9709 ( .C1(n10171), .C2(n8378), .A(n8036), .B(n8035), .ZN(n8037)
         );
  INV_X1 U9710 ( .A(n8037), .ZN(P2_U3171) );
  INV_X1 U9711 ( .A(n8038), .ZN(n8056) );
  OAI222_X1 U9712 ( .A1(n8908), .A2(n8056), .B1(P2_U3151), .B2(n8040), .C1(
        n8039), .C2(n4517), .ZN(P2_U3269) );
  NAND2_X1 U9713 ( .A1(n8041), .A2(n8076), .ZN(n8043) );
  NAND2_X1 U9714 ( .A1(n8043), .A2(n8042), .ZN(n8044) );
  INV_X1 U9715 ( .A(n8044), .ZN(n8045) );
  INV_X1 U9716 ( .A(n8077), .ZN(n8074) );
  OR2_X1 U9717 ( .A1(n8044), .A2(n8077), .ZN(n8181) );
  OAI211_X1 U9718 ( .C1(n8045), .C2(n8074), .A(n10123), .B(n8181), .ZN(n8047)
         );
  AOI22_X1 U9719 ( .A1(n10118), .A2(n8509), .B1(n8507), .B2(n10120), .ZN(n8046) );
  NAND2_X1 U9720 ( .A1(n8047), .A2(n8046), .ZN(n10185) );
  INV_X1 U9721 ( .A(n10185), .ZN(n8055) );
  NAND3_X1 U9722 ( .A1(n8049), .A2(n8048), .A3(n8074), .ZN(n8050) );
  NAND2_X1 U9723 ( .A1(n8051), .A2(n8050), .ZN(n10187) );
  INV_X1 U9724 ( .A(n8098), .ZN(n10184) );
  NOR2_X1 U9725 ( .A1(n10184), .A2(n8735), .ZN(n8053) );
  OAI22_X1 U9726 ( .A1(n8779), .A2(n5487), .B1(n8096), .B2(n8776), .ZN(n8052)
         );
  AOI211_X1 U9727 ( .C1(n10187), .C2(n10132), .A(n8053), .B(n8052), .ZN(n8054)
         );
  OAI21_X1 U9728 ( .B1(n8055), .B2(n10136), .A(n8054), .ZN(P2_U3222) );
  OAI222_X1 U9729 ( .A1(n8057), .A2(P1_U3086), .B1(n9910), .B2(n8056), .C1(
        n10424), .C2(n8225), .ZN(P1_U3329) );
  XNOR2_X1 U9730 ( .A(n10176), .B(n8281), .ZN(n8089) );
  INV_X1 U9731 ( .A(n8058), .ZN(n8060) );
  NAND2_X1 U9732 ( .A1(n8060), .A2(n8510), .ZN(n8061) );
  NAND2_X1 U9733 ( .A1(n8062), .A2(n8061), .ZN(n8072) );
  XNOR2_X1 U9734 ( .A(n8072), .B(n8509), .ZN(n8090) );
  XOR2_X1 U9735 ( .A(n8089), .B(n8090), .Z(n8069) );
  AOI21_X1 U9736 ( .B1(n8493), .B2(n8510), .A(n8063), .ZN(n8065) );
  OR2_X1 U9737 ( .A1(n8488), .A2(n8127), .ZN(n8064) );
  OAI211_X1 U9738 ( .C1(n8490), .C2(n8066), .A(n8065), .B(n8064), .ZN(n8067)
         );
  AOI21_X1 U9739 ( .B1(n10176), .B2(n8378), .A(n8067), .ZN(n8068) );
  OAI21_X1 U9740 ( .B1(n8069), .B2(n8482), .A(n8068), .ZN(P2_U3157) );
  XNOR2_X1 U9741 ( .A(n8077), .B(n7421), .ZN(n8092) );
  OR2_X1 U9742 ( .A1(n8089), .A2(n8509), .ZN(n8070) );
  NAND2_X1 U9743 ( .A1(n8072), .A2(n8071), .ZN(n8082) );
  NOR2_X1 U9744 ( .A1(n8073), .A2(n8281), .ZN(n8075) );
  AOI211_X1 U9745 ( .C1(n8281), .C2(n8508), .A(n8075), .B(n8074), .ZN(n8080)
         );
  NOR2_X1 U9746 ( .A1(n8076), .A2(n7421), .ZN(n8078) );
  AOI211_X1 U9747 ( .C1(n8508), .C2(n7421), .A(n8078), .B(n8077), .ZN(n8079)
         );
  XOR2_X1 U9748 ( .A(n7421), .B(n10194), .Z(n8228) );
  XNOR2_X1 U9749 ( .A(n8228), .B(n8232), .ZN(n8083) );
  XNOR2_X1 U9750 ( .A(n8229), .B(n8083), .ZN(n8088) );
  INV_X1 U9751 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10604) );
  NOR2_X1 U9752 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10604), .ZN(n8111) );
  NOR2_X1 U9753 ( .A1(n8477), .A2(n8127), .ZN(n8084) );
  AOI211_X1 U9754 ( .C1(n8475), .C2(n8506), .A(n8111), .B(n8084), .ZN(n8085)
         );
  OAI21_X1 U9755 ( .B1(n8128), .B2(n8490), .A(n8085), .ZN(n8086) );
  AOI21_X1 U9756 ( .B1(n10194), .B2(n8378), .A(n8086), .ZN(n8087) );
  OAI21_X1 U9757 ( .B1(n8088), .B2(n8482), .A(n8087), .ZN(P2_U3164) );
  OAI22_X1 U9758 ( .A1(n8090), .A2(n8089), .B1(n8509), .B2(n8072), .ZN(n8091)
         );
  XOR2_X1 U9759 ( .A(n8092), .B(n8091), .Z(n8100) );
  AOI21_X1 U9760 ( .B1(n8493), .B2(n8509), .A(n8093), .ZN(n8095) );
  OR2_X1 U9761 ( .A1(n8488), .A2(n8232), .ZN(n8094) );
  OAI211_X1 U9762 ( .C1(n8490), .C2(n8096), .A(n8095), .B(n8094), .ZN(n8097)
         );
  AOI21_X1 U9763 ( .B1(n8098), .B2(n8378), .A(n8097), .ZN(n8099) );
  OAI21_X1 U9764 ( .B1(n8100), .B2(n8482), .A(n8099), .ZN(P2_U3176) );
  INV_X1 U9765 ( .A(n8101), .ZN(n8103) );
  OAI222_X1 U9766 ( .A1(n8908), .A2(n8103), .B1(n5772), .B2(P2_U3151), .C1(
        n8102), .C2(n4517), .ZN(P2_U3267) );
  OAI222_X1 U9767 ( .A1(n8343), .A2(n10569), .B1(P1_U3086), .B2(n9378), .C1(
        n8103), .C2(n9910), .ZN(P1_U3327) );
  AOI21_X1 U9768 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(n8121) );
  INV_X1 U9769 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10248) );
  OAI21_X1 U9770 ( .B1(n8109), .B2(n8108), .A(n8107), .ZN(n8110) );
  NAND2_X1 U9771 ( .A1(n8110), .A2(n10095), .ZN(n8113) );
  INV_X1 U9772 ( .A(n8111), .ZN(n8112) );
  OAI211_X1 U9773 ( .C1(n10248), .C2(n8611), .A(n8113), .B(n8112), .ZN(n8118)
         );
  AOI21_X1 U9774 ( .B1(n4613), .B2(n8115), .A(n8114), .ZN(n8116) );
  NOR2_X1 U9775 ( .A1(n8116), .A2(n10100), .ZN(n8117) );
  AOI211_X1 U9776 ( .C1(n8596), .C2(n8119), .A(n8118), .B(n8117), .ZN(n8120)
         );
  OAI21_X1 U9777 ( .B1(n8121), .B2(n8618), .A(n8120), .ZN(P2_U3194) );
  OAI21_X1 U9778 ( .B1(n5172), .B2(n5747), .A(n8122), .ZN(n10191) );
  NAND2_X1 U9779 ( .A1(n8181), .A2(n8123), .ZN(n8125) );
  XNOR2_X1 U9780 ( .A(n8125), .B(n8124), .ZN(n8126) );
  OAI222_X1 U9781 ( .A1(n8760), .A2(n8226), .B1(n8762), .B2(n8127), .C1(n8757), 
        .C2(n8126), .ZN(n10192) );
  NAND2_X1 U9782 ( .A1(n10192), .A2(n8779), .ZN(n8132) );
  OAI22_X1 U9783 ( .A1(n8779), .A2(n8129), .B1(n8128), .B2(n8776), .ZN(n8130)
         );
  AOI21_X1 U9784 ( .B1(n10194), .B2(n10130), .A(n8130), .ZN(n8131) );
  OAI211_X1 U9785 ( .C1(n8770), .C2(n10191), .A(n8132), .B(n8131), .ZN(
        P2_U3221) );
  INV_X1 U9786 ( .A(n8134), .ZN(n8138) );
  OR2_X1 U9787 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  OAI211_X1 U9788 ( .C1(n8133), .C2(n8138), .A(n10123), .B(n8137), .ZN(n8140)
         );
  AOI22_X1 U9789 ( .A1(n8773), .A2(n10120), .B1(n10118), .B2(n8505), .ZN(n8139) );
  NAND2_X1 U9790 ( .A1(n8140), .A2(n8139), .ZN(n8200) );
  MUX2_X1 U9791 ( .A(n8200), .B(P2_REG1_REG_15__SCAN_IN), .S(n10211), .Z(n8144) );
  XNOR2_X1 U9792 ( .A(n8142), .B(n8141), .ZN(n8203) );
  INV_X1 U9793 ( .A(n8203), .ZN(n8145) );
  NAND2_X1 U9794 ( .A1(n10213), .A2(n10188), .ZN(n8823) );
  INV_X1 U9795 ( .A(n8244), .ZN(n8497) );
  OAI22_X1 U9796 ( .A1(n8145), .A2(n8823), .B1(n8497), .B2(n8829), .ZN(n8143)
         );
  OR2_X1 U9797 ( .A1(n8144), .A2(n8143), .ZN(P2_U3474) );
  MUX2_X1 U9798 ( .A(n8200), .B(P2_REG0_REG_15__SCAN_IN), .S(n10198), .Z(n8147) );
  INV_X1 U9799 ( .A(n10188), .ZN(n10190) );
  OR2_X1 U9800 ( .A1(n10198), .A2(n10190), .ZN(n8895) );
  OAI22_X1 U9801 ( .A1(n8145), .A2(n8895), .B1(n8497), .B2(n8900), .ZN(n8146)
         );
  OR2_X1 U9802 ( .A1(n8147), .A2(n8146), .ZN(P2_U3435) );
  XNOR2_X1 U9803 ( .A(n8148), .B(n8149), .ZN(n8163) );
  INV_X1 U9804 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8152) );
  XNOR2_X1 U9805 ( .A(n8150), .B(n8149), .ZN(n8151) );
  AOI222_X1 U9806 ( .A1(n10123), .A2(n8151), .B1(n8506), .B2(n10118), .C1(
        n8504), .C2(n10120), .ZN(n8158) );
  MUX2_X1 U9807 ( .A(n8152), .B(n8158), .S(n10196), .Z(n8154) );
  NAND2_X1 U9808 ( .A1(n8240), .A2(n8891), .ZN(n8153) );
  OAI211_X1 U9809 ( .C1(n8163), .C2(n8895), .A(n8154), .B(n8153), .ZN(P2_U3432) );
  MUX2_X1 U9810 ( .A(n8155), .B(n8158), .S(n10213), .Z(n8157) );
  NAND2_X1 U9811 ( .A1(n8240), .A2(n6959), .ZN(n8156) );
  OAI211_X1 U9812 ( .C1(n8823), .C2(n8163), .A(n8157), .B(n8156), .ZN(P2_U3473) );
  INV_X1 U9813 ( .A(n8158), .ZN(n8160) );
  OAI22_X1 U9814 ( .A1(n8372), .A2(n8679), .B1(n8367), .B2(n8776), .ZN(n8159)
         );
  OAI21_X1 U9815 ( .B1(n8160), .B2(n8159), .A(n8779), .ZN(n8162) );
  NAND2_X1 U9816 ( .A1(n10136), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8161) );
  OAI211_X1 U9817 ( .C1(n8163), .C2(n8770), .A(n8162), .B(n8161), .ZN(P2_U3219) );
  XNOR2_X1 U9818 ( .A(n8164), .B(n8165), .ZN(n8178) );
  INV_X1 U9819 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8168) );
  XNOR2_X1 U9820 ( .A(n8166), .B(n8165), .ZN(n8167) );
  AOI222_X1 U9821 ( .A1(n10123), .A2(n8167), .B1(n8504), .B2(n10118), .C1(
        n8503), .C2(n10120), .ZN(n8174) );
  MUX2_X1 U9822 ( .A(n8168), .B(n8174), .S(n10196), .Z(n8170) );
  NAND2_X1 U9823 ( .A1(n8414), .A2(n8891), .ZN(n8169) );
  OAI211_X1 U9824 ( .C1(n8178), .C2(n8895), .A(n8170), .B(n8169), .ZN(P2_U3438) );
  MUX2_X1 U9825 ( .A(n8171), .B(n8174), .S(n10213), .Z(n8173) );
  NAND2_X1 U9826 ( .A1(n8414), .A2(n6959), .ZN(n8172) );
  OAI211_X1 U9827 ( .C1(n8178), .C2(n8823), .A(n8173), .B(n8172), .ZN(P2_U3475) );
  MUX2_X1 U9828 ( .A(n8175), .B(n8174), .S(n8779), .Z(n8177) );
  AOI22_X1 U9829 ( .A1(n8414), .A2(n10130), .B1(n10133), .B2(n8421), .ZN(n8176) );
  OAI211_X1 U9830 ( .C1(n8178), .C2(n8770), .A(n8177), .B(n8176), .ZN(P2_U3217) );
  XNOR2_X1 U9831 ( .A(n8179), .B(n8184), .ZN(n8199) );
  INV_X1 U9832 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U9833 ( .A1(n8181), .A2(n8180), .ZN(n8183) );
  AND2_X1 U9834 ( .A1(n8183), .A2(n8182), .ZN(n8185) );
  XNOR2_X1 U9835 ( .A(n8185), .B(n8184), .ZN(n8186) );
  AOI222_X1 U9836 ( .A1(n10123), .A2(n8186), .B1(n8507), .B2(n10118), .C1(
        n8505), .C2(n10120), .ZN(n8193) );
  MUX2_X1 U9837 ( .A(n8187), .B(n8193), .S(n10196), .Z(n8189) );
  NAND2_X1 U9838 ( .A1(n8237), .A2(n8891), .ZN(n8188) );
  OAI211_X1 U9839 ( .C1(n8199), .C2(n8895), .A(n8189), .B(n8188), .ZN(P2_U3429) );
  MUX2_X1 U9840 ( .A(n8190), .B(n8193), .S(n10213), .Z(n8192) );
  NAND2_X1 U9841 ( .A1(n8237), .A2(n6959), .ZN(n8191) );
  OAI211_X1 U9842 ( .C1(n8823), .C2(n8199), .A(n8192), .B(n8191), .ZN(P2_U3472) );
  INV_X1 U9843 ( .A(n8193), .ZN(n8196) );
  OAI22_X1 U9844 ( .A1(n8194), .A2(n8679), .B1(n8235), .B2(n8776), .ZN(n8195)
         );
  OAI21_X1 U9845 ( .B1(n8196), .B2(n8195), .A(n8779), .ZN(n8198) );
  NAND2_X1 U9846 ( .A1(n10136), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8197) );
  OAI211_X1 U9847 ( .C1(n8199), .C2(n8770), .A(n8198), .B(n8197), .ZN(P2_U3220) );
  OAI22_X1 U9848 ( .A1(n8497), .A2(n8735), .B1(n8489), .B2(n8776), .ZN(n8202)
         );
  MUX2_X1 U9849 ( .A(n8200), .B(P2_REG2_REG_15__SCAN_IN), .S(n10136), .Z(n8201) );
  AOI211_X1 U9850 ( .C1(n8203), .C2(n10132), .A(n8202), .B(n8201), .ZN(n8204)
         );
  INV_X1 U9851 ( .A(n8204), .ZN(P2_U3218) );
  INV_X1 U9852 ( .A(n8618), .ZN(n10114) );
  XNOR2_X1 U9853 ( .A(n8205), .B(n5318), .ZN(n8218) );
  INV_X1 U9854 ( .A(n8206), .ZN(n8207) );
  AOI21_X1 U9855 ( .B1(n6634), .B2(n8208), .A(n8207), .ZN(n8210) );
  OAI22_X1 U9856 ( .A1(n10100), .A2(n8210), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8209), .ZN(n8217) );
  INV_X1 U9857 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8215) );
  OAI211_X1 U9858 ( .C1(n8213), .C2(n8212), .A(n8211), .B(n10095), .ZN(n8214)
         );
  OAI21_X1 U9859 ( .B1(n8611), .B2(n8215), .A(n8214), .ZN(n8216) );
  AOI211_X1 U9860 ( .C1(n10114), .C2(n8218), .A(n8217), .B(n8216), .ZN(n8219)
         );
  OAI21_X1 U9861 ( .B1(n6685), .B2(n6680), .A(n8219), .ZN(P2_U3183) );
  INV_X1 U9862 ( .A(n9059), .ZN(n8224) );
  OAI222_X1 U9863 ( .A1(n5285), .A2(P2_U3151), .B1(n8908), .B2(n8224), .C1(
        n4517), .C2(n6851), .ZN(P2_U3265) );
  INV_X1 U9864 ( .A(n8220), .ZN(n8322) );
  OAI222_X1 U9865 ( .A1(n8343), .A2(n10617), .B1(n9910), .B2(n8322), .C1(n9300), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U9866 ( .A1(n4517), .A2(n8222), .B1(n8908), .B2(n8221), .C1(
        P2_U3151), .C2(n10107), .ZN(P2_U3293) );
  INV_X1 U9867 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10402) );
  OAI222_X1 U9868 ( .A1(n8225), .A2(n10402), .B1(n9910), .B2(n8224), .C1(
        P1_U3086), .C2(n8223), .ZN(P1_U3325) );
  XNOR2_X1 U9869 ( .A(n8237), .B(n7421), .ZN(n8227) );
  NAND2_X1 U9870 ( .A1(n8227), .A2(n8226), .ZN(n8241) );
  OAI21_X1 U9871 ( .B1(n8227), .B2(n8226), .A(n8241), .ZN(n8231) );
  AOI21_X1 U9872 ( .B1(n8231), .B2(n8230), .A(n8364), .ZN(n8239) );
  NAND2_X1 U9873 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8529) );
  OAI21_X1 U9874 ( .B1(n8477), .B2(n8232), .A(n8529), .ZN(n8233) );
  AOI21_X1 U9875 ( .B1(n8475), .B2(n8505), .A(n8233), .ZN(n8234) );
  OAI21_X1 U9876 ( .B1(n8235), .B2(n8490), .A(n8234), .ZN(n8236) );
  AOI21_X1 U9877 ( .B1(n8237), .B2(n8378), .A(n8236), .ZN(n8238) );
  OAI21_X1 U9878 ( .B1(n8239), .B2(n8482), .A(n8238), .ZN(P2_U3174) );
  XNOR2_X1 U9879 ( .A(n8809), .B(n7421), .ZN(n8264) );
  INV_X1 U9880 ( .A(n8264), .ZN(n8275) );
  XNOR2_X1 U9881 ( .A(n8240), .B(n7421), .ZN(n8242) );
  INV_X1 U9882 ( .A(n8242), .ZN(n8243) );
  INV_X1 U9883 ( .A(n8241), .ZN(n8363) );
  XNOR2_X1 U9884 ( .A(n8242), .B(n8505), .ZN(n8362) );
  OAI21_X1 U9885 ( .B1(n8243), .B2(n8505), .A(n8361), .ZN(n8484) );
  INV_X1 U9886 ( .A(n8484), .ZN(n8246) );
  XNOR2_X1 U9887 ( .A(n8244), .B(n7421), .ZN(n8248) );
  XNOR2_X1 U9888 ( .A(n8248), .B(n8419), .ZN(n8483) );
  INV_X1 U9889 ( .A(n8483), .ZN(n8245) );
  XNOR2_X1 U9890 ( .A(n8414), .B(n8281), .ZN(n8247) );
  NOR2_X1 U9891 ( .A1(n8247), .A2(n8773), .ZN(n8426) );
  AOI21_X1 U9892 ( .B1(n8247), .B2(n8773), .A(n8426), .ZN(n8415) );
  INV_X1 U9893 ( .A(n8248), .ZN(n8249) );
  NAND2_X1 U9894 ( .A1(n8249), .A2(n8504), .ZN(n8416) );
  XNOR2_X1 U9895 ( .A(n8830), .B(n7421), .ZN(n8251) );
  NAND2_X1 U9896 ( .A1(n8251), .A2(n8761), .ZN(n8468) );
  INV_X1 U9897 ( .A(n8251), .ZN(n8252) );
  NAND2_X1 U9898 ( .A1(n8252), .A2(n8503), .ZN(n8253) );
  NAND2_X1 U9899 ( .A1(n8427), .A2(n8468), .ZN(n8257) );
  XNOR2_X1 U9900 ( .A(n8767), .B(n7421), .ZN(n8254) );
  NAND2_X1 U9901 ( .A1(n8254), .A2(n8744), .ZN(n8382) );
  INV_X1 U9902 ( .A(n8254), .ZN(n8255) );
  NAND2_X1 U9903 ( .A1(n8255), .A2(n8772), .ZN(n8256) );
  AND2_X1 U9904 ( .A1(n8382), .A2(n8256), .ZN(n8469) );
  NAND2_X1 U9905 ( .A1(n8257), .A2(n8469), .ZN(n8381) );
  XNOR2_X1 U9906 ( .A(n8892), .B(n7421), .ZN(n8258) );
  NAND2_X1 U9907 ( .A1(n8258), .A2(n8759), .ZN(n8445) );
  INV_X1 U9908 ( .A(n8258), .ZN(n8259) );
  NAND2_X1 U9909 ( .A1(n8259), .A2(n8728), .ZN(n8260) );
  XNOR2_X1 U9910 ( .A(n8719), .B(n7421), .ZN(n8261) );
  NAND2_X1 U9911 ( .A1(n8261), .A2(n8708), .ZN(n8456) );
  INV_X1 U9912 ( .A(n8261), .ZN(n8262) );
  INV_X1 U9913 ( .A(n8708), .ZN(n8729) );
  NAND2_X1 U9914 ( .A1(n8262), .A2(n8729), .ZN(n8263) );
  XNOR2_X1 U9915 ( .A(n8264), .B(n8501), .ZN(n8457) );
  INV_X1 U9916 ( .A(n8272), .ZN(n8265) );
  XNOR2_X1 U9917 ( .A(n8444), .B(n7421), .ZN(n8269) );
  NAND2_X1 U9918 ( .A1(n8269), .A2(n8745), .ZN(n8394) );
  INV_X1 U9919 ( .A(n8457), .ZN(n8266) );
  INV_X1 U9920 ( .A(n8268), .ZN(n8274) );
  INV_X1 U9921 ( .A(n8269), .ZN(n8270) );
  NAND2_X1 U9922 ( .A1(n8270), .A2(n8502), .ZN(n8271) );
  OAI21_X1 U9923 ( .B1(n8275), .B2(n8501), .A(n8460), .ZN(n8279) );
  INV_X1 U9924 ( .A(n8279), .ZN(n8277) );
  XNOR2_X1 U9925 ( .A(n8872), .B(n7421), .ZN(n8278) );
  INV_X1 U9926 ( .A(n8278), .ZN(n8276) );
  XNOR2_X1 U9927 ( .A(n8680), .B(n8281), .ZN(n8282) );
  NAND2_X1 U9928 ( .A1(n8282), .A2(n8692), .ZN(n8404) );
  INV_X1 U9929 ( .A(n8282), .ZN(n8283) );
  NAND2_X1 U9930 ( .A1(n8283), .A2(n8500), .ZN(n8284) );
  NAND2_X1 U9931 ( .A1(n8403), .A2(n8404), .ZN(n8288) );
  XNOR2_X1 U9932 ( .A(n8860), .B(n7421), .ZN(n8285) );
  NAND2_X1 U9933 ( .A1(n8285), .A2(n8653), .ZN(n8290) );
  INV_X1 U9934 ( .A(n8285), .ZN(n8286) );
  INV_X1 U9935 ( .A(n8653), .ZN(n8676) );
  NAND2_X1 U9936 ( .A1(n8286), .A2(n8676), .ZN(n8287) );
  INV_X1 U9937 ( .A(n8290), .ZN(n8289) );
  XNOR2_X1 U9938 ( .A(n8324), .B(n8664), .ZN(n8292) );
  NOR3_X1 U9939 ( .A1(n8407), .A2(n8289), .A3(n8292), .ZN(n8301) );
  INV_X1 U9940 ( .A(n8292), .ZN(n8291) );
  INV_X1 U9941 ( .A(n8296), .ZN(n8294) );
  AND2_X1 U9942 ( .A1(n8405), .A2(n8292), .ZN(n8293) );
  INV_X1 U9943 ( .A(n8295), .ZN(n8298) );
  AND2_X1 U9944 ( .A1(n8404), .A2(n8296), .ZN(n8297) );
  OAI21_X1 U9945 ( .B1(n8301), .B2(n4914), .A(n8472), .ZN(n8305) );
  INV_X1 U9946 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10602) );
  OAI22_X1 U9947 ( .A1(n8653), .A2(n8477), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10602), .ZN(n8303) );
  NOR2_X1 U9948 ( .A1(n8654), .A2(n8488), .ZN(n8302) );
  AOI211_X1 U9949 ( .C1(n8657), .C2(n8479), .A(n8303), .B(n8302), .ZN(n8304)
         );
  OAI211_X1 U9950 ( .C1(n8856), .C2(n8496), .A(n8305), .B(n8304), .ZN(P2_U3180) );
  AOI22_X1 U9951 ( .A1(n9734), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9977), .B2(
        n8306), .ZN(n8309) );
  NAND2_X1 U9952 ( .A1(n8307), .A2(n4511), .ZN(n8308) );
  OAI211_X1 U9953 ( .C1(n8310), .C2(n9741), .A(n8309), .B(n8308), .ZN(n8311)
         );
  AOI21_X1 U9954 ( .B1(n8312), .B2(n9731), .A(n8311), .ZN(n8313) );
  OAI21_X1 U9955 ( .B1(n8314), .B2(n9991), .A(n8313), .ZN(P1_U3356) );
  OAI222_X1 U9956 ( .A1(n8343), .A2(n8316), .B1(P1_U3086), .B2(n8315), .C1(
        n8319), .C2(n9910), .ZN(P1_U3326) );
  OAI222_X1 U9957 ( .A1(n8323), .A2(n8319), .B1(P2_U3151), .B2(n8318), .C1(
        n8317), .C2(n4517), .ZN(P2_U3266) );
  OAI222_X1 U9958 ( .A1(n8323), .A2(n8322), .B1(n8321), .B2(P2_U3151), .C1(
        n8320), .C2(n4517), .ZN(P2_U3268) );
  INV_X1 U9959 ( .A(n8324), .ZN(n8325) );
  NAND2_X1 U9960 ( .A1(n8327), .A2(n8326), .ZN(n8352) );
  INV_X1 U9961 ( .A(n8352), .ZN(n8329) );
  XNOR2_X1 U9962 ( .A(n8849), .B(n7421), .ZN(n8330) );
  XNOR2_X1 U9963 ( .A(n8330), .B(n8654), .ZN(n8351) );
  NAND2_X1 U9964 ( .A1(n8329), .A2(n8328), .ZN(n8353) );
  INV_X1 U9965 ( .A(n8330), .ZN(n8331) );
  NAND2_X1 U9966 ( .A1(n8331), .A2(n8633), .ZN(n8332) );
  NAND2_X1 U9967 ( .A1(n8353), .A2(n8332), .ZN(n8334) );
  XNOR2_X1 U9968 ( .A(n8334), .B(n8333), .ZN(n8340) );
  INV_X1 U9969 ( .A(n8639), .ZN(n8336) );
  OAI22_X1 U9970 ( .A1(n8336), .A2(n8490), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8335), .ZN(n8338) );
  OAI22_X1 U9971 ( .A1(n8654), .A2(n8477), .B1(n8499), .B2(n8488), .ZN(n8337)
         );
  AOI211_X1 U9972 ( .C1(n8843), .C2(n8378), .A(n8338), .B(n8337), .ZN(n8339)
         );
  OAI21_X1 U9973 ( .B1(n8340), .B2(n8482), .A(n8339), .ZN(P2_U3160) );
  OAI222_X1 U9974 ( .A1(n8343), .A2(n8342), .B1(n9910), .B2(n8341), .C1(
        P1_U3086), .C2(n9340), .ZN(P1_U3336) );
  AOI22_X1 U9975 ( .A1(n8620), .A2(n10133), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10136), .ZN(n8345) );
  NAND2_X1 U9976 ( .A1(n5828), .A2(n10130), .ZN(n8344) );
  OAI211_X1 U9977 ( .C1(n8347), .C2(n8346), .A(n8345), .B(n8344), .ZN(n8348)
         );
  INV_X1 U9978 ( .A(n8348), .ZN(n8349) );
  OAI21_X1 U9979 ( .B1(n8350), .B2(n10136), .A(n8349), .ZN(P2_U3204) );
  AOI21_X1 U9980 ( .B1(n8352), .B2(n8351), .A(n8482), .ZN(n8354) );
  NAND2_X1 U9981 ( .A1(n8354), .A2(n8353), .ZN(n8359) );
  INV_X1 U9982 ( .A(n8648), .ZN(n8356) );
  AOI22_X1 U9983 ( .A1(n8645), .A2(n8493), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8355) );
  OAI21_X1 U9984 ( .B1(n8356), .B2(n8490), .A(n8355), .ZN(n8357) );
  AOI21_X1 U9985 ( .B1(n8646), .B2(n8475), .A(n8357), .ZN(n8358) );
  OAI211_X1 U9986 ( .C1(n8360), .C2(n8496), .A(n8359), .B(n8358), .ZN(P2_U3154) );
  INV_X1 U9987 ( .A(n8361), .ZN(n8366) );
  NOR3_X1 U9988 ( .A1(n8364), .A2(n8363), .A3(n8362), .ZN(n8365) );
  OAI21_X1 U9989 ( .B1(n8366), .B2(n8365), .A(n8472), .ZN(n8371) );
  NAND2_X1 U9990 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8541) );
  OAI21_X1 U9991 ( .B1(n8488), .B2(n8419), .A(n8541), .ZN(n8369) );
  NOR2_X1 U9992 ( .A1(n8490), .A2(n8367), .ZN(n8368) );
  AOI211_X1 U9993 ( .C1(n8493), .C2(n8506), .A(n8369), .B(n8368), .ZN(n8370)
         );
  OAI211_X1 U9994 ( .C1(n8372), .C2(n8496), .A(n8371), .B(n8370), .ZN(P2_U3155) );
  INV_X1 U9995 ( .A(n8373), .ZN(n8437) );
  AOI21_X1 U9996 ( .B1(n8677), .B2(n8374), .A(n8437), .ZN(n8380) );
  AOI22_X1 U9997 ( .A1(n8501), .A2(n8493), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8376) );
  NAND2_X1 U9998 ( .A1(n8479), .A2(n8694), .ZN(n8375) );
  OAI211_X1 U9999 ( .C1(n8692), .C2(n8488), .A(n8376), .B(n8375), .ZN(n8377)
         );
  AOI21_X1 U10000 ( .B1(n8872), .B2(n8378), .A(n8377), .ZN(n8379) );
  OAI21_X1 U10001 ( .B1(n8380), .B2(n8482), .A(n8379), .ZN(P2_U3156) );
  INV_X1 U10002 ( .A(n8892), .ZN(n8390) );
  INV_X1 U10003 ( .A(n8381), .ZN(n8473) );
  NOR3_X1 U10004 ( .A1(n8473), .A2(n4906), .A3(n8383), .ZN(n8384) );
  INV_X1 U10005 ( .A(n8391), .ZN(n8448) );
  OAI21_X1 U10006 ( .B1(n8384), .B2(n8448), .A(n8472), .ZN(n8389) );
  NAND2_X1 U10007 ( .A1(n8493), .A2(n8772), .ZN(n8386) );
  OAI211_X1 U10008 ( .C1(n8745), .C2(n8488), .A(n8386), .B(n8385), .ZN(n8387)
         );
  AOI21_X1 U10009 ( .B1(n8479), .B2(n8750), .A(n8387), .ZN(n8388) );
  OAI211_X1 U10010 ( .C1(n8390), .C2(n8496), .A(n8389), .B(n8388), .ZN(
        P2_U3159) );
  NAND2_X1 U10011 ( .A1(n8391), .A2(n8445), .ZN(n8392) );
  NAND2_X1 U10012 ( .A1(n8392), .A2(n8446), .ZN(n8395) );
  INV_X1 U10013 ( .A(n8395), .ZN(n8449) );
  INV_X1 U10014 ( .A(n8394), .ZN(n8393) );
  NOR3_X1 U10015 ( .A1(n8449), .A2(n8393), .A3(n8396), .ZN(n8398) );
  NAND2_X1 U10016 ( .A1(n8395), .A2(n8394), .ZN(n8397) );
  OAI21_X1 U10017 ( .B1(n8398), .B2(n8459), .A(n8472), .ZN(n8402) );
  NOR2_X1 U10018 ( .A1(n8745), .A2(n8477), .ZN(n8400) );
  OAI22_X1 U10019 ( .A1(n8717), .A2(n8488), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10441), .ZN(n8399) );
  AOI211_X1 U10020 ( .C1(n8718), .C2(n8479), .A(n8400), .B(n8399), .ZN(n8401)
         );
  OAI211_X1 U10021 ( .C1(n8881), .C2(n8496), .A(n8402), .B(n8401), .ZN(
        P2_U3163) );
  INV_X1 U10022 ( .A(n8404), .ZN(n8406) );
  NOR3_X1 U10023 ( .A1(n8438), .A2(n8406), .A3(n8405), .ZN(n8408) );
  OAI21_X1 U10024 ( .B1(n8408), .B2(n8407), .A(n8472), .ZN(n8413) );
  OAI22_X1 U10025 ( .A1(n8692), .A2(n8477), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8409), .ZN(n8411) );
  NOR2_X1 U10026 ( .A1(n8664), .A2(n8488), .ZN(n8410) );
  AOI211_X1 U10027 ( .C1(n8666), .C2(n8479), .A(n8411), .B(n8410), .ZN(n8412)
         );
  OAI211_X1 U10028 ( .C1(n8798), .C2(n8496), .A(n8413), .B(n8412), .ZN(
        P2_U3165) );
  INV_X1 U10029 ( .A(n8414), .ZN(n8424) );
  AOI21_X1 U10030 ( .B1(n8485), .B2(n8416), .A(n8415), .ZN(n8417) );
  OAI21_X1 U10031 ( .B1(n4604), .B2(n8417), .A(n8472), .ZN(n8423) );
  NAND2_X1 U10032 ( .A1(n8475), .A2(n8503), .ZN(n8418) );
  NAND2_X1 U10033 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8574) );
  OAI211_X1 U10034 ( .C1(n8419), .C2(n8477), .A(n8418), .B(n8574), .ZN(n8420)
         );
  AOI21_X1 U10035 ( .B1(n8479), .B2(n8421), .A(n8420), .ZN(n8422) );
  OAI211_X1 U10036 ( .C1(n8424), .C2(n8496), .A(n8423), .B(n8422), .ZN(
        P2_U3166) );
  INV_X1 U10037 ( .A(n8830), .ZN(n8433) );
  NOR3_X1 U10038 ( .A1(n4604), .A2(n8426), .A3(n8425), .ZN(n8428) );
  INV_X1 U10039 ( .A(n8427), .ZN(n8471) );
  OAI21_X1 U10040 ( .B1(n8428), .B2(n8471), .A(n8472), .ZN(n8432) );
  NAND2_X1 U10041 ( .A1(n8475), .A2(n8772), .ZN(n8429) );
  NAND2_X1 U10042 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8595) );
  OAI211_X1 U10043 ( .C1(n8487), .C2(n8477), .A(n8429), .B(n8595), .ZN(n8430)
         );
  AOI21_X1 U10044 ( .B1(n8479), .B2(n8775), .A(n8430), .ZN(n8431) );
  OAI211_X1 U10045 ( .C1(n8433), .C2(n8496), .A(n8432), .B(n8431), .ZN(
        P2_U3168) );
  INV_X1 U10046 ( .A(n8434), .ZN(n8436) );
  NOR3_X1 U10047 ( .A1(n8437), .A2(n8436), .A3(n8435), .ZN(n8439) );
  OAI21_X1 U10048 ( .B1(n8439), .B2(n8438), .A(n8472), .ZN(n8443) );
  AOI22_X1 U10049 ( .A1(n8677), .A2(n8493), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8440) );
  OAI21_X1 U10050 ( .B1(n8653), .B2(n8488), .A(n8440), .ZN(n8441) );
  AOI21_X1 U10051 ( .B1(n8682), .B2(n8479), .A(n8441), .ZN(n8442) );
  OAI211_X1 U10052 ( .C1(n8680), .C2(n8496), .A(n8443), .B(n8442), .ZN(
        P2_U3169) );
  INV_X1 U10053 ( .A(n8444), .ZN(n8888) );
  INV_X1 U10054 ( .A(n8445), .ZN(n8447) );
  NOR3_X1 U10055 ( .A1(n8448), .A2(n8447), .A3(n8446), .ZN(n8450) );
  OAI21_X1 U10056 ( .B1(n8450), .B2(n8449), .A(n8472), .ZN(n8455) );
  NOR2_X1 U10057 ( .A1(n8477), .A2(n8759), .ZN(n8453) );
  OAI22_X1 U10058 ( .A1(n8708), .A2(n8488), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8451), .ZN(n8452) );
  AOI211_X1 U10059 ( .C1(n8479), .C2(n8733), .A(n8453), .B(n8452), .ZN(n8454)
         );
  OAI211_X1 U10060 ( .C1(n8888), .C2(n8496), .A(n8455), .B(n8454), .ZN(
        P2_U3173) );
  INV_X1 U10061 ( .A(n8809), .ZN(n8467) );
  INV_X1 U10062 ( .A(n8456), .ZN(n8458) );
  NOR3_X1 U10063 ( .A1(n8459), .A2(n8458), .A3(n8457), .ZN(n8462) );
  INV_X1 U10064 ( .A(n8460), .ZN(n8461) );
  OAI21_X1 U10065 ( .B1(n8462), .B2(n8461), .A(n8472), .ZN(n8466) );
  AOI22_X1 U10066 ( .A1(n8729), .A2(n8493), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8463) );
  OAI21_X1 U10067 ( .B1(n8707), .B2(n8488), .A(n8463), .ZN(n8464) );
  AOI21_X1 U10068 ( .B1(n8709), .B2(n8479), .A(n8464), .ZN(n8465) );
  OAI211_X1 U10069 ( .C1(n8467), .C2(n8496), .A(n8466), .B(n8465), .ZN(
        P2_U3175) );
  INV_X1 U10070 ( .A(n8767), .ZN(n8901) );
  INV_X1 U10071 ( .A(n8468), .ZN(n8470) );
  NOR3_X1 U10072 ( .A1(n8471), .A2(n8470), .A3(n8469), .ZN(n8474) );
  OAI21_X1 U10073 ( .B1(n8474), .B2(n8473), .A(n8472), .ZN(n8481) );
  NAND2_X1 U10074 ( .A1(n8475), .A2(n8728), .ZN(n8476) );
  NAND2_X1 U10075 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8609) );
  OAI211_X1 U10076 ( .C1(n8761), .C2(n8477), .A(n8476), .B(n8609), .ZN(n8478)
         );
  AOI21_X1 U10077 ( .B1(n8479), .B2(n8763), .A(n8478), .ZN(n8480) );
  OAI211_X1 U10078 ( .C1(n8901), .C2(n8496), .A(n8481), .B(n8480), .ZN(
        P2_U3178) );
  AOI21_X1 U10079 ( .B1(n8484), .B2(n8483), .A(n8482), .ZN(n8486) );
  NAND2_X1 U10080 ( .A1(n8486), .A2(n8485), .ZN(n8495) );
  NAND2_X1 U10081 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8557) );
  OAI21_X1 U10082 ( .B1(n8488), .B2(n8487), .A(n8557), .ZN(n8492) );
  NOR2_X1 U10083 ( .A1(n8490), .A2(n8489), .ZN(n8491) );
  AOI211_X1 U10084 ( .C1(n8493), .C2(n8505), .A(n8492), .B(n8491), .ZN(n8494)
         );
  OAI211_X1 U10085 ( .C1(n8497), .C2(n8496), .A(n8495), .B(n8494), .ZN(
        P2_U3181) );
  MUX2_X1 U10086 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8498), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10087 ( .A(n8499), .ZN(n8632) );
  MUX2_X1 U10088 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8632), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10089 ( .A(n8646), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8606), .Z(
        P2_U3519) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8633), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10091 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8645), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10092 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8676), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10093 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8500), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10094 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8501), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10095 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8729), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10096 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8502), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10097 ( .A(n8728), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8606), .Z(
        P2_U3510) );
  MUX2_X1 U10098 ( .A(n8772), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8606), .Z(
        P2_U3509) );
  MUX2_X1 U10099 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8503), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10100 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8773), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10101 ( .A(n8504), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8606), .Z(
        P2_U3506) );
  MUX2_X1 U10102 ( .A(n8505), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8606), .Z(
        P2_U3505) );
  MUX2_X1 U10103 ( .A(n8506), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8606), .Z(
        P2_U3504) );
  MUX2_X1 U10104 ( .A(n8507), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8606), .Z(
        P2_U3503) );
  MUX2_X1 U10105 ( .A(n8508), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8606), .Z(
        P2_U3502) );
  MUX2_X1 U10106 ( .A(n8509), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8606), .Z(
        P2_U3501) );
  MUX2_X1 U10107 ( .A(n8510), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8606), .Z(
        P2_U3500) );
  MUX2_X1 U10108 ( .A(n8511), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8606), .Z(
        P2_U3499) );
  MUX2_X1 U10109 ( .A(n10121), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8606), .Z(
        P2_U3498) );
  MUX2_X1 U10110 ( .A(n8512), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8606), .Z(
        P2_U3497) );
  MUX2_X1 U10111 ( .A(n10119), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8606), .Z(
        P2_U3496) );
  MUX2_X1 U10112 ( .A(n8513), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8606), .Z(
        P2_U3494) );
  MUX2_X1 U10113 ( .A(n8514), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8606), .Z(
        P2_U3493) );
  MUX2_X1 U10114 ( .A(n8515), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8606), .Z(
        P2_U3492) );
  MUX2_X1 U10115 ( .A(n8516), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8606), .Z(
        P2_U3491) );
  AOI21_X1 U10116 ( .B1(n8519), .B2(n8518), .A(n8517), .ZN(n8534) );
  INV_X1 U10117 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10252) );
  INV_X1 U10118 ( .A(n8520), .ZN(n8523) );
  INV_X1 U10119 ( .A(n8521), .ZN(n8522) );
  OAI21_X1 U10120 ( .B1(n8523), .B2(P2_REG1_REG_13__SCAN_IN), .A(n8522), .ZN(
        n8528) );
  OAI21_X1 U10121 ( .B1(n8526), .B2(n8525), .A(n8524), .ZN(n8527) );
  AOI22_X1 U10122 ( .A1(n10114), .A2(n8528), .B1(n8527), .B2(n10095), .ZN(
        n8530) );
  OAI211_X1 U10123 ( .C1(n10252), .C2(n8611), .A(n8530), .B(n8529), .ZN(n8531)
         );
  AOI21_X1 U10124 ( .B1(n8532), .B2(n8596), .A(n8531), .ZN(n8533) );
  OAI21_X1 U10125 ( .B1(n8534), .B2(n10100), .A(n8533), .ZN(P2_U3195) );
  AOI21_X1 U10126 ( .B1(n4610), .B2(n8536), .A(n8535), .ZN(n8551) );
  INV_X1 U10127 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10256) );
  OAI21_X1 U10128 ( .B1(n8539), .B2(n8538), .A(n8537), .ZN(n8540) );
  NAND2_X1 U10129 ( .A1(n8540), .A2(n10095), .ZN(n8542) );
  OAI211_X1 U10130 ( .C1(n8611), .C2(n10256), .A(n8542), .B(n8541), .ZN(n8548)
         );
  AOI21_X1 U10131 ( .B1(n8545), .B2(n8544), .A(n8543), .ZN(n8546) );
  NOR2_X1 U10132 ( .A1(n8546), .A2(n10100), .ZN(n8547) );
  AOI211_X1 U10133 ( .C1(n8596), .C2(n8549), .A(n8548), .B(n8547), .ZN(n8550)
         );
  OAI21_X1 U10134 ( .B1(n8551), .B2(n8618), .A(n8550), .ZN(P2_U3196) );
  AOI21_X1 U10135 ( .B1(n6614), .B2(n8553), .A(n8552), .ZN(n8567) );
  OAI21_X1 U10136 ( .B1(n8556), .B2(n8555), .A(n8554), .ZN(n8565) );
  INV_X1 U10137 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10260) );
  OAI21_X1 U10138 ( .B1(n8611), .B2(n10260), .A(n8557), .ZN(n8564) );
  AOI21_X1 U10139 ( .B1(n8560), .B2(n8559), .A(n8558), .ZN(n8561) );
  OAI22_X1 U10140 ( .A1(n6680), .A2(n8562), .B1(n8561), .B2(n8618), .ZN(n8563)
         );
  AOI211_X1 U10141 ( .C1(n10095), .C2(n8565), .A(n8564), .B(n8563), .ZN(n8566)
         );
  OAI21_X1 U10142 ( .B1(n8567), .B2(n10100), .A(n8566), .ZN(P2_U3197) );
  AOI21_X1 U10143 ( .B1(n4574), .B2(n8569), .A(n8568), .ZN(n8584) );
  INV_X1 U10144 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10264) );
  OAI21_X1 U10145 ( .B1(n8572), .B2(n8571), .A(n8570), .ZN(n8573) );
  NAND2_X1 U10146 ( .A1(n8573), .A2(n10095), .ZN(n8575) );
  OAI211_X1 U10147 ( .C1(n10264), .C2(n8611), .A(n8575), .B(n8574), .ZN(n8581)
         );
  AOI21_X1 U10148 ( .B1(n8578), .B2(n8577), .A(n8576), .ZN(n8579) );
  NOR2_X1 U10149 ( .A1(n8579), .A2(n10100), .ZN(n8580) );
  AOI211_X1 U10150 ( .C1(n8596), .C2(n8582), .A(n8581), .B(n8580), .ZN(n8583)
         );
  OAI21_X1 U10151 ( .B1(n8584), .B2(n8618), .A(n8583), .ZN(P2_U3198) );
  AOI21_X1 U10152 ( .B1(n8778), .B2(n8586), .A(n8585), .ZN(n8599) );
  INV_X1 U10153 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10267) );
  OAI21_X1 U10154 ( .B1(n8589), .B2(n8588), .A(n8587), .ZN(n8594) );
  INV_X1 U10155 ( .A(n8590), .ZN(n8593) );
  INV_X1 U10156 ( .A(n8591), .ZN(n8592) );
  OAI21_X1 U10157 ( .B1(n8599), .B2(n10100), .A(n8598), .ZN(P2_U3199) );
  AOI21_X1 U10158 ( .B1(n8602), .B2(n8601), .A(n8600), .ZN(n8619) );
  INV_X1 U10159 ( .A(n8603), .ZN(n8605) );
  NAND2_X1 U10160 ( .A1(n8605), .A2(n8604), .ZN(n8608) );
  OAI21_X1 U10161 ( .B1(n8608), .B2(n8606), .A(n6680), .ZN(n8616) );
  INV_X1 U10162 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10271) );
  NAND3_X1 U10163 ( .A1(n8608), .A2(n10095), .A3(n8607), .ZN(n8610) );
  OAI211_X1 U10164 ( .C1(n10271), .C2(n8611), .A(n8610), .B(n8609), .ZN(n8615)
         );
  NAND2_X1 U10165 ( .A1(n8620), .A2(n10133), .ZN(n8623) );
  NAND2_X1 U10166 ( .A1(n8622), .A2(n8621), .ZN(n8835) );
  AOI21_X1 U10167 ( .B1(n8623), .B2(n8835), .A(n10136), .ZN(n8626) );
  AOI21_X1 U10168 ( .B1(n10136), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8626), .ZN(
        n8624) );
  OAI21_X1 U10169 ( .B1(n8625), .B2(n8735), .A(n8624), .ZN(P2_U3202) );
  AOI21_X1 U10170 ( .B1(n10136), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8626), .ZN(
        n8627) );
  OAI21_X1 U10171 ( .B1(n8628), .B2(n8735), .A(n8627), .ZN(P2_U3203) );
  INV_X1 U10172 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U10173 ( .A1(n8632), .A2(n10120), .ZN(n8635) );
  MUX2_X1 U10174 ( .A(n8638), .B(n8841), .S(n8779), .Z(n8641) );
  AOI22_X1 U10175 ( .A1(n8843), .A2(n10130), .B1(n10133), .B2(n8639), .ZN(
        n8640) );
  OAI211_X1 U10176 ( .C1(n8846), .C2(n8770), .A(n8641), .B(n8640), .ZN(
        P2_U3205) );
  INV_X1 U10177 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8647) );
  MUX2_X1 U10178 ( .A(n8647), .B(n8847), .S(n8779), .Z(n8650) );
  AOI22_X1 U10179 ( .A1(n8849), .A2(n10130), .B1(n10133), .B2(n8648), .ZN(
        n8649) );
  OAI211_X1 U10180 ( .C1(n8852), .C2(n8770), .A(n8650), .B(n8649), .ZN(
        P2_U3206) );
  XOR2_X1 U10181 ( .A(n8656), .B(n8651), .Z(n8652) );
  OAI222_X1 U10182 ( .A1(n8760), .A2(n8654), .B1(n8762), .B2(n8653), .C1(n8652), .C2(n8757), .ZN(n8794) );
  INV_X1 U10183 ( .A(n8794), .ZN(n8661) );
  XOR2_X1 U10184 ( .A(n8656), .B(n8655), .Z(n8795) );
  AOI22_X1 U10185 ( .A1(n8657), .A2(n10133), .B1(n10136), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8658) );
  OAI21_X1 U10186 ( .B1(n8856), .B2(n8735), .A(n8658), .ZN(n8659) );
  AOI21_X1 U10187 ( .B1(n8795), .B2(n10132), .A(n8659), .ZN(n8660) );
  OAI21_X1 U10188 ( .B1(n8661), .B2(n10136), .A(n8660), .ZN(P2_U3207) );
  NOR2_X1 U10189 ( .A1(n8798), .A2(n8679), .ZN(n8665) );
  XOR2_X1 U10190 ( .A(n8667), .B(n8662), .Z(n8663) );
  OAI222_X1 U10191 ( .A1(n8762), .A2(n8692), .B1(n8760), .B2(n8664), .C1(n8757), .C2(n8663), .ZN(n8857) );
  AOI211_X1 U10192 ( .C1(n10133), .C2(n8666), .A(n8665), .B(n8857), .ZN(n8671)
         );
  XOR2_X1 U10193 ( .A(n8668), .B(n8667), .Z(n8863) );
  INV_X1 U10194 ( .A(n8863), .ZN(n8669) );
  AOI22_X1 U10195 ( .A1(n8669), .A2(n10132), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10136), .ZN(n8670) );
  OAI21_X1 U10196 ( .B1(n8671), .B2(n10136), .A(n8670), .ZN(P2_U3208) );
  XNOR2_X1 U10197 ( .A(n8672), .B(n8674), .ZN(n8869) );
  XNOR2_X1 U10198 ( .A(n8675), .B(n8674), .ZN(n8678) );
  AOI222_X1 U10199 ( .A1(n10123), .A2(n8678), .B1(n8677), .B2(n10118), .C1(
        n8676), .C2(n10120), .ZN(n8864) );
  OAI21_X1 U10200 ( .B1(n8680), .B2(n8679), .A(n8864), .ZN(n8681) );
  NAND2_X1 U10201 ( .A1(n8681), .A2(n8779), .ZN(n8684) );
  AOI22_X1 U10202 ( .A1(n8682), .A2(n10133), .B1(n10136), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8683) );
  OAI211_X1 U10203 ( .C1(n8869), .C2(n8770), .A(n8684), .B(n8683), .ZN(
        P2_U3209) );
  NAND2_X1 U10204 ( .A1(n8698), .A2(n8685), .ZN(n8687) );
  NAND2_X1 U10205 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  XNOR2_X1 U10206 ( .A(n8688), .B(n8689), .ZN(n8875) );
  INV_X1 U10207 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8693) );
  XNOR2_X1 U10208 ( .A(n8690), .B(n8689), .ZN(n8691) );
  OAI222_X1 U10209 ( .A1(n8762), .A2(n8717), .B1(n8760), .B2(n8692), .C1(n8757), .C2(n8691), .ZN(n8804) );
  INV_X1 U10210 ( .A(n8804), .ZN(n8870) );
  MUX2_X1 U10211 ( .A(n8693), .B(n8870), .S(n8779), .Z(n8696) );
  AOI22_X1 U10212 ( .A1(n8872), .A2(n10130), .B1(n10133), .B2(n8694), .ZN(
        n8695) );
  OAI211_X1 U10213 ( .C1(n8875), .C2(n8770), .A(n8696), .B(n8695), .ZN(
        P2_U3210) );
  NAND2_X1 U10214 ( .A1(n8698), .A2(n8697), .ZN(n8732) );
  NAND2_X1 U10215 ( .A1(n8732), .A2(n8699), .ZN(n8721) );
  NAND2_X1 U10216 ( .A1(n8721), .A2(n8700), .ZN(n8702) );
  NAND2_X1 U10217 ( .A1(n8702), .A2(n8701), .ZN(n8703) );
  XNOR2_X1 U10218 ( .A(n8703), .B(n8705), .ZN(n8879) );
  XOR2_X1 U10219 ( .A(n8705), .B(n8704), .Z(n8706) );
  OAI222_X1 U10220 ( .A1(n8762), .A2(n8708), .B1(n8760), .B2(n8707), .C1(n8757), .C2(n8706), .ZN(n8808) );
  NAND2_X1 U10221 ( .A1(n8808), .A2(n8779), .ZN(n8714) );
  INV_X1 U10222 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8711) );
  INV_X1 U10223 ( .A(n8709), .ZN(n8710) );
  OAI22_X1 U10224 ( .A1(n8779), .A2(n8711), .B1(n8710), .B2(n8776), .ZN(n8712)
         );
  AOI21_X1 U10225 ( .B1(n8809), .B2(n10130), .A(n8712), .ZN(n8713) );
  OAI211_X1 U10226 ( .C1(n8879), .C2(n8770), .A(n8714), .B(n8713), .ZN(
        P2_U3211) );
  XNOR2_X1 U10227 ( .A(n8715), .B(n8722), .ZN(n8716) );
  OAI222_X1 U10228 ( .A1(n8762), .A2(n8745), .B1(n8760), .B2(n8717), .C1(n8757), .C2(n8716), .ZN(n8880) );
  AOI21_X1 U10229 ( .B1(n10133), .B2(n8718), .A(n8880), .ZN(n8726) );
  AOI22_X1 U10230 ( .A1(n8719), .A2(n10130), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n10136), .ZN(n8725) );
  NAND2_X1 U10231 ( .A1(n8721), .A2(n8720), .ZN(n8723) );
  XNOR2_X1 U10232 ( .A(n8723), .B(n8722), .ZN(n8812) );
  NAND2_X1 U10233 ( .A1(n8812), .A2(n10132), .ZN(n8724) );
  OAI211_X1 U10234 ( .C1(n8726), .C2(n10136), .A(n8725), .B(n8724), .ZN(
        P2_U3212) );
  OAI21_X1 U10235 ( .B1(n4611), .B2(n8731), .A(n8727), .ZN(n8730) );
  AOI222_X1 U10236 ( .A1(n10123), .A2(n8730), .B1(n8729), .B2(n10120), .C1(
        n8728), .C2(n10118), .ZN(n8815) );
  XOR2_X1 U10237 ( .A(n8732), .B(n8731), .Z(n8817) );
  AOI22_X1 U10238 ( .A1(n10136), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n10133), 
        .B2(n8733), .ZN(n8734) );
  OAI21_X1 U10239 ( .B1(n8888), .B2(n8735), .A(n8734), .ZN(n8736) );
  AOI21_X1 U10240 ( .B1(n8817), .B2(n10132), .A(n8736), .ZN(n8737) );
  OAI21_X1 U10241 ( .B1(n8815), .B2(n10136), .A(n8737), .ZN(P2_U3213) );
  XNOR2_X1 U10242 ( .A(n8738), .B(n8739), .ZN(n8896) );
  NAND2_X1 U10243 ( .A1(n8740), .A2(n8739), .ZN(n8741) );
  NAND2_X1 U10244 ( .A1(n8741), .A2(n10123), .ZN(n8742) );
  OR2_X1 U10245 ( .A1(n8743), .A2(n8742), .ZN(n8748) );
  OAI22_X1 U10246 ( .A1(n8745), .A2(n8760), .B1(n8744), .B2(n8762), .ZN(n8746)
         );
  INV_X1 U10247 ( .A(n8746), .ZN(n8747) );
  MUX2_X1 U10248 ( .A(n8890), .B(n8749), .S(n10136), .Z(n8752) );
  AOI22_X1 U10249 ( .A1(n8892), .A2(n10130), .B1(n10133), .B2(n8750), .ZN(
        n8751) );
  OAI211_X1 U10250 ( .C1(n8896), .C2(n8770), .A(n8752), .B(n8751), .ZN(
        P2_U3214) );
  OAI21_X1 U10251 ( .B1(n8754), .B2(n8755), .A(n8753), .ZN(n8824) );
  XOR2_X1 U10252 ( .A(n8756), .B(n8755), .Z(n8758) );
  OAI222_X1 U10253 ( .A1(n8762), .A2(n8761), .B1(n8760), .B2(n8759), .C1(n8758), .C2(n8757), .ZN(n8825) );
  NAND2_X1 U10254 ( .A1(n8825), .A2(n8779), .ZN(n8769) );
  INV_X1 U10255 ( .A(n8763), .ZN(n8764) );
  OAI22_X1 U10256 ( .A1(n8779), .A2(n8765), .B1(n8764), .B2(n8776), .ZN(n8766)
         );
  AOI21_X1 U10257 ( .B1(n8767), .B2(n10130), .A(n8766), .ZN(n8768) );
  OAI211_X1 U10258 ( .C1(n8824), .C2(n8770), .A(n8769), .B(n8768), .ZN(
        P2_U3215) );
  XOR2_X1 U10259 ( .A(n8771), .B(n8781), .Z(n8774) );
  AOI222_X1 U10260 ( .A1(n10123), .A2(n8774), .B1(n8773), .B2(n10118), .C1(
        n8772), .C2(n10120), .ZN(n8833) );
  INV_X1 U10261 ( .A(n8775), .ZN(n8777) );
  OAI22_X1 U10262 ( .A1(n8779), .A2(n8778), .B1(n8777), .B2(n8776), .ZN(n8780)
         );
  AOI21_X1 U10263 ( .B1(n8830), .B2(n10130), .A(n8780), .ZN(n8784) );
  XNOR2_X1 U10264 ( .A(n8782), .B(n8781), .ZN(n8831) );
  NAND2_X1 U10265 ( .A1(n8831), .A2(n10132), .ZN(n8783) );
  OAI211_X1 U10266 ( .C1(n8833), .C2(n10136), .A(n8784), .B(n8783), .ZN(
        P2_U3216) );
  NAND2_X1 U10267 ( .A1(n8834), .A2(n6959), .ZN(n8786) );
  INV_X1 U10268 ( .A(n8835), .ZN(n8785) );
  NAND2_X1 U10269 ( .A1(n8785), .A2(n10213), .ZN(n8787) );
  OAI211_X1 U10270 ( .C1(n10213), .C2(n6880), .A(n8786), .B(n8787), .ZN(
        P2_U3490) );
  INV_X1 U10271 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U10272 ( .A1(n8838), .A2(n6959), .ZN(n8788) );
  OAI211_X1 U10273 ( .C1(n10213), .C2(n8789), .A(n8788), .B(n8787), .ZN(
        P2_U3489) );
  INV_X1 U10274 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8790) );
  MUX2_X1 U10275 ( .A(n8790), .B(n8841), .S(n10213), .Z(n8792) );
  NAND2_X1 U10276 ( .A1(n8843), .A2(n6959), .ZN(n8791) );
  OAI211_X1 U10277 ( .C1(n8846), .C2(n8823), .A(n8792), .B(n8791), .ZN(
        P2_U3487) );
  INV_X1 U10278 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8793) );
  INV_X1 U10279 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8796) );
  AOI21_X1 U10280 ( .B1(n8795), .B2(n10188), .A(n8794), .ZN(n8853) );
  OAI21_X1 U10281 ( .B1(n8856), .B2(n8829), .A(n8797), .ZN(P2_U3485) );
  MUX2_X1 U10282 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8857), .S(n10213), .Z(
        n8800) );
  OAI22_X1 U10283 ( .A1(n8863), .A2(n8823), .B1(n8798), .B2(n8829), .ZN(n8799)
         );
  OR2_X1 U10284 ( .A1(n8800), .A2(n8799), .ZN(P2_U3484) );
  INV_X1 U10285 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8801) );
  MUX2_X1 U10286 ( .A(n8801), .B(n8864), .S(n10213), .Z(n8803) );
  NAND2_X1 U10287 ( .A1(n8866), .A2(n6959), .ZN(n8802) );
  OAI211_X1 U10288 ( .C1(n8823), .C2(n8869), .A(n8803), .B(n8802), .ZN(
        P2_U3483) );
  MUX2_X1 U10289 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8804), .S(n10213), .Z(
        n8807) );
  OAI22_X1 U10290 ( .A1(n8875), .A2(n8823), .B1(n8805), .B2(n8829), .ZN(n8806)
         );
  OR2_X1 U10291 ( .A1(n8807), .A2(n8806), .ZN(P2_U3482) );
  INV_X1 U10292 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8810) );
  AOI21_X1 U10293 ( .B1(n10195), .B2(n8809), .A(n8808), .ZN(n8876) );
  MUX2_X1 U10294 ( .A(n8810), .B(n8876), .S(n10213), .Z(n8811) );
  OAI21_X1 U10295 ( .B1(n8879), .B2(n8823), .A(n8811), .ZN(P2_U3481) );
  MUX2_X1 U10296 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8880), .S(n10213), .Z(
        n8814) );
  INV_X1 U10297 ( .A(n8812), .ZN(n8882) );
  OAI22_X1 U10298 ( .A1(n8882), .A2(n8823), .B1(n8881), .B2(n8829), .ZN(n8813)
         );
  OR2_X1 U10299 ( .A1(n8814), .A2(n8813), .ZN(P2_U3480) );
  INV_X1 U10300 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8818) );
  INV_X1 U10301 ( .A(n8815), .ZN(n8816) );
  AOI21_X1 U10302 ( .B1(n8817), .B2(n10188), .A(n8816), .ZN(n8885) );
  MUX2_X1 U10303 ( .A(n8818), .B(n8885), .S(n10213), .Z(n8819) );
  OAI21_X1 U10304 ( .B1(n8888), .B2(n8829), .A(n8819), .ZN(P2_U3479) );
  MUX2_X1 U10305 ( .A(n8890), .B(n8820), .S(n10211), .Z(n8822) );
  NAND2_X1 U10306 ( .A1(n8892), .A2(n6959), .ZN(n8821) );
  OAI211_X1 U10307 ( .C1(n8896), .C2(n8823), .A(n8822), .B(n8821), .ZN(
        P2_U3478) );
  INV_X1 U10308 ( .A(n8824), .ZN(n8826) );
  AOI21_X1 U10309 ( .B1(n8826), .B2(n10188), .A(n8825), .ZN(n8897) );
  MUX2_X1 U10310 ( .A(n8827), .B(n8897), .S(n10213), .Z(n8828) );
  OAI21_X1 U10311 ( .B1(n8901), .B2(n8829), .A(n8828), .ZN(P2_U3477) );
  AOI22_X1 U10312 ( .A1(n8831), .A2(n10188), .B1(n10195), .B2(n8830), .ZN(
        n8832) );
  NAND2_X1 U10313 ( .A1(n8833), .A2(n8832), .ZN(n8902) );
  MUX2_X1 U10314 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8902), .S(n10213), .Z(
        P2_U3476) );
  INV_X1 U10315 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U10316 ( .A1(n8834), .A2(n8891), .ZN(n8836) );
  OR2_X1 U10317 ( .A1(n8835), .A2(n10198), .ZN(n8839) );
  OAI211_X1 U10318 ( .C1(n8837), .C2(n10196), .A(n8836), .B(n8839), .ZN(
        P2_U3458) );
  NAND2_X1 U10319 ( .A1(n8838), .A2(n8891), .ZN(n8840) );
  OAI211_X1 U10320 ( .C1(n5779), .C2(n10196), .A(n8840), .B(n8839), .ZN(
        P2_U3457) );
  MUX2_X1 U10321 ( .A(n8842), .B(n8841), .S(n10196), .Z(n8845) );
  NAND2_X1 U10322 ( .A1(n8843), .A2(n8891), .ZN(n8844) );
  OAI211_X1 U10323 ( .C1(n8846), .C2(n8895), .A(n8845), .B(n8844), .ZN(
        P2_U3455) );
  MUX2_X1 U10324 ( .A(n8848), .B(n8847), .S(n10196), .Z(n8851) );
  NAND2_X1 U10325 ( .A1(n8849), .A2(n8891), .ZN(n8850) );
  OAI211_X1 U10326 ( .C1(n8852), .C2(n8895), .A(n8851), .B(n8850), .ZN(
        P2_U3454) );
  OAI21_X1 U10327 ( .B1(n8856), .B2(n8900), .A(n8855), .ZN(P2_U3453) );
  INV_X1 U10328 ( .A(n8857), .ZN(n8858) );
  MUX2_X1 U10329 ( .A(n8859), .B(n8858), .S(n10196), .Z(n8862) );
  NAND2_X1 U10330 ( .A1(n8860), .A2(n8891), .ZN(n8861) );
  OAI211_X1 U10331 ( .C1(n8863), .C2(n8895), .A(n8862), .B(n8861), .ZN(
        P2_U3452) );
  MUX2_X1 U10332 ( .A(n8865), .B(n8864), .S(n10196), .Z(n8868) );
  NAND2_X1 U10333 ( .A1(n8866), .A2(n8891), .ZN(n8867) );
  OAI211_X1 U10334 ( .C1(n8869), .C2(n8895), .A(n8868), .B(n8867), .ZN(
        P2_U3451) );
  MUX2_X1 U10335 ( .A(n8871), .B(n8870), .S(n10196), .Z(n8874) );
  NAND2_X1 U10336 ( .A1(n8872), .A2(n8891), .ZN(n8873) );
  OAI211_X1 U10337 ( .C1(n8875), .C2(n8895), .A(n8874), .B(n8873), .ZN(
        P2_U3450) );
  MUX2_X1 U10338 ( .A(n8877), .B(n8876), .S(n10196), .Z(n8878) );
  OAI21_X1 U10339 ( .B1(n8879), .B2(n8895), .A(n8878), .ZN(P2_U3449) );
  MUX2_X1 U10340 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8880), .S(n10196), .Z(
        n8884) );
  OAI22_X1 U10341 ( .A1(n8882), .A2(n8895), .B1(n8881), .B2(n8900), .ZN(n8883)
         );
  OR2_X1 U10342 ( .A1(n8884), .A2(n8883), .ZN(P2_U3448) );
  INV_X1 U10343 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8886) );
  MUX2_X1 U10344 ( .A(n8886), .B(n8885), .S(n10196), .Z(n8887) );
  OAI21_X1 U10345 ( .B1(n8888), .B2(n8900), .A(n8887), .ZN(P2_U3447) );
  INV_X1 U10346 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8889) );
  MUX2_X1 U10347 ( .A(n8890), .B(n8889), .S(n10198), .Z(n8894) );
  NAND2_X1 U10348 ( .A1(n8892), .A2(n8891), .ZN(n8893) );
  OAI211_X1 U10349 ( .C1(n8896), .C2(n8895), .A(n8894), .B(n8893), .ZN(
        P2_U3446) );
  MUX2_X1 U10350 ( .A(n8898), .B(n8897), .S(n10196), .Z(n8899) );
  OAI21_X1 U10351 ( .B1(n8901), .B2(n8900), .A(n8899), .ZN(P2_U3444) );
  MUX2_X1 U10352 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8902), .S(n10196), .Z(
        P2_U3441) );
  INV_X1 U10353 ( .A(n9053), .ZN(n9911) );
  NAND3_X1 U10354 ( .A1(n8903), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8904) );
  OAI22_X1 U10355 ( .A1(n8905), .A2(n8904), .B1(n6872), .B2(n4517), .ZN(n8906)
         );
  INV_X1 U10356 ( .A(n8906), .ZN(n8907) );
  OAI21_X1 U10357 ( .B1(n9911), .B2(n8908), .A(n8907), .ZN(P2_U3264) );
  NAND2_X1 U10358 ( .A1(n8911), .A2(n8910), .ZN(n8913) );
  XNOR2_X1 U10359 ( .A(n8913), .B(n8912), .ZN(n8920) );
  AND2_X1 U10360 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9459) );
  OAI22_X1 U10361 ( .A1(n8915), .A2(n9028), .B1(n9029), .B2(n8914), .ZN(n8916)
         );
  AOI211_X1 U10362 ( .C1(n9033), .C2(n8917), .A(n9459), .B(n8916), .ZN(n8919)
         );
  NAND2_X1 U10363 ( .A1(n9111), .A2(n9051), .ZN(n8918) );
  OAI211_X1 U10364 ( .C1(n8920), .C2(n9046), .A(n8919), .B(n8918), .ZN(
        P1_U3215) );
  INV_X1 U10365 ( .A(n9656), .ZN(n9888) );
  INV_X1 U10366 ( .A(n8921), .ZN(n8925) );
  AOI21_X1 U10367 ( .B1(n8922), .B2(n9002), .A(n8923), .ZN(n8924) );
  OAI21_X1 U10368 ( .B1(n8925), .B2(n8924), .A(n9025), .ZN(n8930) );
  INV_X1 U10369 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8926) );
  NOR2_X1 U10370 ( .A1(n8926), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8928) );
  OAI22_X1 U10371 ( .A1(n9651), .A2(n9028), .B1(n9029), .B2(n9682), .ZN(n8927)
         );
  AOI211_X1 U10372 ( .C1(n9033), .C2(n9648), .A(n8928), .B(n8927), .ZN(n8929)
         );
  OAI211_X1 U10373 ( .C1(n9888), .C2(n9036), .A(n8930), .B(n8929), .ZN(
        P1_U3216) );
  XNOR2_X1 U10374 ( .A(n8932), .B(n8931), .ZN(n8937) );
  AND2_X1 U10375 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9556) );
  OAI22_X1 U10376 ( .A1(n8933), .A2(n9029), .B1(n8944), .B2(n9028), .ZN(n8934)
         );
  AOI211_X1 U10377 ( .C1(n9033), .C2(n9716), .A(n9556), .B(n8934), .ZN(n8936)
         );
  NAND2_X1 U10378 ( .A1(n9843), .A2(n9051), .ZN(n8935) );
  OAI211_X1 U10379 ( .C1(n8937), .C2(n9046), .A(n8936), .B(n8935), .ZN(
        P1_U3219) );
  XNOR2_X1 U10380 ( .A(n8939), .B(n8938), .ZN(n8940) );
  XNOR2_X1 U10381 ( .A(n8941), .B(n8940), .ZN(n8948) );
  INV_X1 U10382 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8942) );
  OAI22_X1 U10383 ( .A1(n9041), .A2(n8943), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8942), .ZN(n8946) );
  OAI22_X1 U10384 ( .A1(n8944), .A2(n9029), .B1(n9028), .B2(n9682), .ZN(n8945)
         );
  AOI211_X1 U10385 ( .C1(n9688), .C2(n9051), .A(n8946), .B(n8945), .ZN(n8947)
         );
  OAI21_X1 U10386 ( .B1(n8948), .B2(n9046), .A(n8947), .ZN(P1_U3223) );
  AOI21_X1 U10387 ( .B1(n8950), .B2(n8949), .A(n9023), .ZN(n8956) );
  INV_X1 U10388 ( .A(n9624), .ZN(n8952) );
  OAI22_X1 U10389 ( .A1(n9041), .A2(n8952), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8951), .ZN(n8954) );
  OAI22_X1 U10390 ( .A1(n9651), .A2(n9029), .B1(n9028), .B2(n9195), .ZN(n8953)
         );
  AOI211_X1 U10391 ( .C1(n9878), .C2(n9051), .A(n8954), .B(n8953), .ZN(n8955)
         );
  OAI21_X1 U10392 ( .B1(n8956), .B2(n9046), .A(n8955), .ZN(P1_U3225) );
  NOR2_X1 U10393 ( .A1(n8958), .A2(n5079), .ZN(n8959) );
  XNOR2_X1 U10394 ( .A(n8960), .B(n8959), .ZN(n8966) );
  AOI22_X1 U10395 ( .A1(n9037), .A2(n9918), .B1(n9038), .B2(n10065), .ZN(n8961) );
  NAND2_X1 U10396 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9502) );
  OAI211_X1 U10397 ( .C1(n9041), .C2(n8962), .A(n8961), .B(n9502), .ZN(n8963)
         );
  AOI21_X1 U10398 ( .B1(n8964), .B2(n9051), .A(n8963), .ZN(n8965) );
  OAI21_X1 U10399 ( .B1(n8966), .B2(n9046), .A(n8965), .ZN(P1_U3226) );
  XNOR2_X1 U10400 ( .A(n8968), .B(n8967), .ZN(n8969) );
  XNOR2_X1 U10401 ( .A(n8970), .B(n8969), .ZN(n8980) );
  NOR3_X1 U10402 ( .A1(n9041), .A2(P1_REG3_REG_17__SCAN_IN), .A3(n8971), .ZN(
        n8976) );
  AOI21_X1 U10403 ( .B1(n8972), .B2(n8971), .A(P1_U3086), .ZN(n8974) );
  OAI22_X1 U10404 ( .A1(n8974), .A2(n6275), .B1(n8973), .B2(n9029), .ZN(n8975)
         );
  AOI211_X1 U10405 ( .C1(n9037), .C2(n9711), .A(n8976), .B(n8975), .ZN(n8979)
         );
  NAND2_X1 U10406 ( .A1(n8977), .A2(n9051), .ZN(n8978) );
  OAI211_X1 U10407 ( .C1(n8980), .C2(n9046), .A(n8979), .B(n8978), .ZN(
        P1_U3228) );
  AOI22_X1 U10408 ( .A1(n9033), .A2(n9637), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8986) );
  AOI22_X1 U10409 ( .A1(n9038), .A2(n9816), .B1(n9037), .B2(n9784), .ZN(n8985)
         );
  NAND2_X1 U10410 ( .A1(n9636), .A2(n9051), .ZN(n8984) );
  NAND4_X1 U10411 ( .A1(n8987), .A2(n8986), .A3(n8985), .A4(n8984), .ZN(
        P1_U3229) );
  NOR2_X1 U10412 ( .A1(n8989), .A2(n4755), .ZN(n8990) );
  XNOR2_X1 U10413 ( .A(n8991), .B(n8990), .ZN(n8997) );
  INV_X1 U10414 ( .A(n9699), .ZN(n8993) );
  INV_X1 U10415 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8992) );
  OAI22_X1 U10416 ( .A1(n9041), .A2(n8993), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8992), .ZN(n8995) );
  OAI22_X1 U10417 ( .A1(n9737), .A2(n9029), .B1(n9028), .B2(n9184), .ZN(n8994)
         );
  AOI211_X1 U10418 ( .C1(n9698), .C2(n9051), .A(n8995), .B(n8994), .ZN(n8996)
         );
  OAI21_X1 U10419 ( .B1(n8997), .B2(n9046), .A(n8996), .ZN(P1_U3233) );
  XNOR2_X1 U10420 ( .A(n8999), .B(n8998), .ZN(n9001) );
  INV_X1 U10421 ( .A(n9003), .ZN(n9000) );
  NAND2_X1 U10422 ( .A1(n9001), .A2(n9000), .ZN(n9005) );
  INV_X1 U10423 ( .A(n9002), .ZN(n9004) );
  AOI22_X1 U10424 ( .A1(n9005), .A2(n8922), .B1(n9004), .B2(n9003), .ZN(n9011)
         );
  INV_X1 U10425 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9006) );
  OAI22_X1 U10426 ( .A1(n9041), .A2(n9007), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9006), .ZN(n9009) );
  OAI22_X1 U10427 ( .A1(n9184), .A2(n9029), .B1(n9028), .B2(n9666), .ZN(n9008)
         );
  AOI211_X1 U10428 ( .C1(n9670), .C2(n9051), .A(n9009), .B(n9008), .ZN(n9010)
         );
  OAI21_X1 U10429 ( .B1(n9011), .B2(n9046), .A(n9010), .ZN(P1_U3235) );
  XNOR2_X1 U10430 ( .A(n9013), .B(n9012), .ZN(n9014) );
  XNOR2_X1 U10431 ( .A(n9015), .B(n9014), .ZN(n9016) );
  NAND2_X1 U10432 ( .A1(n9016), .A2(n9025), .ZN(n9020) );
  AND2_X1 U10433 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9531) );
  OAI22_X1 U10434 ( .A1(n9017), .A2(n9029), .B1(n9737), .B2(n9028), .ZN(n9018)
         );
  AOI211_X1 U10435 ( .C1(n9033), .C2(n9733), .A(n9531), .B(n9018), .ZN(n9019)
         );
  OAI211_X1 U10436 ( .C1(n9905), .C2(n9036), .A(n9020), .B(n9019), .ZN(
        P1_U3238) );
  INV_X1 U10437 ( .A(n9613), .ZN(n9875) );
  OAI21_X1 U10438 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(n9024) );
  NAND3_X1 U10439 ( .A1(n9026), .A2(n9025), .A3(n9024), .ZN(n9035) );
  NOR2_X1 U10440 ( .A1(n9027), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9032) );
  OAI22_X1 U10441 ( .A1(n9030), .A2(n9029), .B1(n9028), .B2(n9608), .ZN(n9031)
         );
  AOI211_X1 U10442 ( .C1(n9033), .C2(n9605), .A(n9032), .B(n9031), .ZN(n9034)
         );
  OAI211_X1 U10443 ( .C1(n9875), .C2(n9036), .A(n9035), .B(n9034), .ZN(
        P1_U3240) );
  AOI22_X1 U10444 ( .A1(n9038), .A2(n9346), .B1(n9037), .B2(n9345), .ZN(n9039)
         );
  NAND2_X1 U10445 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9477) );
  OAI211_X1 U10446 ( .C1(n9041), .C2(n9040), .A(n9039), .B(n9477), .ZN(n9050)
         );
  INV_X1 U10447 ( .A(n9042), .ZN(n9048) );
  AOI21_X1 U10448 ( .B1(n9047), .B2(n9044), .A(n9043), .ZN(n9045) );
  AOI211_X1 U10449 ( .C1(n9048), .C2(n9047), .A(n9046), .B(n9045), .ZN(n9049)
         );
  AOI211_X1 U10450 ( .C1(n9927), .C2(n9051), .A(n9050), .B(n9049), .ZN(n9052)
         );
  INV_X1 U10451 ( .A(n9052), .ZN(P1_U3241) );
  NAND2_X1 U10452 ( .A1(n9053), .A2(n9058), .ZN(n9055) );
  OR2_X1 U10453 ( .A1(n9060), .A2(n10455), .ZN(n9054) );
  INV_X1 U10454 ( .A(n9860), .ZN(n9056) );
  INV_X1 U10455 ( .A(n9057), .ZN(n9559) );
  AND2_X1 U10456 ( .A1(n9860), .A2(n9057), .ZN(n9098) );
  INV_X1 U10457 ( .A(n9098), .ZN(n9339) );
  NAND2_X1 U10458 ( .A1(n9059), .A2(n9058), .ZN(n9062) );
  OR2_X1 U10459 ( .A1(n9060), .A2(n10402), .ZN(n9061) );
  OR2_X1 U10460 ( .A1(n9564), .A2(n9099), .ZN(n9321) );
  NAND2_X1 U10461 ( .A1(n9564), .A2(n9099), .ZN(n9292) );
  INV_X1 U10462 ( .A(n9064), .ZN(n9067) );
  NAND4_X1 U10463 ( .A1(n9755), .A2(n9067), .A3(n9066), .A4(n9065), .ZN(n9070)
         );
  NOR3_X1 U10464 ( .A1(n9070), .A2(n9069), .A3(n9068), .ZN(n9071) );
  AND4_X1 U10465 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(n9075)
         );
  NAND3_X1 U10466 ( .A1(n9077), .A2(n9076), .A3(n9075), .ZN(n9078) );
  NOR2_X1 U10467 ( .A1(n9079), .A2(n9078), .ZN(n9080) );
  NAND3_X1 U10468 ( .A1(n9081), .A2(n5059), .A3(n9080), .ZN(n9082) );
  NOR2_X1 U10469 ( .A1(n9083), .A2(n9082), .ZN(n9084) );
  NAND4_X1 U10470 ( .A1(n9085), .A2(n4552), .A3(n9084), .A4(n9161), .ZN(n9086)
         );
  OR3_X1 U10471 ( .A1(n9729), .A2(n9087), .A3(n9086), .ZN(n9088) );
  NOR2_X1 U10472 ( .A1(n9707), .A2(n9088), .ZN(n9089) );
  AND2_X1 U10473 ( .A1(n9695), .A2(n9089), .ZN(n9090) );
  NAND4_X1 U10474 ( .A1(n9646), .A2(n9090), .A3(n9661), .A4(n9677), .ZN(n9091)
         );
  NOR2_X1 U10475 ( .A1(n9640), .A2(n9091), .ZN(n9093) );
  INV_X1 U10476 ( .A(n9614), .ZN(n9092) );
  AND4_X1 U10477 ( .A1(n9589), .A2(n9628), .A3(n9093), .A4(n9092), .ZN(n9094)
         );
  AND2_X1 U10478 ( .A1(n9576), .A2(n9094), .ZN(n9095) );
  AND4_X1 U10479 ( .A1(n9321), .A2(n9096), .A3(n9292), .A4(n9095), .ZN(n9097)
         );
  NAND2_X1 U10480 ( .A1(n9339), .A2(n9097), .ZN(n9325) );
  NOR2_X1 U10481 ( .A1(n9099), .A2(n9559), .ZN(n9213) );
  NOR2_X1 U10482 ( .A1(n9098), .A2(n9213), .ZN(n9101) );
  NOR2_X1 U10483 ( .A1(n9860), .A2(n9099), .ZN(n9100) );
  MUX2_X1 U10484 ( .A(n9101), .B(n9100), .S(n9564), .Z(n9218) );
  OR2_X1 U10485 ( .A1(n9670), .A2(n9682), .ZN(n9102) );
  NAND2_X1 U10486 ( .A1(n9190), .A2(n9102), .ZN(n9225) );
  NAND2_X1 U10487 ( .A1(n9224), .A2(n9103), .ZN(n9231) );
  MUX2_X1 U10488 ( .A(n9225), .B(n9231), .S(n9215), .Z(n9192) );
  INV_X1 U10489 ( .A(n9276), .ZN(n9104) );
  NAND2_X1 U10490 ( .A1(n9280), .A2(n9104), .ZN(n9105) );
  NAND2_X1 U10491 ( .A1(n9105), .A2(n9277), .ZN(n9109) );
  INV_X1 U10492 ( .A(n9164), .ZN(n9106) );
  NAND2_X1 U10493 ( .A1(n9277), .A2(n9106), .ZN(n9107) );
  NAND2_X1 U10494 ( .A1(n9107), .A2(n9280), .ZN(n9108) );
  MUX2_X1 U10495 ( .A(n9109), .B(n9108), .S(n9215), .Z(n9168) );
  OR2_X1 U10496 ( .A1(n9111), .A2(n9110), .ZN(n9275) );
  AND2_X1 U10497 ( .A1(n9275), .A2(n9215), .ZN(n9112) );
  AND2_X1 U10498 ( .A1(n9276), .A2(n9112), .ZN(n9162) );
  INV_X1 U10499 ( .A(n9255), .ZN(n9115) );
  OAI211_X1 U10500 ( .C1(n9116), .C2(n9115), .A(n9114), .B(n9113), .ZN(n9117)
         );
  MUX2_X1 U10501 ( .A(n9118), .B(n9117), .S(n9215), .Z(n9137) );
  INV_X1 U10502 ( .A(n9136), .ZN(n9120) );
  AND2_X1 U10503 ( .A1(n9119), .A2(n9258), .ZN(n9138) );
  OAI21_X1 U10504 ( .B1(n9137), .B2(n9120), .A(n9138), .ZN(n9121) );
  NAND2_X1 U10505 ( .A1(n9121), .A2(n9261), .ZN(n9123) );
  INV_X1 U10506 ( .A(n9215), .ZN(n9207) );
  NAND4_X1 U10507 ( .A1(n9123), .A2(n9207), .A3(n9124), .A4(n9122), .ZN(n9147)
         );
  OR2_X1 U10508 ( .A1(n9140), .A2(n9207), .ZN(n9127) );
  INV_X1 U10509 ( .A(n9124), .ZN(n9125) );
  NAND2_X1 U10510 ( .A1(n9125), .A2(n9207), .ZN(n9126) );
  NAND4_X1 U10511 ( .A1(n9129), .A2(n9128), .A3(n9127), .A4(n9126), .ZN(n9134)
         );
  AND2_X1 U10512 ( .A1(n9215), .A2(n9351), .ZN(n9132) );
  OAI21_X1 U10513 ( .B1(n9351), .B2(n9215), .A(n9131), .ZN(n9130) );
  OAI21_X1 U10514 ( .B1(n9132), .B2(n9131), .A(n9130), .ZN(n9133) );
  AND3_X1 U10515 ( .A1(n9134), .A2(n9148), .A3(n9133), .ZN(n9146) );
  AND2_X1 U10516 ( .A1(n9136), .A2(n9135), .ZN(n9257) );
  NAND2_X1 U10517 ( .A1(n9137), .A2(n9257), .ZN(n9139) );
  NAND2_X1 U10518 ( .A1(n9139), .A2(n9138), .ZN(n9144) );
  AND4_X1 U10519 ( .A1(n9141), .A2(n9215), .A3(n9140), .A4(n9261), .ZN(n9143)
         );
  INV_X1 U10520 ( .A(n9151), .ZN(n9142) );
  AOI21_X1 U10521 ( .B1(n9144), .B2(n9143), .A(n9142), .ZN(n9145) );
  NAND3_X1 U10522 ( .A1(n9147), .A2(n9146), .A3(n9145), .ZN(n9152) );
  NAND2_X1 U10523 ( .A1(n9152), .A2(n9148), .ZN(n9149) );
  NAND2_X1 U10524 ( .A1(n9155), .A2(n9153), .ZN(n9246) );
  AOI21_X1 U10525 ( .B1(n9149), .B2(n9263), .A(n9246), .ZN(n9150) );
  NAND2_X1 U10526 ( .A1(n9156), .A2(n9154), .ZN(n9271) );
  OAI21_X1 U10527 ( .B1(n9150), .B2(n9271), .A(n9269), .ZN(n9159) );
  NAND2_X1 U10528 ( .A1(n9157), .A2(n9156), .ZN(n9158) );
  MUX2_X1 U10529 ( .A(n9159), .B(n9158), .S(n9207), .Z(n9160) );
  INV_X1 U10530 ( .A(n9162), .ZN(n9165) );
  NAND2_X1 U10531 ( .A1(n9164), .A2(n9163), .ZN(n9278) );
  OAI21_X1 U10532 ( .B1(n9168), .B2(n9167), .A(n9166), .ZN(n9176) );
  NAND3_X1 U10533 ( .A1(n9176), .A2(n9170), .A3(n9724), .ZN(n9169) );
  AND3_X1 U10534 ( .A1(n9169), .A2(n9173), .A3(n9172), .ZN(n9179) );
  AND2_X1 U10535 ( .A1(n9180), .A2(n9170), .ZN(n9283) );
  INV_X1 U10536 ( .A(n9283), .ZN(n9177) );
  NAND2_X1 U10537 ( .A1(n9172), .A2(n9171), .ZN(n9175) );
  INV_X1 U10538 ( .A(n9173), .ZN(n9174) );
  AOI21_X1 U10539 ( .B1(n9283), .B2(n9175), .A(n9174), .ZN(n9285) );
  OAI211_X1 U10540 ( .C1(n9177), .C2(n9176), .A(n9285), .B(n9183), .ZN(n9178)
         );
  MUX2_X1 U10541 ( .A(n9179), .B(n9178), .S(n9215), .Z(n9182) );
  AOI21_X1 U10542 ( .B1(n9185), .B2(n9180), .A(n9215), .ZN(n9181) );
  NOR2_X1 U10543 ( .A1(n9182), .A2(n9181), .ZN(n9189) );
  NAND2_X1 U10544 ( .A1(n9186), .A2(n9183), .ZN(n9230) );
  OR2_X1 U10545 ( .A1(n9688), .A2(n9184), .ZN(n9229) );
  NAND2_X1 U10546 ( .A1(n9229), .A2(n9185), .ZN(n9242) );
  MUX2_X1 U10547 ( .A(n9230), .B(n9242), .S(n9215), .Z(n9188) );
  MUX2_X1 U10548 ( .A(n9186), .B(n9229), .S(n9207), .Z(n9187) );
  MUX2_X1 U10549 ( .A(n9224), .B(n9190), .S(n9215), .Z(n9191) );
  MUX2_X1 U10550 ( .A(n9233), .B(n9227), .S(n9207), .Z(n9193) );
  INV_X1 U10551 ( .A(n9245), .ZN(n9194) );
  OAI211_X1 U10552 ( .C1(n9198), .C2(n9194), .A(n9308), .B(n9237), .ZN(n9196)
         );
  NOR2_X1 U10553 ( .A1(n9613), .A2(n9195), .ZN(n9199) );
  INV_X1 U10554 ( .A(n9199), .ZN(n9222) );
  NAND2_X1 U10555 ( .A1(n9196), .A2(n9222), .ZN(n9202) );
  INV_X1 U10556 ( .A(n9237), .ZN(n9197) );
  AOI21_X1 U10557 ( .B1(n9198), .B2(n9245), .A(n9197), .ZN(n9200) );
  OAI21_X1 U10558 ( .B1(n9200), .B2(n9199), .A(n9308), .ZN(n9201) );
  MUX2_X1 U10559 ( .A(n9202), .B(n9201), .S(n9215), .Z(n9204) );
  INV_X1 U10560 ( .A(n9223), .ZN(n9203) );
  NOR2_X1 U10561 ( .A1(n9204), .A2(n9203), .ZN(n9208) );
  NAND2_X1 U10562 ( .A1(n9206), .A2(n9205), .ZN(n9241) );
  MUX2_X1 U10563 ( .A(n9208), .B(n9207), .S(n9241), .Z(n9210) );
  OAI21_X1 U10564 ( .B1(n9241), .B2(n9223), .A(n9290), .ZN(n9209) );
  MUX2_X1 U10565 ( .A(n9316), .B(n9291), .S(n9215), .Z(n9211) );
  INV_X1 U10566 ( .A(n9213), .ZN(n9214) );
  AND2_X1 U10567 ( .A1(n9564), .A2(n9214), .ZN(n9315) );
  NOR2_X1 U10568 ( .A1(n9860), .A2(n9321), .ZN(n9216) );
  MUX2_X1 U10569 ( .A(n9315), .B(n9216), .S(n9215), .Z(n9217) );
  OAI21_X1 U10570 ( .B1(n9331), .B2(n9299), .A(n9249), .ZN(n9221) );
  NOR3_X1 U10571 ( .A1(n9336), .A2(n9340), .A3(n9219), .ZN(n9220) );
  OAI211_X1 U10572 ( .C1(n9296), .C2(n9325), .A(n9221), .B(n9220), .ZN(n9344)
         );
  NAND2_X1 U10573 ( .A1(n9223), .A2(n9222), .ZN(n9312) );
  NAND2_X1 U10574 ( .A1(n9225), .A2(n9224), .ZN(n9226) );
  NAND2_X1 U10575 ( .A1(n9227), .A2(n9226), .ZN(n9228) );
  NAND2_X1 U10576 ( .A1(n9228), .A2(n9233), .ZN(n9244) );
  INV_X1 U10577 ( .A(n9229), .ZN(n9235) );
  INV_X1 U10578 ( .A(n9230), .ZN(n9234) );
  INV_X1 U10579 ( .A(n9231), .ZN(n9232) );
  OAI211_X1 U10580 ( .C1(n9235), .C2(n9234), .A(n9233), .B(n9232), .ZN(n9236)
         );
  NAND3_X1 U10581 ( .A1(n9245), .A2(n9244), .A3(n9236), .ZN(n9238) );
  AND2_X1 U10582 ( .A1(n9238), .A2(n9237), .ZN(n9239) );
  NOR2_X1 U10583 ( .A1(n9312), .A2(n9239), .ZN(n9240) );
  OR2_X1 U10584 ( .A1(n9241), .A2(n9240), .ZN(n9314) );
  INV_X1 U10585 ( .A(n9242), .ZN(n9243) );
  NAND3_X1 U10586 ( .A1(n9245), .A2(n9244), .A3(n9243), .ZN(n9309) );
  INV_X1 U10587 ( .A(n9246), .ZN(n9268) );
  INV_X1 U10588 ( .A(n9247), .ZN(n9250) );
  NAND2_X1 U10589 ( .A1(n10001), .A2(n9750), .ZN(n9248) );
  AND3_X1 U10590 ( .A1(n9250), .A2(n9249), .A3(n9248), .ZN(n9252) );
  OAI21_X1 U10591 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(n9256) );
  AOI21_X1 U10592 ( .B1(n9256), .B2(n9255), .A(n9254), .ZN(n9260) );
  INV_X1 U10593 ( .A(n9257), .ZN(n9259) );
  OAI21_X1 U10594 ( .B1(n9260), .B2(n9259), .A(n9258), .ZN(n9262) );
  NAND2_X1 U10595 ( .A1(n9262), .A2(n9261), .ZN(n9265) );
  OAI211_X1 U10596 ( .C1(n9266), .C2(n9265), .A(n9264), .B(n9263), .ZN(n9267)
         );
  AND2_X1 U10597 ( .A1(n9268), .A2(n9267), .ZN(n9272) );
  OAI211_X1 U10598 ( .C1(n9272), .C2(n9271), .A(n9270), .B(n9269), .ZN(n9273)
         );
  AND3_X1 U10599 ( .A1(n9275), .A2(n9274), .A3(n9273), .ZN(n9279) );
  OAI211_X1 U10600 ( .C1(n9279), .C2(n9278), .A(n9277), .B(n9276), .ZN(n9281)
         );
  NAND2_X1 U10601 ( .A1(n9281), .A2(n9280), .ZN(n9282) );
  NAND3_X1 U10602 ( .A1(n9283), .A2(n9724), .A3(n9282), .ZN(n9284) );
  AND2_X1 U10603 ( .A1(n9285), .A2(n9284), .ZN(n9286) );
  OAI21_X1 U10604 ( .B1(n9309), .B2(n9286), .A(n9308), .ZN(n9287) );
  INV_X1 U10605 ( .A(n9287), .ZN(n9288) );
  NOR2_X1 U10606 ( .A1(n9312), .A2(n9288), .ZN(n9289) );
  NOR2_X1 U10607 ( .A1(n9314), .A2(n9289), .ZN(n9293) );
  NAND2_X1 U10608 ( .A1(n9291), .A2(n9290), .ZN(n9318) );
  OAI211_X1 U10609 ( .C1(n9293), .C2(n9318), .A(n9292), .B(n9316), .ZN(n9294)
         );
  NAND2_X1 U10610 ( .A1(n9294), .A2(n9321), .ZN(n9295) );
  NAND2_X1 U10611 ( .A1(n9339), .A2(n9295), .ZN(n9297) );
  INV_X1 U10612 ( .A(n9296), .ZN(n9333) );
  AND2_X1 U10613 ( .A1(n9297), .A2(n9333), .ZN(n9328) );
  INV_X1 U10614 ( .A(n9328), .ZN(n9305) );
  NOR3_X1 U10615 ( .A1(n9336), .A2(n9340), .A3(n9306), .ZN(n9304) );
  INV_X1 U10616 ( .A(n9336), .ZN(n9307) );
  AOI21_X1 U10617 ( .B1(n9307), .B2(n9299), .A(n9298), .ZN(n9303) );
  INV_X1 U10618 ( .A(n9300), .ZN(n9941) );
  NAND4_X1 U10619 ( .A1(n9301), .A2(n9941), .A3(n9995), .A4(n10063), .ZN(n9302) );
  AOI22_X1 U10620 ( .A1(n9305), .A2(n9304), .B1(n9303), .B2(n9302), .ZN(n9343)
         );
  AND4_X1 U10621 ( .A1(n9333), .A2(n9307), .A3(n9306), .A4(n9340), .ZN(n9330)
         );
  OAI21_X1 U10622 ( .B1(n9309), .B2(n9692), .A(n9308), .ZN(n9310) );
  INV_X1 U10623 ( .A(n9310), .ZN(n9311) );
  NOR2_X1 U10624 ( .A1(n9312), .A2(n9311), .ZN(n9313) );
  NOR2_X1 U10625 ( .A1(n9314), .A2(n9313), .ZN(n9319) );
  INV_X1 U10626 ( .A(n9315), .ZN(n9317) );
  OAI211_X1 U10627 ( .C1(n9319), .C2(n9318), .A(n9317), .B(n9316), .ZN(n9320)
         );
  OAI21_X1 U10628 ( .B1(n9321), .B2(n9559), .A(n9320), .ZN(n9322) );
  NAND2_X1 U10629 ( .A1(n9322), .A2(n9339), .ZN(n9324) );
  NAND2_X1 U10630 ( .A1(n9324), .A2(n9323), .ZN(n9326) );
  NAND2_X1 U10631 ( .A1(n9326), .A2(n9325), .ZN(n9329) );
  NOR2_X1 U10632 ( .A1(n6465), .A2(n9336), .ZN(n9327) );
  AOI22_X1 U10633 ( .A1(n9330), .A2(n9329), .B1(n9328), .B2(n9327), .ZN(n9342)
         );
  OAI21_X1 U10634 ( .B1(n9333), .B2(n9340), .A(n9332), .ZN(n9338) );
  NOR3_X1 U10635 ( .A1(n9336), .A2(n9335), .A3(n9334), .ZN(n9337) );
  OAI211_X1 U10636 ( .C1(n9340), .C2(n9339), .A(n9338), .B(n9337), .ZN(n9341)
         );
  NAND4_X1 U10637 ( .A1(n9344), .A2(n9343), .A3(n9342), .A4(n9341), .ZN(
        P1_U3242) );
  MUX2_X1 U10638 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9573), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10639 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9776), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10640 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9783), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10641 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9775), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10642 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9784), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10643 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9806), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10644 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9827), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10645 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9817), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10646 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9828), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10647 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9846), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10648 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9711), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10649 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9918), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10650 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9345), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10651 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10065), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10652 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9346), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10653 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n10062), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10654 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9347), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10655 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9348), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10656 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9349), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10657 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9350), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10658 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9351), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10659 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9352), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10660 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n10029), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10661 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9353), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10662 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9354), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10663 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9355), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10664 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9997), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10665 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9998), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10666 ( .C1(n9356), .C2(n9380), .A(n9528), .B(n9948), .ZN(n9364)
         );
  OAI211_X1 U10667 ( .C1(n9359), .C2(n9358), .A(n9551), .B(n9357), .ZN(n9363)
         );
  AOI22_X1 U10668 ( .A1(n9946), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9362) );
  NAND2_X1 U10669 ( .A1(n9958), .A2(n9360), .ZN(n9361) );
  NAND4_X1 U10670 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(
        P1_U3244) );
  NOR2_X1 U10671 ( .A1(n9457), .A2(n9365), .ZN(n9366) );
  AOI211_X1 U10672 ( .C1(n9946), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9367), .B(
        n9366), .ZN(n9377) );
  OAI211_X1 U10673 ( .C1(n9370), .C2(n9369), .A(n9528), .B(n9368), .ZN(n9376)
         );
  INV_X1 U10674 ( .A(n9396), .ZN(n9374) );
  NAND3_X1 U10675 ( .A1(n9953), .A2(n9372), .A3(n9371), .ZN(n9373) );
  NAND3_X1 U10676 ( .A1(n9551), .A2(n9374), .A3(n9373), .ZN(n9375) );
  NAND3_X1 U10677 ( .A1(n9377), .A2(n9376), .A3(n9375), .ZN(P1_U3246) );
  INV_X1 U10678 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9379) );
  AOI21_X1 U10679 ( .B1(n9941), .B2(n9379), .A(n9378), .ZN(n9940) );
  MUX2_X1 U10680 ( .A(n9381), .B(n9380), .S(n9941), .Z(n9383) );
  NAND2_X1 U10681 ( .A1(n9383), .A2(n9382), .ZN(n9384) );
  OAI211_X1 U10682 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9940), .A(n9384), .B(
        P1_U3973), .ZN(n9964) );
  NOR2_X1 U10683 ( .A1(n9457), .A2(n9385), .ZN(n9386) );
  AOI211_X1 U10684 ( .C1(n9946), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9387), .B(
        n9386), .ZN(n9399) );
  OAI211_X1 U10685 ( .C1(n9390), .C2(n9389), .A(n9528), .B(n9388), .ZN(n9398)
         );
  MUX2_X1 U10686 ( .A(n7031), .B(P1_REG1_REG_4__SCAN_IN), .S(n9391), .Z(n9394)
         );
  INV_X1 U10687 ( .A(n9392), .ZN(n9393) );
  NAND2_X1 U10688 ( .A1(n9394), .A2(n9393), .ZN(n9395) );
  OAI211_X1 U10689 ( .C1(n9396), .C2(n9395), .A(n9551), .B(n9404), .ZN(n9397)
         );
  NAND4_X1 U10690 ( .A1(n9964), .A2(n9399), .A3(n9398), .A4(n9397), .ZN(
        P1_U3247) );
  OAI211_X1 U10691 ( .C1(n9401), .C2(n9400), .A(n9528), .B(n4770), .ZN(n9412)
         );
  NAND3_X1 U10692 ( .A1(n9404), .A2(n9403), .A3(n9402), .ZN(n9405) );
  NAND3_X1 U10693 ( .A1(n9551), .A2(n9406), .A3(n9405), .ZN(n9411) );
  AOI21_X1 U10694 ( .B1(n9946), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9407), .ZN(
        n9410) );
  NAND2_X1 U10695 ( .A1(n9958), .A2(n9408), .ZN(n9409) );
  NAND4_X1 U10696 ( .A1(n9412), .A2(n9411), .A3(n9410), .A4(n9409), .ZN(
        P1_U3248) );
  OAI21_X1 U10697 ( .B1(n9415), .B2(n9414), .A(n9413), .ZN(n9416) );
  NAND2_X1 U10698 ( .A1(n9416), .A2(n9528), .ZN(n9426) );
  AOI21_X1 U10699 ( .B1(n9946), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9417), .ZN(
        n9425) );
  OAI21_X1 U10700 ( .B1(n9420), .B2(n9419), .A(n9418), .ZN(n9421) );
  NAND2_X1 U10701 ( .A1(n9421), .A2(n9551), .ZN(n9424) );
  NAND2_X1 U10702 ( .A1(n9958), .A2(n9422), .ZN(n9423) );
  NAND4_X1 U10703 ( .A1(n9426), .A2(n9425), .A3(n9424), .A4(n9423), .ZN(
        P1_U3252) );
  OAI211_X1 U10704 ( .C1(n9429), .C2(n9428), .A(n9427), .B(n9551), .ZN(n9440)
         );
  AOI21_X1 U10705 ( .B1(n9946), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n9430), .ZN(
        n9439) );
  INV_X1 U10706 ( .A(n9431), .ZN(n9432) );
  OAI21_X1 U10707 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9435) );
  OR2_X1 U10708 ( .A1(n9962), .A2(n9435), .ZN(n9438) );
  NAND2_X1 U10709 ( .A1(n9958), .A2(n9436), .ZN(n9437) );
  NAND4_X1 U10710 ( .A1(n9440), .A2(n9439), .A3(n9438), .A4(n9437), .ZN(
        P1_U3254) );
  AOI21_X1 U10711 ( .B1(n7311), .B2(n9442), .A(n9441), .ZN(n9445) );
  INV_X1 U10712 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9443) );
  MUX2_X1 U10713 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9443), .S(n9462), .Z(n9444) );
  NAND2_X1 U10714 ( .A1(n9444), .A2(n9445), .ZN(n9467) );
  OAI211_X1 U10715 ( .C1(n9445), .C2(n9444), .A(n9551), .B(n9467), .ZN(n9456)
         );
  AOI21_X1 U10716 ( .B1(n9946), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9446), .ZN(
        n9455) );
  OAI21_X1 U10717 ( .B1(n9448), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9447), .ZN(
        n9451) );
  INV_X1 U10718 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9449) );
  AOI22_X1 U10719 ( .A1(n9462), .A2(n9449), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n9468), .ZN(n9450) );
  NOR2_X1 U10720 ( .A1(n9450), .A2(n9451), .ZN(n9461) );
  AOI21_X1 U10721 ( .B1(n9451), .B2(n9450), .A(n9461), .ZN(n9452) );
  NAND2_X1 U10722 ( .A1(n9528), .A2(n9452), .ZN(n9454) );
  NAND2_X1 U10723 ( .A1(n9958), .A2(n9462), .ZN(n9453) );
  NAND4_X1 U10724 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(n9453), .ZN(
        P1_U3256) );
  NOR2_X1 U10725 ( .A1(n9457), .A2(n9475), .ZN(n9458) );
  AOI211_X1 U10726 ( .C1(n9946), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9459), .B(
        n9458), .ZN(n9473) );
  INV_X1 U10727 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9460) );
  MUX2_X1 U10728 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n9460), .S(n9480), .Z(n9465) );
  AOI21_X1 U10729 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9462), .A(n9461), .ZN(
        n9463) );
  OAI211_X1 U10730 ( .C1(n9465), .C2(n9464), .A(n9528), .B(n9479), .ZN(n9472)
         );
  INV_X1 U10731 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9466) );
  MUX2_X1 U10732 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9466), .S(n9480), .Z(n9470) );
  OAI21_X1 U10733 ( .B1(n9468), .B2(n9443), .A(n9467), .ZN(n9469) );
  NAND2_X1 U10734 ( .A1(n9469), .A2(n9470), .ZN(n9474) );
  OAI211_X1 U10735 ( .C1(n9470), .C2(n9469), .A(n9551), .B(n9474), .ZN(n9471)
         );
  NAND3_X1 U10736 ( .A1(n9473), .A2(n9472), .A3(n9471), .ZN(P1_U3257) );
  OAI21_X1 U10737 ( .B1(n9466), .B2(n9475), .A(n9474), .ZN(n9487) );
  XNOR2_X1 U10738 ( .A(n9487), .B(n9494), .ZN(n9476) );
  NAND2_X1 U10739 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9476), .ZN(n9489) );
  OAI211_X1 U10740 ( .C1(n9476), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9551), .B(
        n9489), .ZN(n9486) );
  INV_X1 U10741 ( .A(n9477), .ZN(n9478) );
  AOI21_X1 U10742 ( .B1(n9946), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9478), .ZN(
        n9485) );
  XNOR2_X1 U10743 ( .A(n9495), .B(n9494), .ZN(n9481) );
  NOR2_X1 U10744 ( .A1(n6217), .A2(n9481), .ZN(n9496) );
  AOI21_X1 U10745 ( .B1(n6217), .B2(n9481), .A(n9496), .ZN(n9482) );
  NAND2_X1 U10746 ( .A1(n9528), .A2(n9482), .ZN(n9484) );
  NAND2_X1 U10747 ( .A1(n9958), .A2(n9488), .ZN(n9483) );
  NAND4_X1 U10748 ( .A1(n9486), .A2(n9485), .A3(n9484), .A4(n9483), .ZN(
        P1_U3258) );
  NAND2_X1 U10749 ( .A1(n9488), .A2(n9487), .ZN(n9490) );
  NAND2_X1 U10750 ( .A1(n9490), .A2(n9489), .ZN(n9493) );
  INV_X1 U10751 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9491) );
  MUX2_X1 U10752 ( .A(n9491), .B(P1_REG1_REG_16__SCAN_IN), .S(n9515), .Z(n9492) );
  NOR2_X1 U10753 ( .A1(n9492), .A2(n9493), .ZN(n9508) );
  AOI21_X1 U10754 ( .B1(n9493), .B2(n9492), .A(n9508), .ZN(n9507) );
  NOR2_X1 U10755 ( .A1(n9495), .A2(n9494), .ZN(n9497) );
  NOR2_X1 U10756 ( .A1(n9497), .A2(n9496), .ZN(n9500) );
  NAND2_X1 U10757 ( .A1(n9515), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9498) );
  OAI21_X1 U10758 ( .B1(n9515), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9498), .ZN(
        n9499) );
  NOR2_X1 U10759 ( .A1(n9500), .A2(n9499), .ZN(n9514) );
  AOI211_X1 U10760 ( .C1(n9500), .C2(n9499), .A(n9514), .B(n9962), .ZN(n9501)
         );
  INV_X1 U10761 ( .A(n9501), .ZN(n9506) );
  INV_X1 U10762 ( .A(n9946), .ZN(n9520) );
  INV_X1 U10763 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9503) );
  OAI21_X1 U10764 ( .B1(n9520), .B2(n9503), .A(n9502), .ZN(n9504) );
  AOI21_X1 U10765 ( .B1(n9515), .B2(n9958), .A(n9504), .ZN(n9505) );
  OAI211_X1 U10766 ( .C1(n9507), .C2(n9957), .A(n9506), .B(n9505), .ZN(
        P1_U3259) );
  AOI21_X1 U10767 ( .B1(n9509), .B2(n9491), .A(n9508), .ZN(n9512) );
  AOI22_X1 U10768 ( .A1(n9532), .A2(n6255), .B1(P1_REG1_REG_17__SCAN_IN), .B2(
        n9510), .ZN(n9511) );
  NOR2_X1 U10769 ( .A1(n9512), .A2(n9511), .ZN(n9536) );
  AOI21_X1 U10770 ( .B1(n9512), .B2(n9511), .A(n9536), .ZN(n9524) );
  NOR2_X1 U10771 ( .A1(n9532), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9513) );
  AOI21_X1 U10772 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9532), .A(n9513), .ZN(
        n9517) );
  AOI21_X1 U10773 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9515), .A(n9514), .ZN(
        n9516) );
  NAND2_X1 U10774 ( .A1(n9517), .A2(n9516), .ZN(n9525) );
  OAI21_X1 U10775 ( .B1(n9517), .B2(n9516), .A(n9525), .ZN(n9518) );
  NAND2_X1 U10776 ( .A1(n9518), .A2(n9528), .ZN(n9523) );
  INV_X1 U10777 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9519) );
  OAI22_X1 U10778 ( .A1(n9520), .A2(n9519), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6275), .ZN(n9521) );
  AOI21_X1 U10779 ( .B1(n9958), .B2(n9532), .A(n9521), .ZN(n9522) );
  OAI211_X1 U10780 ( .C1(n9524), .C2(n9957), .A(n9523), .B(n9522), .ZN(
        P1_U3260) );
  OAI21_X1 U10781 ( .B1(n9532), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9525), .ZN(
        n9526) );
  INV_X1 U10782 ( .A(n9526), .ZN(n9530) );
  INV_X1 U10783 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9527) );
  MUX2_X1 U10784 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9527), .S(n9546), .Z(n9529) );
  NAND2_X1 U10785 ( .A1(n9530), .A2(n9529), .ZN(n9544) );
  OAI211_X1 U10786 ( .C1(n9530), .C2(n9529), .A(n9544), .B(n9528), .ZN(n9542)
         );
  AOI21_X1 U10787 ( .B1(n9946), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9531), .ZN(
        n9541) );
  OR2_X1 U10788 ( .A1(n9532), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9534) );
  INV_X1 U10789 ( .A(n9534), .ZN(n9533) );
  NOR2_X1 U10790 ( .A1(n9536), .A2(n9533), .ZN(n9538) );
  XNOR2_X1 U10791 ( .A(n9546), .B(n9853), .ZN(n9537) );
  NAND2_X1 U10792 ( .A1(n9537), .A2(n9534), .ZN(n9535) );
  OR2_X1 U10793 ( .A1(n9536), .A2(n9535), .ZN(n9548) );
  OAI211_X1 U10794 ( .C1(n9538), .C2(n9537), .A(n9551), .B(n9548), .ZN(n9540)
         );
  NAND2_X1 U10795 ( .A1(n9958), .A2(n9546), .ZN(n9539) );
  NAND4_X1 U10796 ( .A1(n9542), .A2(n9541), .A3(n9540), .A4(n9539), .ZN(
        P1_U3261) );
  NAND2_X1 U10797 ( .A1(n9546), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U10798 ( .A1(n9544), .A2(n9543), .ZN(n9545) );
  XNOR2_X1 U10799 ( .A(n9545), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9550) );
  NAND2_X1 U10800 ( .A1(n9546), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U10801 ( .A1(n9548), .A2(n9547), .ZN(n9549) );
  XNOR2_X1 U10802 ( .A(n9549), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9552) );
  INV_X1 U10803 ( .A(n9550), .ZN(n9554) );
  AOI21_X1 U10804 ( .B1(n9552), .B2(n9551), .A(n9958), .ZN(n9553) );
  NAND2_X1 U10805 ( .A1(n9762), .A2(n9987), .ZN(n9562) );
  NOR2_X1 U10806 ( .A1(n9559), .A2(n9558), .ZN(n9765) );
  INV_X1 U10807 ( .A(n9765), .ZN(n9560) );
  NOR2_X1 U10808 ( .A1(n9991), .A2(n9560), .ZN(n9566) );
  AOI21_X1 U10809 ( .B1(n9734), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9566), .ZN(
        n9561) );
  OAI211_X1 U10810 ( .C1(n9860), .C2(n9719), .A(n9562), .B(n9561), .ZN(
        P1_U3263) );
  INV_X1 U10811 ( .A(n9564), .ZN(n9864) );
  XNOR2_X1 U10812 ( .A(n9564), .B(n9563), .ZN(n9565) );
  NAND2_X1 U10813 ( .A1(n9766), .A2(n9987), .ZN(n9568) );
  AOI21_X1 U10814 ( .B1(n9734), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9566), .ZN(
        n9567) );
  OAI211_X1 U10815 ( .C1(n9864), .C2(n9719), .A(n9568), .B(n9567), .ZN(
        P1_U3264) );
  NAND2_X1 U10816 ( .A1(n9570), .A2(n9569), .ZN(n9571) );
  NAND3_X1 U10817 ( .A1(n9572), .A2(n10075), .A3(n9571), .ZN(n9575) );
  AOI22_X1 U10818 ( .A1(n10063), .A2(n9783), .B1(n9573), .B2(n10030), .ZN(
        n9574) );
  AND2_X2 U10819 ( .A1(n9575), .A2(n9574), .ZN(n9770) );
  NAND2_X1 U10820 ( .A1(n9577), .A2(n9576), .ZN(n9578) );
  NAND2_X1 U10821 ( .A1(n9579), .A2(n9578), .ZN(n9771) );
  INV_X1 U10822 ( .A(n9771), .ZN(n9586) );
  OAI211_X1 U10823 ( .C1(n9581), .C2(n9593), .A(n9983), .B(n9580), .ZN(n9769)
         );
  AOI22_X1 U10824 ( .A1(n9734), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9977), .B2(
        n9582), .ZN(n9584) );
  NAND2_X1 U10825 ( .A1(n9867), .A2(n4511), .ZN(n9583) );
  OAI211_X1 U10826 ( .C1(n9769), .C2(n9741), .A(n9584), .B(n9583), .ZN(n9585)
         );
  AOI21_X1 U10827 ( .B1(n9586), .B2(n9731), .A(n9585), .ZN(n9587) );
  OAI21_X1 U10828 ( .B1(n9734), .B2(n9770), .A(n9587), .ZN(P1_U3265) );
  XNOR2_X1 U10829 ( .A(n9588), .B(n5052), .ZN(n9781) );
  XNOR2_X1 U10830 ( .A(n9590), .B(n9589), .ZN(n9774) );
  NAND2_X1 U10831 ( .A1(n9871), .A2(n9609), .ZN(n9591) );
  NAND2_X1 U10832 ( .A1(n9591), .A2(n9983), .ZN(n9592) );
  OR2_X1 U10833 ( .A1(n9593), .A2(n9592), .ZN(n9778) );
  NAND2_X1 U10834 ( .A1(n9732), .A2(n9775), .ZN(n9596) );
  AOI22_X1 U10835 ( .A1(n9991), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9977), .B2(
        n9594), .ZN(n9595) );
  OAI211_X1 U10836 ( .C1(n9738), .C2(n9597), .A(n9596), .B(n9595), .ZN(n9598)
         );
  AOI21_X1 U10837 ( .B1(n9871), .B2(n4511), .A(n9598), .ZN(n9599) );
  OAI21_X1 U10838 ( .B1(n9778), .B2(n9741), .A(n9599), .ZN(n9600) );
  AOI21_X1 U10839 ( .B1(n9774), .B2(n9731), .A(n9600), .ZN(n9601) );
  OAI21_X1 U10840 ( .B1(n9781), .B2(n9747), .A(n9601), .ZN(P1_U3266) );
  INV_X1 U10841 ( .A(n9602), .ZN(n9603) );
  AOI21_X1 U10842 ( .B1(n9614), .B2(n9604), .A(n9603), .ZN(n9787) );
  NAND2_X1 U10843 ( .A1(n9732), .A2(n9784), .ZN(n9607) );
  AOI22_X1 U10844 ( .A1(n9991), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9977), .B2(
        n9605), .ZN(n9606) );
  OAI211_X1 U10845 ( .C1(n9738), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9612)
         );
  INV_X1 U10846 ( .A(n9623), .ZN(n9610) );
  OAI211_X1 U10847 ( .C1(n9875), .C2(n9610), .A(n9609), .B(n9983), .ZN(n9785)
         );
  NOR2_X1 U10848 ( .A1(n9785), .A2(n9741), .ZN(n9611) );
  AOI211_X1 U10849 ( .C1(n4511), .C2(n9613), .A(n9612), .B(n9611), .ZN(n9617)
         );
  XNOR2_X1 U10850 ( .A(n9615), .B(n9614), .ZN(n9789) );
  NAND2_X1 U10851 ( .A1(n9789), .A2(n9731), .ZN(n9616) );
  OAI211_X1 U10852 ( .C1(n9787), .C2(n9747), .A(n9617), .B(n9616), .ZN(
        P1_U3267) );
  OAI211_X1 U10853 ( .C1(n9619), .C2(n9628), .A(n9618), .B(n10075), .ZN(n9621)
         );
  AOI22_X1 U10854 ( .A1(n10063), .A2(n9806), .B1(n9775), .B2(n10030), .ZN(
        n9620) );
  NAND2_X1 U10855 ( .A1(n9621), .A2(n9620), .ZN(n9793) );
  INV_X1 U10856 ( .A(n9793), .ZN(n9632) );
  OR2_X1 U10857 ( .A1(n9626), .A2(n4558), .ZN(n9622) );
  AND3_X1 U10858 ( .A1(n9623), .A2(n9622), .A3(n9983), .ZN(n9792) );
  AOI22_X1 U10859 ( .A1(n9734), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9977), .B2(
        n9624), .ZN(n9625) );
  OAI21_X1 U10860 ( .B1(n9626), .B2(n9719), .A(n9625), .ZN(n9627) );
  AOI21_X1 U10861 ( .B1(n9792), .B2(n9987), .A(n9627), .ZN(n9631) );
  XNOR2_X1 U10862 ( .A(n9629), .B(n9628), .ZN(n9794) );
  NAND2_X1 U10863 ( .A1(n9794), .A2(n9731), .ZN(n9630) );
  OAI211_X1 U10864 ( .C1(n9632), .C2(n9991), .A(n9631), .B(n9630), .ZN(
        P1_U3268) );
  OAI211_X1 U10865 ( .C1(n4576), .C2(n5047), .A(n9633), .B(n10075), .ZN(n9635)
         );
  AOI22_X1 U10866 ( .A1(n10063), .A2(n9816), .B1(n9784), .B2(n10030), .ZN(
        n9634) );
  NAND2_X1 U10867 ( .A1(n9635), .A2(n9634), .ZN(n9800) );
  INV_X1 U10868 ( .A(n9800), .ZN(n9644) );
  AOI211_X1 U10869 ( .C1(n9636), .C2(n9652), .A(n9715), .B(n4558), .ZN(n9801)
         );
  INV_X1 U10870 ( .A(n9636), .ZN(n9884) );
  AOI22_X1 U10871 ( .A1(n9734), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9977), .B2(
        n9637), .ZN(n9638) );
  OAI21_X1 U10872 ( .B1(n9884), .B2(n9719), .A(n9638), .ZN(n9639) );
  AOI21_X1 U10873 ( .B1(n9801), .B2(n9987), .A(n9639), .ZN(n9643) );
  XNOR2_X1 U10874 ( .A(n9641), .B(n9640), .ZN(n9802) );
  NAND2_X1 U10875 ( .A1(n9802), .A2(n9731), .ZN(n9642) );
  OAI211_X1 U10876 ( .C1(n9644), .C2(n9991), .A(n9643), .B(n9642), .ZN(
        P1_U3269) );
  XNOR2_X1 U10877 ( .A(n9645), .B(n9646), .ZN(n9810) );
  INV_X1 U10878 ( .A(n9810), .ZN(n9659) );
  XNOR2_X1 U10879 ( .A(n9647), .B(n9646), .ZN(n9805) );
  NAND2_X1 U10880 ( .A1(n9805), .A2(n9731), .ZN(n9658) );
  NAND2_X1 U10881 ( .A1(n9732), .A2(n9827), .ZN(n9650) );
  AOI22_X1 U10882 ( .A1(n9734), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9977), .B2(
        n9648), .ZN(n9649) );
  OAI211_X1 U10883 ( .C1(n9738), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9655)
         );
  AOI21_X1 U10884 ( .B1(n9667), .B2(n9656), .A(n9715), .ZN(n9653) );
  NAND2_X1 U10885 ( .A1(n9653), .A2(n9652), .ZN(n9808) );
  NOR2_X1 U10886 ( .A1(n9808), .A2(n9741), .ZN(n9654) );
  AOI211_X1 U10887 ( .C1(n4511), .C2(n9656), .A(n9655), .B(n9654), .ZN(n9657)
         );
  OAI211_X1 U10888 ( .C1(n9659), .C2(n9747), .A(n9658), .B(n9657), .ZN(
        P1_U3270) );
  XNOR2_X1 U10889 ( .A(n9660), .B(n9661), .ZN(n9822) );
  INV_X1 U10890 ( .A(n9822), .ZN(n9673) );
  XNOR2_X1 U10891 ( .A(n9662), .B(n9661), .ZN(n9815) );
  NAND2_X1 U10892 ( .A1(n9815), .A2(n9731), .ZN(n9672) );
  NAND2_X1 U10893 ( .A1(n9732), .A2(n9817), .ZN(n9665) );
  AOI22_X1 U10894 ( .A1(n9991), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9977), .B2(
        n9663), .ZN(n9664) );
  OAI211_X1 U10895 ( .C1(n9738), .C2(n9666), .A(n9665), .B(n9664), .ZN(n9669)
         );
  OAI211_X1 U10896 ( .C1(n9892), .C2(n9684), .A(n9983), .B(n9667), .ZN(n9819)
         );
  NOR2_X1 U10897 ( .A1(n9819), .A2(n9741), .ZN(n9668) );
  AOI211_X1 U10898 ( .C1(n4511), .C2(n9670), .A(n9669), .B(n9668), .ZN(n9671)
         );
  OAI211_X1 U10899 ( .C1(n9673), .C2(n9747), .A(n9672), .B(n9671), .ZN(
        P1_U3271) );
  OAI21_X1 U10900 ( .B1(n9675), .B2(n9677), .A(n9674), .ZN(n9676) );
  INV_X1 U10901 ( .A(n9676), .ZN(n9831) );
  XOR2_X1 U10902 ( .A(n9678), .B(n9677), .Z(n9833) );
  NAND2_X1 U10903 ( .A1(n9833), .A2(n9731), .ZN(n9690) );
  NAND2_X1 U10904 ( .A1(n9732), .A2(n9828), .ZN(n9681) );
  AOI22_X1 U10905 ( .A1(n9734), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9977), .B2(
        n9679), .ZN(n9680) );
  OAI211_X1 U10906 ( .C1(n9738), .C2(n9682), .A(n9681), .B(n9680), .ZN(n9687)
         );
  INV_X1 U10907 ( .A(n9683), .ZN(n9697) );
  INV_X1 U10908 ( .A(n9684), .ZN(n9685) );
  OAI211_X1 U10909 ( .C1(n9896), .C2(n9697), .A(n9685), .B(n9983), .ZN(n9829)
         );
  NOR2_X1 U10910 ( .A1(n9829), .A2(n9741), .ZN(n9686) );
  AOI211_X1 U10911 ( .C1(n4511), .C2(n9688), .A(n9687), .B(n9686), .ZN(n9689)
         );
  OAI211_X1 U10912 ( .C1(n9831), .C2(n9747), .A(n9690), .B(n9689), .ZN(
        P1_U3272) );
  OAI211_X1 U10913 ( .C1(n9695), .C2(n9692), .A(n9691), .B(n10075), .ZN(n9694)
         );
  AOI22_X1 U10914 ( .A1(n10063), .A2(n9846), .B1(n9817), .B2(n10030), .ZN(
        n9693) );
  NAND2_X1 U10915 ( .A1(n9694), .A2(n9693), .ZN(n9836) );
  INV_X1 U10916 ( .A(n9836), .ZN(n9704) );
  XNOR2_X1 U10917 ( .A(n4636), .B(n9695), .ZN(n9838) );
  NAND2_X1 U10918 ( .A1(n9838), .A2(n9731), .ZN(n9703) );
  AOI211_X1 U10919 ( .C1(n9698), .C2(n9714), .A(n9715), .B(n9697), .ZN(n9837)
         );
  AOI22_X1 U10920 ( .A1(n9734), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9977), .B2(
        n9699), .ZN(n9700) );
  OAI21_X1 U10921 ( .B1(n4966), .B2(n9719), .A(n9700), .ZN(n9701) );
  AOI21_X1 U10922 ( .B1(n9837), .B2(n9987), .A(n9701), .ZN(n9702) );
  OAI211_X1 U10923 ( .C1(n9991), .C2(n9704), .A(n9703), .B(n9702), .ZN(
        P1_U3273) );
  XOR2_X1 U10924 ( .A(n9705), .B(n9707), .Z(n9845) );
  INV_X1 U10925 ( .A(n9706), .ZN(n9710) );
  INV_X1 U10926 ( .A(n9707), .ZN(n9709) );
  OAI211_X1 U10927 ( .C1(n9710), .C2(n9709), .A(n10075), .B(n9708), .ZN(n9713)
         );
  AOI22_X1 U10928 ( .A1(n9711), .A2(n10063), .B1(n10030), .B2(n9828), .ZN(
        n9712) );
  NAND2_X1 U10929 ( .A1(n9713), .A2(n9712), .ZN(n9841) );
  AOI211_X1 U10930 ( .C1(n9843), .C2(n9739), .A(n9715), .B(n4967), .ZN(n9842)
         );
  NAND2_X1 U10931 ( .A1(n9842), .A2(n9987), .ZN(n9718) );
  AOI22_X1 U10932 ( .A1(n9734), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9977), .B2(
        n9716), .ZN(n9717) );
  OAI211_X1 U10933 ( .C1(n9720), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9721)
         );
  AOI21_X1 U10934 ( .B1(n9757), .B2(n9841), .A(n9721), .ZN(n9722) );
  OAI21_X1 U10935 ( .B1(n9845), .B2(n9723), .A(n9722), .ZN(P1_U3274) );
  NAND2_X1 U10936 ( .A1(n9725), .A2(n9724), .ZN(n9728) );
  INV_X1 U10937 ( .A(n9726), .ZN(n9727) );
  AOI21_X1 U10938 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9850) );
  XOR2_X1 U10939 ( .A(n9730), .B(n9729), .Z(n9852) );
  NAND2_X1 U10940 ( .A1(n9852), .A2(n9731), .ZN(n9746) );
  NAND2_X1 U10941 ( .A1(n9732), .A2(n9918), .ZN(n9736) );
  AOI22_X1 U10942 ( .A1(n9734), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9977), .B2(
        n9733), .ZN(n9735) );
  OAI211_X1 U10943 ( .C1(n9738), .C2(n9737), .A(n9736), .B(n9735), .ZN(n9743)
         );
  OAI211_X1 U10944 ( .C1(n9905), .C2(n9740), .A(n9983), .B(n9739), .ZN(n9847)
         );
  NOR2_X1 U10945 ( .A1(n9847), .A2(n9741), .ZN(n9742) );
  AOI211_X1 U10946 ( .C1(n4511), .C2(n9744), .A(n9743), .B(n9742), .ZN(n9745)
         );
  OAI211_X1 U10947 ( .C1(n9850), .C2(n9747), .A(n9746), .B(n9745), .ZN(
        P1_U3275) );
  OAI21_X1 U10948 ( .B1(n9749), .B2(n4511), .A(n9748), .ZN(n9761) );
  NAND2_X1 U10949 ( .A1(n9751), .A2(n9750), .ZN(n9760) );
  INV_X1 U10950 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9752) );
  OAI22_X1 U10951 ( .A1(n9755), .A2(n9754), .B1(n9753), .B2(n9752), .ZN(n9756)
         );
  NAND2_X1 U10952 ( .A1(n9757), .A2(n9756), .ZN(n9759) );
  NAND2_X1 U10953 ( .A1(n9991), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9758) );
  NAND4_X1 U10954 ( .A1(n9761), .A2(n9760), .A3(n9759), .A4(n9758), .ZN(
        P1_U3293) );
  INV_X1 U10955 ( .A(n9798), .ZN(n9855) );
  INV_X1 U10956 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9763) );
  NOR2_X1 U10957 ( .A1(n9762), .A2(n9765), .ZN(n9857) );
  MUX2_X1 U10958 ( .A(n9763), .B(n9857), .S(n10094), .Z(n9764) );
  OAI21_X1 U10959 ( .B1(n9860), .B2(n9855), .A(n9764), .ZN(P1_U3553) );
  INV_X1 U10960 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9767) );
  NOR2_X1 U10961 ( .A1(n9766), .A2(n9765), .ZN(n9861) );
  MUX2_X1 U10962 ( .A(n9767), .B(n9861), .S(n10094), .Z(n9768) );
  OAI21_X1 U10963 ( .B1(n9864), .B2(n9855), .A(n9768), .ZN(P1_U3552) );
  AOI21_X1 U10964 ( .B1(n9798), .B2(n9867), .A(n9772), .ZN(n9773) );
  INV_X1 U10965 ( .A(n9773), .ZN(P1_U3550) );
  NAND2_X1 U10966 ( .A1(n9774), .A2(n10060), .ZN(n9780) );
  AOI22_X1 U10967 ( .A1(n9776), .A2(n10064), .B1(n10063), .B2(n9775), .ZN(
        n9777) );
  AND2_X1 U10968 ( .A1(n9778), .A2(n9777), .ZN(n9779) );
  OAI211_X1 U10969 ( .C1(n9849), .C2(n9781), .A(n9779), .B(n9780), .ZN(n9869)
         );
  INV_X1 U10970 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9790) );
  AOI22_X1 U10971 ( .A1(n10063), .A2(n9784), .B1(n9783), .B2(n10030), .ZN(
        n9786) );
  OAI211_X1 U10972 ( .C1(n9787), .C2(n9849), .A(n9786), .B(n9785), .ZN(n9788)
         );
  AOI21_X1 U10973 ( .B1(n9789), .B2(n10060), .A(n9788), .ZN(n9872) );
  MUX2_X1 U10974 ( .A(n9790), .B(n9872), .S(n10094), .Z(n9791) );
  OAI21_X1 U10975 ( .B1(n9875), .B2(n9855), .A(n9791), .ZN(P1_U3548) );
  NOR2_X1 U10976 ( .A1(n9793), .A2(n9792), .ZN(n9796) );
  NAND2_X1 U10977 ( .A1(n9794), .A2(n10060), .ZN(n9795) );
  NAND2_X1 U10978 ( .A1(n9796), .A2(n9795), .ZN(n9876) );
  MUX2_X1 U10979 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9876), .S(n10094), .Z(
        n9797) );
  AOI21_X1 U10980 ( .B1(n9798), .B2(n9878), .A(n9797), .ZN(n9799) );
  INV_X1 U10981 ( .A(n9799), .ZN(P1_U3547) );
  INV_X1 U10982 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9803) );
  AOI211_X1 U10983 ( .C1(n10060), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9881)
         );
  MUX2_X1 U10984 ( .A(n9803), .B(n9881), .S(n10094), .Z(n9804) );
  OAI21_X1 U10985 ( .B1(n9884), .B2(n9855), .A(n9804), .ZN(P1_U3546) );
  INV_X1 U10986 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U10987 ( .A1(n9805), .A2(n10060), .ZN(n9812) );
  AOI22_X1 U10988 ( .A1(n10064), .A2(n9806), .B1(n9827), .B2(n10063), .ZN(
        n9807) );
  NAND2_X1 U10989 ( .A1(n9808), .A2(n9807), .ZN(n9809) );
  AOI21_X1 U10990 ( .B1(n9810), .B2(n9821), .A(n9809), .ZN(n9811) );
  AND2_X1 U10991 ( .A1(n9812), .A2(n9811), .ZN(n9885) );
  MUX2_X1 U10992 ( .A(n9813), .B(n9885), .S(n10094), .Z(n9814) );
  OAI21_X1 U10993 ( .B1(n9888), .B2(n9855), .A(n9814), .ZN(P1_U3545) );
  INV_X1 U10994 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U10995 ( .A1(n9815), .A2(n10060), .ZN(n9824) );
  AOI22_X1 U10996 ( .A1(n10063), .A2(n9817), .B1(n9816), .B2(n10030), .ZN(
        n9818) );
  NAND2_X1 U10997 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  AOI21_X1 U10998 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9823) );
  AND2_X1 U10999 ( .A1(n9824), .A2(n9823), .ZN(n9889) );
  MUX2_X1 U11000 ( .A(n9825), .B(n9889), .S(n10094), .Z(n9826) );
  OAI21_X1 U11001 ( .B1(n9892), .B2(n9855), .A(n9826), .ZN(P1_U3544) );
  INV_X1 U11002 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9834) );
  AOI22_X1 U11003 ( .A1(n10063), .A2(n9828), .B1(n9827), .B2(n10030), .ZN(
        n9830) );
  OAI211_X1 U11004 ( .C1(n9831), .C2(n9849), .A(n9830), .B(n9829), .ZN(n9832)
         );
  AOI21_X1 U11005 ( .B1(n9833), .B2(n10060), .A(n9832), .ZN(n9893) );
  MUX2_X1 U11006 ( .A(n9834), .B(n9893), .S(n10094), .Z(n9835) );
  OAI21_X1 U11007 ( .B1(n9896), .B2(n9855), .A(n9835), .ZN(P1_U3543) );
  INV_X1 U11008 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9839) );
  AOI211_X1 U11009 ( .C1(n9838), .C2(n10060), .A(n9837), .B(n9836), .ZN(n9897)
         );
  MUX2_X1 U11010 ( .A(n9839), .B(n9897), .S(n10094), .Z(n9840) );
  OAI21_X1 U11011 ( .B1(n4966), .B2(n9855), .A(n9840), .ZN(P1_U3542) );
  AOI211_X1 U11012 ( .C1(n10042), .C2(n9843), .A(n9842), .B(n9841), .ZN(n9844)
         );
  OAI21_X1 U11013 ( .B1(n10070), .B2(n9845), .A(n9844), .ZN(n9900) );
  MUX2_X1 U11014 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9900), .S(n10094), .Z(
        P1_U3541) );
  AOI22_X1 U11015 ( .A1(n9918), .A2(n10063), .B1(n10030), .B2(n9846), .ZN(
        n9848) );
  OAI211_X1 U11016 ( .C1(n9850), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9851)
         );
  AOI21_X1 U11017 ( .B1(n9852), .B2(n10060), .A(n9851), .ZN(n9901) );
  MUX2_X1 U11018 ( .A(n9853), .B(n9901), .S(n10094), .Z(n9854) );
  OAI21_X1 U11019 ( .B1(n9905), .B2(n9855), .A(n9854), .ZN(P1_U3540) );
  MUX2_X1 U11020 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9856), .S(n10094), .Z(
        P1_U3522) );
  INV_X1 U11021 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9858) );
  MUX2_X1 U11022 ( .A(n9858), .B(n9857), .S(n10078), .Z(n9859) );
  OAI21_X1 U11023 ( .B1(n9860), .B2(n9904), .A(n9859), .ZN(P1_U3521) );
  INV_X1 U11024 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9862) );
  MUX2_X1 U11025 ( .A(n9862), .B(n9861), .S(n10078), .Z(n9863) );
  OAI21_X1 U11026 ( .B1(n9864), .B2(n9904), .A(n9863), .ZN(P1_U3520) );
  AOI21_X1 U11027 ( .B1(n9879), .B2(n9867), .A(n9866), .ZN(n9868) );
  INV_X1 U11028 ( .A(n9868), .ZN(P1_U3518) );
  INV_X1 U11029 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9873) );
  MUX2_X1 U11030 ( .A(n9873), .B(n9872), .S(n10078), .Z(n9874) );
  OAI21_X1 U11031 ( .B1(n9875), .B2(n9904), .A(n9874), .ZN(P1_U3516) );
  MUX2_X1 U11032 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9876), .S(n10078), .Z(
        n9877) );
  AOI21_X1 U11033 ( .B1(n9879), .B2(n9878), .A(n9877), .ZN(n9880) );
  INV_X1 U11034 ( .A(n9880), .ZN(P1_U3515) );
  INV_X1 U11035 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9882) );
  MUX2_X1 U11036 ( .A(n9882), .B(n9881), .S(n10078), .Z(n9883) );
  OAI21_X1 U11037 ( .B1(n9884), .B2(n9904), .A(n9883), .ZN(P1_U3514) );
  INV_X1 U11038 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9886) );
  MUX2_X1 U11039 ( .A(n9886), .B(n9885), .S(n10078), .Z(n9887) );
  OAI21_X1 U11040 ( .B1(n9888), .B2(n9904), .A(n9887), .ZN(P1_U3513) );
  INV_X1 U11041 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9890) );
  MUX2_X1 U11042 ( .A(n9890), .B(n9889), .S(n10078), .Z(n9891) );
  OAI21_X1 U11043 ( .B1(n9892), .B2(n9904), .A(n9891), .ZN(P1_U3512) );
  INV_X1 U11044 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9894) );
  MUX2_X1 U11045 ( .A(n9894), .B(n9893), .S(n10078), .Z(n9895) );
  OAI21_X1 U11046 ( .B1(n9896), .B2(n9904), .A(n9895), .ZN(P1_U3511) );
  INV_X1 U11047 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9898) );
  MUX2_X1 U11048 ( .A(n9898), .B(n9897), .S(n10078), .Z(n9899) );
  OAI21_X1 U11049 ( .B1(n4966), .B2(n9904), .A(n9899), .ZN(P1_U3510) );
  MUX2_X1 U11050 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9900), .S(n10078), .Z(
        P1_U3509) );
  INV_X1 U11051 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9902) );
  MUX2_X1 U11052 ( .A(n9902), .B(n9901), .S(n10078), .Z(n9903) );
  OAI21_X1 U11053 ( .B1(n9905), .B2(n9904), .A(n9903), .ZN(P1_U3507) );
  NOR4_X1 U11054 ( .A1(n9906), .A2(P1_IR_REG_30__SCAN_IN), .A3(n6130), .A4(
        P1_U3086), .ZN(n9907) );
  AOI21_X1 U11055 ( .B1(n9908), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9907), .ZN(
        n9909) );
  OAI21_X1 U11056 ( .B1(n9911), .B2(n9910), .A(n9909), .ZN(P1_U3324) );
  MUX2_X1 U11057 ( .A(n9912), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U11058 ( .B1(n9914), .B2(n10068), .A(n9913), .ZN(n9916) );
  AOI211_X1 U11059 ( .C1(n9917), .C2(n10060), .A(n9916), .B(n9915), .ZN(n9935)
         );
  AOI22_X1 U11060 ( .A1(n10094), .A2(n9935), .B1(n6255), .B2(n10092), .ZN(
        P1_U3539) );
  AOI22_X1 U11061 ( .A1(n9918), .A2(n10064), .B1(n10063), .B2(n10065), .ZN(
        n9919) );
  OAI211_X1 U11062 ( .C1(n9921), .C2(n10068), .A(n9920), .B(n9919), .ZN(n9925)
         );
  AND3_X1 U11063 ( .A1(n9923), .A2(n10060), .A3(n9922), .ZN(n9924) );
  AOI211_X1 U11064 ( .C1(n10075), .C2(n9926), .A(n9925), .B(n9924), .ZN(n9937)
         );
  AOI22_X1 U11065 ( .A1(n10094), .A2(n9937), .B1(n9491), .B2(n10092), .ZN(
        P1_U3538) );
  INV_X1 U11066 ( .A(n9927), .ZN(n9929) );
  OAI21_X1 U11067 ( .B1(n9929), .B2(n10068), .A(n9928), .ZN(n9931) );
  AOI211_X1 U11068 ( .C1(n9932), .C2(n10060), .A(n9931), .B(n9930), .ZN(n9939)
         );
  INV_X1 U11069 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9933) );
  AOI22_X1 U11070 ( .A1(n10094), .A2(n9939), .B1(n9933), .B2(n10092), .ZN(
        P1_U3537) );
  INV_X1 U11071 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9934) );
  AOI22_X1 U11072 ( .A1(n10078), .A2(n9935), .B1(n9934), .B2(n10076), .ZN(
        P1_U3504) );
  INV_X1 U11073 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9936) );
  AOI22_X1 U11074 ( .A1(n10078), .A2(n9937), .B1(n9936), .B2(n10076), .ZN(
        P1_U3501) );
  INV_X1 U11075 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U11076 ( .A1(n10078), .A2(n9939), .B1(n9938), .B2(n10076), .ZN(
        P1_U3498) );
  XNOR2_X1 U11077 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11078 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11079 ( .B1(n9941), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9940), .ZN(
        n9942) );
  XOR2_X1 U11080 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9942), .Z(n9945) );
  AOI22_X1 U11081 ( .A1(n9946), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9943) );
  OAI21_X1 U11082 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(P1_U3243) );
  AOI22_X1 U11083 ( .A1(n9946), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9966) );
  INV_X1 U11084 ( .A(n9947), .ZN(n9950) );
  NAND3_X1 U11085 ( .A1(n9950), .A2(n9949), .A3(n9948), .ZN(n9952) );
  NAND2_X1 U11086 ( .A1(n9952), .A2(n9951), .ZN(n9961) );
  OAI21_X1 U11087 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(n9956) );
  OR2_X1 U11088 ( .A1(n9957), .A2(n9956), .ZN(n9960) );
  NAND2_X1 U11089 ( .A1(n9958), .A2(n4647), .ZN(n9959) );
  OAI211_X1 U11090 ( .C1(n9962), .C2(n9961), .A(n9960), .B(n9959), .ZN(n9963)
         );
  INV_X1 U11091 ( .A(n9963), .ZN(n9965) );
  NAND3_X1 U11092 ( .A1(n9966), .A2(n9965), .A3(n9964), .ZN(P1_U3245) );
  XNOR2_X1 U11093 ( .A(n9967), .B(n9973), .ZN(n9976) );
  OAI22_X1 U11094 ( .A1(n9971), .A2(n9970), .B1(n9969), .B2(n9968), .ZN(n9975)
         );
  XNOR2_X1 U11095 ( .A(n9972), .B(n9973), .ZN(n9981) );
  NOR2_X1 U11096 ( .A1(n9981), .A2(n9996), .ZN(n9974) );
  AOI211_X1 U11097 ( .C1(n10075), .C2(n9976), .A(n9975), .B(n9974), .ZN(n10050) );
  AOI222_X1 U11098 ( .A1(n9980), .A2(n4511), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9991), .C1(n9978), .C2(n9977), .ZN(n9990) );
  INV_X1 U11099 ( .A(n9981), .ZN(n10053) );
  NOR2_X1 U11100 ( .A1(n9991), .A2(n9982), .ZN(n9988) );
  OAI211_X1 U11101 ( .C1(n9985), .C2(n10049), .A(n9984), .B(n9983), .ZN(n10048) );
  INV_X1 U11102 ( .A(n10048), .ZN(n9986) );
  AOI22_X1 U11103 ( .A1(n10053), .A2(n9988), .B1(n9987), .B2(n9986), .ZN(n9989) );
  OAI211_X1 U11104 ( .C1(n9991), .C2(n10050), .A(n9990), .B(n9989), .ZN(
        P1_U3286) );
  AND2_X1 U11105 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9992), .ZN(P1_U3294) );
  AND2_X1 U11106 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9992), .ZN(P1_U3295) );
  AND2_X1 U11107 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9992), .ZN(P1_U3296) );
  AND2_X1 U11108 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9992), .ZN(P1_U3297) );
  AND2_X1 U11109 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9992), .ZN(P1_U3298) );
  AND2_X1 U11110 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9992), .ZN(P1_U3299) );
  AND2_X1 U11111 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9992), .ZN(P1_U3300) );
  AND2_X1 U11112 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9992), .ZN(P1_U3301) );
  AND2_X1 U11113 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9992), .ZN(P1_U3302) );
  AND2_X1 U11114 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9992), .ZN(P1_U3303) );
  AND2_X1 U11115 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9992), .ZN(P1_U3304) );
  AND2_X1 U11116 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9992), .ZN(P1_U3305) );
  AND2_X1 U11117 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9992), .ZN(P1_U3306) );
  AND2_X1 U11118 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9992), .ZN(P1_U3307) );
  AND2_X1 U11119 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9992), .ZN(P1_U3308) );
  AND2_X1 U11120 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9992), .ZN(P1_U3309) );
  AND2_X1 U11121 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9992), .ZN(P1_U3310) );
  AND2_X1 U11122 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9992), .ZN(P1_U3311) );
  AND2_X1 U11123 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9992), .ZN(P1_U3312) );
  AND2_X1 U11124 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9992), .ZN(P1_U3313) );
  AND2_X1 U11125 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9992), .ZN(P1_U3314) );
  AND2_X1 U11126 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9992), .ZN(P1_U3315) );
  AND2_X1 U11127 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9992), .ZN(P1_U3316) );
  AND2_X1 U11128 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9992), .ZN(P1_U3317) );
  AND2_X1 U11129 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9992), .ZN(P1_U3318) );
  AND2_X1 U11130 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9992), .ZN(P1_U3319) );
  INV_X1 U11131 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10576) );
  NOR2_X1 U11132 ( .A1(n9993), .A2(n10576), .ZN(P1_U3320) );
  INV_X1 U11133 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10367) );
  NOR2_X1 U11134 ( .A1(n9993), .A2(n10367), .ZN(P1_U3321) );
  AND2_X1 U11135 ( .A1(n9992), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3322) );
  INV_X1 U11136 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10404) );
  NOR2_X1 U11137 ( .A1(n9993), .A2(n10404), .ZN(P1_U3323) );
  OAI21_X1 U11138 ( .B1(n9995), .B2(n10601), .A(n9994), .ZN(P1_U3439) );
  INV_X1 U11139 ( .A(n9996), .ZN(n10009) );
  INV_X1 U11140 ( .A(n10008), .ZN(n10006) );
  AOI22_X1 U11141 ( .A1(n10063), .A2(n9998), .B1(n9997), .B2(n10030), .ZN(
        n10000) );
  OAI211_X1 U11142 ( .C1(n10001), .C2(n10068), .A(n10000), .B(n9999), .ZN(
        n10002) );
  INV_X1 U11143 ( .A(n10002), .ZN(n10004) );
  OAI211_X1 U11144 ( .C1(n10006), .C2(n10005), .A(n10004), .B(n10003), .ZN(
        n10007) );
  AOI21_X1 U11145 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(n10080) );
  INV_X1 U11146 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U11147 ( .A1(n10078), .A2(n10080), .B1(n10010), .B2(n10076), .ZN(
        P1_U3456) );
  OAI21_X1 U11148 ( .B1(n10012), .B2(n10068), .A(n10011), .ZN(n10014) );
  AOI211_X1 U11149 ( .C1(n10060), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10081) );
  INV_X1 U11150 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10016) );
  AOI22_X1 U11151 ( .A1(n10078), .A2(n10081), .B1(n10016), .B2(n10076), .ZN(
        P1_U3459) );
  OAI211_X1 U11152 ( .C1(n10019), .C2(n10068), .A(n10018), .B(n10017), .ZN(
        n10020) );
  AOI21_X1 U11153 ( .B1(n10060), .B2(n10021), .A(n10020), .ZN(n10083) );
  INV_X1 U11154 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10022) );
  AOI22_X1 U11155 ( .A1(n10078), .A2(n10083), .B1(n10022), .B2(n10076), .ZN(
        P1_U3462) );
  OAI21_X1 U11156 ( .B1(n10024), .B2(n10068), .A(n10023), .ZN(n10026) );
  AOI211_X1 U11157 ( .C1(n10060), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10084) );
  INV_X1 U11158 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10028) );
  AOI22_X1 U11159 ( .A1(n10078), .A2(n10084), .B1(n10028), .B2(n10076), .ZN(
        P1_U3465) );
  AOI22_X1 U11160 ( .A1(n10031), .A2(n10042), .B1(n10030), .B2(n10029), .ZN(
        n10032) );
  NAND2_X1 U11161 ( .A1(n10033), .A2(n10032), .ZN(n10034) );
  NOR2_X1 U11162 ( .A1(n10035), .A2(n10034), .ZN(n10038) );
  NAND2_X1 U11163 ( .A1(n10036), .A2(n10060), .ZN(n10037) );
  AND2_X1 U11164 ( .A1(n10038), .A2(n10037), .ZN(n10086) );
  INV_X1 U11165 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10039) );
  AOI22_X1 U11166 ( .A1(n10078), .A2(n10086), .B1(n10039), .B2(n10076), .ZN(
        P1_U3468) );
  AOI21_X1 U11167 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n10043) );
  OAI211_X1 U11168 ( .C1(n10070), .C2(n10045), .A(n10044), .B(n10043), .ZN(
        n10046) );
  INV_X1 U11169 ( .A(n10046), .ZN(n10088) );
  INV_X1 U11170 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U11171 ( .A1(n10078), .A2(n10088), .B1(n10047), .B2(n10076), .ZN(
        P1_U3471) );
  OAI21_X1 U11172 ( .B1(n10049), .B2(n10068), .A(n10048), .ZN(n10052) );
  INV_X1 U11173 ( .A(n10050), .ZN(n10051) );
  AOI211_X1 U11174 ( .C1(n10054), .C2(n10053), .A(n10052), .B(n10051), .ZN(
        n10090) );
  INV_X1 U11175 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11176 ( .A1(n10078), .A2(n10090), .B1(n10055), .B2(n10076), .ZN(
        P1_U3474) );
  OAI21_X1 U11177 ( .B1(n4974), .B2(n10068), .A(n10056), .ZN(n10058) );
  AOI211_X1 U11178 ( .C1(n10060), .C2(n10059), .A(n10058), .B(n10057), .ZN(
        n10091) );
  INV_X1 U11179 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10061) );
  AOI22_X1 U11180 ( .A1(n10078), .A2(n10091), .B1(n10061), .B2(n10076), .ZN(
        P1_U3492) );
  AOI22_X1 U11181 ( .A1(n10065), .A2(n10064), .B1(n10063), .B2(n10062), .ZN(
        n10066) );
  OAI211_X1 U11182 ( .C1(n10069), .C2(n10068), .A(n10067), .B(n10066), .ZN(
        n10073) );
  NOR2_X1 U11183 ( .A1(n10071), .A2(n10070), .ZN(n10072) );
  AOI211_X1 U11184 ( .C1(n10075), .C2(n10074), .A(n10073), .B(n10072), .ZN(
        n10093) );
  INV_X1 U11185 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10077) );
  AOI22_X1 U11186 ( .A1(n10078), .A2(n10093), .B1(n10077), .B2(n10076), .ZN(
        P1_U3495) );
  AOI22_X1 U11187 ( .A1(n10094), .A2(n10080), .B1(n10079), .B2(n10092), .ZN(
        P1_U3523) );
  AOI22_X1 U11188 ( .A1(n10094), .A2(n10081), .B1(n7027), .B2(n10092), .ZN(
        P1_U3524) );
  AOI22_X1 U11189 ( .A1(n10094), .A2(n10083), .B1(n10082), .B2(n10092), .ZN(
        P1_U3525) );
  AOI22_X1 U11190 ( .A1(n10094), .A2(n10084), .B1(n7031), .B2(n10092), .ZN(
        P1_U3526) );
  AOI22_X1 U11191 ( .A1(n10094), .A2(n10086), .B1(n10085), .B2(n10092), .ZN(
        P1_U3527) );
  AOI22_X1 U11192 ( .A1(n10094), .A2(n10088), .B1(n10087), .B2(n10092), .ZN(
        P1_U3528) );
  AOI22_X1 U11193 ( .A1(n10094), .A2(n10090), .B1(n10089), .B2(n10092), .ZN(
        P1_U3529) );
  AOI22_X1 U11194 ( .A1(n10094), .A2(n10091), .B1(n9443), .B2(n10092), .ZN(
        P1_U3535) );
  AOI22_X1 U11195 ( .A1(n10094), .A2(n10093), .B1(n9466), .B2(n10092), .ZN(
        P1_U3536) );
  OAI211_X1 U11196 ( .C1(n10098), .C2(n10097), .A(n10096), .B(n10095), .ZN(
        n10099) );
  INV_X1 U11197 ( .A(n10099), .ZN(n10109) );
  OAI21_X1 U11198 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(n10104) );
  AOI22_X1 U11199 ( .A1(n10105), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n6720), .B2(
        n10104), .ZN(n10106) );
  OAI21_X1 U11200 ( .B1(n6680), .B2(n10107), .A(n10106), .ZN(n10108) );
  NOR2_X1 U11201 ( .A1(n10109), .A2(n10108), .ZN(n10116) );
  OAI21_X1 U11202 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(n10113) );
  NAND2_X1 U11203 ( .A1(n10114), .A2(n10113), .ZN(n10115) );
  OAI211_X1 U11204 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7276), .A(n10116), .B(
        n10115), .ZN(P2_U3184) );
  XOR2_X1 U11205 ( .A(n10117), .B(n10128), .Z(n10122) );
  AOI222_X1 U11206 ( .A1(n10123), .A2(n10122), .B1(n10121), .B2(n10120), .C1(
        n10119), .C2(n10118), .ZN(n10156) );
  INV_X1 U11207 ( .A(n10124), .ZN(n10134) );
  OAI21_X1 U11208 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(n10129) );
  XNOR2_X1 U11209 ( .A(n10129), .B(n10128), .ZN(n10159) );
  AOI222_X1 U11210 ( .A1(n10134), .A2(n10133), .B1(n10159), .B2(n10132), .C1(
        n10131), .C2(n10130), .ZN(n10135) );
  OAI221_X1 U11211 ( .B1(n10136), .B2(n10156), .C1(n8779), .C2(n6631), .A(
        n10135), .ZN(P2_U3227) );
  INV_X1 U11212 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U11213 ( .A1(n10137), .A2(n10183), .ZN(n10139) );
  AOI211_X1 U11214 ( .C1(n10181), .C2(n10140), .A(n10139), .B(n10138), .ZN(
        n10199) );
  AOI22_X1 U11215 ( .A1(n10198), .A2(n10141), .B1(n10199), .B2(n10196), .ZN(
        P2_U3393) );
  OAI22_X1 U11216 ( .A1(n10143), .A2(n10162), .B1(n10142), .B2(n10183), .ZN(
        n10145) );
  NOR2_X1 U11217 ( .A1(n10145), .A2(n10144), .ZN(n10201) );
  AOI22_X1 U11218 ( .A1(n10198), .A2(n5342), .B1(n10201), .B2(n10196), .ZN(
        P2_U3396) );
  INV_X1 U11219 ( .A(n10146), .ZN(n10150) );
  OAI22_X1 U11220 ( .A1(n10148), .A2(n10190), .B1(n10147), .B2(n10183), .ZN(
        n10149) );
  NOR2_X1 U11221 ( .A1(n10150), .A2(n10149), .ZN(n10202) );
  AOI22_X1 U11222 ( .A1(n10198), .A2(n5371), .B1(n10202), .B2(n10196), .ZN(
        P2_U3402) );
  INV_X1 U11223 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11224 ( .A1(n10152), .A2(n10181), .B1(n10195), .B2(n10151), .ZN(
        n10153) );
  AND2_X1 U11225 ( .A1(n10154), .A2(n10153), .ZN(n10203) );
  AOI22_X1 U11226 ( .A1(n10198), .A2(n10155), .B1(n10203), .B2(n10196), .ZN(
        P2_U3405) );
  OAI21_X1 U11227 ( .B1(n10157), .B2(n10183), .A(n10156), .ZN(n10158) );
  AOI21_X1 U11228 ( .B1(n10159), .B2(n10188), .A(n10158), .ZN(n10204) );
  AOI22_X1 U11229 ( .A1(n10198), .A2(n5401), .B1(n10204), .B2(n10196), .ZN(
        P2_U3408) );
  INV_X1 U11230 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10166) );
  INV_X1 U11231 ( .A(n10160), .ZN(n10165) );
  OAI22_X1 U11232 ( .A1(n10163), .A2(n10162), .B1(n10161), .B2(n10183), .ZN(
        n10164) );
  NOR2_X1 U11233 ( .A1(n10165), .A2(n10164), .ZN(n10205) );
  AOI22_X1 U11234 ( .A1(n10198), .A2(n10166), .B1(n10205), .B2(n10196), .ZN(
        P2_U3411) );
  AOI22_X1 U11235 ( .A1(n10168), .A2(n10188), .B1(n10195), .B2(n10167), .ZN(
        n10169) );
  AND2_X1 U11236 ( .A1(n10170), .A2(n10169), .ZN(n10206) );
  AOI22_X1 U11237 ( .A1(n10198), .A2(n5436), .B1(n10206), .B2(n10196), .ZN(
        P2_U3414) );
  INV_X1 U11238 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U11239 ( .A1(n10172), .A2(n10181), .B1(n10195), .B2(n10171), .ZN(
        n10173) );
  AND2_X1 U11240 ( .A1(n10174), .A2(n10173), .ZN(n10207) );
  AOI22_X1 U11241 ( .A1(n10198), .A2(n10175), .B1(n10207), .B2(n10196), .ZN(
        P2_U3417) );
  INV_X1 U11242 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10182) );
  INV_X1 U11243 ( .A(n10176), .ZN(n10177) );
  NOR2_X1 U11244 ( .A1(n10177), .A2(n10183), .ZN(n10179) );
  AOI211_X1 U11245 ( .C1(n10181), .C2(n10180), .A(n10179), .B(n10178), .ZN(
        n10209) );
  AOI22_X1 U11246 ( .A1(n10198), .A2(n10182), .B1(n10209), .B2(n10196), .ZN(
        P2_U3420) );
  INV_X1 U11247 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10189) );
  NOR2_X1 U11248 ( .A1(n10184), .A2(n10183), .ZN(n10186) );
  AOI211_X1 U11249 ( .C1(n10188), .C2(n10187), .A(n10186), .B(n10185), .ZN(
        n10210) );
  AOI22_X1 U11250 ( .A1(n10198), .A2(n10189), .B1(n10210), .B2(n10196), .ZN(
        P2_U3423) );
  INV_X1 U11251 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10197) );
  NOR2_X1 U11252 ( .A1(n10191), .A2(n10190), .ZN(n10193) );
  AOI211_X1 U11253 ( .C1(n10195), .C2(n10194), .A(n10193), .B(n10192), .ZN(
        n10212) );
  AOI22_X1 U11254 ( .A1(n10198), .A2(n10197), .B1(n10212), .B2(n10196), .ZN(
        P2_U3426) );
  AOI22_X1 U11255 ( .A1(n10213), .A2(n10199), .B1(n5318), .B2(n10211), .ZN(
        P2_U3460) );
  AOI22_X1 U11256 ( .A1(n10213), .A2(n10201), .B1(n10200), .B2(n10211), .ZN(
        P2_U3461) );
  AOI22_X1 U11257 ( .A1(n10213), .A2(n10202), .B1(n6585), .B2(n10211), .ZN(
        P2_U3463) );
  AOI22_X1 U11258 ( .A1(n10213), .A2(n10203), .B1(n5383), .B2(n10211), .ZN(
        P2_U3464) );
  AOI22_X1 U11259 ( .A1(n10213), .A2(n10204), .B1(n5404), .B2(n10211), .ZN(
        P2_U3465) );
  AOI22_X1 U11260 ( .A1(n10213), .A2(n10205), .B1(n5418), .B2(n10211), .ZN(
        P2_U3466) );
  AOI22_X1 U11261 ( .A1(n10213), .A2(n10206), .B1(n6593), .B2(n10211), .ZN(
        P2_U3467) );
  AOI22_X1 U11262 ( .A1(n10213), .A2(n10207), .B1(n5445), .B2(n10211), .ZN(
        P2_U3468) );
  INV_X1 U11263 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U11264 ( .A1(n10213), .A2(n10209), .B1(n10208), .B2(n10211), .ZN(
        P2_U3469) );
  AOI22_X1 U11265 ( .A1(n10213), .A2(n10210), .B1(n5486), .B2(n10211), .ZN(
        P2_U3470) );
  AOI22_X1 U11266 ( .A1(n10213), .A2(n10212), .B1(n6624), .B2(n10211), .ZN(
        P2_U3471) );
  INV_X1 U11267 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10215) );
  NAND2_X1 U11268 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10214) );
  NOR2_X1 U11269 ( .A1(n10215), .A2(n10214), .ZN(n10217) );
  AOI21_X1 U11270 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U11271 ( .A1(n10217), .A2(n10219), .ZN(n10216) );
  XOR2_X1 U11272 ( .A(n10216), .B(P2_ADDR_REG_1__SCAN_IN), .Z(ADD_1068_U5) );
  XOR2_X1 U11273 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11274 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10269) );
  NOR2_X1 U11275 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10266) );
  NOR2_X1 U11276 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10263) );
  NOR2_X1 U11277 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10259) );
  NOR2_X1 U11278 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10255) );
  NOR2_X1 U11279 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10251) );
  NOR2_X1 U11280 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10247) );
  NOR2_X1 U11281 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10243) );
  NOR2_X1 U11282 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10239) );
  NOR2_X1 U11283 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10235) );
  NOR2_X1 U11284 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10231) );
  NOR2_X1 U11285 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10229) );
  NOR2_X1 U11286 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10227) );
  NOR2_X1 U11287 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10225) );
  NAND2_X1 U11288 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10223) );
  XOR2_X1 U11289 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10682) );
  NAND2_X1 U11290 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10221) );
  NOR2_X1 U11291 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10217), .ZN(n10218) );
  NOR2_X1 U11292 ( .A1(n10219), .A2(n10218), .ZN(n10672) );
  XOR2_X1 U11293 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10671) );
  NAND2_X1 U11294 ( .A1(n10672), .A2(n10671), .ZN(n10220) );
  NAND2_X1 U11295 ( .A1(n10221), .A2(n10220), .ZN(n10681) );
  NAND2_X1 U11296 ( .A1(n10682), .A2(n10681), .ZN(n10222) );
  NAND2_X1 U11297 ( .A1(n10223), .A2(n10222), .ZN(n10684) );
  XNOR2_X1 U11298 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10683) );
  NOR2_X1 U11299 ( .A1(n10684), .A2(n10683), .ZN(n10224) );
  NOR2_X1 U11300 ( .A1(n10225), .A2(n10224), .ZN(n10674) );
  XNOR2_X1 U11301 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10673) );
  NOR2_X1 U11302 ( .A1(n10674), .A2(n10673), .ZN(n10226) );
  NOR2_X1 U11303 ( .A1(n10227), .A2(n10226), .ZN(n10680) );
  XNOR2_X1 U11304 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10679) );
  NOR2_X1 U11305 ( .A1(n10680), .A2(n10679), .ZN(n10228) );
  NOR2_X1 U11306 ( .A1(n10229), .A2(n10228), .ZN(n10676) );
  XNOR2_X1 U11307 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10675) );
  NOR2_X1 U11308 ( .A1(n10676), .A2(n10675), .ZN(n10230) );
  NOR2_X1 U11309 ( .A1(n10231), .A2(n10230), .ZN(n10678) );
  INV_X1 U11310 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U11311 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10233), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10232), .ZN(n10677) );
  NOR2_X1 U11312 ( .A1(n10678), .A2(n10677), .ZN(n10234) );
  NOR2_X1 U11313 ( .A1(n10235), .A2(n10234), .ZN(n10670) );
  INV_X1 U11314 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U11315 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10237), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10236), .ZN(n10669) );
  NOR2_X1 U11316 ( .A1(n10670), .A2(n10669), .ZN(n10238) );
  NOR2_X1 U11317 ( .A1(n10239), .A2(n10238), .ZN(n10288) );
  INV_X1 U11318 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U11319 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10241), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10240), .ZN(n10287) );
  NOR2_X1 U11320 ( .A1(n10288), .A2(n10287), .ZN(n10242) );
  NOR2_X1 U11321 ( .A1(n10243), .A2(n10242), .ZN(n10286) );
  INV_X1 U11322 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10245) );
  INV_X1 U11323 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U11324 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10245), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10244), .ZN(n10285) );
  NOR2_X1 U11325 ( .A1(n10286), .A2(n10285), .ZN(n10246) );
  NOR2_X1 U11326 ( .A1(n10247), .A2(n10246), .ZN(n10284) );
  INV_X1 U11327 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U11328 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10249), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10248), .ZN(n10283) );
  NOR2_X1 U11329 ( .A1(n10284), .A2(n10283), .ZN(n10250) );
  NOR2_X1 U11330 ( .A1(n10251), .A2(n10250), .ZN(n10282) );
  INV_X1 U11331 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U11332 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10253), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10252), .ZN(n10281) );
  NOR2_X1 U11333 ( .A1(n10282), .A2(n10281), .ZN(n10254) );
  NOR2_X1 U11334 ( .A1(n10255), .A2(n10254), .ZN(n10280) );
  INV_X1 U11335 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U11336 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n10257), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n10256), .ZN(n10279) );
  NOR2_X1 U11337 ( .A1(n10280), .A2(n10279), .ZN(n10258) );
  NOR2_X1 U11338 ( .A1(n10259), .A2(n10258), .ZN(n10278) );
  INV_X1 U11339 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U11340 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n10261), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10260), .ZN(n10277) );
  NOR2_X1 U11341 ( .A1(n10278), .A2(n10277), .ZN(n10262) );
  NOR2_X1 U11342 ( .A1(n10263), .A2(n10262), .ZN(n10276) );
  AOI22_X1 U11343 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9503), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n10264), .ZN(n10275) );
  NOR2_X1 U11344 ( .A1(n10276), .A2(n10275), .ZN(n10265) );
  NOR2_X1 U11345 ( .A1(n10266), .A2(n10265), .ZN(n10274) );
  AOI22_X1 U11346 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9519), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10267), .ZN(n10273) );
  NOR2_X1 U11347 ( .A1(n10274), .A2(n10273), .ZN(n10268) );
  NOR2_X1 U11348 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  AND2_X1 U11349 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10270), .ZN(n10289) );
  NOR2_X1 U11350 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10270), .ZN(n10291) );
  NOR2_X1 U11351 ( .A1(n10289), .A2(n10291), .ZN(n10272) );
  XNOR2_X1 U11352 ( .A(n10272), .B(n10271), .ZN(ADD_1068_U55) );
  XNOR2_X1 U11353 ( .A(n10274), .B(n10273), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11354 ( .A(n10276), .B(n10275), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11355 ( .A(n10278), .B(n10277), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11356 ( .A(n10280), .B(n10279), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11357 ( .A(n10282), .B(n10281), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11358 ( .A(n10284), .B(n10283), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11359 ( .A(n10286), .B(n10285), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11360 ( .A(n10288), .B(n10287), .ZN(ADD_1068_U63) );
  NOR2_X1 U11361 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10289), .ZN(n10290) );
  NOR2_X1 U11362 ( .A1(n10291), .A2(n10290), .ZN(n10668) );
  XNOR2_X1 U11363 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10666) );
  INV_X1 U11364 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10664) );
  XNOR2_X1 U11365 ( .A(keyinput_g43), .B(n10566), .ZN(n10298) );
  AOI22_X1 U11366 ( .A1(SI_31_), .A2(keyinput_g1), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .ZN(n10292) );
  OAI221_X1 U11367 ( .B1(SI_31_), .B2(keyinput_g1), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_g82), .A(n10292), .ZN(n10297)
         );
  AOI22_X1 U11368 ( .A1(SI_15_), .A2(keyinput_g17), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n10293) );
  OAI221_X1 U11369 ( .B1(SI_15_), .B2(keyinput_g17), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n10293), .ZN(n10296)
         );
  AOI22_X1 U11370 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_g118), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_g106), .ZN(n10294) );
  OAI221_X1 U11371 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_g118), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_g106), .A(n10294), .ZN(n10295) );
  NOR4_X1 U11372 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10326) );
  AOI22_X1 U11373 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        SI_22_), .B2(keyinput_g10), .ZN(n10299) );
  OAI221_X1 U11374 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        SI_22_), .C2(keyinput_g10), .A(n10299), .ZN(n10306) );
  AOI22_X1 U11375 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n10300) );
  OAI221_X1 U11376 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n10300), .ZN(n10305)
         );
  AOI22_X1 U11377 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n10301) );
  OAI221_X1 U11378 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n10301), .ZN(n10304)
         );
  AOI22_X1 U11379 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .ZN(n10302) );
  OAI221_X1 U11380 ( .B1(SI_4_), .B2(keyinput_g28), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput_g87), .A(n10302), .ZN(n10303)
         );
  NOR4_X1 U11381 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10325) );
  AOI22_X1 U11382 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_g90), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_g101), .ZN(n10307) );
  OAI221_X1 U11383 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_g90), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_g101), .A(n10307), .ZN(n10314) );
  AOI22_X1 U11384 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_g102), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .ZN(n10308) );
  OAI221_X1 U11385 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_g102), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput_g67), .A(n10308), .ZN(n10313)
         );
  AOI22_X1 U11386 ( .A1(SI_21_), .A2(keyinput_g11), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n10309) );
  OAI221_X1 U11387 ( .B1(SI_21_), .B2(keyinput_g11), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n10309), .ZN(n10312)
         );
  AOI22_X1 U11388 ( .A1(SI_18_), .A2(keyinput_g14), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_g73), .ZN(n10310) );
  OAI221_X1 U11389 ( .B1(SI_18_), .B2(keyinput_g14), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput_g73), .A(n10310), .ZN(n10311)
         );
  NOR4_X1 U11390 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10324) );
  AOI22_X1 U11391 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput_g127), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_g94), .ZN(n10315) );
  OAI221_X1 U11392 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput_g127), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_g94), .A(n10315), .ZN(n10322) );
  AOI22_X1 U11393 ( .A1(SI_2_), .A2(keyinput_g30), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .ZN(n10316) );
  OAI221_X1 U11394 ( .B1(SI_2_), .B2(keyinput_g30), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n10316), .ZN(n10321)
         );
  AOI22_X1 U11395 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput_g77), .B1(
        SI_20_), .B2(keyinput_g12), .ZN(n10317) );
  OAI221_X1 U11396 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_g77), .C1(
        SI_20_), .C2(keyinput_g12), .A(n10317), .ZN(n10320) );
  AOI22_X1 U11397 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(SI_16_), 
        .B2(keyinput_g16), .ZN(n10318) );
  OAI221_X1 U11398 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(SI_16_), 
        .C2(keyinput_g16), .A(n10318), .ZN(n10319) );
  NOR4_X1 U11399 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10323) );
  NAND4_X1 U11400 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10471) );
  AOI22_X1 U11401 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g93), .B1(SI_10_), 
        .B2(keyinput_g22), .ZN(n10327) );
  OAI221_X1 U11402 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g93), .C1(SI_10_), 
        .C2(keyinput_g22), .A(n10327), .ZN(n10334) );
  AOI22_X1 U11403 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_g96), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .ZN(n10328) );
  OAI221_X1 U11404 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_g96), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_g84), .A(n10328), .ZN(n10333)
         );
  AOI22_X1 U11405 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_g120), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n10329) );
  OAI221_X1 U11406 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_g120), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n10329), .ZN(n10332)
         );
  AOI22_X1 U11407 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_g107), .B1(SI_24_), .B2(keyinput_g8), .ZN(n10330) );
  OAI221_X1 U11408 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_g107), .C1(
        SI_24_), .C2(keyinput_g8), .A(n10330), .ZN(n10331) );
  NOR4_X1 U11409 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10363) );
  AOI22_X1 U11410 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_g125), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_g104), .ZN(n10335) );
  OAI221_X1 U11411 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_g125), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_g104), .A(n10335), .ZN(n10342) );
  AOI22_X1 U11412 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n10336) );
  OAI221_X1 U11413 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n10336), .ZN(n10341) );
  AOI22_X1 U11414 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_g95), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput_g99), .ZN(n10337) );
  OAI221_X1 U11415 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_g95), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_g99), .A(n10337), .ZN(n10340) );
  AOI22_X1 U11416 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g92), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n10338) );
  OAI221_X1 U11417 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g92), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n10338), .ZN(n10339)
         );
  NOR4_X1 U11418 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10362) );
  AOI22_X1 U11419 ( .A1(SI_23_), .A2(keyinput_g9), .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n10343) );
  OAI221_X1 U11420 ( .B1(SI_23_), .B2(keyinput_g9), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n10343), .ZN(n10350)
         );
  AOI22_X1 U11421 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_g117), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n10344) );
  OAI221_X1 U11422 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_g117), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n10344), .ZN(n10349)
         );
  AOI22_X1 U11423 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_g115), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .ZN(n10345) );
  OAI221_X1 U11424 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_g115), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_g76), .A(n10345), .ZN(n10348)
         );
  AOI22_X1 U11425 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_g121), .B1(SI_17_), .B2(keyinput_g15), .ZN(n10346) );
  OAI221_X1 U11426 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_g121), .C1(
        SI_17_), .C2(keyinput_g15), .A(n10346), .ZN(n10347) );
  NOR4_X1 U11427 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10361) );
  AOI22_X1 U11428 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n10351) );
  OAI221_X1 U11429 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n10351), .ZN(n10359)
         );
  AOI22_X1 U11430 ( .A1(SI_3_), .A2(keyinput_g29), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_g53), .ZN(n10352) );
  OAI221_X1 U11431 ( .B1(SI_3_), .B2(keyinput_g29), .C1(P2_REG3_REG_9__SCAN_IN), .C2(keyinput_g53), .A(n10352), .ZN(n10358) );
  AOI22_X1 U11432 ( .A1(SI_9_), .A2(keyinput_g23), .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n10353) );
  OAI221_X1 U11433 ( .B1(SI_9_), .B2(keyinput_g23), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n10353), .ZN(n10357)
         );
  XNOR2_X1 U11434 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g110), .ZN(n10355)
         );
  XNOR2_X1 U11435 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_g52), .ZN(n10354)
         );
  NAND2_X1 U11436 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  NOR4_X1 U11437 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10360) );
  NAND4_X1 U11438 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10470) );
  AOI22_X1 U11439 ( .A1(n10366), .A2(keyinput_g79), .B1(keyinput_g25), .B2(
        n10365), .ZN(n10364) );
  OAI221_X1 U11440 ( .B1(n10366), .B2(keyinput_g79), .C1(n10365), .C2(
        keyinput_g25), .A(n10364), .ZN(n10370) );
  XNOR2_X1 U11441 ( .A(n10367), .B(keyinput_g126), .ZN(n10369) );
  XOR2_X1 U11442 ( .A(SI_0_), .B(keyinput_g32), .Z(n10368) );
  OR3_X1 U11443 ( .A1(n10370), .A2(n10369), .A3(n10368), .ZN(n10377) );
  INV_X1 U11444 ( .A(SI_30_), .ZN(n10372) );
  AOI22_X1 U11445 ( .A1(n10372), .A2(keyinput_g2), .B1(n5218), .B2(
        keyinput_g20), .ZN(n10371) );
  OAI221_X1 U11446 ( .B1(n10372), .B2(keyinput_g2), .C1(n5218), .C2(
        keyinput_g20), .A(n10371), .ZN(n10376) );
  AOI22_X1 U11447 ( .A1(n10374), .A2(keyinput_g80), .B1(n8409), .B2(
        keyinput_g47), .ZN(n10373) );
  OAI221_X1 U11448 ( .B1(n10374), .B2(keyinput_g80), .C1(n8409), .C2(
        keyinput_g47), .A(n10373), .ZN(n10375) );
  NOR3_X1 U11449 ( .A1(n10377), .A2(n10376), .A3(n10375), .ZN(n10416) );
  INV_X1 U11450 ( .A(SI_13_), .ZN(n10581) );
  AOI22_X1 U11451 ( .A1(n10379), .A2(keyinput_g78), .B1(keyinput_g19), .B2(
        n10581), .ZN(n10378) );
  OAI221_X1 U11452 ( .B1(n10379), .B2(keyinput_g78), .C1(n10581), .C2(
        keyinput_g19), .A(n10378), .ZN(n10388) );
  INV_X1 U11453 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U11454 ( .A1(n5858), .A2(keyinput_g109), .B1(n10381), .B2(
        keyinput_g38), .ZN(n10380) );
  OAI221_X1 U11455 ( .B1(n5858), .B2(keyinput_g109), .C1(n10381), .C2(
        keyinput_g38), .A(n10380), .ZN(n10387) );
  XNOR2_X1 U11456 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_g68), .ZN(n10385) );
  XNOR2_X1 U11457 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_g100), .ZN(n10384)
         );
  XNOR2_X1 U11458 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g91), .ZN(n10383) );
  XNOR2_X1 U11459 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n10382)
         );
  NAND4_X1 U11460 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10386) );
  NOR3_X1 U11461 ( .A1(n10388), .A2(n10387), .A3(n10386), .ZN(n10415) );
  AOI22_X1 U11462 ( .A1(n10390), .A2(keyinput_g39), .B1(keyinput_g111), .B2(
        n5868), .ZN(n10389) );
  INV_X1 U11463 ( .A(SI_14_), .ZN(n10392) );
  AOI22_X1 U11464 ( .A1(n10392), .A2(keyinput_g18), .B1(n10584), .B2(
        keyinput_g71), .ZN(n10391) );
  OAI221_X1 U11465 ( .B1(n10392), .B2(keyinput_g18), .C1(n10584), .C2(
        keyinput_g71), .A(n10391), .ZN(n10399) );
  INV_X1 U11466 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U11467 ( .A1(n10565), .A2(keyinput_g98), .B1(n10394), .B2(
        keyinput_g81), .ZN(n10393) );
  OAI221_X1 U11468 ( .B1(n10565), .B2(keyinput_g98), .C1(n10394), .C2(
        keyinput_g81), .A(n10393), .ZN(n10398) );
  INV_X1 U11469 ( .A(P2_B_REG_SCAN_IN), .ZN(n10396) );
  AOI22_X1 U11470 ( .A1(n6447), .A2(keyinput_g113), .B1(n10396), .B2(
        keyinput_g64), .ZN(n10395) );
  OAI221_X1 U11471 ( .B1(n6447), .B2(keyinput_g113), .C1(n10396), .C2(
        keyinput_g64), .A(n10395), .ZN(n10397) );
  NOR4_X1 U11472 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10414) );
  INV_X1 U11473 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U11474 ( .A1(n10402), .A2(keyinput_g66), .B1(n10559), .B2(
        keyinput_g103), .ZN(n10401) );
  OAI221_X1 U11475 ( .B1(n10402), .B2(keyinput_g66), .C1(n10559), .C2(
        keyinput_g103), .A(n10401), .ZN(n10412) );
  AOI22_X1 U11476 ( .A1(n6444), .A2(keyinput_g112), .B1(keyinput_g124), .B2(
        n10404), .ZN(n10403) );
  OAI221_X1 U11477 ( .B1(n6444), .B2(keyinput_g112), .C1(n10404), .C2(
        keyinput_g124), .A(n10403), .ZN(n10411) );
  INV_X1 U11478 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U11479 ( .A1(n10555), .A2(keyinput_g116), .B1(n10617), .B2(
        keyinput_g69), .ZN(n10405) );
  OAI221_X1 U11480 ( .B1(n10555), .B2(keyinput_g116), .C1(n10617), .C2(
        keyinput_g69), .A(n10405), .ZN(n10410) );
  AOI22_X1 U11481 ( .A1(n10408), .A2(keyinput_g21), .B1(keyinput_g89), .B2(
        n10407), .ZN(n10406) );
  OAI221_X1 U11482 ( .B1(n10408), .B2(keyinput_g21), .C1(n10407), .C2(
        keyinput_g89), .A(n10406), .ZN(n10409) );
  NOR4_X1 U11483 ( .A1(n10412), .A2(n10411), .A3(n10410), .A4(n10409), .ZN(
        n10413) );
  NAND4_X1 U11484 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10469) );
  AOI22_X1 U11485 ( .A1(n10575), .A2(keyinput_g13), .B1(n10418), .B2(
        keyinput_g72), .ZN(n10417) );
  OAI221_X1 U11486 ( .B1(n10575), .B2(keyinput_g13), .C1(n10418), .C2(
        keyinput_g72), .A(n10417), .ZN(n10428) );
  AOI22_X1 U11487 ( .A1(n10421), .A2(keyinput_g6), .B1(n10420), .B2(
        keyinput_g4), .ZN(n10419) );
  OAI221_X1 U11488 ( .B1(n10421), .B2(keyinput_g6), .C1(n10420), .C2(
        keyinput_g4), .A(n10419), .ZN(n10427) );
  AOI22_X1 U11489 ( .A1(n10611), .A2(keyinput_g123), .B1(n5385), .B2(
        keyinput_g49), .ZN(n10422) );
  OAI221_X1 U11490 ( .B1(n10611), .B2(keyinput_g123), .C1(n5385), .C2(
        keyinput_g49), .A(n10422), .ZN(n10426) );
  AOI22_X1 U11491 ( .A1(n10601), .A2(keyinput_g122), .B1(n10424), .B2(
        keyinput_g70), .ZN(n10423) );
  OAI221_X1 U11492 ( .B1(n10601), .B2(keyinput_g122), .C1(n10424), .C2(
        keyinput_g70), .A(n10423), .ZN(n10425) );
  NOR4_X1 U11493 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .ZN(
        n10467) );
  AOI22_X1 U11494 ( .A1(n10605), .A2(keyinput_g83), .B1(keyinput_g44), .B2(
        n8209), .ZN(n10429) );
  OAI221_X1 U11495 ( .B1(n10605), .B2(keyinput_g83), .C1(n8209), .C2(
        keyinput_g44), .A(n10429), .ZN(n10438) );
  INV_X1 U11496 ( .A(SI_5_), .ZN(n10558) );
  AOI22_X1 U11497 ( .A1(n10431), .A2(keyinput_g5), .B1(keyinput_g27), .B2(
        n10558), .ZN(n10430) );
  OAI221_X1 U11498 ( .B1(n10431), .B2(keyinput_g5), .C1(n10558), .C2(
        keyinput_g27), .A(n10430), .ZN(n10437) );
  XNOR2_X1 U11499 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_g51), .ZN(n10435)
         );
  XNOR2_X1 U11500 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g108), .ZN(n10434)
         );
  XNOR2_X1 U11501 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10433) );
  XNOR2_X1 U11502 ( .A(SI_8_), .B(keyinput_g24), .ZN(n10432) );
  NAND4_X1 U11503 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        n10436) );
  NOR3_X1 U11504 ( .A1(n10438), .A2(n10437), .A3(n10436), .ZN(n10466) );
  AOI22_X1 U11505 ( .A1(n10441), .A2(keyinput_g45), .B1(keyinput_g33), .B2(
        n10440), .ZN(n10439) );
  OAI221_X1 U11506 ( .B1(n10441), .B2(keyinput_g45), .C1(n10440), .C2(
        keyinput_g33), .A(n10439), .ZN(n10450) );
  AOI22_X1 U11507 ( .A1(n5902), .A2(keyinput_g119), .B1(n10443), .B2(
        keyinput_g35), .ZN(n10442) );
  OAI221_X1 U11508 ( .B1(n5902), .B2(keyinput_g119), .C1(n10443), .C2(
        keyinput_g35), .A(n10442), .ZN(n10449) );
  AOI22_X1 U11509 ( .A1(n7276), .A2(keyinput_g59), .B1(n5717), .B2(keyinput_g3), .ZN(n10444) );
  OAI221_X1 U11510 ( .B1(n7276), .B2(keyinput_g59), .C1(n5717), .C2(
        keyinput_g3), .A(n10444), .ZN(n10448) );
  XNOR2_X1 U11511 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_g114), .ZN(n10446)
         );
  XNOR2_X1 U11512 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_g74), .ZN(n10445) );
  NAND2_X1 U11513 ( .A1(n10446), .A2(n10445), .ZN(n10447) );
  NOR4_X1 U11514 ( .A1(n10450), .A2(n10449), .A3(n10448), .A4(n10447), .ZN(
        n10465) );
  AOI22_X1 U11515 ( .A1(n10633), .A2(keyinput_g40), .B1(n10452), .B2(
        keyinput_g50), .ZN(n10451) );
  OAI221_X1 U11516 ( .B1(n10633), .B2(keyinput_g40), .C1(n10452), .C2(
        keyinput_g50), .A(n10451), .ZN(n10463) );
  AOI22_X1 U11517 ( .A1(n10455), .A2(keyinput_g65), .B1(n10454), .B2(
        keyinput_g26), .ZN(n10453) );
  OAI221_X1 U11518 ( .B1(n10455), .B2(keyinput_g65), .C1(n10454), .C2(
        keyinput_g26), .A(n10453), .ZN(n10462) );
  AOI22_X1 U11519 ( .A1(n10457), .A2(keyinput_g85), .B1(n10602), .B2(
        keyinput_g62), .ZN(n10456) );
  OAI221_X1 U11520 ( .B1(n10457), .B2(keyinput_g85), .C1(n10602), .C2(
        keyinput_g62), .A(n10456), .ZN(n10461) );
  XNOR2_X1 U11521 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g97), .ZN(n10459) );
  XNOR2_X1 U11522 ( .A(SI_25_), .B(keyinput_g7), .ZN(n10458) );
  NAND2_X1 U11523 ( .A1(n10459), .A2(n10458), .ZN(n10460) );
  NOR4_X1 U11524 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10464) );
  NAND4_X1 U11525 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n10468) );
  NOR4_X1 U11526 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .ZN(
        n10663) );
  XOR2_X1 U11527 ( .A(SI_1_), .B(keyinput_f31), .Z(n10478) );
  AOI22_X1 U11528 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_f89), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .ZN(n10472) );
  OAI221_X1 U11529 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n10472), .ZN(n10477) );
  AOI22_X1 U11530 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_f113), .B1(SI_2_), 
        .B2(keyinput_f30), .ZN(n10473) );
  OAI221_X1 U11531 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_f113), .C1(SI_2_), .C2(keyinput_f30), .A(n10473), .ZN(n10476) );
  AOI22_X1 U11532 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_f124), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .ZN(n10474) );
  OAI221_X1 U11533 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_f124), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_f77), .A(n10474), .ZN(n10475)
         );
  NOR4_X1 U11534 ( .A1(n10478), .A2(n10477), .A3(n10476), .A4(n10475), .ZN(
        n10506) );
  AOI22_X1 U11535 ( .A1(SI_6_), .A2(keyinput_f26), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_f81), .ZN(n10479) );
  OAI221_X1 U11536 ( .B1(SI_6_), .B2(keyinput_f26), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_f81), .A(n10479), .ZN(n10486)
         );
  AOI22_X1 U11537 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_f112), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n10480) );
  OAI221_X1 U11538 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_f112), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n10480), .ZN(n10485)
         );
  AOI22_X1 U11539 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_f109), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n10481) );
  OAI221_X1 U11540 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_f109), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n10481), .ZN(n10484)
         );
  AOI22_X1 U11541 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_f125), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n10482) );
  OAI221_X1 U11542 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_f125), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_f56), .A(n10482), .ZN(n10483)
         );
  NOR4_X1 U11543 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10505) );
  AOI22_X1 U11544 ( .A1(SI_30_), .A2(keyinput_f2), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .ZN(n10487) );
  OAI221_X1 U11545 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput_f73), .A(n10487), .ZN(n10494)
         );
  AOI22_X1 U11546 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_f97), .B1(
        P2_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n10488) );
  OAI221_X1 U11547 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_f97), .C1(
        P2_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n10488), .ZN(n10493) );
  AOI22_X1 U11548 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_f99), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .ZN(n10489) );
  OAI221_X1 U11549 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_f99), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_f70), .A(n10489), .ZN(n10492)
         );
  AOI22_X1 U11550 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_f114), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput_f121), .ZN(n10490) );
  OAI221_X1 U11551 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_f114), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput_f121), .A(n10490), .ZN(n10491) );
  NOR4_X1 U11552 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10504) );
  AOI22_X1 U11553 ( .A1(SI_0_), .A2(keyinput_f32), .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n10495) );
  OAI221_X1 U11554 ( .B1(SI_0_), .B2(keyinput_f32), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n10495), .ZN(n10502)
         );
  AOI22_X1 U11555 ( .A1(SI_27_), .A2(keyinput_f5), .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n10496) );
  OAI221_X1 U11556 ( .B1(SI_27_), .B2(keyinput_f5), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n10496), .ZN(n10501)
         );
  AOI22_X1 U11557 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_f95), .B1(SI_29_), 
        .B2(keyinput_f3), .ZN(n10497) );
  OAI221_X1 U11558 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_f95), .C1(SI_29_), 
        .C2(keyinput_f3), .A(n10497), .ZN(n10500) );
  AOI22_X1 U11559 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_f106), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput_f96), .ZN(n10498) );
  OAI221_X1 U11560 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_f106), .C1(
        P1_IR_REG_6__SCAN_IN), .C2(keyinput_f96), .A(n10498), .ZN(n10499) );
  NOR4_X1 U11561 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10503) );
  NAND4_X1 U11562 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10659) );
  AOI22_X1 U11563 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f118), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n10507) );
  OAI221_X1 U11564 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f118), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n10507), .ZN(n10514)
         );
  AOI22_X1 U11565 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_f80), .B1(
        SI_18_), .B2(keyinput_f14), .ZN(n10508) );
  OAI221_X1 U11566 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .C1(
        SI_18_), .C2(keyinput_f14), .A(n10508), .ZN(n10513) );
  AOI22_X1 U11567 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_f67), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n10509) );
  OAI221_X1 U11568 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n10509), .ZN(n10512) );
  AOI22_X1 U11569 ( .A1(SI_11_), .A2(keyinput_f21), .B1(SI_15_), .B2(
        keyinput_f17), .ZN(n10510) );
  OAI221_X1 U11570 ( .B1(SI_11_), .B2(keyinput_f21), .C1(SI_15_), .C2(
        keyinput_f17), .A(n10510), .ZN(n10511) );
  NOR4_X1 U11571 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n10542) );
  AOI22_X1 U11572 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f101), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n10515) );
  OAI221_X1 U11573 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f101), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n10515), .ZN(n10522) );
  AOI22_X1 U11574 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n10516) );
  OAI221_X1 U11575 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n10516), .ZN(n10521)
         );
  AOI22_X1 U11576 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_f90), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n10517) );
  OAI221_X1 U11577 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_f90), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n10517), .ZN(n10520)
         );
  AOI22_X1 U11578 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_f87), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .ZN(n10518) );
  OAI221_X1 U11579 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n10518), .ZN(n10519) );
  NOR4_X1 U11580 ( .A1(n10522), .A2(n10521), .A3(n10520), .A4(n10519), .ZN(
        n10541) );
  AOI22_X1 U11581 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_f126), .B1(SI_26_), 
        .B2(keyinput_f6), .ZN(n10523) );
  OAI221_X1 U11582 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_f126), .C1(SI_26_), 
        .C2(keyinput_f6), .A(n10523), .ZN(n10530) );
  AOI22_X1 U11583 ( .A1(SI_14_), .A2(keyinput_f18), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .ZN(n10524) );
  OAI221_X1 U11584 ( .B1(SI_14_), .B2(keyinput_f18), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput_f72), .A(n10524), .ZN(n10529)
         );
  AOI22_X1 U11585 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .ZN(n10525) );
  OAI221_X1 U11586 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_f85), .A(n10525), .ZN(n10528)
         );
  AOI22_X1 U11587 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_f111), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .ZN(n10526) );
  OAI221_X1 U11588 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_f111), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_f84), .A(n10526), .ZN(n10527)
         );
  NOR4_X1 U11589 ( .A1(n10530), .A2(n10529), .A3(n10528), .A4(n10527), .ZN(
        n10540) );
  AOI22_X1 U11590 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_f79), .ZN(n10531) );
  OAI221_X1 U11591 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_f79), .A(n10531), .ZN(n10538)
         );
  AOI22_X1 U11592 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_f86), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n10532) );
  OAI221_X1 U11593 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n10532), .ZN(n10537)
         );
  AOI22_X1 U11594 ( .A1(SI_12_), .A2(keyinput_f20), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_f78), .ZN(n10533) );
  OAI221_X1 U11595 ( .B1(SI_12_), .B2(keyinput_f20), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput_f78), .A(n10533), .ZN(n10536)
         );
  AOI22_X1 U11596 ( .A1(SI_28_), .A2(keyinput_f4), .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n10534) );
  OAI221_X1 U11597 ( .B1(SI_28_), .B2(keyinput_f4), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n10534), .ZN(n10535)
         );
  NOR4_X1 U11598 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10539) );
  NAND4_X1 U11599 ( .A1(n10542), .A2(n10541), .A3(n10540), .A4(n10539), .ZN(
        n10658) );
  AOI22_X1 U11600 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .ZN(n10543) );
  OAI221_X1 U11601 ( .B1(SI_31_), .B2(keyinput_f1), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n10543), .ZN(n10550)
         );
  AOI22_X1 U11602 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_f104), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_f102), .ZN(n10544) );
  OAI221_X1 U11603 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_f104), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_f102), .A(n10544), .ZN(n10549) );
  AOI22_X1 U11604 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_f94), .B1(SI_25_), 
        .B2(keyinput_f7), .ZN(n10545) );
  OAI221_X1 U11605 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_f94), .C1(SI_25_), 
        .C2(keyinput_f7), .A(n10545), .ZN(n10548) );
  AOI22_X1 U11606 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P2_STATE_REG_SCAN_IN), 
        .B2(keyinput_f34), .ZN(n10546) );
  OAI221_X1 U11607 ( .B1(SI_7_), .B2(keyinput_f25), .C1(P2_STATE_REG_SCAN_IN), 
        .C2(keyinput_f34), .A(n10546), .ZN(n10547) );
  NOR4_X1 U11608 ( .A1(n10550), .A2(n10549), .A3(n10548), .A4(n10547), .ZN(
        n10596) );
  AOI22_X1 U11609 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .ZN(n10551) );
  OAI221_X1 U11610 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_f76), .A(n10551), .ZN(n10563)
         );
  AOI22_X1 U11611 ( .A1(SI_10_), .A2(keyinput_f22), .B1(n10553), .B2(
        keyinput_f8), .ZN(n10552) );
  OAI221_X1 U11612 ( .B1(SI_10_), .B2(keyinput_f22), .C1(n10553), .C2(
        keyinput_f8), .A(n10552), .ZN(n10562) );
  INV_X1 U11613 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U11614 ( .A1(n10556), .A2(keyinput_f37), .B1(keyinput_f116), .B2(
        n10555), .ZN(n10554) );
  OAI221_X1 U11615 ( .B1(n10556), .B2(keyinput_f37), .C1(n10555), .C2(
        keyinput_f116), .A(n10554), .ZN(n10561) );
  AOI22_X1 U11616 ( .A1(n10559), .A2(keyinput_f103), .B1(n10558), .B2(
        keyinput_f27), .ZN(n10557) );
  OAI221_X1 U11617 ( .B1(n10559), .B2(keyinput_f103), .C1(n10558), .C2(
        keyinput_f27), .A(n10557), .ZN(n10560) );
  NOR4_X1 U11618 ( .A1(n10563), .A2(n10562), .A3(n10561), .A4(n10560), .ZN(
        n10595) );
  AOI22_X1 U11619 ( .A1(n10566), .A2(keyinput_f43), .B1(keyinput_f98), .B2(
        n10565), .ZN(n10564) );
  OAI221_X1 U11620 ( .B1(n10566), .B2(keyinput_f43), .C1(n10565), .C2(
        keyinput_f98), .A(n10564), .ZN(n10573) );
  AOI22_X1 U11621 ( .A1(n10569), .A2(keyinput_f68), .B1(keyinput_f15), .B2(
        n10568), .ZN(n10567) );
  OAI221_X1 U11622 ( .B1(n10569), .B2(keyinput_f68), .C1(n10568), .C2(
        keyinput_f15), .A(n10567), .ZN(n10572) );
  XNOR2_X1 U11623 ( .A(n10570), .B(keyinput_f29), .ZN(n10571) );
  OR3_X1 U11624 ( .A1(n10573), .A2(n10572), .A3(n10571), .ZN(n10579) );
  AOI22_X1 U11625 ( .A1(n10575), .A2(keyinput_f13), .B1(keyinput_f59), .B2(
        n7276), .ZN(n10574) );
  OAI221_X1 U11626 ( .B1(n10575), .B2(keyinput_f13), .C1(n7276), .C2(
        keyinput_f59), .A(n10574), .ZN(n10578) );
  XNOR2_X1 U11627 ( .A(n10576), .B(keyinput_f127), .ZN(n10577) );
  NOR3_X1 U11628 ( .A1(n10579), .A2(n10578), .A3(n10577), .ZN(n10594) );
  INV_X1 U11629 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U11630 ( .A1(n10582), .A2(keyinput_f51), .B1(keyinput_f19), .B2(
        n10581), .ZN(n10580) );
  OAI221_X1 U11631 ( .B1(n10582), .B2(keyinput_f51), .C1(n10581), .C2(
        keyinput_f19), .A(n10580), .ZN(n10592) );
  AOI22_X1 U11632 ( .A1(n10585), .A2(keyinput_f9), .B1(n10584), .B2(
        keyinput_f71), .ZN(n10583) );
  OAI221_X1 U11633 ( .B1(n10585), .B2(keyinput_f9), .C1(n10584), .C2(
        keyinput_f71), .A(n10583), .ZN(n10591) );
  XOR2_X1 U11634 ( .A(n10440), .B(keyinput_f33), .Z(n10589) );
  XNOR2_X1 U11635 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_f88), .ZN(n10588)
         );
  XNOR2_X1 U11636 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_f92), .ZN(n10587) );
  XNOR2_X1 U11637 ( .A(SI_4_), .B(keyinput_f28), .ZN(n10586) );
  NAND4_X1 U11638 ( .A1(n10589), .A2(n10588), .A3(n10587), .A4(n10586), .ZN(
        n10590) );
  NOR3_X1 U11639 ( .A1(n10592), .A2(n10591), .A3(n10590), .ZN(n10593) );
  NAND4_X1 U11640 ( .A1(n10596), .A2(n10595), .A3(n10594), .A4(n10593), .ZN(
        n10657) );
  INV_X1 U11641 ( .A(SI_21_), .ZN(n10598) );
  AOI22_X1 U11642 ( .A1(n10599), .A2(keyinput_f12), .B1(n10598), .B2(
        keyinput_f11), .ZN(n10597) );
  OAI221_X1 U11643 ( .B1(n10599), .B2(keyinput_f12), .C1(n10598), .C2(
        keyinput_f11), .A(n10597), .ZN(n10610) );
  AOI22_X1 U11644 ( .A1(n10602), .A2(keyinput_f62), .B1(keyinput_f122), .B2(
        n10601), .ZN(n10600) );
  OAI221_X1 U11645 ( .B1(n10602), .B2(keyinput_f62), .C1(n10601), .C2(
        keyinput_f122), .A(n10600), .ZN(n10609) );
  AOI22_X1 U11646 ( .A1(n10605), .A2(keyinput_f83), .B1(n10604), .B2(
        keyinput_f46), .ZN(n10603) );
  OAI221_X1 U11647 ( .B1(n10605), .B2(keyinput_f83), .C1(n10604), .C2(
        keyinput_f46), .A(n10603), .ZN(n10608) );
  XNOR2_X1 U11648 ( .A(n10606), .B(keyinput_f110), .ZN(n10607) );
  NOR4_X1 U11649 ( .A1(n10610), .A2(n10609), .A3(n10608), .A4(n10607), .ZN(
        n10613) );
  XOR2_X1 U11650 ( .A(keyinput_f123), .B(n10611), .Z(n10612) );
  AND2_X1 U11651 ( .A1(n10613), .A2(n10612), .ZN(n10655) );
  AOI22_X1 U11652 ( .A1(n10615), .A2(keyinput_f82), .B1(keyinput_f119), .B2(
        n5902), .ZN(n10614) );
  OAI221_X1 U11653 ( .B1(n10615), .B2(keyinput_f82), .C1(n5902), .C2(
        keyinput_f119), .A(n10614), .ZN(n10625) );
  AOI22_X1 U11654 ( .A1(n10618), .A2(keyinput_f23), .B1(n10617), .B2(
        keyinput_f69), .ZN(n10616) );
  OAI221_X1 U11655 ( .B1(n10618), .B2(keyinput_f23), .C1(n10617), .C2(
        keyinput_f69), .A(n10616), .ZN(n10624) );
  XNOR2_X1 U11656 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_f100), .ZN(n10622)
         );
  XNOR2_X1 U11657 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_f107), .ZN(n10621)
         );
  XNOR2_X1 U11658 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_f93), .ZN(n10620) );
  XNOR2_X1 U11659 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_f48), .ZN(n10619)
         );
  NAND4_X1 U11660 ( .A1(n10622), .A2(n10621), .A3(n10620), .A4(n10619), .ZN(
        n10623) );
  NOR3_X1 U11661 ( .A1(n10625), .A2(n10624), .A3(n10623), .ZN(n10654) );
  INV_X1 U11662 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U11663 ( .A1(n10627), .A2(keyinput_f36), .B1(n8335), .B2(
        keyinput_f42), .ZN(n10626) );
  OAI221_X1 U11664 ( .B1(n10627), .B2(keyinput_f36), .C1(n8335), .C2(
        keyinput_f42), .A(n10626), .ZN(n10639) );
  INV_X1 U11665 ( .A(keyinput_f0), .ZN(n10629) );
  AOI22_X1 U11666 ( .A1(n10630), .A2(keyinput_f54), .B1(P2_WR_REG_SCAN_IN), 
        .B2(n10629), .ZN(n10628) );
  OAI221_X1 U11667 ( .B1(n10630), .B2(keyinput_f54), .C1(n10629), .C2(
        P2_WR_REG_SCAN_IN), .A(n10628), .ZN(n10638) );
  AOI22_X1 U11668 ( .A1(n10633), .A2(keyinput_f40), .B1(keyinput_f24), .B2(
        n10632), .ZN(n10631) );
  OAI221_X1 U11669 ( .B1(n10633), .B2(keyinput_f40), .C1(n10632), .C2(
        keyinput_f24), .A(n10631), .ZN(n10637) );
  XNOR2_X1 U11670 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_f115), .ZN(n10635)
         );
  XNOR2_X1 U11671 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_f41), .ZN(n10634)
         );
  NAND2_X1 U11672 ( .A1(n10635), .A2(n10634), .ZN(n10636) );
  NOR4_X1 U11673 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10653) );
  INV_X1 U11674 ( .A(SI_16_), .ZN(n10641) );
  AOI22_X1 U11675 ( .A1(n10642), .A2(keyinput_f74), .B1(keyinput_f16), .B2(
        n10641), .ZN(n10640) );
  OAI221_X1 U11676 ( .B1(n10642), .B2(keyinput_f74), .C1(n10641), .C2(
        keyinput_f16), .A(n10640), .ZN(n10651) );
  XOR2_X1 U11677 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f91), .Z(n10650) );
  XNOR2_X1 U11678 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_f60), .ZN(n10646)
         );
  XNOR2_X1 U11679 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_f117), .ZN(n10645)
         );
  XNOR2_X1 U11680 ( .A(SI_22_), .B(keyinput_f10), .ZN(n10644) );
  XNOR2_X1 U11681 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_f108), .ZN(n10643)
         );
  NAND4_X1 U11682 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .ZN(
        n10649) );
  INV_X1 U11683 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10647) );
  XNOR2_X1 U11684 ( .A(keyinput_f120), .B(n10647), .ZN(n10648) );
  NOR4_X1 U11685 ( .A1(n10651), .A2(n10650), .A3(n10649), .A4(n10648), .ZN(
        n10652) );
  NAND4_X1 U11686 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(
        n10656) );
  NOR4_X1 U11687 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n10661) );
  XNOR2_X1 U11688 ( .A(n10664), .B(keyinput_f105), .ZN(n10660) );
  OAI22_X1 U11689 ( .A1(n10661), .A2(n10660), .B1(n10664), .B2(keyinput_g105), 
        .ZN(n10662) );
  AOI211_X1 U11690 ( .C1(keyinput_g105), .C2(n10664), .A(n10663), .B(n10662), 
        .ZN(n10665) );
  XOR2_X1 U11691 ( .A(n10666), .B(n10665), .Z(n10667) );
  XNOR2_X1 U11692 ( .A(n10668), .B(n10667), .ZN(ADD_1068_U4) );
  XNOR2_X1 U11693 ( .A(n10670), .B(n10669), .ZN(ADD_1068_U47) );
  XOR2_X1 U11694 ( .A(n10672), .B(n10671), .Z(ADD_1068_U54) );
  XNOR2_X1 U11695 ( .A(n10674), .B(n10673), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11696 ( .A(n10676), .B(n10675), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11697 ( .A(n10678), .B(n10677), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11698 ( .A(n10680), .B(n10679), .ZN(ADD_1068_U50) );
  XOR2_X1 U11699 ( .A(n10682), .B(n10681), .Z(ADD_1068_U53) );
  XNOR2_X1 U11700 ( .A(n10684), .B(n10683), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U5024 ( .A(n5943), .Z(n6387) );
  CLKBUF_X1 U5021 ( .A(n5948), .Z(n6535) );
  OAI211_X1 U5022 ( .C1(n9771), .C2(n10070), .A(n9770), .B(n9769), .ZN(n9865)
         );
  INV_X1 U5027 ( .A(n5339), .ZN(n5776) );
  CLKBUF_X2 U5036 ( .A(n6440), .Z(n6422) );
  CLKBUF_X1 U5056 ( .A(n5886), .Z(n5880) );
  XNOR2_X1 U5176 ( .A(n5281), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8318) );
endmodule

