

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650;

  INV_X2 U4894 ( .A(n8861), .ZN(P2_U3966) );
  INV_X2 U4896 ( .A(n6950), .ZN(n8760) );
  INV_X1 U4897 ( .A(n5633), .ZN(n6535) );
  INV_X1 U4898 ( .A(n9345), .ZN(n8280) );
  CLKBUF_X1 U4899 ( .A(n6584), .Z(n4830) );
  NAND2_X1 U4900 ( .A1(n5586), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5588) );
  XNOR2_X1 U4901 ( .A(n5603), .B(n5602), .ZN(n5604) );
  INV_X1 U4902 ( .A(n8587), .ZN(n8580) );
  INV_X2 U4903 ( .A(n6127), .ZN(n6129) );
  OR2_X1 U4904 ( .A1(n7573), .A2(n10612), .ZN(n7601) );
  NOR2_X1 U4905 ( .A1(n6301), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6261) );
  OR2_X1 U4906 ( .A1(n8809), .A2(n8812), .ZN(n8810) );
  NAND2_X1 U4907 ( .A1(n10449), .A2(n8890), .ZN(n8434) );
  INV_X2 U4908 ( .A(n5720), .ZN(n6536) );
  INV_X1 U4910 ( .A(n6768), .ZN(n10378) );
  OAI22_X1 U4911 ( .A1(n8760), .A2(n6788), .B1(n10413), .B2(n8763), .ZN(n6789)
         );
  AND2_X2 U4912 ( .A1(n8241), .A2(n6522), .ZN(n4874) );
  INV_X1 U4913 ( .A(n8761), .ZN(n4854) );
  NAND2_X1 U4914 ( .A1(n6646), .A2(n7388), .ZN(n7110) );
  NAND2_X1 U4915 ( .A1(n5585), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6144) );
  NOR2_X1 U4916 ( .A1(n9256), .A2(n4888), .ZN(n9199) );
  AOI21_X1 U4917 ( .B1(n8940), .B2(n6192), .A(n6126), .ZN(n8958) );
  NAND2_X1 U4918 ( .A1(n6791), .A2(n6790), .ZN(n4829) );
  OAI21_X2 U4919 ( .B1(n7805), .B2(n5255), .A(n5253), .ZN(n8104) );
  OAI21_X2 U4920 ( .B1(n7706), .B2(n7705), .A(n7704), .ZN(n7805) );
  INV_X8 U4921 ( .A(n4832), .ZN(n8257) );
  NOR2_X2 U4922 ( .A1(n8048), .A2(n8620), .ZN(n8047) );
  OAI22_X2 U4923 ( .A1(n8021), .A2(n8618), .B1(n10637), .B2(n8020), .ZN(n8048)
         );
  XNOR2_X2 U4924 ( .A(n5588), .B(n5587), .ZN(n5610) );
  AND2_X1 U4925 ( .A1(n5605), .A2(n5604), .ZN(n6584) );
  XNOR2_X2 U4926 ( .A(n6144), .B(n6143), .ZN(n6173) );
  XNOR2_X2 U4927 ( .A(n5011), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10292) );
  NAND2_X1 U4928 ( .A1(n4847), .A2(n4834), .ZN(n9196) );
  NAND2_X1 U4929 ( .A1(n4840), .A2(n9268), .ZN(n9208) );
  NAND2_X1 U4930 ( .A1(n5352), .A2(n5350), .ZN(n7936) );
  NAND2_X1 U4931 ( .A1(n7741), .A2(n7742), .ZN(n7740) );
  AND2_X1 U4932 ( .A1(n7782), .A2(n7781), .ZN(n7783) );
  INV_X1 U4933 ( .A(n9289), .ZN(n4834) );
  INV_X1 U4934 ( .A(n7125), .ZN(n4835) );
  AND3_X1 U4935 ( .A1(n5669), .A2(n5668), .A3(n5667), .ZN(n10451) );
  INV_X1 U4936 ( .A(n6779), .ZN(n6788) );
  CLKBUF_X3 U4937 ( .A(n6951), .Z(n8752) );
  NAND2_X1 U4938 ( .A1(n8598), .A2(n8636), .ZN(n8433) );
  INV_X1 U4939 ( .A(n5610), .ZN(n8598) );
  OAI21_X1 U4941 ( .B1(n6519), .B2(P1_IR_REG_29__SCAN_IN), .A(n6520), .ZN(
        n6523) );
  INV_X2 U4942 ( .A(n5491), .ZN(n4832) );
  OAI21_X1 U4943 ( .B1(n5112), .B2(n4936), .A(n5111), .ZN(n5110) );
  OR2_X1 U4944 ( .A1(n8639), .A2(n8638), .ZN(n5112) );
  OAI21_X1 U4945 ( .B1(n9191), .B2(n4849), .A(n4848), .ZN(n4847) );
  NAND2_X1 U4946 ( .A1(n9191), .A2(n9190), .ZN(n4848) );
  NAND2_X1 U4947 ( .A1(n5090), .A2(n8591), .ZN(n8637) );
  NAND2_X1 U4948 ( .A1(n4940), .A2(n4938), .ZN(n9191) );
  AND2_X1 U4949 ( .A1(n8810), .A2(n6077), .ZN(n8847) );
  NAND2_X1 U4950 ( .A1(n4850), .A2(n9197), .ZN(n8732) );
  OR2_X1 U4951 ( .A1(n6054), .A2(n6053), .ZN(n5476) );
  OR2_X1 U4952 ( .A1(n9199), .A2(n5462), .ZN(n8733) );
  NAND2_X1 U4953 ( .A1(n9199), .A2(n5462), .ZN(n4850) );
  NAND2_X1 U4954 ( .A1(n5389), .A2(n5388), .ZN(n8998) );
  INV_X1 U4955 ( .A(n5236), .ZN(n4849) );
  AOI21_X1 U4956 ( .B1(n5422), .B2(n9595), .A(n9292), .ZN(n5421) );
  NOR2_X1 U4957 ( .A1(n9258), .A2(n9257), .ZN(n9256) );
  OAI21_X1 U4958 ( .B1(n9208), .B2(n5239), .A(n5237), .ZN(n5247) );
  NAND2_X1 U4959 ( .A1(n4839), .A2(n4838), .ZN(n4840) );
  NAND2_X1 U4960 ( .A1(n4842), .A2(n4841), .ZN(n9267) );
  OR2_X1 U4961 ( .A1(n8704), .A2(n4837), .ZN(n9268) );
  OR2_X1 U4962 ( .A1(n8704), .A2(n8703), .ZN(n4842) );
  NAND2_X1 U4963 ( .A1(n8704), .A2(n4841), .ZN(n4839) );
  OR2_X1 U4964 ( .A1(n9741), .A2(n8383), .ZN(n8385) );
  NAND3_X1 U4965 ( .A1(n4853), .A2(n8109), .A3(n8110), .ZN(n8172) );
  NAND2_X1 U4966 ( .A1(n4853), .A2(n8120), .ZN(n8121) );
  AOI21_X2 U4967 ( .B1(n7936), .B2(n7932), .A(n7934), .ZN(n8137) );
  NAND2_X1 U4968 ( .A1(n8702), .A2(n8706), .ZN(n4837) );
  AOI21_X1 U4969 ( .B1(n4841), .B2(n8703), .A(n9269), .ZN(n4838) );
  NOR2_X1 U4970 ( .A1(n7880), .A2(n7881), .ZN(n7954) );
  NAND2_X1 U4971 ( .A1(n8339), .A2(n8338), .ZN(n9812) );
  AND2_X1 U4972 ( .A1(n5213), .A2(n5211), .ZN(n7674) );
  NAND2_X1 U4973 ( .A1(n7325), .A2(n7324), .ZN(n7307) );
  NAND2_X1 U4974 ( .A1(n7809), .A2(n7808), .ZN(n9434) );
  NAND2_X1 U4975 ( .A1(n4851), .A2(n7302), .ZN(n7325) );
  NAND2_X1 U4976 ( .A1(n7301), .A2(n7300), .ZN(n4851) );
  NAND2_X1 U4977 ( .A1(n7031), .A2(n7032), .ZN(n7301) );
  NAND2_X1 U4978 ( .A1(n7710), .A2(n7709), .ZN(n9871) );
  INV_X1 U4979 ( .A(n7601), .ZN(n5136) );
  NAND2_X1 U4980 ( .A1(n4852), .A2(n4872), .ZN(n7030) );
  INV_X2 U4981 ( .A(n10469), .ZN(n4833) );
  NAND2_X1 U4982 ( .A1(n7485), .A2(n7484), .ZN(n7728) );
  NAND2_X1 U4983 ( .A1(n4973), .A2(n5754), .ZN(n10596) );
  NAND2_X1 U4984 ( .A1(n6794), .A2(n6793), .ZN(n6847) );
  NOR2_X2 U4985 ( .A1(n9745), .A2(n6731), .ZN(n9262) );
  INV_X2 U4986 ( .A(n10539), .ZN(n10498) );
  OAI21_X1 U4987 ( .B1(n5740), .B2(n5739), .A(n5509), .ZN(n5767) );
  NAND2_X1 U4988 ( .A1(n4845), .A2(n4844), .ZN(n4843) );
  INV_X1 U4989 ( .A(n6890), .ZN(n4844) );
  INV_X2 U4990 ( .A(n8434), .ZN(n6911) );
  NAND2_X1 U4991 ( .A1(n8466), .A2(n7084), .ZN(n7356) );
  INV_X1 U4992 ( .A(n7074), .ZN(n10440) );
  NAND4_X1 U4993 ( .A1(n5673), .A2(n5672), .A3(n5671), .A4(n5670), .ZN(n8860)
         );
  INV_X1 U4994 ( .A(n8761), .ZN(n4836) );
  AND4_X1 U4995 ( .A1(n5729), .A2(n5728), .A3(n5727), .A4(n5726), .ZN(n7403)
         );
  AND4_X1 U4996 ( .A1(n5738), .A2(n5737), .A3(n5736), .A4(n5735), .ZN(n7397)
         );
  NAND2_X1 U4997 ( .A1(n4881), .A2(n5609), .ZN(n7074) );
  AND4_X1 U4998 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n7118)
         );
  AND4_X1 U4999 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n7240)
         );
  AND2_X1 U5000 ( .A1(n4855), .A2(n6649), .ZN(n6950) );
  NAND4_X1 U5001 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n6779)
         );
  NAND4_X1 U5002 ( .A1(n6527), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(n10355)
         );
  OR2_X2 U5003 ( .A1(n7110), .A2(n6647), .ZN(n8763) );
  INV_X1 U5004 ( .A(n6171), .ZN(n10340) );
  INV_X1 U5005 ( .A(n4855), .ZN(n8764) );
  INV_X1 U5006 ( .A(n7366), .ZN(n10405) );
  AND2_X2 U5007 ( .A1(n7110), .A2(n6815), .ZN(n4856) );
  AND3_X2 U5008 ( .A1(n6707), .A2(n6706), .A3(n6705), .ZN(n10351) );
  INV_X1 U5009 ( .A(n7097), .ZN(n10350) );
  NAND2_X1 U5010 ( .A1(n6173), .A2(n8423), .ZN(n6171) );
  XNOR2_X1 U5011 ( .A(n6232), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6698) );
  INV_X2 U5012 ( .A(n6806), .ZN(n6944) );
  NAND2_X1 U5013 ( .A1(n6231), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6232) );
  AND2_X2 U5014 ( .A1(n6522), .A2(n6523), .ZN(n6800) );
  INV_X1 U5015 ( .A(n5605), .ZN(n8249) );
  INV_X1 U5016 ( .A(n6521), .ZN(n6522) );
  INV_X1 U5017 ( .A(n6523), .ZN(n8241) );
  XNOR2_X1 U5018 ( .A(n5590), .B(n5589), .ZN(n8423) );
  NAND2_X1 U5019 ( .A1(n8263), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5600) );
  INV_X1 U5020 ( .A(n5604), .ZN(n8227) );
  NAND2_X1 U5021 ( .A1(n5575), .A2(n5574), .ZN(n8902) );
  NAND2_X1 U5022 ( .A1(n5299), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5590) );
  NOR2_X1 U5023 ( .A1(n5299), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6133) );
  XNOR2_X1 U5024 ( .A(n6219), .B(n6218), .ZN(n7749) );
  NAND2_X2 U5025 ( .A1(n4832), .A2(P2_U3152), .ZN(n7619) );
  NAND2_X1 U5026 ( .A1(n6244), .A2(n6228), .ZN(n6307) );
  NAND2_X1 U5027 ( .A1(n5574), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5572) );
  NAND2_X2 U5028 ( .A1(n5088), .A2(n5087), .ZN(n5491) );
  AND3_X2 U5029 ( .A1(n5880), .A2(n5678), .A3(n5566), .ZN(n5883) );
  NOR2_X1 U5030 ( .A1(n5570), .A2(n5569), .ZN(n5571) );
  NOR2_X2 U5031 ( .A1(n5665), .A2(n5559), .ZN(n5678) );
  AND2_X1 U5032 ( .A1(n6212), .A2(n5263), .ZN(n5267) );
  AND2_X1 U5033 ( .A1(n6221), .A2(n6218), .ZN(n5413) );
  AND4_X1 U5034 ( .A1(n6252), .A2(n6226), .A3(n6262), .A4(n6209), .ZN(n6212)
         );
  AND4_X1 U5035 ( .A1(n6206), .A2(n6204), .A3(n6205), .A4(n10200), .ZN(n5171)
         );
  AND3_X1 U5036 ( .A1(n6268), .A2(n6286), .A3(n6207), .ZN(n6208) );
  INV_X1 U5037 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6226) );
  NOR2_X1 U5038 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5560) );
  INV_X1 U5039 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6616) );
  INV_X1 U5040 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5589) );
  NOR2_X1 U5041 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5591) );
  INV_X1 U5042 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6169) );
  OR2_X1 U5043 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5559) );
  INV_X1 U5044 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5842) );
  INV_X1 U5045 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6221) );
  NOR2_X1 U5046 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6210) );
  NOR2_X1 U5047 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6211) );
  INV_X4 U5048 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5049 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5587) );
  INV_X1 U5050 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6230) );
  INV_X1 U5051 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6218) );
  NOR2_X1 U5052 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6268) );
  NOR2_X1 U5053 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5558) );
  INV_X1 U5054 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6238) );
  INV_X1 U5055 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6252) );
  INV_X4 U5056 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X2 U5057 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U5058 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6205) );
  NOR2_X1 U5059 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n6204) );
  INV_X1 U5060 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5795) );
  INV_X1 U5061 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6143) );
  INV_X1 U5062 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6147) );
  INV_X1 U5063 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5743) );
  INV_X1 U5064 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5716) );
  NOR2_X1 U5065 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5561) );
  INV_X1 U5066 ( .A(n8706), .ZN(n4841) );
  NAND3_X1 U5067 ( .A1(n6847), .A2(n6845), .A3(n6846), .ZN(n6848) );
  NAND2_X1 U5068 ( .A1(n4846), .A2(n4843), .ZN(n6794) );
  INV_X1 U5069 ( .A(n6892), .ZN(n4845) );
  NAND2_X1 U5070 ( .A1(n6889), .A2(n6714), .ZN(n4846) );
  NAND3_X1 U5071 ( .A1(n8732), .A2(n5227), .A3(n8733), .ZN(n5223) );
  OAI21_X2 U5072 ( .B1(n6307), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6617) );
  AND2_X2 U5073 ( .A1(n6261), .A2(n6224), .ZN(n6244) );
  NAND2_X1 U5074 ( .A1(n4852), .A2(n5261), .ZN(n6964) );
  NAND2_X1 U5075 ( .A1(n6961), .A2(n5262), .ZN(n4852) );
  AOI21_X1 U5076 ( .B1(n4853), .B2(n8109), .A(n8110), .ZN(n8111) );
  OAI211_X2 U5077 ( .C1(n8108), .C2(n5252), .A(n8107), .B(n4941), .ZN(n4853)
         );
  INV_X4 U5078 ( .A(n5173), .ZN(n6801) );
  NOR2_X2 U5079 ( .A1(n9821), .A2(n9682), .ZN(n9662) );
  AND2_X2 U5080 ( .A1(n7110), .A2(n6815), .ZN(n4855) );
  INV_X2 U5081 ( .A(n6697), .ZN(n10385) );
  OAI21_X2 U5082 ( .B1(n9013), .B2(n9005), .A(n8998), .ZN(n8978) );
  NAND2_X1 U5083 ( .A1(n10449), .A2(n8890), .ZN(n4857) );
  NAND2_X1 U5084 ( .A1(n10449), .A2(n8890), .ZN(n4858) );
  NAND2_X2 U5085 ( .A1(n8249), .A2(n8227), .ZN(n5620) );
  XNOR2_X2 U5086 ( .A(n5572), .B(n5597), .ZN(n6184) );
  AOI21_X2 U5087 ( .B1(n8137), .B2(n8138), .A(n8139), .ZN(n8131) );
  NAND2_X2 U5088 ( .A1(n8439), .A2(n6173), .ZN(n8587) );
  INV_X1 U5089 ( .A(n5945), .ZN(n4859) );
  NAND2_X1 U5090 ( .A1(n6382), .A2(n8257), .ZN(n5945) );
  OAI21_X1 U5091 ( .B1(n6080), .B2(n6079), .A(n6078), .ZN(n6100) );
  NAND2_X1 U5092 ( .A1(n5544), .A2(n5543), .ZN(n5879) );
  OAI21_X1 U5093 ( .B1(n5822), .B2(n5118), .A(n5115), .ZN(n5544) );
  INV_X1 U5094 ( .A(n5119), .ZN(n5118) );
  AND2_X1 U5095 ( .A1(n5116), .A2(n5542), .ZN(n5115) );
  NAND2_X1 U5096 ( .A1(n5822), .A2(n5470), .ZN(n5121) );
  NAND2_X1 U5097 ( .A1(n5222), .A2(n5221), .ZN(n5220) );
  NAND2_X1 U5098 ( .A1(n8241), .A2(n6521), .ZN(n5173) );
  INV_X1 U5099 ( .A(SI_10_), .ZN(n10082) );
  INV_X1 U5100 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6207) );
  AND2_X1 U5101 ( .A1(n5471), .A2(n5770), .ZN(n5517) );
  NAND2_X1 U5102 ( .A1(n5514), .A2(n10082), .ZN(n5519) );
  NAND2_X1 U5103 ( .A1(n5506), .A2(n10039), .ZN(n5509) );
  OR2_X1 U5104 ( .A1(n9110), .A2(n8970), .ZN(n8573) );
  OR2_X1 U5105 ( .A1(n9005), .A2(n8813), .ZN(n8563) );
  NAND2_X1 U5106 ( .A1(n5432), .A2(n8442), .ZN(n5431) );
  NAND2_X1 U5107 ( .A1(n9015), .A2(n4885), .ZN(n5432) );
  OR2_X1 U5108 ( .A1(n9155), .A2(n8913), .ZN(n8535) );
  NAND2_X1 U5109 ( .A1(n9077), .A2(n8234), .ZN(n5371) );
  NAND2_X1 U5110 ( .A1(n10630), .A2(n7956), .ZN(n5401) );
  OR2_X1 U5111 ( .A1(n10596), .A2(n7446), .ZN(n8502) );
  NOR2_X1 U5112 ( .A1(n9015), .A2(n5393), .ZN(n5392) );
  INV_X1 U5113 ( .A(n5395), .ZN(n5393) );
  NOR2_X1 U5114 ( .A1(n8004), .A2(n7827), .ZN(n6167) );
  NAND2_X1 U5115 ( .A1(n5883), .A2(n5576), .ZN(n5584) );
  INV_X1 U5116 ( .A(n5257), .ZN(n5256) );
  OAI21_X1 U5117 ( .B1(n4878), .B2(n8105), .A(n8106), .ZN(n5257) );
  NOR2_X1 U5118 ( .A1(n9493), .A2(n5295), .ZN(n9371) );
  INV_X1 U5119 ( .A(n9530), .ZN(n5296) );
  OR2_X1 U5120 ( .A1(n9790), .A2(n9598), .ZN(n9308) );
  AND2_X1 U5121 ( .A1(n4979), .A2(n9595), .ZN(n4977) );
  NAND2_X1 U5122 ( .A1(n9594), .A2(n5161), .ZN(n5160) );
  NOR2_X1 U5123 ( .A1(n8663), .A2(n8662), .ZN(n5473) );
  OR2_X1 U5124 ( .A1(n9801), .A2(n9597), .ZN(n9377) );
  OR2_X1 U5125 ( .A1(n9855), .A2(n9744), .ZN(n9389) );
  OR2_X1 U5126 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  OR2_X1 U5127 ( .A1(n9434), .A2(n9430), .ZN(n9422) );
  NAND2_X1 U5128 ( .A1(n7335), .A2(n7334), .ZN(n4999) );
  OAI21_X1 U5129 ( .B1(n6055), .B2(n5289), .A(n6059), .ZN(n6080) );
  INV_X1 U5130 ( .A(n6056), .ZN(n5289) );
  NOR2_X1 U5131 ( .A1(n5979), .A2(n5126), .ZN(n5125) );
  INV_X1 U5132 ( .A(n5962), .ZN(n5126) );
  NAND2_X1 U5133 ( .A1(n5961), .A2(n5960), .ZN(n5268) );
  INV_X1 U5134 ( .A(SI_12_), .ZN(n5282) );
  OAI21_X1 U5135 ( .B1(n6173), .B2(n8973), .A(n8423), .ZN(n5327) );
  NAND2_X1 U5136 ( .A1(n5921), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5932) );
  AND2_X1 U5137 ( .A1(n6166), .A2(n7145), .ZN(n6193) );
  INV_X1 U5138 ( .A(n6089), .ZN(n6192) );
  NAND2_X2 U5139 ( .A1(n8249), .A2(n5604), .ZN(n5633) );
  NAND2_X1 U5140 ( .A1(n5377), .A2(n5376), .ZN(n8937) );
  AOI21_X1 U5141 ( .B1(n5379), .B2(n5382), .A(n4900), .ZN(n5376) );
  OR2_X1 U5142 ( .A1(n9122), .A2(n8997), .ZN(n8966) );
  OR2_X1 U5143 ( .A1(n9138), .A2(n9049), .ZN(n5395) );
  NAND2_X1 U5144 ( .A1(n7587), .A2(n4964), .ZN(n4963) );
  INV_X1 U5145 ( .A(n10441), .ZN(n9082) );
  INV_X1 U5146 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U5147 ( .A1(n5883), .A2(n5133), .ZN(n5574) );
  AND2_X1 U5148 ( .A1(n5571), .A2(n5461), .ZN(n5133) );
  NAND2_X1 U5149 ( .A1(n5215), .A2(n7509), .ZN(n5214) );
  OR2_X1 U5150 ( .A1(n9345), .A2(n6919), .ZN(n6695) );
  INV_X1 U5151 ( .A(n6965), .ZN(n6962) );
  OR2_X1 U5152 ( .A1(n9778), .A2(n9351), .ZN(n9533) );
  INV_X1 U5153 ( .A(n6823), .ZN(n8672) );
  NAND2_X1 U5154 ( .A1(n5205), .A2(n5204), .ZN(n5203) );
  INV_X1 U5155 ( .A(n8330), .ZN(n5204) );
  AND2_X1 U5156 ( .A1(n9377), .A2(n9376), .ZN(n9475) );
  OR2_X1 U5157 ( .A1(n9816), .A2(n9239), .ZN(n9626) );
  NAND2_X1 U5158 ( .A1(n5206), .A2(n5205), .ZN(n9639) );
  OR2_X1 U5159 ( .A1(n8078), .A2(n8077), .ZN(n8177) );
  INV_X1 U5160 ( .A(n7917), .ZN(n5191) );
  NAND2_X1 U5161 ( .A1(n7124), .A2(n9356), .ZN(n7243) );
  NAND2_X1 U5162 ( .A1(n4982), .A2(n9572), .ZN(n9571) );
  INV_X1 U5163 ( .A(n9569), .ZN(n4982) );
  XNOR2_X1 U5164 ( .A(n8261), .B(n8260), .ZN(n9344) );
  NAND2_X1 U5165 ( .A1(n8256), .A2(n8255), .ZN(n8261) );
  AND2_X1 U5166 ( .A1(n5038), .A2(n5039), .ZN(n5037) );
  NAND2_X1 U5167 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(n6277), .ZN(n5039) );
  NAND2_X1 U5168 ( .A1(n6220), .A2(n5207), .ZN(n5208) );
  NOR2_X1 U5169 ( .A1(n5334), .A2(n5330), .ZN(n5329) );
  NOR2_X1 U5170 ( .A1(n6181), .A2(n6114), .ZN(n5334) );
  INV_X1 U5171 ( .A(n5332), .ZN(n5330) );
  INV_X1 U5172 ( .A(n9789), .ZN(n5407) );
  INV_X1 U5173 ( .A(n9395), .ZN(n5014) );
  NAND2_X1 U5174 ( .A1(n5017), .A2(n5016), .ZN(n5015) );
  NAND2_X1 U5175 ( .A1(n9392), .A2(n9488), .ZN(n5017) );
  NAND2_X1 U5176 ( .A1(n10520), .A2(n9492), .ZN(n5016) );
  NOR2_X1 U5177 ( .A1(n5049), .A2(n5045), .ZN(n5044) );
  NOR2_X1 U5178 ( .A1(n5051), .A2(n9421), .ZN(n5045) );
  NOR2_X1 U5179 ( .A1(n5054), .A2(n5050), .ZN(n5049) );
  OAI21_X1 U5180 ( .B1(n5033), .B2(n5032), .A(n5031), .ZN(n9420) );
  NAND2_X1 U5181 ( .A1(n4879), .A2(n5047), .ZN(n5046) );
  NAND2_X1 U5182 ( .A1(n5048), .A2(n5051), .ZN(n5047) );
  OR2_X1 U5183 ( .A1(n5054), .A2(n5053), .ZN(n5048) );
  NAND2_X1 U5184 ( .A1(n9484), .A2(n9491), .ZN(n5030) );
  AND2_X1 U5185 ( .A1(n9778), .A2(n9351), .ZN(n9493) );
  NOR2_X1 U5186 ( .A1(n7253), .A2(n5428), .ZN(n5427) );
  INV_X1 U5187 ( .A(n9517), .ZN(n5428) );
  INV_X1 U5188 ( .A(n5273), .ZN(n5272) );
  OAI21_X1 U5189 ( .B1(n6115), .B2(n5274), .A(n8223), .ZN(n5273) );
  INV_X1 U5190 ( .A(n6117), .ZN(n5274) );
  INV_X1 U5191 ( .A(n5940), .ZN(n5099) );
  NOR2_X1 U5192 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .ZN(
        n5478) );
  NAND2_X1 U5193 ( .A1(n5280), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5279) );
  INV_X1 U5194 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5280) );
  OAI21_X1 U5195 ( .B1(n8131), .B2(n8129), .A(n5307), .ZN(n5306) );
  AND2_X1 U5196 ( .A1(n5977), .A2(n5308), .ZN(n5307) );
  NAND2_X1 U5197 ( .A1(n5310), .A2(n5309), .ZN(n5308) );
  NAND2_X1 U5198 ( .A1(n8586), .A2(n5092), .ZN(n5091) );
  NOR2_X1 U5199 ( .A1(n5094), .A2(n5093), .ZN(n5092) );
  INV_X1 U5200 ( .A(n8583), .ZN(n5093) );
  INV_X1 U5201 ( .A(n8592), .ZN(n5095) );
  NAND2_X1 U5202 ( .A1(n5148), .A2(n5147), .ZN(n5146) );
  NOR2_X1 U5203 ( .A1(n5448), .A2(n5444), .ZN(n5443) );
  INV_X1 U5204 ( .A(n8440), .ZN(n5444) );
  INV_X1 U5205 ( .A(n5449), .ZN(n5448) );
  NOR2_X1 U5206 ( .A1(n8942), .A2(n5450), .ZN(n5449) );
  INV_X1 U5207 ( .A(n8573), .ZN(n5450) );
  INV_X1 U5208 ( .A(n5451), .ZN(n5447) );
  AND2_X1 U5209 ( .A1(n8948), .A2(n8595), .ZN(n5451) );
  OR2_X1 U5210 ( .A1(n9117), .A2(n8957), .ZN(n8596) );
  NAND2_X1 U5211 ( .A1(n5114), .A2(n4867), .ZN(n8552) );
  NOR2_X1 U5212 ( .A1(n9155), .A2(n9158), .ZN(n5142) );
  AND2_X1 U5213 ( .A1(n5401), .A2(n8616), .ZN(n5399) );
  AND2_X1 U5214 ( .A1(n5134), .A2(n10630), .ZN(n5137) );
  INV_X1 U5215 ( .A(n5138), .ZN(n5134) );
  NOR2_X1 U5216 ( .A1(n7175), .A2(n5457), .ZN(n5456) );
  INV_X1 U5217 ( .A(n7085), .ZN(n5457) );
  NAND2_X1 U5218 ( .A1(n10440), .A2(n7237), .ZN(n8472) );
  NOR2_X1 U5219 ( .A1(n7601), .A2(n10149), .ZN(n7778) );
  NAND2_X1 U5220 ( .A1(n7410), .A2(n7409), .ZN(n5375) );
  NOR2_X1 U5221 ( .A1(n8720), .A2(n5246), .ZN(n5245) );
  OAI22_X1 U5222 ( .A1(n8720), .A2(n5244), .B1(n8718), .B2(n8719), .ZN(n5243)
         );
  NAND2_X1 U5223 ( .A1(n9206), .A2(n9205), .ZN(n5244) );
  INV_X1 U5224 ( .A(n5254), .ZN(n5253) );
  OAI21_X1 U5225 ( .B1(n4877), .B2(n5255), .A(n8092), .ZN(n5254) );
  INV_X1 U5226 ( .A(n5260), .ZN(n5255) );
  OR2_X1 U5227 ( .A1(n5253), .A2(n5251), .ZN(n5250) );
  AND2_X1 U5228 ( .A1(n4877), .A2(n5252), .ZN(n5251) );
  INV_X1 U5229 ( .A(n8092), .ZN(n5258) );
  NAND2_X1 U5230 ( .A1(n6327), .A2(n6326), .ZN(n10317) );
  INV_X1 U5231 ( .A(n9463), .ZN(n5419) );
  AND2_X1 U5232 ( .A1(n8392), .A2(n9667), .ZN(n5418) );
  NAND2_X1 U5233 ( .A1(n8272), .A2(n9390), .ZN(n5201) );
  NAND2_X1 U5234 ( .A1(n4983), .A2(n9367), .ZN(n8206) );
  INV_X1 U5235 ( .A(n8208), .ZN(n4983) );
  INV_X1 U5236 ( .A(n4991), .ZN(n4985) );
  NAND2_X1 U5237 ( .A1(n6922), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7527) );
  OR2_X1 U5238 ( .A1(n7313), .A2(n7312), .ZN(n7491) );
  AND2_X1 U5239 ( .A1(n7248), .A2(n7242), .ZN(n4974) );
  NAND2_X1 U5240 ( .A1(n10515), .A2(n10486), .ZN(n9519) );
  NOR2_X1 U5241 ( .A1(n8291), .A2(n4998), .ZN(n4997) );
  INV_X1 U5242 ( .A(n8278), .ZN(n4998) );
  OR2_X1 U5243 ( .A1(n9837), .A2(n9723), .ZN(n5188) );
  OR2_X1 U5244 ( .A1(n5404), .A2(n5041), .ZN(n5038) );
  NAND2_X1 U5245 ( .A1(n8248), .A2(n8247), .ZN(n8252) );
  OAI21_X1 U5246 ( .B1(n4862), .B2(n6277), .A(n6240), .ZN(n5151) );
  AND2_X1 U5247 ( .A1(n6211), .A2(n6210), .ZN(n5263) );
  NAND2_X1 U5248 ( .A1(n6229), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6233) );
  AND2_X1 U5249 ( .A1(n5548), .A2(n5547), .ZN(n5878) );
  NOR2_X1 U5250 ( .A1(n5535), .A2(n5120), .ZN(n5119) );
  INV_X1 U5251 ( .A(n5533), .ZN(n5120) );
  INV_X1 U5252 ( .A(n5837), .ZN(n5535) );
  NAND2_X1 U5253 ( .A1(n5171), .A2(n6208), .ZN(n6301) );
  XNOR2_X1 U5254 ( .A(n5522), .B(n10080), .ZN(n5793) );
  NAND2_X1 U5255 ( .A1(n5521), .A2(n5463), .ZN(n5794) );
  AND2_X1 U5256 ( .A1(n5520), .A2(n5519), .ZN(n5463) );
  OR2_X1 U5257 ( .A1(n5518), .A2(n5768), .ZN(n5520) );
  NAND2_X1 U5258 ( .A1(n5085), .A2(n5500), .ZN(n5715) );
  INV_X1 U5259 ( .A(n5698), .ZN(n5086) );
  NAND2_X1 U5260 ( .A1(n8332), .A2(n5657), .ZN(n5114) );
  INV_X1 U5261 ( .A(n7167), .ZN(n5340) );
  NOR2_X1 U5262 ( .A1(n5340), .A2(n5344), .ZN(n5337) );
  NAND2_X1 U5263 ( .A1(n5721), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5733) );
  INV_X1 U5264 ( .A(n5723), .ZN(n5721) );
  AOI21_X1 U5265 ( .B1(n7390), .B2(n7389), .A(n5469), .ZN(n7623) );
  NOR2_X1 U5266 ( .A1(n7831), .A2(n5356), .ZN(n5355) );
  INV_X1 U5267 ( .A(n7754), .ZN(n5356) );
  NOR2_X1 U5268 ( .A1(n5897), .A2(n5354), .ZN(n5353) );
  INV_X1 U5269 ( .A(n5358), .ZN(n5354) );
  INV_X1 U5270 ( .A(n5355), .ZN(n5351) );
  OR2_X1 U5271 ( .A1(n5757), .A2(n5756), .ZN(n5776) );
  AND2_X1 U5272 ( .A1(n7046), .A2(n5347), .ZN(n5346) );
  NAND2_X1 U5273 ( .A1(n7004), .A2(n5349), .ZN(n5347) );
  NAND2_X1 U5274 ( .A1(n5938), .A2(n5310), .ZN(n5315) );
  INV_X1 U5275 ( .A(n5320), .ZN(n5319) );
  XNOR2_X1 U5276 ( .A(n8637), .B(n5089), .ZN(n8594) );
  INV_X1 U5277 ( .A(n8593), .ZN(n5089) );
  OR2_X1 U5278 ( .A1(n7752), .A2(n6168), .ZN(n6367) );
  NOR2_X1 U5279 ( .A1(n6429), .A2(n6428), .ZN(n6427) );
  NOR2_X1 U5280 ( .A1(n6427), .A2(n5002), .ZN(n6392) );
  NOR2_X1 U5281 ( .A1(n5004), .A2(n5003), .ZN(n5002) );
  OR2_X1 U5282 ( .A1(n6392), .A2(n6391), .ZN(n5001) );
  NOR2_X1 U5283 ( .A1(n6413), .A2(n4922), .ZN(n6416) );
  OR2_X1 U5284 ( .A1(n6416), .A2(n6415), .ZN(n5008) );
  INV_X1 U5285 ( .A(n5146), .ZN(n5145) );
  AND2_X1 U5286 ( .A1(n6122), .A2(n6186), .ZN(n8940) );
  NOR2_X1 U5287 ( .A1(n8967), .A2(n5384), .ZN(n5383) );
  AND2_X1 U5288 ( .A1(n8596), .A2(n8595), .ZN(n8967) );
  INV_X1 U5289 ( .A(n6044), .ZN(n6043) );
  NOR2_X1 U5290 ( .A1(n5390), .A2(n8993), .ZN(n5388) );
  NAND2_X1 U5291 ( .A1(n8414), .A2(n9056), .ZN(n8415) );
  OR2_X1 U5292 ( .A1(n4875), .A2(n4951), .ZN(n4950) );
  INV_X1 U5293 ( .A(n5431), .ZN(n4951) );
  NAND2_X1 U5294 ( .A1(n4949), .A2(n5431), .ZN(n8994) );
  NAND2_X1 U5295 ( .A1(n8416), .A2(n4875), .ZN(n4949) );
  OR2_X1 U5296 ( .A1(n9024), .A2(n8918), .ZN(n5394) );
  AND2_X1 U5297 ( .A1(n8552), .A2(n8442), .ZN(n9015) );
  OR2_X1 U5298 ( .A1(n9031), .A2(n9033), .ZN(n5434) );
  NOR2_X1 U5299 ( .A1(n9041), .A2(n8917), .ZN(n9024) );
  AOI21_X1 U5300 ( .B1(n5367), .B2(n8624), .A(n4899), .ZN(n5366) );
  OR2_X1 U5301 ( .A1(n5932), .A2(n5931), .ZN(n5950) );
  INV_X1 U5302 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5582) );
  AND2_X1 U5303 ( .A1(n4952), .A2(n4914), .ZN(n4957) );
  NAND2_X1 U5304 ( .A1(n9078), .A2(n8447), .ZN(n4956) );
  AND2_X1 U5305 ( .A1(n5371), .A2(n5372), .ZN(n5370) );
  NAND2_X1 U5306 ( .A1(n9067), .A2(n5371), .ZN(n5368) );
  NAND2_X1 U5307 ( .A1(n4861), .A2(n5441), .ZN(n4952) );
  NAND2_X1 U5308 ( .A1(n8028), .A2(n8229), .ZN(n5372) );
  INV_X1 U5309 ( .A(n7954), .ZN(n5440) );
  NAND2_X1 U5310 ( .A1(n8450), .A2(n4869), .ZN(n5437) );
  OR2_X1 U5311 ( .A1(n10637), .A2(n7952), .ZN(n8451) );
  AND2_X1 U5312 ( .A1(n8453), .A2(n8454), .ZN(n8619) );
  NOR2_X1 U5313 ( .A1(n8619), .A2(n5403), .ZN(n5400) );
  AND4_X1 U5314 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n7956)
         );
  AND2_X1 U5315 ( .A1(n4963), .A2(n8457), .ZN(n7773) );
  AND4_X1 U5316 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n7882)
         );
  NAND2_X1 U5317 ( .A1(n8457), .A2(n8456), .ZN(n7599) );
  OAI21_X1 U5318 ( .B1(n5459), .B2(n7427), .A(n4966), .ZN(n7569) );
  INV_X1 U5319 ( .A(n5460), .ZN(n5459) );
  AOI21_X1 U5320 ( .B1(n5460), .B2(n4967), .A(n5458), .ZN(n4966) );
  AND4_X1 U5321 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n7627)
         );
  AND2_X1 U5322 ( .A1(n7210), .A2(n8487), .ZN(n7211) );
  OR2_X1 U5323 ( .A1(n7209), .A2(n8486), .ZN(n7210) );
  AND2_X1 U5324 ( .A1(n8433), .A2(n8593), .ZN(n10437) );
  OR2_X1 U5325 ( .A1(n6761), .A2(n6185), .ZN(n10441) );
  INV_X1 U5326 ( .A(n10437), .ZN(n9085) );
  NAND2_X1 U5327 ( .A1(n6107), .A2(n6106), .ZN(n9110) );
  INV_X1 U5328 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5566) );
  AND2_X1 U5329 ( .A1(n5862), .A2(n5844), .ZN(n7973) );
  NAND2_X1 U5330 ( .A1(n7804), .A2(n7803), .ZN(n5260) );
  NAND2_X1 U5331 ( .A1(n6929), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8340) );
  INV_X1 U5332 ( .A(n8323), .ZN(n6929) );
  NAND2_X1 U5333 ( .A1(n9208), .A2(n5245), .ZN(n5242) );
  INV_X1 U5334 ( .A(n5243), .ZN(n5240) );
  INV_X1 U5335 ( .A(n7035), .ZN(n6921) );
  NAND2_X1 U5336 ( .A1(n6923), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7688) );
  INV_X1 U5337 ( .A(n7527), .ZN(n6923) );
  INV_X1 U5338 ( .A(n5245), .ZN(n5238) );
  NOR2_X1 U5339 ( .A1(n5243), .A2(n9216), .ZN(n5241) );
  NOR2_X1 U5340 ( .A1(n5222), .A2(n5221), .ZN(n5219) );
  INV_X1 U5341 ( .A(n7520), .ZN(n5217) );
  OAI21_X1 U5342 ( .B1(n7249), .B2(n8763), .A(n6948), .ZN(n6949) );
  INV_X1 U5343 ( .A(n8740), .ZN(n5228) );
  INV_X1 U5344 ( .A(n9237), .ZN(n5226) );
  NAND2_X1 U5345 ( .A1(n10317), .A2(n5076), .ZN(n5075) );
  NAND2_X1 U5346 ( .A1(n6328), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U5347 ( .A1(n5077), .A2(n5075), .ZN(n6570) );
  INV_X1 U5348 ( .A(n6572), .ZN(n5077) );
  INV_X1 U5349 ( .A(n6331), .ZN(n5062) );
  AOI21_X1 U5350 ( .B1(n6668), .B2(n5062), .A(n10260), .ZN(n5061) );
  NAND2_X1 U5351 ( .A1(n6607), .A2(n5073), .ZN(n5072) );
  INV_X1 U5352 ( .A(n6340), .ZN(n5073) );
  INV_X1 U5353 ( .A(n5072), .ZN(n5071) );
  OR2_X1 U5354 ( .A1(n7379), .A2(n7378), .ZN(n5067) );
  NAND2_X1 U5355 ( .A1(n5067), .A2(n5066), .ZN(n5065) );
  NAND2_X1 U5356 ( .A1(n7708), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5066) );
  AND2_X1 U5357 ( .A1(n5065), .A2(n5064), .ZN(n7607) );
  INV_X1 U5358 ( .A(n7608), .ZN(n5064) );
  NOR2_X1 U5359 ( .A1(n7607), .A2(n5063), .ZN(n6348) );
  AND2_X1 U5360 ( .A1(n7807), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5063) );
  OR2_X1 U5361 ( .A1(n7943), .A2(n7942), .ZN(n5056) );
  INV_X1 U5362 ( .A(n5160), .ZN(n5157) );
  NAND2_X1 U5363 ( .A1(n9600), .A2(n5422), .ZN(n9575) );
  NAND2_X1 U5364 ( .A1(n9600), .A2(n9375), .ZN(n9573) );
  NOR2_X1 U5365 ( .A1(n4894), .A2(n4980), .ZN(n4979) );
  NOR2_X1 U5366 ( .A1(n4981), .A2(n5205), .ZN(n4980) );
  NAND2_X1 U5367 ( .A1(n8394), .A2(n10473), .ZN(n8403) );
  NAND2_X1 U5368 ( .A1(n6927), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8297) );
  INV_X1 U5369 ( .A(n8284), .ZN(n6927) );
  AND2_X1 U5370 ( .A1(n9676), .A2(n9295), .ZN(n9694) );
  NAND2_X1 U5371 ( .A1(n5197), .A2(n5196), .ZN(n9721) );
  NAND2_X1 U5372 ( .A1(n5200), .A2(n8274), .ZN(n5196) );
  NAND2_X1 U5373 ( .A1(n8272), .A2(n5198), .ZN(n5197) );
  AND2_X1 U5374 ( .A1(n8274), .A2(n9390), .ZN(n5198) );
  OAI21_X1 U5375 ( .B1(n8085), .B2(n5412), .A(n5410), .ZN(n8382) );
  INV_X1 U5376 ( .A(n5411), .ZN(n5410) );
  OAI21_X1 U5377 ( .B1(n4863), .B2(n5412), .A(n9389), .ZN(n5411) );
  NAND2_X1 U5378 ( .A1(n6925), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8078) );
  INV_X1 U5379 ( .A(n8067), .ZN(n6925) );
  AND3_X1 U5380 ( .A1(n8082), .A2(n8081), .A3(n8080), .ZN(n9271) );
  AND4_X1 U5381 ( .A1(n7820), .A2(n7819), .A3(n7818), .A4(n7817), .ZN(n8094)
         );
  NAND2_X1 U5382 ( .A1(n8085), .A2(n4863), .ZN(n8211) );
  INV_X1 U5383 ( .A(n7916), .ZN(n5190) );
  NAND2_X1 U5384 ( .A1(n7901), .A2(n7900), .ZN(n7917) );
  OR2_X1 U5385 ( .A1(n7486), .A2(n9555), .ZN(n4991) );
  NOR2_X1 U5386 ( .A1(n9409), .A2(n4988), .ZN(n4987) );
  INV_X1 U5387 ( .A(n4990), .ZN(n4988) );
  NAND2_X1 U5388 ( .A1(n7486), .A2(n9555), .ZN(n4990) );
  NAND2_X1 U5389 ( .A1(n7466), .A2(n7465), .ZN(n7487) );
  AND2_X1 U5390 ( .A1(n9402), .A2(n9403), .ZN(n9401) );
  NAND2_X1 U5391 ( .A1(n6857), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6967) );
  AND2_X1 U5392 ( .A1(n7388), .A2(n9697), .ZN(n7105) );
  NAND2_X1 U5393 ( .A1(n9761), .A2(n7099), .ZN(n7124) );
  AND2_X1 U5394 ( .A1(n10346), .A2(n7098), .ZN(n9763) );
  NAND2_X1 U5395 ( .A1(n8671), .A2(n8670), .ZN(n9785) );
  NAND2_X1 U5396 ( .A1(n8060), .A2(n8059), .ZN(n9858) );
  XNOR2_X1 U5397 ( .A(n8252), .B(n8251), .ZN(n9339) );
  NAND2_X1 U5398 ( .A1(n6102), .A2(n6101), .ZN(n6116) );
  XNOR2_X1 U5399 ( .A(n6213), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6495) );
  INV_X1 U5400 ( .A(n6301), .ZN(n5170) );
  NAND2_X1 U5401 ( .A1(n5123), .A2(n5122), .ZN(n6000) );
  NAND2_X1 U5402 ( .A1(n5128), .A2(n6036), .ZN(n5122) );
  AND2_X1 U5403 ( .A1(n5125), .A2(n6036), .ZN(n5124) );
  NAND2_X1 U5404 ( .A1(n5100), .A2(n5104), .ZN(n5941) );
  NAND2_X1 U5405 ( .A1(n5102), .A2(n5101), .ZN(n5100) );
  NAND2_X1 U5406 ( .A1(n5121), .A2(n5533), .ZN(n5838) );
  NAND2_X1 U5407 ( .A1(n5528), .A2(n5527), .ZN(n5805) );
  NAND2_X1 U5408 ( .A1(n5361), .A2(n5360), .ZN(n8784) );
  AOI21_X1 U5409 ( .B1(n5362), .B2(n8812), .A(n6098), .ZN(n5360) );
  AND2_X1 U5410 ( .A1(n5333), .A2(n6180), .ZN(n5332) );
  NAND2_X1 U5411 ( .A1(n6114), .A2(n6178), .ZN(n5333) );
  INV_X1 U5412 ( .A(n6178), .ZN(n5335) );
  NAND2_X1 U5413 ( .A1(n6042), .A2(n6041), .ZN(n9005) );
  NAND2_X1 U5414 ( .A1(n5987), .A2(n5986), .ZN(n9138) );
  AND4_X1 U5415 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n8032)
         );
  NOR2_X1 U5416 ( .A1(n5435), .A2(n8644), .ZN(n5111) );
  AND2_X1 U5417 ( .A1(n6072), .A2(n6071), .ZN(n8997) );
  INV_X1 U5418 ( .A(n8813), .ZN(n9013) );
  AND3_X1 U5419 ( .A1(n5926), .A2(n5925), .A3(n5924), .ZN(n8234) );
  AND2_X1 U5420 ( .A1(n6371), .A2(n6369), .ZN(n8896) );
  NAND2_X1 U5421 ( .A1(n8429), .A2(n8428), .ZN(n9090) );
  OR2_X1 U5422 ( .A1(n5945), .A2(n5642), .ZN(n5647) );
  INV_X1 U5423 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U5424 ( .A1(n8335), .A2(n8334), .ZN(n9816) );
  NAND2_X1 U5425 ( .A1(n8750), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U5426 ( .A1(n9279), .A2(n9278), .ZN(n4940) );
  INV_X1 U5427 ( .A(n8751), .ZN(n4939) );
  AND4_X1 U5428 ( .A1(n6972), .A2(n6971), .A3(n6970), .A4(n6969), .ZN(n7342)
         );
  XNOR2_X1 U5429 ( .A(n6711), .B(n8761), .ZN(n6892) );
  XNOR2_X1 U5430 ( .A(n8739), .B(n8737), .ZN(n9237) );
  NAND2_X1 U5431 ( .A1(n8320), .A2(n8319), .ZN(n9821) );
  NAND2_X1 U5432 ( .A1(n8277), .A2(n8276), .ZN(n9843) );
  OR2_X1 U5433 ( .A1(n6960), .A2(n6959), .ZN(n5262) );
  NAND2_X1 U5434 ( .A1(n6960), .A2(n6959), .ZN(n5261) );
  AND2_X1 U5435 ( .A1(n8362), .A2(n8361), .ZN(n9285) );
  OR2_X1 U5436 ( .A1(n9230), .A2(n8672), .ZN(n8362) );
  AND2_X1 U5437 ( .A1(n5019), .A2(n5286), .ZN(n5018) );
  INV_X1 U5438 ( .A(n9542), .ZN(n5286) );
  OR2_X1 U5439 ( .A1(n4866), .A2(n9538), .ZN(n5019) );
  OR2_X1 U5440 ( .A1(n9499), .A2(n9697), .ZN(n5287) );
  AND2_X1 U5441 ( .A1(n5288), .A2(n9538), .ZN(n5022) );
  INV_X1 U5442 ( .A(n9718), .ZN(n5406) );
  NAND2_X1 U5443 ( .A1(n9571), .A2(n9570), .ZN(n9793) );
  XNOR2_X1 U5444 ( .A(n8380), .B(n9475), .ZN(n9805) );
  AOI21_X1 U5445 ( .B1(n9639), .B2(n8660), .A(n8366), .ZN(n8380) );
  OR2_X1 U5446 ( .A1(n10552), .A2(n6725), .ZN(n10488) );
  AND2_X1 U5447 ( .A1(n5409), .A2(n4930), .ZN(n9788) );
  NAND2_X1 U5448 ( .A1(n8694), .A2(n10473), .ZN(n5409) );
  NAND2_X1 U5449 ( .A1(n5179), .A2(n5178), .ZN(n9789) );
  OR2_X1 U5450 ( .A1(n9571), .A2(n5182), .ZN(n5178) );
  OAI21_X1 U5451 ( .B1(n5015), .B2(n10519), .A(n9521), .ZN(n9393) );
  OAI21_X1 U5452 ( .B1(n5015), .B2(n9396), .A(n5013), .ZN(n9398) );
  NOR2_X1 U5453 ( .A1(n5014), .A2(n7253), .ZN(n5013) );
  AOI21_X1 U5454 ( .B1(n5036), .B2(n5035), .A(n5034), .ZN(n5033) );
  NAND2_X1 U5455 ( .A1(n9405), .A2(n9404), .ZN(n5034) );
  NAND2_X1 U5456 ( .A1(n9399), .A2(n9488), .ZN(n5036) );
  AOI21_X1 U5457 ( .B1(n9400), .B2(n9492), .A(n7338), .ZN(n5035) );
  AND2_X1 U5458 ( .A1(n9414), .A2(n9413), .ZN(n5031) );
  NAND2_X1 U5459 ( .A1(n9408), .A2(n9409), .ZN(n5032) );
  NAND2_X1 U5460 ( .A1(n9425), .A2(n9492), .ZN(n5053) );
  NAND2_X1 U5461 ( .A1(n9422), .A2(n5052), .ZN(n5051) );
  AND2_X1 U5462 ( .A1(n9438), .A2(n9488), .ZN(n5052) );
  NOR2_X1 U5463 ( .A1(n9424), .A2(n5046), .ZN(n5042) );
  NAND2_X1 U5464 ( .A1(n4904), .A2(n5044), .ZN(n5043) );
  NOR2_X1 U5465 ( .A1(n9678), .A2(n5027), .ZN(n5026) );
  INV_X1 U5466 ( .A(n9694), .ZN(n5027) );
  AOI21_X1 U5467 ( .B1(n5025), .B2(n5024), .A(n5023), .ZN(n9469) );
  NAND2_X1 U5468 ( .A1(n9464), .A2(n9651), .ZN(n5023) );
  NOR2_X1 U5469 ( .A1(n9465), .A2(n9660), .ZN(n5024) );
  NAND2_X1 U5470 ( .A1(n9461), .A2(n5026), .ZN(n5025) );
  INV_X1 U5471 ( .A(n8129), .ZN(n5309) );
  NAND2_X1 U5472 ( .A1(n8585), .A2(n8584), .ZN(n5094) );
  NAND2_X1 U5473 ( .A1(n7070), .A2(n10405), .ZN(n8466) );
  NOR2_X1 U5474 ( .A1(n9352), .A2(n5298), .ZN(n5297) );
  NAND2_X1 U5475 ( .A1(n5429), .A2(n9517), .ZN(n10520) );
  NAND2_X1 U5476 ( .A1(n9391), .A2(n10471), .ZN(n5429) );
  INV_X1 U5477 ( .A(n5551), .ZN(n5291) );
  INV_X1 U5478 ( .A(n5878), .ZN(n5107) );
  NAND2_X1 U5479 ( .A1(n5119), .A2(n5117), .ZN(n5116) );
  INV_X1 U5480 ( .A(n5470), .ZN(n5117) );
  OAI21_X1 U5481 ( .B1(n5794), .B2(n5524), .A(n5523), .ZN(n5526) );
  INV_X1 U5482 ( .A(SI_11_), .ZN(n10080) );
  AND2_X1 U5483 ( .A1(n5313), .A2(n6008), .ZN(n5311) );
  NOR2_X1 U5484 ( .A1(n7753), .A2(n5856), .ZN(n5358) );
  NOR2_X1 U5485 ( .A1(n5974), .A2(n5973), .ZN(n6014) );
  AND2_X1 U5486 ( .A1(n7070), .A2(n4858), .ZN(n5649) );
  OR2_X1 U5487 ( .A1(n8929), .A2(n8419), .ZN(n8581) );
  OR2_X1 U5488 ( .A1(n9105), .A2(n8958), .ZN(n8576) );
  OR2_X1 U5489 ( .A1(n6121), .A2(n6120), .ZN(n6186) );
  AOI21_X1 U5490 ( .B1(n5381), .B2(n5380), .A(n8948), .ZN(n5379) );
  INV_X1 U5491 ( .A(n5383), .ZN(n5380) );
  INV_X1 U5492 ( .A(n5465), .ZN(n5430) );
  NAND2_X1 U5493 ( .A1(n8442), .A2(n8918), .ZN(n5433) );
  OR2_X1 U5494 ( .A1(n9143), .A2(n9056), .ZN(n8626) );
  NOR2_X1 U5495 ( .A1(n8534), .A2(n5365), .ZN(n5364) );
  INV_X1 U5496 ( .A(n5370), .ZN(n5365) );
  INV_X1 U5497 ( .A(n5368), .ZN(n5367) );
  NAND2_X1 U5498 ( .A1(n5847), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U5499 ( .A1(n10622), .A2(n5139), .ZN(n5138) );
  INV_X1 U5500 ( .A(n7599), .ZN(n8614) );
  NAND2_X1 U5501 ( .A1(n5784), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5812) );
  INV_X1 U5502 ( .A(n5786), .ZN(n5784) );
  INV_X1 U5503 ( .A(n7426), .ZN(n4967) );
  INV_X1 U5504 ( .A(n8505), .ZN(n5458) );
  AND2_X1 U5505 ( .A1(n8613), .A2(n8502), .ZN(n5460) );
  NOR2_X1 U5506 ( .A1(n8609), .A2(n7425), .ZN(n7426) );
  NOR2_X1 U5507 ( .A1(n7218), .A2(n7411), .ZN(n5132) );
  OR2_X1 U5508 ( .A1(n5741), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5742) );
  NOR2_X1 U5509 ( .A1(n5742), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5773) );
  AOI21_X1 U5510 ( .B1(n5029), .B2(n5028), .A(n9495), .ZN(n9501) );
  AND2_X1 U5511 ( .A1(n9496), .A2(n4865), .ZN(n5028) );
  NAND2_X1 U5512 ( .A1(n5030), .A2(n9485), .ZN(n5029) );
  INV_X1 U5513 ( .A(n9493), .ZN(n9536) );
  OR2_X1 U5514 ( .A1(n9796), .A2(n8771), .ZN(n9375) );
  INV_X1 U5515 ( .A(n4997), .ZN(n4993) );
  AND2_X1 U5516 ( .A1(n9694), .A2(n9458), .ZN(n5414) );
  AND2_X1 U5517 ( .A1(n5168), .A2(n5167), .ZN(n5166) );
  NOR2_X1 U5518 ( .A1(n9843), .A2(n9848), .ZN(n5168) );
  NAND2_X1 U5519 ( .A1(n8056), .A2(n8055), .ZN(n8208) );
  INV_X1 U5520 ( .A(n5427), .ZN(n5426) );
  AOI21_X1 U5521 ( .B1(n7248), .B2(n5427), .A(n5425), .ZN(n5424) );
  INV_X1 U5522 ( .A(n9762), .ZN(n9353) );
  NAND2_X1 U5523 ( .A1(n10356), .A2(n10385), .ZN(n9510) );
  NAND2_X1 U5524 ( .A1(n10348), .A2(n10347), .ZN(n10346) );
  OR2_X1 U5525 ( .A1(n9785), .A2(n9578), .ZN(n9482) );
  NAND2_X1 U5526 ( .A1(n9790), .A2(n5187), .ZN(n5186) );
  OR2_X1 U5527 ( .A1(n7467), .A2(n7486), .ZN(n7500) );
  NAND2_X1 U5528 ( .A1(n5429), .A2(n5427), .ZN(n10523) );
  NOR2_X1 U5529 ( .A1(n9771), .A2(n7104), .ZN(n7129) );
  NAND2_X1 U5530 ( .A1(n5149), .A2(n10385), .ZN(n9771) );
  INV_X1 U5531 ( .A(n10349), .ZN(n5149) );
  OR2_X1 U5532 ( .A1(n6722), .A2(n6716), .ZN(n7100) );
  NAND2_X1 U5533 ( .A1(n8266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5041) );
  AND2_X1 U5534 ( .A1(n4862), .A2(n5209), .ZN(n5207) );
  AND2_X1 U5535 ( .A1(n6517), .A2(n6239), .ZN(n5209) );
  NAND2_X1 U5536 ( .A1(n5270), .A2(n5269), .ZN(n8244) );
  AOI21_X1 U5537 ( .B1(n5272), .B2(n5274), .A(n4932), .ZN(n5269) );
  AOI21_X1 U5538 ( .B1(n6040), .B2(n6039), .A(n6038), .ZN(n6055) );
  INV_X1 U5539 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U5540 ( .A1(n5130), .A2(n5127), .ZN(n6040) );
  INV_X1 U5541 ( .A(n5995), .ZN(n5129) );
  NAND2_X1 U5542 ( .A1(n5096), .A2(n5097), .ZN(n5961) );
  AOI21_X1 U5543 ( .B1(n4860), .B2(n5108), .A(n5098), .ZN(n5097) );
  INV_X1 U5544 ( .A(n5939), .ZN(n5098) );
  AND2_X1 U5545 ( .A1(n5962), .A2(n5944), .ZN(n5960) );
  INV_X1 U5546 ( .A(n5105), .ZN(n5104) );
  OAI21_X1 U5547 ( .B1(n5293), .B2(n5106), .A(n5290), .ZN(n5105) );
  NAND2_X1 U5548 ( .A1(n5107), .A2(n5548), .ZN(n5106) );
  AOI21_X1 U5549 ( .B1(n5292), .B2(n5291), .A(n4903), .ZN(n5290) );
  INV_X1 U5550 ( .A(n5879), .ZN(n5102) );
  NAND2_X1 U5551 ( .A1(n5103), .A2(n5548), .ZN(n5899) );
  OR2_X1 U5552 ( .A1(n5526), .A2(n5525), .ZN(n5528) );
  AND2_X1 U5553 ( .A1(n5519), .A2(n5516), .ZN(n5770) );
  NAND2_X1 U5554 ( .A1(n5511), .A2(n10086), .ZN(n5768) );
  NAND2_X1 U5555 ( .A1(n5504), .A2(n5503), .ZN(n5740) );
  INV_X1 U5556 ( .A(n5714), .ZN(n5501) );
  NAND2_X1 U5557 ( .A1(n5509), .A2(n5508), .ZN(n5739) );
  XNOR2_X1 U5558 ( .A(n5502), .B(SI_7_), .ZN(n5714) );
  OR2_X1 U5559 ( .A1(n6273), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6275) );
  XNOR2_X1 U5560 ( .A(n5499), .B(SI_6_), .ZN(n5698) );
  NAND2_X1 U5561 ( .A1(n5498), .A2(n5497), .ZN(n5699) );
  NAND2_X1 U5562 ( .A1(n5277), .A2(n5276), .ZN(n5479) );
  NAND2_X1 U5563 ( .A1(n5279), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U5564 ( .A1(n5275), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5088) );
  INV_X1 U5565 ( .A(n5279), .ZN(n5275) );
  OR2_X1 U5566 ( .A1(n5776), .A2(n10105), .ZN(n5786) );
  INV_X1 U5567 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10105) );
  OR2_X1 U5568 ( .A1(n5731), .A2(n5730), .ZN(n5349) );
  NAND2_X1 U5569 ( .A1(n7740), .A2(n5358), .ZN(n5357) );
  INV_X1 U5570 ( .A(n5324), .ZN(n5323) );
  NAND2_X1 U5571 ( .A1(n6024), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6044) );
  INV_X1 U5572 ( .A(n6026), .ZN(n6024) );
  NAND2_X1 U5573 ( .A1(n5655), .A2(n5325), .ZN(n5324) );
  INV_X1 U5574 ( .A(n5656), .ZN(n5325) );
  NAND2_X1 U5575 ( .A1(n5732), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5757) );
  INV_X1 U5576 ( .A(n5733), .ZN(n5732) );
  NAND2_X1 U5577 ( .A1(n5825), .A2(n5824), .ZN(n7771) );
  NAND2_X1 U5578 ( .A1(n5304), .A2(n5302), .ZN(n8799) );
  NOR2_X1 U5579 ( .A1(n5464), .A2(n5937), .ZN(n5303) );
  INV_X1 U5580 ( .A(n6073), .ZN(n6076) );
  AND2_X1 U5581 ( .A1(n8846), .A2(n6077), .ZN(n5362) );
  AND2_X1 U5582 ( .A1(n8430), .A2(n8584), .ZN(n8435) );
  NAND2_X1 U5583 ( .A1(n5095), .A2(n5091), .ZN(n5090) );
  NAND2_X1 U5584 ( .A1(n6376), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5000) );
  AND2_X1 U5585 ( .A1(n5008), .A2(n5007), .ZN(n6442) );
  NAND2_X1 U5586 ( .A1(n6444), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5007) );
  NOR2_X1 U5587 ( .A1(n6442), .A2(n6441), .ZN(n6453) );
  NOR2_X1 U5588 ( .A1(n8950), .A2(n5146), .ZN(n8928) );
  AND2_X1 U5589 ( .A1(n8581), .A2(n8582), .ZN(n8921) );
  NAND2_X1 U5590 ( .A1(n5442), .A2(n5445), .ZN(n8924) );
  AOI21_X1 U5591 ( .B1(n5447), .B2(n5449), .A(n5446), .ZN(n5445) );
  INV_X1 U5592 ( .A(n8577), .ZN(n5446) );
  NAND2_X1 U5593 ( .A1(n8960), .A2(n8573), .ZN(n4972) );
  NAND2_X1 U5594 ( .A1(n8944), .A2(n9080), .ZN(n4970) );
  NAND2_X1 U5595 ( .A1(n8576), .A2(n8577), .ZN(n8942) );
  OR2_X1 U5596 ( .A1(n8950), .A2(n9105), .ZN(n8938) );
  INV_X1 U5597 ( .A(n8942), .ZN(n8936) );
  NAND2_X1 U5598 ( .A1(n5452), .A2(n5451), .ZN(n8960) );
  AOI21_X1 U5599 ( .B1(n8953), .B2(n6192), .A(n6111), .ZN(n8970) );
  AOI21_X1 U5600 ( .B1(n4876), .B2(n4951), .A(n4948), .ZN(n4947) );
  INV_X1 U5601 ( .A(n8563), .ZN(n4948) );
  NAND2_X1 U5602 ( .A1(n8980), .A2(n5384), .ZN(n8979) );
  NOR2_X1 U5603 ( .A1(n9132), .A2(n9025), .ZN(n9002) );
  OR2_X1 U5604 ( .A1(n9138), .A2(n9043), .ZN(n9025) );
  AND2_X1 U5605 ( .A1(n5142), .A2(n5141), .ZN(n5140) );
  INV_X1 U5606 ( .A(n5950), .ZN(n5948) );
  AND2_X1 U5607 ( .A1(n8541), .A2(n8916), .ZN(n9062) );
  OAI211_X1 U5608 ( .C1(n4959), .C2(n4955), .A(n4954), .B(n8535), .ZN(n9055)
         );
  OR2_X1 U5609 ( .A1(n4957), .A2(n4955), .ZN(n4954) );
  NAND2_X1 U5610 ( .A1(n4956), .A2(n8534), .ZN(n4955) );
  NAND2_X1 U5611 ( .A1(n9069), .A2(n9077), .ZN(n9070) );
  AND2_X1 U5612 ( .A1(n8028), .A2(n8043), .ZN(n9069) );
  OR2_X1 U5613 ( .A1(n5869), .A2(n5868), .ZN(n5888) );
  NAND2_X1 U5614 ( .A1(n5887), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5905) );
  INV_X1 U5615 ( .A(n5888), .ZN(n5887) );
  NAND2_X1 U5616 ( .A1(n5136), .A2(n4868), .ZN(n8040) );
  AND2_X1 U5617 ( .A1(n8450), .A2(n8449), .ZN(n8620) );
  NAND2_X1 U5618 ( .A1(n5398), .A2(n5401), .ZN(n5397) );
  INV_X1 U5619 ( .A(n5400), .ZN(n5398) );
  AND2_X1 U5620 ( .A1(n8451), .A2(n8452), .ZN(n8618) );
  NAND2_X1 U5621 ( .A1(n5136), .A2(n5137), .ZN(n8024) );
  NOR2_X1 U5622 ( .A1(n7601), .A2(n5138), .ZN(n7885) );
  AND4_X1 U5623 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n7952)
         );
  OAI211_X1 U5624 ( .C1(n7587), .C2(n4962), .A(n8517), .B(n4960), .ZN(n7880)
         );
  NAND2_X1 U5625 ( .A1(n4965), .A2(n4961), .ZN(n4960) );
  NAND2_X1 U5626 ( .A1(n5811), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5827) );
  INV_X1 U5627 ( .A(n5812), .ZN(n5811) );
  OR2_X1 U5628 ( .A1(n5827), .A2(n5826), .ZN(n5848) );
  NAND2_X1 U5629 ( .A1(n7454), .A2(n10604), .ZN(n7573) );
  NAND2_X1 U5630 ( .A1(n7445), .A2(n5460), .ZN(n7570) );
  NAND2_X1 U5631 ( .A1(n7427), .A2(n7426), .ZN(n7445) );
  NAND2_X1 U5632 ( .A1(n5132), .A2(n5131), .ZN(n7432) );
  INV_X1 U5633 ( .A(n5132), .ZN(n7404) );
  AND4_X1 U5634 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n7446)
         );
  NAND2_X1 U5635 ( .A1(n5703), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5723) );
  AOI21_X1 U5636 ( .B1(n10438), .B2(n5456), .A(n5455), .ZN(n5453) );
  INV_X1 U5637 ( .A(n8482), .ZN(n5455) );
  NAND2_X1 U5638 ( .A1(n10444), .A2(n7085), .ZN(n7177) );
  AND2_X1 U5639 ( .A1(n10448), .A2(n10501), .ZN(n7217) );
  NOR2_X1 U5640 ( .A1(n10446), .A2(n10465), .ZN(n10448) );
  OR2_X1 U5641 ( .A1(n10436), .A2(n10438), .ZN(n10444) );
  INV_X1 U5642 ( .A(n8475), .ZN(n8602) );
  NAND2_X1 U5643 ( .A1(n5475), .A2(n7083), .ZN(n7357) );
  NOR2_X1 U5644 ( .A1(n6768), .A2(n10339), .ZN(n7361) );
  NAND2_X1 U5645 ( .A1(n6912), .A2(n10339), .ZN(n8599) );
  NAND2_X1 U5646 ( .A1(n5326), .A2(n8890), .ZN(n6763) );
  OAI21_X1 U5647 ( .B1(n8423), .B2(n8598), .A(n6173), .ZN(n5326) );
  NAND2_X1 U5648 ( .A1(n6064), .A2(n6063), .ZN(n9122) );
  AND2_X1 U5649 ( .A1(n5394), .A2(n5392), .ZN(n9137) );
  NAND2_X1 U5650 ( .A1(n5809), .A2(n5808), .ZN(n10149) );
  NOR2_X1 U5651 ( .A1(n8607), .A2(n5374), .ZN(n5373) );
  INV_X1 U5652 ( .A(n7413), .ZN(n5374) );
  AND2_X1 U5653 ( .A1(n7147), .A2(n6173), .ZN(n10609) );
  INV_X1 U5654 ( .A(n10644), .ZN(n10620) );
  AND2_X1 U5655 ( .A1(n6774), .A2(n6759), .ZN(n7154) );
  AND2_X1 U5656 ( .A1(n7152), .A2(n6755), .ZN(n6776) );
  NOR2_X1 U5657 ( .A1(n6167), .A2(n6150), .ZN(n9937) );
  NAND2_X1 U5658 ( .A1(n5300), .A2(n4887), .ZN(n5299) );
  NOR2_X1 U5659 ( .A1(n5565), .A2(n5564), .ZN(n5880) );
  OR3_X1 U5660 ( .A1(n5806), .A2(P2_IR_REG_11__SCAN_IN), .A3(
        P2_IR_REG_10__SCAN_IN), .ZN(n5823) );
  XNOR2_X1 U5661 ( .A(n6241), .B(n6239), .ZN(n6313) );
  NAND2_X1 U5662 ( .A1(n6516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6241) );
  INV_X1 U5663 ( .A(n9190), .ZN(n5236) );
  NAND2_X1 U5664 ( .A1(n6920), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7035) );
  INV_X1 U5665 ( .A(n6967), .ZN(n6920) );
  OR2_X1 U5666 ( .A1(n8739), .A2(n8738), .ZN(n8740) );
  INV_X1 U5667 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7284) );
  OR2_X1 U5668 ( .A1(n8309), .A2(n8308), .ZN(n8321) );
  NAND2_X1 U5669 ( .A1(n6928), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8323) );
  INV_X1 U5670 ( .A(n8321), .ZN(n6928) );
  OAI22_X1 U5671 ( .A1(n7118), .A2(n8763), .B1(n10385), .B2(n8764), .ZN(n6700)
         );
  NAND2_X1 U5672 ( .A1(n5249), .A2(n4893), .ZN(n8120) );
  NAND2_X1 U5673 ( .A1(n5253), .A2(n5255), .ZN(n5248) );
  NAND2_X1 U5674 ( .A1(n5259), .A2(n4878), .ZN(n4941) );
  OR2_X1 U5675 ( .A1(n9500), .A2(n10493), .ZN(n5288) );
  AND2_X1 U5676 ( .A1(n6937), .A2(n6936), .ZN(n9239) );
  NOR2_X1 U5677 ( .A1(n6669), .A2(n6668), .ZN(n6667) );
  OR2_X1 U5678 ( .A1(n6677), .A2(n6300), .ZN(n10232) );
  OAI21_X1 U5679 ( .B1(n9661), .B2(n4976), .A(n4975), .ZN(n9569) );
  AOI21_X1 U5680 ( .B1(n4977), .B2(n4981), .A(n4905), .ZN(n4975) );
  INV_X1 U5681 ( .A(n4977), .ZN(n4976) );
  OR2_X1 U5682 ( .A1(n9584), .A2(n8672), .ZN(n8658) );
  OR2_X1 U5683 ( .A1(n8365), .A2(n8364), .ZN(n8662) );
  NAND2_X1 U5684 ( .A1(n5417), .A2(n5416), .ZN(n9616) );
  NAND2_X1 U5685 ( .A1(n4906), .A2(n8392), .ZN(n5416) );
  NAND2_X1 U5686 ( .A1(n5420), .A2(n9463), .ZN(n9649) );
  NAND2_X1 U5687 ( .A1(n9668), .A2(n9667), .ZN(n5420) );
  OAI21_X1 U5688 ( .B1(n9719), .B2(n4994), .A(n4992), .ZN(n9674) );
  INV_X1 U5689 ( .A(n4995), .ZN(n4994) );
  AOI21_X1 U5690 ( .B1(n4993), .B2(n4995), .A(n4925), .ZN(n4992) );
  AND2_X1 U5691 ( .A1(n5188), .A2(n4928), .ZN(n4995) );
  NAND2_X1 U5692 ( .A1(n9749), .A2(n5164), .ZN(n9690) );
  NOR2_X1 U5693 ( .A1(n9833), .A2(n5165), .ZN(n5164) );
  INV_X1 U5694 ( .A(n5166), .ZN(n5165) );
  NAND2_X1 U5695 ( .A1(n6926), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8284) );
  OR2_X1 U5696 ( .A1(n9848), .A2(n9271), .ZN(n9724) );
  NAND2_X1 U5697 ( .A1(n9749), .A2(n5168), .ZN(n9730) );
  NAND2_X1 U5698 ( .A1(n9749), .A2(n9755), .ZN(n9750) );
  NAND2_X1 U5699 ( .A1(n5201), .A2(n5199), .ZN(n9738) );
  OR2_X1 U5700 ( .A1(n7815), .A2(n7814), .ZN(n8067) );
  AND2_X1 U5701 ( .A1(n8119), .A2(n8214), .ZN(n9749) );
  NAND2_X1 U5702 ( .A1(n8206), .A2(n8061), .ZN(n8272) );
  NOR2_X1 U5703 ( .A1(n8215), .A2(n9858), .ZN(n8214) );
  AND3_X1 U5704 ( .A1(n8071), .A2(n8070), .A3(n8069), .ZN(n9744) );
  NAND2_X1 U5705 ( .A1(n8085), .A2(n9422), .ZN(n8209) );
  OR2_X1 U5706 ( .A1(n7993), .A2(n9434), .ZN(n8215) );
  OAI21_X1 U5707 ( .B1(n7901), .B2(n5193), .A(n5189), .ZN(n7918) );
  AOI21_X1 U5708 ( .B1(n5192), .B2(n9418), .A(n4898), .ZN(n5189) );
  OR2_X1 U5709 ( .A1(n7995), .A2(n9871), .ZN(n7993) );
  NAND2_X1 U5710 ( .A1(n7907), .A2(n7912), .ZN(n7995) );
  OAI21_X1 U5711 ( .B1(n7487), .B2(n4986), .A(n4984), .ZN(n7729) );
  AOI21_X1 U5712 ( .B1(n4987), .B2(n4985), .A(n4897), .ZN(n4984) );
  INV_X1 U5713 ( .A(n4987), .ZN(n4986) );
  NOR2_X1 U5714 ( .A1(n7500), .A2(n7728), .ZN(n7733) );
  AND4_X1 U5715 ( .A1(n7496), .A2(n7495), .A3(n7494), .A4(n7493), .ZN(n7896)
         );
  NAND2_X1 U5716 ( .A1(n7347), .A2(n10564), .ZN(n7467) );
  NAND2_X1 U5717 ( .A1(n4999), .A2(n7336), .ZN(n7339) );
  AND2_X1 U5718 ( .A1(n7262), .A2(n7266), .ZN(n7347) );
  AND2_X1 U5719 ( .A1(n5195), .A2(n5194), .ZN(n10509) );
  NAND2_X1 U5720 ( .A1(n7243), .A2(n4974), .ZN(n5195) );
  NAND2_X1 U5721 ( .A1(n7129), .A2(n4835), .ZN(n10476) );
  OR2_X1 U5722 ( .A1(n10476), .A2(n7259), .ZN(n10510) );
  AND4_X1 U5723 ( .A1(n6830), .A2(n6829), .A3(n6828), .A4(n6827), .ZN(n7247)
         );
  NAND2_X1 U5724 ( .A1(n9763), .A2(n9762), .ZN(n9761) );
  AND2_X1 U5725 ( .A1(n9498), .A2(n6727), .ZN(n10516) );
  NAND2_X1 U5726 ( .A1(n5187), .A2(n10516), .ZN(n8693) );
  INV_X1 U5727 ( .A(n5186), .ZN(n5181) );
  NAND2_X1 U5728 ( .A1(n9482), .A2(n9489), .ZN(n9352) );
  INV_X1 U5729 ( .A(n9352), .ZN(n5182) );
  AND2_X1 U5730 ( .A1(n5182), .A2(n5186), .ZN(n5180) );
  NAND2_X1 U5731 ( .A1(n4996), .A2(n5188), .ZN(n9692) );
  NAND2_X1 U5732 ( .A1(n9719), .A2(n4997), .ZN(n4996) );
  NAND2_X1 U5733 ( .A1(n8065), .A2(n8064), .ZN(n9855) );
  AND2_X1 U5734 ( .A1(n7261), .A2(n9540), .ZN(n10549) );
  INV_X1 U5735 ( .A(n10477), .ZN(n10565) );
  NAND2_X1 U5736 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  OR2_X1 U5737 ( .A1(n9345), .A2(n6701), .ZN(n6707) );
  AND2_X1 U5738 ( .A1(n9502), .A2(n7462), .ZN(n7261) );
  NOR2_X1 U5739 ( .A1(n4870), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5404) );
  XNOR2_X1 U5740 ( .A(n8244), .B(n8243), .ZN(n8668) );
  NAND2_X1 U5741 ( .A1(n5152), .A2(n5150), .ZN(n6242) );
  INV_X1 U5742 ( .A(n5151), .ZN(n5150) );
  CLKBUF_X1 U5743 ( .A(n6313), .Z(n10220) );
  NAND2_X1 U5744 ( .A1(n6220), .A2(n5413), .ZN(n6236) );
  NAND2_X1 U5745 ( .A1(n5130), .A2(n5982), .ZN(n5996) );
  CLKBUF_X1 U5746 ( .A(n6646), .Z(n6234) );
  AND2_X1 U5747 ( .A1(n6245), .A2(n6227), .ZN(n6228) );
  XNOR2_X1 U5748 ( .A(n5861), .B(n5860), .ZN(n8057) );
  NAND2_X1 U5749 ( .A1(n5121), .A2(n5119), .ZN(n5859) );
  NAND2_X1 U5750 ( .A1(n5074), .A2(n6279), .ZN(n6282) );
  OR2_X1 U5751 ( .A1(n6278), .A2(n6277), .ZN(n5074) );
  NAND2_X1 U5752 ( .A1(n5074), .A2(n6288), .ZN(n6287) );
  AND2_X1 U5753 ( .A1(n6095), .A2(n6094), .ZN(n8957) );
  OR2_X1 U5754 ( .A1(n8972), .A2(n6089), .ZN(n6095) );
  NAND2_X1 U5755 ( .A1(n5114), .A2(n6006), .ZN(n9132) );
  NAND2_X1 U5756 ( .A1(n5336), .A2(n5338), .ZN(n7371) );
  INV_X1 U5757 ( .A(n5339), .ZN(n5338) );
  OAI21_X1 U5758 ( .B1(n5341), .B2(n5340), .A(n5766), .ZN(n5339) );
  NAND2_X1 U5759 ( .A1(n5345), .A2(n5349), .ZN(n7047) );
  OR2_X1 U5760 ( .A1(n7003), .A2(n7004), .ZN(n5345) );
  AND2_X1 U5761 ( .A1(n6193), .A2(n6182), .ZN(n8815) );
  AND2_X1 U5762 ( .A1(n8815), .A2(n9080), .ZN(n8804) );
  NAND2_X1 U5763 ( .A1(n5357), .A2(n7754), .ZN(n7830) );
  NAND2_X1 U5764 ( .A1(n5886), .A2(n5885), .ZN(n9169) );
  NAND2_X1 U5765 ( .A1(n5318), .A2(n7010), .ZN(n6994) );
  NAND2_X1 U5766 ( .A1(n6885), .A2(n5322), .ZN(n5318) );
  OAI21_X1 U5767 ( .B1(n6885), .B2(n5321), .A(n5319), .ZN(n6993) );
  NAND2_X1 U5768 ( .A1(n5351), .A2(n5359), .ZN(n5350) );
  NAND2_X1 U5769 ( .A1(n7740), .A2(n5353), .ZN(n5352) );
  NAND2_X1 U5770 ( .A1(n6885), .A2(n5324), .ZN(n7013) );
  AND4_X1 U5771 ( .A1(n5781), .A2(n5780), .A3(n5779), .A4(n5778), .ZN(n7442)
         );
  NAND2_X1 U5772 ( .A1(n7168), .A2(n7167), .ZN(n7166) );
  NAND2_X1 U5773 ( .A1(n5342), .A2(n5341), .ZN(n7168) );
  NAND2_X1 U5774 ( .A1(n7003), .A2(n5343), .ZN(n5342) );
  INV_X1 U5775 ( .A(n5305), .ZN(n5314) );
  AOI21_X1 U5776 ( .B1(n8131), .B2(n5937), .A(n8129), .ZN(n5305) );
  NOR2_X1 U5777 ( .A1(n8837), .A2(n8838), .ZN(n8836) );
  AND2_X1 U5778 ( .A1(n8815), .A2(n9082), .ZN(n8802) );
  NAND2_X1 U5779 ( .A1(n5319), .A2(n5321), .ZN(n5316) );
  NAND2_X1 U5780 ( .A1(n6885), .A2(n5319), .ZN(n5317) );
  AND2_X1 U5781 ( .A1(n6174), .A2(n10373), .ZN(n10399) );
  INV_X1 U5782 ( .A(n8820), .ZN(n8848) );
  INV_X1 U5783 ( .A(n8804), .ZN(n10393) );
  NAND2_X1 U5784 ( .A1(n8810), .A2(n5362), .ZN(n8845) );
  INV_X1 U5785 ( .A(n8802), .ZN(n10394) );
  NAND2_X1 U5786 ( .A1(n7740), .A2(n5857), .ZN(n7757) );
  INV_X1 U5787 ( .A(n10399), .ZN(n8851) );
  NAND2_X1 U5788 ( .A1(n6203), .A2(n10274), .ZN(n8861) );
  INV_X1 U5789 ( .A(n5001), .ZN(n6390) );
  INV_X1 U5790 ( .A(n5008), .ZN(n6439) );
  NOR2_X1 U5791 ( .A1(n6467), .A2(n5010), .ZN(n6470) );
  AND2_X1 U5792 ( .A1(n6472), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5010) );
  NOR2_X1 U5793 ( .A1(n6470), .A2(n6469), .ZN(n7189) );
  NOR2_X1 U5794 ( .A1(n7189), .A2(n5009), .ZN(n7190) );
  AND2_X1 U5795 ( .A1(n7195), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U5796 ( .A1(n7190), .A2(n7191), .ZN(n7539) );
  NOR2_X1 U5797 ( .A1(n7562), .A2(n5006), .ZN(n7542) );
  AND2_X1 U5798 ( .A1(n7567), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U5799 ( .A1(n7542), .A2(n7541), .ZN(n7644) );
  NAND2_X1 U5800 ( .A1(n7644), .A2(n5005), .ZN(n7647) );
  OR2_X1 U5801 ( .A1(n7650), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U5802 ( .A1(n7647), .A2(n7646), .ZN(n7972) );
  XNOR2_X1 U5803 ( .A(n8900), .B(n9090), .ZN(n9092) );
  NOR2_X1 U5804 ( .A1(n9094), .A2(n5144), .ZN(n5143) );
  NAND2_X1 U5805 ( .A1(n5145), .A2(n8955), .ZN(n5144) );
  AOI21_X1 U5806 ( .B1(n4971), .B2(n9085), .A(n4968), .ZN(n9108) );
  NAND2_X1 U5807 ( .A1(n4970), .A2(n4969), .ZN(n4968) );
  XNOR2_X1 U5808 ( .A(n4972), .B(n8942), .ZN(n4971) );
  NAND2_X1 U5809 ( .A1(n8943), .A2(n9082), .ZN(n4969) );
  NAND2_X1 U5810 ( .A1(n5378), .A2(n5381), .ZN(n8949) );
  NAND2_X1 U5811 ( .A1(n8978), .A2(n5383), .ZN(n5378) );
  NAND2_X1 U5812 ( .A1(n6085), .A2(n6084), .ZN(n9117) );
  AOI21_X1 U5813 ( .B1(n8978), .B2(n8919), .A(n5385), .ZN(n8965) );
  AND2_X1 U5814 ( .A1(n6087), .A2(n6066), .ZN(n8986) );
  AND2_X1 U5815 ( .A1(n5389), .A2(n5391), .ZN(n9000) );
  OAI21_X1 U5816 ( .B1(n8416), .B2(n4951), .A(n4876), .ZN(n8992) );
  NAND2_X1 U5817 ( .A1(n5394), .A2(n5395), .ZN(n9016) );
  AND2_X1 U5818 ( .A1(n5434), .A2(n4885), .ZN(n9012) );
  INV_X1 U5819 ( .A(n5434), .ZN(n9032) );
  NAND2_X1 U5820 ( .A1(n5581), .A2(n5580), .ZN(n9155) );
  NAND2_X1 U5821 ( .A1(n4953), .A2(n4956), .ZN(n8413) );
  NAND2_X1 U5822 ( .A1(n4957), .A2(n4959), .ZN(n4953) );
  NAND2_X1 U5823 ( .A1(n8231), .A2(n8624), .ZN(n8915) );
  NAND2_X1 U5824 ( .A1(n5369), .A2(n5368), .ZN(n8231) );
  NAND2_X1 U5825 ( .A1(n8230), .A2(n5370), .ZN(n5369) );
  NAND2_X1 U5826 ( .A1(n4959), .A2(n4958), .ZN(n9079) );
  AND2_X1 U5827 ( .A1(n4952), .A2(n8528), .ZN(n4958) );
  NAND2_X1 U5828 ( .A1(n8230), .A2(n5372), .ZN(n9068) );
  NAND2_X1 U5829 ( .A1(n5438), .A2(n5437), .ZN(n8232) );
  NAND2_X1 U5830 ( .A1(n5440), .A2(n5439), .ZN(n5438) );
  NAND2_X1 U5831 ( .A1(n5846), .A2(n5845), .ZN(n7889) );
  NAND2_X1 U5832 ( .A1(n7877), .A2(n5402), .ZN(n7878) );
  NAND2_X1 U5833 ( .A1(n4963), .A2(n4961), .ZN(n7879) );
  AND2_X1 U5834 ( .A1(n7587), .A2(n8506), .ZN(n7772) );
  NAND2_X1 U5835 ( .A1(n5800), .A2(n5799), .ZN(n10612) );
  NAND2_X1 U5836 ( .A1(n7270), .A2(n5657), .ZN(n4973) );
  NAND2_X1 U5837 ( .A1(n5387), .A2(n7080), .ZN(n7204) );
  OR2_X1 U5838 ( .A1(n6383), .A2(n6755), .ZN(n10373) );
  INV_X1 U5839 ( .A(n9076), .ZN(n10466) );
  INV_X1 U5840 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6512) );
  AND2_X1 U5841 ( .A1(n5645), .A2(n5644), .ZN(n10307) );
  NAND2_X1 U5842 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5011) );
  AND4_X1 U5843 ( .A1(n6863), .A2(n6862), .A3(n6861), .A4(n6860), .ZN(n7249)
         );
  NAND2_X1 U5844 ( .A1(n5259), .A2(n5260), .ZN(n8093) );
  NAND2_X1 U5845 ( .A1(n7507), .A2(n5219), .ZN(n7519) );
  INV_X1 U5846 ( .A(n8759), .ZN(n5231) );
  NAND2_X1 U5847 ( .A1(n5242), .A2(n5240), .ZN(n9215) );
  AND4_X1 U5848 ( .A1(n7693), .A2(n7692), .A3(n7691), .A4(n7690), .ZN(n9428)
         );
  NAND2_X1 U5849 ( .A1(n7678), .A2(n7677), .ZN(n9877) );
  NAND2_X1 U5850 ( .A1(n5224), .A2(n8740), .ZN(n9229) );
  NAND2_X1 U5851 ( .A1(n9236), .A2(n9237), .ZN(n5224) );
  NAND2_X1 U5852 ( .A1(n8352), .A2(n8351), .ZN(n9806) );
  AND4_X1 U5853 ( .A1(n7040), .A2(n7039), .A3(n7038), .A4(n7037), .ZN(n7337)
         );
  OAI21_X1 U5854 ( .B1(n9208), .B2(n9206), .A(n9205), .ZN(n9249) );
  AND4_X1 U5855 ( .A1(n7532), .A2(n7531), .A3(n7530), .A4(n7529), .ZN(n7985)
         );
  INV_X1 U5856 ( .A(n5241), .ZN(n5239) );
  AOI21_X1 U5857 ( .B1(n5241), .B2(n5238), .A(n9218), .ZN(n5237) );
  AND4_X1 U5858 ( .A1(n7318), .A2(n7317), .A3(n7316), .A4(n7315), .ZN(n7535)
         );
  NAND2_X1 U5859 ( .A1(n5216), .A2(n5212), .ZN(n5211) );
  INV_X1 U5860 ( .A(n5219), .ZN(n5212) );
  AND2_X1 U5861 ( .A1(n6822), .A2(n6821), .ZN(n9274) );
  AOI21_X1 U5862 ( .B1(n5227), .B2(n5226), .A(n4902), .ZN(n5225) );
  NAND2_X1 U5863 ( .A1(n8367), .A2(n6944), .ZN(n8370) );
  AND4_X1 U5864 ( .A1(n7719), .A2(n7718), .A3(n7717), .A4(n7716), .ZN(n9430)
         );
  NAND2_X1 U5865 ( .A1(n4873), .A2(P1_B_REG_SCAN_IN), .ZN(n5284) );
  NAND2_X1 U5866 ( .A1(n8379), .A2(n8378), .ZN(n9618) );
  INV_X1 U5867 ( .A(n9285), .ZN(n9631) );
  INV_X1 U5868 ( .A(n7337), .ZN(n9556) );
  INV_X1 U5869 ( .A(n7342), .ZN(n10513) );
  INV_X1 U5870 ( .A(n7249), .ZN(n10474) );
  INV_X1 U5871 ( .A(n7247), .ZN(n10515) );
  NAND2_X1 U5872 ( .A1(n6823), .A2(n6877), .ZN(n6734) );
  NAND2_X1 U5873 ( .A1(n4880), .A2(n8241), .ZN(n5172) );
  INV_X1 U5874 ( .A(n5075), .ZN(n6573) );
  NOR2_X1 U5875 ( .A1(n6667), .A2(n6331), .ZN(n10261) );
  NAND2_X1 U5876 ( .A1(n6669), .A2(n5062), .ZN(n5058) );
  NAND2_X1 U5877 ( .A1(n5060), .A2(n4920), .ZN(n5059) );
  INV_X1 U5878 ( .A(n5061), .ZN(n5060) );
  NOR2_X1 U5879 ( .A1(n6592), .A2(n6591), .ZN(n6590) );
  OR2_X1 U5880 ( .A1(n6590), .A2(n5072), .ZN(n6606) );
  NOR2_X1 U5881 ( .A1(n6590), .A2(n6340), .ZN(n6608) );
  INV_X1 U5882 ( .A(n5070), .ZN(n5069) );
  OAI21_X1 U5883 ( .B1(n5072), .B2(n6339), .A(n6341), .ZN(n5070) );
  INV_X1 U5884 ( .A(n5067), .ZN(n7377) );
  INV_X1 U5885 ( .A(n5065), .ZN(n7609) );
  NOR2_X1 U5886 ( .A1(n7796), .A2(n6349), .ZN(n7943) );
  INV_X1 U5887 ( .A(n5056), .ZN(n7941) );
  NOR2_X1 U5888 ( .A1(n8157), .A2(n8156), .ZN(n8155) );
  AND2_X1 U5889 ( .A1(n5056), .A2(n5055), .ZN(n8157) );
  NAND2_X1 U5890 ( .A1(n8063), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5055) );
  NOR2_X1 U5891 ( .A1(n10245), .A2(n5082), .ZN(n5081) );
  AND2_X1 U5892 ( .A1(n10250), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5082) );
  INV_X1 U5893 ( .A(n6355), .ZN(n5080) );
  OR2_X1 U5894 ( .A1(n6357), .A2(n6358), .ZN(n5084) );
  NAND2_X1 U5895 ( .A1(n9347), .A2(n9346), .ZN(n9778) );
  AOI21_X1 U5896 ( .B1(n9339), .B2(n6944), .A(n9338), .ZN(n9564) );
  AND2_X1 U5897 ( .A1(n9583), .A2(n9582), .ZN(n9791) );
  OAI21_X1 U5898 ( .B1(n9793), .B2(n10526), .A(n9581), .ZN(n9795) );
  NAND2_X1 U5899 ( .A1(n4978), .A2(n4979), .ZN(n9591) );
  NAND2_X1 U5900 ( .A1(n9661), .A2(n5202), .ZN(n4978) );
  AOI21_X1 U5901 ( .B1(n8405), .B2(n9764), .A(n8404), .ZN(n9804) );
  INV_X1 U5902 ( .A(n9805), .ZN(n8405) );
  NAND2_X1 U5903 ( .A1(n8403), .A2(n8402), .ZN(n8404) );
  INV_X1 U5904 ( .A(n9816), .ZN(n9648) );
  NAND2_X1 U5905 ( .A1(n5206), .A2(n8331), .ZN(n9641) );
  NAND2_X1 U5906 ( .A1(n8307), .A2(n8306), .ZN(n9828) );
  NAND2_X1 U5907 ( .A1(n9719), .A2(n8278), .ZN(n9706) );
  NAND2_X1 U5908 ( .A1(n8211), .A2(n9444), .ZN(n8381) );
  NAND2_X1 U5909 ( .A1(n7917), .A2(n5192), .ZN(n7986) );
  NOR2_X1 U5910 ( .A1(n5191), .A2(n5190), .ZN(n7988) );
  NAND2_X1 U5911 ( .A1(n4989), .A2(n4990), .ZN(n7488) );
  NAND2_X1 U5912 ( .A1(n7487), .A2(n4991), .ZN(n4989) );
  AOI21_X1 U5913 ( .B1(n7243), .B2(n7242), .A(n4864), .ZN(n10470) );
  OAI21_X1 U5914 ( .B1(n9788), .B2(n10592), .A(n5184), .ZN(n5177) );
  INV_X1 U5915 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5185) );
  AOI21_X1 U5916 ( .B1(n9786), .B2(n10477), .A(n5156), .ZN(n9787) );
  AND2_X1 U5917 ( .A1(n9785), .A2(n10549), .ZN(n5156) );
  NAND2_X1 U5918 ( .A1(n6518), .A2(n5404), .ZN(n8268) );
  XNOR2_X1 U5919 ( .A(n8224), .B(n8223), .ZN(n8778) );
  NAND2_X1 U5920 ( .A1(n5271), .A2(n6117), .ZN(n8224) );
  XNOR2_X1 U5921 ( .A(n6116), .B(n6115), .ZN(n8664) );
  AND3_X1 U5922 ( .A1(n6211), .A2(n6210), .A3(n6221), .ZN(n5264) );
  NAND2_X1 U5923 ( .A1(n6005), .A2(n6004), .ZN(n8332) );
  INV_X1 U5924 ( .A(n6698), .ZN(n9502) );
  OAI21_X1 U5925 ( .B1(n6288), .B2(n5074), .A(n6287), .ZN(n10319) );
  NAND2_X1 U5926 ( .A1(n5332), .A2(n5335), .ZN(n5331) );
  NAND2_X1 U5927 ( .A1(n5112), .A2(n5436), .ZN(n5109) );
  OAI21_X1 U5928 ( .B1(n9543), .B2(n5285), .A(n5283), .ZN(P1_U3240) );
  OR2_X1 U5929 ( .A1(n9544), .A2(n5284), .ZN(n5283) );
  NAND2_X1 U5930 ( .A1(n5020), .A2(n5018), .ZN(n5285) );
  NAND2_X1 U5931 ( .A1(n5083), .A2(n5078), .ZN(P1_U3260) );
  NAND2_X1 U5932 ( .A1(n5079), .A2(n10226), .ZN(n5078) );
  NOR2_X1 U5933 ( .A1(n6359), .A2(n5084), .ZN(n5083) );
  XNOR2_X1 U5934 ( .A(n5081), .B(n5080), .ZN(n5079) );
  OAI211_X1 U5935 ( .C1(n9788), .C2(n10498), .A(n5408), .B(n5405), .ZN(
        P1_U3355) );
  AOI21_X1 U5936 ( .B1(n9786), .B2(n10534), .A(n8695), .ZN(n5408) );
  NAND2_X1 U5937 ( .A1(n5407), .A2(n5406), .ZN(n5405) );
  NAND2_X1 U5938 ( .A1(n5154), .A2(n5153), .ZN(P1_U3552) );
  OR2_X1 U5939 ( .A1(n10591), .A2(n8675), .ZN(n5153) );
  NAND2_X1 U5940 ( .A1(n5155), .A2(n10591), .ZN(n5154) );
  OAI211_X1 U5941 ( .C1(n9863), .C2(n9789), .A(n9788), .B(n9787), .ZN(n5155)
         );
  OAI211_X1 U5942 ( .C1(n9789), .C2(n5183), .A(n5176), .B(n5175), .ZN(P1_U3520) );
  NAND2_X1 U5943 ( .A1(n10595), .A2(n10480), .ZN(n5183) );
  OR2_X1 U5944 ( .A1(n9787), .A2(n10592), .ZN(n5175) );
  INV_X1 U5945 ( .A(n5177), .ZN(n5176) );
  OR2_X1 U5946 ( .A1(n9169), .A2(n8032), .ZN(n8450) );
  AND2_X1 U5947 ( .A1(n8661), .A2(n5203), .ZN(n5202) );
  INV_X1 U5948 ( .A(n5202), .ZN(n4981) );
  AND2_X1 U5949 ( .A1(n5104), .A2(n5099), .ZN(n4860) );
  AND2_X1 U5950 ( .A1(n5437), .A2(n8526), .ZN(n4861) );
  INV_X1 U5951 ( .A(n8105), .ZN(n5252) );
  INV_X1 U5952 ( .A(n5464), .ZN(n5313) );
  AND2_X1 U5953 ( .A1(n4907), .A2(n5413), .ZN(n4862) );
  AND2_X1 U5954 ( .A1(n9443), .A2(n9422), .ZN(n4863) );
  NOR2_X1 U5955 ( .A1(n7246), .A2(n7245), .ZN(n4864) );
  OR2_X1 U5956 ( .A1(n9158), .A2(n8234), .ZN(n8447) );
  OR2_X1 U5957 ( .A1(n9485), .A2(n9492), .ZN(n4865) );
  INV_X1 U5958 ( .A(n5382), .ZN(n5381) );
  OAI22_X1 U5959 ( .A1(n8967), .A2(n5386), .B1(n8920), .B2(n9117), .ZN(n5382)
         );
  OR2_X1 U5960 ( .A1(n9539), .A2(n9697), .ZN(n4866) );
  AND2_X1 U5961 ( .A1(n9423), .A2(n9421), .ZN(n9418) );
  AND2_X1 U5962 ( .A1(n5113), .A2(n6006), .ZN(n4867) );
  AND2_X1 U5963 ( .A1(n5135), .A2(n5137), .ZN(n4868) );
  OR2_X1 U5964 ( .A1(n8030), .A2(n8035), .ZN(n4869) );
  NOR2_X1 U5965 ( .A1(n9609), .A2(n9801), .ZN(n5158) );
  NOR2_X1 U5966 ( .A1(n9609), .A2(n5160), .ZN(n5159) );
  OR2_X1 U5967 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4870) );
  INV_X1 U5968 ( .A(n7248), .ZN(n10471) );
  NAND2_X1 U5969 ( .A1(n9519), .A2(n9517), .ZN(n7248) );
  AND2_X1 U5970 ( .A1(n9625), .A2(n8331), .ZN(n5205) );
  NAND2_X1 U5971 ( .A1(n5903), .A2(n5902), .ZN(n9165) );
  NAND2_X1 U5972 ( .A1(n8667), .A2(n8666), .ZN(n9796) );
  NOR2_X1 U5973 ( .A1(n8614), .A2(n7596), .ZN(n4871) );
  AND2_X1 U5974 ( .A1(n9724), .A2(n9451), .ZN(n9449) );
  INV_X1 U5975 ( .A(n9449), .ZN(n9742) );
  AND2_X1 U5976 ( .A1(n6962), .A2(n5261), .ZN(n4872) );
  NAND2_X1 U5977 ( .A1(n8647), .A2(n8646), .ZN(n9790) );
  NAND2_X1 U5978 ( .A1(n6119), .A2(n6118), .ZN(n9105) );
  INV_X1 U5979 ( .A(n9105), .ZN(n5148) );
  OR2_X1 U5980 ( .A1(n6698), .A2(n9542), .ZN(n4873) );
  NAND3_X1 U5981 ( .A1(n6784), .A2(n6783), .A3(n6782), .ZN(n7104) );
  INV_X2 U5982 ( .A(n8763), .ZN(n6951) );
  NOR2_X1 U5983 ( .A1(n5433), .A2(n5430), .ZN(n4875) );
  AND2_X1 U5984 ( .A1(n4950), .A2(n8993), .ZN(n4876) );
  INV_X1 U5985 ( .A(n5937), .ZN(n5310) );
  OR2_X1 U5986 ( .A1(n7804), .A2(n7803), .ZN(n4877) );
  AND2_X1 U5987 ( .A1(n5260), .A2(n5258), .ZN(n4878) );
  NAND2_X1 U5988 ( .A1(n5294), .A2(n5552), .ZN(n5293) );
  OAI211_X1 U5989 ( .C1(n6694), .C2(n10319), .A(n6696), .B(n6695), .ZN(n6697)
         );
  AND2_X1 U5990 ( .A1(n9446), .A2(n9447), .ZN(n4879) );
  AND2_X1 U5991 ( .A1(n6521), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4880) );
  AND3_X1 U5992 ( .A1(n5608), .A2(n5607), .A3(n5606), .ZN(n4881) );
  NAND2_X1 U5993 ( .A1(n7206), .A2(n7205), .ZN(n4882) );
  AND4_X1 U5994 ( .A1(n6616), .A2(n6230), .A3(n6249), .A4(n6306), .ZN(n4883)
         );
  AND3_X1 U5995 ( .A1(n6638), .A2(n5174), .A3(n5172), .ZN(n4884) );
  NAND2_X1 U5996 ( .A1(n8733), .A2(n8732), .ZN(n9236) );
  OR2_X1 U5997 ( .A1(n9165), .A2(n8229), .ZN(n8528) );
  OR2_X1 U5998 ( .A1(n10149), .A2(n7776), .ZN(n8457) );
  XNOR2_X1 U5999 ( .A(n8860), .B(n10451), .ZN(n10438) );
  XNOR2_X1 U6000 ( .A(n9765), .B(n10351), .ZN(n10348) );
  INV_X1 U6001 ( .A(n10348), .ZN(n10353) );
  NAND2_X1 U6002 ( .A1(n5920), .A2(n5919), .ZN(n9158) );
  OR2_X1 U6003 ( .A1(n9138), .A2(n8551), .ZN(n4885) );
  INV_X1 U6004 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6306) );
  INV_X1 U6005 ( .A(n7506), .ZN(n5221) );
  AND4_X1 U6006 ( .A1(n5637), .A2(n5636), .A3(n5635), .A4(n5634), .ZN(n7071)
         );
  NAND2_X1 U6007 ( .A1(n5210), .A2(n6495), .ZN(n6815) );
  INV_X1 U6008 ( .A(n6815), .ZN(n6647) );
  AND2_X1 U6009 ( .A1(n8400), .A2(n8399), .ZN(n8771) );
  NAND2_X1 U6010 ( .A1(n8416), .A2(n5465), .ZN(n9031) );
  NAND2_X1 U6011 ( .A1(n8823), .A2(n5476), .ZN(n8809) );
  AND2_X1 U6012 ( .A1(n5001), .A2(n5000), .ZN(n4886) );
  INV_X1 U6013 ( .A(n7509), .ZN(n5222) );
  AND3_X1 U6014 ( .A1(n5583), .A2(n5582), .A3(n5587), .ZN(n4887) );
  INV_X1 U6015 ( .A(n8973), .ZN(n8890) );
  AND2_X1 U6016 ( .A1(n5586), .A2(n5579), .ZN(n8973) );
  AND2_X1 U6017 ( .A1(n8507), .A2(n8505), .ZN(n8613) );
  NAND2_X1 U6018 ( .A1(n8966), .A2(n8561), .ZN(n8919) );
  INV_X1 U6019 ( .A(n8919), .ZN(n5384) );
  OR2_X1 U6020 ( .A1(n7889), .A2(n7956), .ZN(n8453) );
  NAND2_X1 U6021 ( .A1(n8164), .A2(n8163), .ZN(n9848) );
  NAND2_X1 U6022 ( .A1(n8295), .A2(n8294), .ZN(n9833) );
  AND2_X1 U6023 ( .A1(n8728), .A2(n8729), .ZN(n4888) );
  AND2_X1 U6024 ( .A1(n9725), .A2(n9300), .ZN(n4889) );
  NAND2_X1 U6025 ( .A1(n8422), .A2(n8421), .ZN(n9094) );
  INV_X1 U6026 ( .A(n5158), .ZN(n5163) );
  AND2_X1 U6027 ( .A1(n5415), .A2(n9300), .ZN(n4890) );
  INV_X1 U6028 ( .A(n5108), .ZN(n5101) );
  NAND2_X1 U6029 ( .A1(n5292), .A2(n5548), .ZN(n5108) );
  AND2_X1 U6030 ( .A1(n5314), .A2(n5315), .ZN(n4891) );
  AND2_X1 U6031 ( .A1(n9462), .A2(n9463), .ZN(n9667) );
  INV_X1 U6032 ( .A(n5403), .ZN(n5402) );
  NAND2_X1 U6033 ( .A1(n5242), .A2(n5241), .ZN(n4892) );
  INV_X1 U6034 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6277) );
  AND2_X1 U6035 ( .A1(n5256), .A2(n5248), .ZN(n4893) );
  XNOR2_X1 U6036 ( .A(n5486), .B(n5485), .ZN(n5640) );
  AND2_X1 U6037 ( .A1(n8497), .A2(n8495), .ZN(n8607) );
  INV_X1 U6038 ( .A(n5159), .ZN(n5162) );
  OR2_X1 U6039 ( .A1(n5473), .A2(n5472), .ZN(n4894) );
  NAND2_X1 U6040 ( .A1(n5452), .A2(n8595), .ZN(n4895) );
  AND2_X1 U6041 ( .A1(n9132), .A2(n5113), .ZN(n4896) );
  NOR2_X1 U6042 ( .A1(n7728), .A2(n9554), .ZN(n4897) );
  NOR2_X1 U6043 ( .A1(n9871), .A2(n9551), .ZN(n4898) );
  NOR2_X1 U6044 ( .A1(n8914), .A2(n8913), .ZN(n4899) );
  NOR2_X1 U6045 ( .A1(n9110), .A2(n8944), .ZN(n4900) );
  INV_X1 U6046 ( .A(n5441), .ZN(n5439) );
  NAND2_X1 U6047 ( .A1(n8450), .A2(n4901), .ZN(n5441) );
  NAND2_X1 U6048 ( .A1(n8573), .A2(n8572), .ZN(n8956) );
  AND2_X1 U6049 ( .A1(n8451), .A2(n8453), .ZN(n4901) );
  INV_X1 U6050 ( .A(n4830), .ZN(n6190) );
  INV_X1 U6051 ( .A(n5386), .ZN(n5385) );
  NAND2_X1 U6052 ( .A1(n8989), .A2(n8997), .ZN(n5386) );
  NOR2_X1 U6053 ( .A1(n8748), .A2(n8747), .ZN(n4902) );
  INV_X1 U6054 ( .A(n5344), .ZN(n5343) );
  NAND2_X1 U6055 ( .A1(n5348), .A2(n5349), .ZN(n5344) );
  AND2_X1 U6056 ( .A1(n5553), .A2(SI_18_), .ZN(n4903) );
  AND2_X1 U6057 ( .A1(n6033), .A2(n6032), .ZN(n9035) );
  INV_X1 U6058 ( .A(n9035), .ZN(n5113) );
  INV_X1 U6059 ( .A(n5193), .ZN(n5192) );
  NAND2_X1 U6060 ( .A1(n7987), .A2(n7916), .ZN(n5193) );
  AND2_X1 U6061 ( .A1(n9445), .A2(n9444), .ZN(n9443) );
  AND2_X1 U6062 ( .A1(n9443), .A2(n9442), .ZN(n4904) );
  NAND2_X1 U6063 ( .A1(n5208), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6519) );
  INV_X1 U6064 ( .A(n9568), .ZN(n9572) );
  AND2_X1 U6065 ( .A1(n9308), .A2(n9481), .ZN(n9568) );
  AND2_X1 U6066 ( .A1(n8726), .A2(n8725), .ZN(n9218) );
  AND2_X1 U6067 ( .A1(n8771), .A2(n9594), .ZN(n4905) );
  INV_X1 U6068 ( .A(n4962), .ZN(n4961) );
  NAND2_X1 U6069 ( .A1(n8515), .A2(n8457), .ZN(n4962) );
  INV_X1 U6070 ( .A(n4965), .ZN(n4964) );
  NAND2_X1 U6071 ( .A1(n8614), .A2(n8506), .ZN(n4965) );
  INV_X1 U6072 ( .A(n5293), .ZN(n5292) );
  INV_X1 U6073 ( .A(n5200), .ZN(n5199) );
  NAND2_X1 U6074 ( .A1(n9742), .A2(n8273), .ZN(n5200) );
  INV_X1 U6075 ( .A(n5216), .ZN(n5215) );
  NAND2_X1 U6076 ( .A1(n5220), .A2(n5217), .ZN(n5216) );
  OR2_X1 U6077 ( .A1(n8390), .A2(n5419), .ZN(n4906) );
  AND2_X1 U6078 ( .A1(n6238), .A2(n6237), .ZN(n4907) );
  AND3_X1 U6079 ( .A1(n9587), .A2(n9614), .A3(n5157), .ZN(n4908) );
  AND2_X1 U6080 ( .A1(n5404), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4909) );
  AND2_X1 U6081 ( .A1(n9626), .A2(n9378), .ZN(n9651) );
  AND2_X1 U6082 ( .A1(n9375), .A2(n9374), .ZN(n9478) );
  INV_X1 U6083 ( .A(n9478), .ZN(n9595) );
  AND2_X1 U6084 ( .A1(n6522), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4910) );
  AND2_X1 U6085 ( .A1(n7338), .A2(n7336), .ZN(n4911) );
  AND2_X1 U6086 ( .A1(n9711), .A2(n9458), .ZN(n4912) );
  NOR2_X1 U6087 ( .A1(n5228), .A2(n8749), .ZN(n5227) );
  AND2_X1 U6088 ( .A1(n4882), .A2(n7080), .ZN(n4913) );
  AND2_X1 U6089 ( .A1(n8447), .A2(n8528), .ZN(n4914) );
  AND2_X1 U6090 ( .A1(n5181), .A2(n9352), .ZN(n4915) );
  AND2_X1 U6091 ( .A1(n4879), .A2(n5043), .ZN(n4916) );
  NAND2_X1 U6092 ( .A1(n5660), .A2(n5494), .ZN(n4917) );
  INV_X1 U6093 ( .A(n5468), .ZN(n5348) );
  INV_X1 U6094 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5461) );
  INV_X1 U6095 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6239) );
  AND2_X1 U6096 ( .A1(n5461), .A2(n5597), .ZN(n4918) );
  INV_X1 U6097 ( .A(n9143), .ZN(n8414) );
  NAND2_X1 U6098 ( .A1(n5964), .A2(n5963), .ZN(n9143) );
  INV_X1 U6099 ( .A(n5423), .ZN(n5422) );
  NAND2_X1 U6100 ( .A1(n9568), .A2(n9375), .ZN(n5423) );
  AND2_X1 U6101 ( .A1(n10515), .A2(n7259), .ZN(n4919) );
  OR2_X1 U6102 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10258), .ZN(n4920) );
  AND2_X1 U6103 ( .A1(n9069), .A2(n5142), .ZN(n4921) );
  NAND2_X1 U6104 ( .A1(n7783), .A2(n8616), .ZN(n7877) );
  NAND2_X1 U6105 ( .A1(n5947), .A2(n5946), .ZN(n9148) );
  INV_X1 U6106 ( .A(n9148), .ZN(n5141) );
  AND2_X1 U6107 ( .A1(n6418), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4922) );
  INV_X1 U6108 ( .A(n9205), .ZN(n5246) );
  INV_X1 U6109 ( .A(n9444), .ZN(n5412) );
  INV_X1 U6110 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U6111 ( .A1(n8370), .A2(n8369), .ZN(n9801) );
  INV_X1 U6112 ( .A(n9801), .ZN(n5161) );
  NAND2_X1 U6113 ( .A1(n8418), .A2(n8417), .ZN(n8929) );
  INV_X1 U6114 ( .A(n8929), .ZN(n5147) );
  AND2_X1 U6115 ( .A1(n8658), .A2(n8657), .ZN(n9598) );
  INV_X1 U6116 ( .A(n9598), .ZN(n5187) );
  NAND2_X1 U6117 ( .A1(n9749), .A2(n5166), .ZN(n5169) );
  AND3_X1 U6118 ( .A1(n5911), .A2(n5910), .A3(n5909), .ZN(n8229) );
  AND2_X1 U6119 ( .A1(n5201), .A2(n8273), .ZN(n4923) );
  NAND2_X1 U6120 ( .A1(n9069), .A2(n5140), .ZN(n4924) );
  AND2_X1 U6121 ( .A1(n9833), .A2(n9713), .ZN(n4925) );
  AND2_X1 U6122 ( .A1(n5357), .A2(n5355), .ZN(n4926) );
  AND2_X1 U6123 ( .A1(n7877), .A2(n5400), .ZN(n4927) );
  INV_X1 U6124 ( .A(n5128), .ZN(n5127) );
  NAND2_X1 U6125 ( .A1(n5129), .A2(n5982), .ZN(n5128) );
  OR2_X1 U6126 ( .A1(n9833), .A2(n9713), .ZN(n4928) );
  INV_X1 U6127 ( .A(n5391), .ZN(n5390) );
  AOI21_X1 U6128 ( .B1(n5392), .B2(n8918), .A(n4896), .ZN(n5391) );
  AND2_X1 U6129 ( .A1(n4920), .A2(n5062), .ZN(n4929) );
  AND2_X1 U6130 ( .A1(n8693), .A2(n8692), .ZN(n4930) );
  NAND2_X1 U6131 ( .A1(n5012), .A2(n7114), .ZN(n9504) );
  INV_X1 U6132 ( .A(n10149), .ZN(n5139) );
  INV_X1 U6133 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U6134 ( .A1(n8282), .A2(n8281), .ZN(n9837) );
  INV_X1 U6135 ( .A(n9837), .ZN(n5167) );
  NAND2_X1 U6136 ( .A1(n5867), .A2(n5866), .ZN(n10637) );
  INV_X1 U6137 ( .A(n10637), .ZN(n5135) );
  NAND2_X1 U6138 ( .A1(n7307), .A2(n7306), .ZN(n7507) );
  INV_X1 U6139 ( .A(n5266), .ZN(n6220) );
  NAND2_X1 U6140 ( .A1(n5375), .A2(n7413), .ZN(n7414) );
  INV_X1 U6141 ( .A(n9521), .ZN(n5425) );
  AND2_X1 U6142 ( .A1(n4989), .A2(n4987), .ZN(n4931) );
  AND2_X1 U6143 ( .A1(n8226), .A2(n10058), .ZN(n4932) );
  AND2_X1 U6144 ( .A1(n5218), .A2(n5220), .ZN(n4933) );
  AND2_X1 U6145 ( .A1(n7445), .A2(n8502), .ZN(n4934) );
  NAND2_X1 U6146 ( .A1(n9502), .A2(n10493), .ZN(n9488) );
  INV_X1 U6147 ( .A(n7419), .ZN(n5131) );
  INV_X1 U6148 ( .A(n7010), .ZN(n5321) );
  AND2_X2 U6149 ( .A1(n10340), .A2(n5610), .ZN(n10449) );
  AND2_X1 U6150 ( .A1(n5058), .A2(n5061), .ZN(n4935) );
  NAND2_X1 U6151 ( .A1(n8434), .A2(n8433), .ZN(n4936) );
  OR2_X1 U6152 ( .A1(n8643), .A2(n8642), .ZN(n4937) );
  AND2_X1 U6153 ( .A1(n5666), .A2(n5679), .ZN(n6430) );
  INV_X1 U6154 ( .A(n6430), .ZN(n5004) );
  INV_X1 U6155 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5003) );
  INV_X1 U6156 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6157 ( .A1(n5312), .A2(n5311), .ZN(n6021) );
  INV_X1 U6158 ( .A(n5584), .ZN(n5300) );
  NAND2_X1 U6159 ( .A1(n6883), .A2(n6882), .ZN(n6885) );
  NAND2_X1 U6160 ( .A1(n5488), .A2(n5487), .ZN(n5489) );
  NAND2_X1 U6161 ( .A1(n4944), .A2(n4942), .ZN(n5684) );
  NAND2_X1 U6162 ( .A1(n4943), .A2(n4917), .ZN(n4942) );
  NAND2_X1 U6163 ( .A1(n5662), .A2(n5494), .ZN(n4943) );
  NAND4_X1 U6164 ( .A1(n5658), .A2(n5490), .A3(n4945), .A4(n5489), .ZN(n4944)
         );
  INV_X1 U6165 ( .A(n5662), .ZN(n4945) );
  NAND2_X1 U6166 ( .A1(n5684), .A2(n5495), .ZN(n5498) );
  NAND2_X1 U6167 ( .A1(n8416), .A2(n4876), .ZN(n4946) );
  NAND2_X1 U6168 ( .A1(n4947), .A2(n4946), .ZN(n8980) );
  NAND2_X1 U6169 ( .A1(n4861), .A2(n7954), .ZN(n4959) );
  XNOR2_X1 U6170 ( .A(n5767), .B(n5471), .ZN(n7270) );
  NAND2_X1 U6171 ( .A1(n9674), .A2(n9678), .ZN(n8316) );
  NAND2_X1 U6172 ( .A1(n4999), .A2(n4911), .ZN(n7466) );
  OAI211_X2 U6173 ( .C1(n6518), .C2(n5041), .A(n5040), .B(n5037), .ZN(n6521)
         );
  NAND2_X1 U6174 ( .A1(n10353), .A2(n10352), .ZN(n5012) );
  NAND2_X1 U6175 ( .A1(n9353), .A2(n9504), .ZN(n7115) );
  NAND2_X1 U6176 ( .A1(n9510), .A2(n9509), .ZN(n9762) );
  NAND3_X1 U6177 ( .A1(n5287), .A2(n5022), .A3(n5021), .ZN(n5020) );
  NAND4_X1 U6178 ( .A1(n9503), .A2(n9533), .A3(n9502), .A4(n6234), .ZN(n5021)
         );
  NAND2_X1 U6179 ( .A1(n6518), .A2(n4909), .ZN(n5040) );
  NOR2_X1 U6180 ( .A1(n5042), .A2(n4916), .ZN(n9448) );
  OR2_X1 U6181 ( .A1(n5053), .A2(n9423), .ZN(n5050) );
  INV_X1 U6182 ( .A(n9426), .ZN(n5054) );
  NAND2_X1 U6183 ( .A1(n6669), .A2(n4929), .ZN(n5057) );
  NAND2_X1 U6184 ( .A1(n5057), .A2(n5059), .ZN(n10211) );
  NAND2_X1 U6185 ( .A1(n6592), .A2(n5071), .ZN(n5068) );
  NAND2_X1 U6186 ( .A1(n5068), .A2(n5069), .ZN(n6685) );
  NAND2_X1 U6187 ( .A1(n5715), .A2(n5501), .ZN(n5504) );
  NAND2_X1 U6188 ( .A1(n5699), .A2(n5086), .ZN(n5085) );
  MUX2_X1 U6189 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5491), .Z(n5486) );
  NAND2_X1 U6190 ( .A1(n5478), .A2(n5278), .ZN(n5087) );
  NAND2_X1 U6191 ( .A1(n5879), .A2(n4860), .ZN(n5096) );
  NAND2_X1 U6192 ( .A1(n5879), .A2(n5878), .ZN(n5103) );
  NAND3_X1 U6193 ( .A1(n5110), .A2(n4937), .A3(n5109), .ZN(P2_U3244) );
  NAND2_X1 U6194 ( .A1(n4885), .A2(n8552), .ZN(n8553) );
  NAND2_X1 U6195 ( .A1(n5268), .A2(n5124), .ZN(n5123) );
  NAND2_X1 U6196 ( .A1(n5268), .A2(n5125), .ZN(n5130) );
  NAND2_X1 U6197 ( .A1(n5268), .A2(n5962), .ZN(n5980) );
  INV_X2 U6198 ( .A(n6382), .ZN(n5917) );
  NAND2_X2 U6199 ( .A1(n6184), .A2(n8902), .ZN(n6382) );
  NOR2_X2 U6200 ( .A1(n7432), .A2(n10596), .ZN(n7454) );
  NAND2_X1 U6201 ( .A1(n5883), .A2(n5571), .ZN(n6136) );
  NAND3_X1 U6202 ( .A1(n9069), .A2(n8414), .A3(n5140), .ZN(n9043) );
  NAND2_X1 U6203 ( .A1(n8971), .A2(n5143), .ZN(n8900) );
  NAND2_X1 U6204 ( .A1(n8971), .A2(n8955), .ZN(n8950) );
  NAND2_X1 U6205 ( .A1(n5266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6206 ( .A1(n6220), .A2(n4862), .ZN(n6516) );
  NAND2_X1 U6207 ( .A1(n9633), .A2(n4908), .ZN(n9583) );
  NAND2_X1 U6208 ( .A1(n9633), .A2(n9614), .ZN(n9609) );
  INV_X1 U6209 ( .A(n5169), .ZN(n9707) );
  NAND4_X1 U6210 ( .A1(n5267), .A2(n5171), .A3(n6208), .A4(n4883), .ZN(n5266)
         );
  NAND3_X1 U6211 ( .A1(n5170), .A2(n5265), .A3(n5264), .ZN(n6217) );
  NAND2_X1 U6212 ( .A1(n8241), .A2(n4910), .ZN(n5174) );
  AOI21_X1 U6213 ( .B1(n9571), .B2(n5180), .A(n4915), .ZN(n5179) );
  OR2_X1 U6214 ( .A1(n10595), .A2(n5185), .ZN(n5184) );
  AOI21_X1 U6215 ( .B1(n7248), .B2(n4864), .A(n4919), .ZN(n5194) );
  NAND2_X1 U6216 ( .A1(n9661), .A2(n8330), .ZN(n5206) );
  INV_X2 U6217 ( .A(n6516), .ZN(n6518) );
  NOR2_X1 U6218 ( .A1(n7749), .A2(n6490), .ZN(n5210) );
  XNOR2_X1 U6219 ( .A(n6233), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6646) );
  NAND3_X1 U6220 ( .A1(n7307), .A2(n7306), .A3(n5222), .ZN(n5218) );
  NAND3_X1 U6221 ( .A1(n7307), .A2(n7306), .A3(n5214), .ZN(n5213) );
  NAND2_X1 U6222 ( .A1(n5223), .A2(n5225), .ZN(n9279) );
  OAI211_X1 U6223 ( .C1(n9191), .C2(n5235), .A(n5232), .B(n5229), .ZN(n8774)
         );
  NAND2_X1 U6224 ( .A1(n9191), .A2(n5230), .ZN(n5229) );
  NOR2_X1 U6225 ( .A1(n8767), .A2(n5231), .ZN(n5230) );
  OAI21_X1 U6226 ( .B1(n8767), .B2(n5234), .A(n5233), .ZN(n5232) );
  NAND2_X1 U6227 ( .A1(n8767), .A2(n8759), .ZN(n5233) );
  AND2_X1 U6228 ( .A1(n9190), .A2(n8759), .ZN(n5234) );
  NAND2_X1 U6229 ( .A1(n8767), .A2(n5236), .ZN(n5235) );
  INV_X1 U6230 ( .A(n5247), .ZN(n9258) );
  NAND2_X1 U6231 ( .A1(n7805), .A2(n4877), .ZN(n5259) );
  NAND2_X1 U6232 ( .A1(n7805), .A2(n5250), .ZN(n5249) );
  AND2_X1 U6233 ( .A1(n4883), .A2(n6212), .ZN(n5265) );
  AND2_X1 U6234 ( .A1(n5490), .A2(n5489), .ZN(n5659) );
  NAND2_X1 U6235 ( .A1(n6116), .A2(n5272), .ZN(n5270) );
  NAND2_X1 U6236 ( .A1(n6116), .A2(n6115), .ZN(n5271) );
  OR2_X1 U6237 ( .A1(n5478), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6238 ( .A1(n5527), .A2(n5282), .ZN(n5281) );
  NAND2_X1 U6239 ( .A1(n5528), .A2(n5281), .ZN(n5822) );
  OAI21_X1 U6240 ( .B1(n5899), .B2(n5549), .A(n5551), .ZN(n5915) );
  NAND2_X1 U6241 ( .A1(n5549), .A2(n5551), .ZN(n5294) );
  NAND3_X1 U6242 ( .A1(n9343), .A2(n5297), .A3(n5296), .ZN(n5295) );
  NAND3_X1 U6243 ( .A1(n9568), .A2(n5474), .A3(n9478), .ZN(n5298) );
  NAND2_X1 U6244 ( .A1(n5301), .A2(n5315), .ZN(n5312) );
  INV_X1 U6245 ( .A(n5306), .ZN(n5301) );
  NAND2_X1 U6246 ( .A1(n5938), .A2(n5303), .ZN(n5302) );
  NAND2_X1 U6247 ( .A1(n5306), .A2(n5313), .ZN(n5304) );
  NAND3_X1 U6248 ( .A1(n5317), .A2(n5316), .A3(n5697), .ZN(n6984) );
  OAI21_X1 U6249 ( .B1(n5322), .B2(n5321), .A(n6995), .ZN(n5320) );
  NOR2_X1 U6250 ( .A1(n7011), .A2(n5323), .ZN(n5322) );
  NAND2_X4 U6251 ( .A1(n5327), .A2(n8433), .ZN(n6127) );
  OAI211_X1 U6252 ( .C1(n8782), .C2(n5331), .A(n5328), .B(n6202), .ZN(P2_U3222) );
  NAND2_X1 U6253 ( .A1(n8782), .A2(n5329), .ZN(n5328) );
  NAND2_X1 U6254 ( .A1(n7003), .A2(n5337), .ZN(n5336) );
  OR2_X1 U6255 ( .A1(n5346), .A2(n5468), .ZN(n5341) );
  INV_X1 U6256 ( .A(n5897), .ZN(n5359) );
  NAND2_X1 U6257 ( .A1(n8809), .A2(n5362), .ZN(n5361) );
  NAND2_X1 U6258 ( .A1(n8230), .A2(n5364), .ZN(n5363) );
  NAND2_X1 U6259 ( .A1(n5363), .A2(n5366), .ZN(n9063) );
  NAND2_X2 U6260 ( .A1(n5375), .A2(n5373), .ZN(n10574) );
  NAND2_X1 U6261 ( .A1(n8978), .A2(n5379), .ZN(n5377) );
  NAND2_X1 U6262 ( .A1(n5387), .A2(n4913), .ZN(n7208) );
  NAND2_X1 U6263 ( .A1(n7079), .A2(n5477), .ZN(n5387) );
  NAND2_X1 U6264 ( .A1(n9024), .A2(n5392), .ZN(n5389) );
  NAND2_X1 U6265 ( .A1(n7783), .A2(n5399), .ZN(n5396) );
  NAND2_X1 U6266 ( .A1(n5396), .A2(n5397), .ZN(n8021) );
  NOR2_X1 U6267 ( .A1(n10622), .A2(n7882), .ZN(n5403) );
  INV_X1 U6268 ( .A(n9765), .ZN(n7113) );
  NAND2_X1 U6269 ( .A1(n9765), .A2(n6951), .ZN(n6710) );
  NAND2_X2 U6270 ( .A1(n4884), .A2(n6639), .ZN(n9765) );
  NAND2_X1 U6271 ( .A1(n9711), .A2(n5414), .ZN(n9675) );
  NAND2_X2 U6272 ( .A1(n9725), .A2(n4890), .ZN(n9711) );
  INV_X1 U6273 ( .A(n9705), .ZN(n5415) );
  NAND2_X1 U6274 ( .A1(n9668), .A2(n5418), .ZN(n5417) );
  OAI21_X1 U6275 ( .B1(n8686), .B2(n5423), .A(n5421), .ZN(n8687) );
  NAND2_X1 U6276 ( .A1(n8686), .A2(n9478), .ZN(n9600) );
  OAI21_X2 U6277 ( .B1(n9391), .B2(n5426), .A(n5424), .ZN(n9328) );
  XNOR2_X1 U6278 ( .A(n8432), .B(n8973), .ZN(n5435) );
  INV_X1 U6279 ( .A(n8644), .ZN(n5436) );
  NOR2_X1 U6280 ( .A1(n7954), .A2(n7953), .ZN(n8036) );
  NAND2_X1 U6281 ( .A1(n8979), .A2(n8440), .ZN(n5452) );
  NAND2_X1 U6282 ( .A1(n8979), .A2(n5443), .ZN(n5442) );
  NAND2_X1 U6283 ( .A1(n10436), .A2(n5456), .ZN(n5454) );
  NAND2_X1 U6284 ( .A1(n5454), .A2(n5453), .ZN(n7209) );
  INV_X1 U6285 ( .A(n5601), .ZN(n5598) );
  NAND3_X1 U6286 ( .A1(n5883), .A2(n4918), .A3(n5571), .ZN(n5601) );
  NAND2_X1 U6287 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  XNOR2_X1 U6288 ( .A(n6100), .B(n6099), .ZN(n8367) );
  MUX2_X1 U6289 ( .A(n9884), .B(P1_REG1_REG_28__SCAN_IN), .S(n10589), .Z(
        P1_U3551) );
  MUX2_X1 U6290 ( .A(n9884), .B(P1_REG0_REG_28__SCAN_IN), .S(n10592), .Z(
        P1_U3519) );
  AOI21_X2 U6291 ( .B1(n7674), .B2(n7673), .A(n7672), .ZN(n7706) );
  INV_X1 U6292 ( .A(n9596), .ZN(n8686) );
  INV_X1 U6293 ( .A(n10392), .ZN(n6760) );
  AOI21_X1 U6294 ( .B1(n8431), .B2(n8435), .A(n8436), .ZN(n8432) );
  AOI21_X2 U6295 ( .B1(n8172), .B2(n8174), .A(n8173), .ZN(n8704) );
  XNOR2_X1 U6296 ( .A(n8761), .B(n8730), .ZN(n5462) );
  NOR2_X1 U6297 ( .A1(n5976), .A2(n8798), .ZN(n5464) );
  OR2_X1 U6298 ( .A1(n8414), .A2(n9056), .ZN(n5465) );
  AND2_X1 U6299 ( .A1(n5148), .A2(n8958), .ZN(n5466) );
  OR2_X1 U6300 ( .A1(n5147), .A2(n10638), .ZN(n5467) );
  AND2_X1 U6301 ( .A1(n5752), .A2(n5751), .ZN(n5468) );
  AND2_X1 U6302 ( .A1(n5804), .A2(n5803), .ZN(n5469) );
  AND2_X1 U6303 ( .A1(n5533), .A2(n5532), .ZN(n5470) );
  AND2_X1 U6304 ( .A1(n5768), .A2(n5513), .ZN(n5471) );
  AND2_X1 U6305 ( .A1(n9801), .A2(n9618), .ZN(n5472) );
  AND4_X1 U6306 ( .A1(n9475), .A2(n9617), .A3(n9370), .A4(n9629), .ZN(n5474)
         );
  INV_X1 U6307 ( .A(n7356), .ZN(n7083) );
  AND2_X1 U6308 ( .A1(n7082), .A2(n7081), .ZN(n5475) );
  OR2_X1 U6309 ( .A1(n7086), .A2(n7185), .ZN(n5477) );
  NAND2_X1 U6310 ( .A1(n6958), .A2(n7029), .ZN(n6965) );
  INV_X1 U6311 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U6312 ( .A1(n7074), .A2(n10420), .ZN(n8471) );
  NAND2_X1 U6313 ( .A1(n6647), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6653) );
  INV_X1 U6314 ( .A(n8355), .ZN(n8353) );
  INV_X1 U6315 ( .A(n7491), .ZN(n6922) );
  INV_X1 U6316 ( .A(n5793), .ZN(n5524) );
  INV_X1 U6317 ( .A(n5848), .ZN(n5847) );
  INV_X1 U6318 ( .A(n5922), .ZN(n5921) );
  OR2_X1 U6319 ( .A1(n5905), .A2(n5904), .ZN(n5922) );
  INV_X1 U6320 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U6321 ( .A1(n8353), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8372) );
  INV_X1 U6322 ( .A(n8177), .ZN(n6926) );
  INV_X1 U6323 ( .A(n9401), .ZN(n7338) );
  AND2_X1 U6324 ( .A1(n5541), .A2(n5858), .ZN(n5542) );
  INV_X1 U6325 ( .A(SI_8_), .ZN(n10039) );
  INV_X1 U6326 ( .A(n6087), .ZN(n6086) );
  NAND2_X1 U6327 ( .A1(n6043), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6065) );
  OR2_X1 U6328 ( .A1(n5965), .A2(n10112), .ZN(n5988) );
  NAND2_X1 U6329 ( .A1(n4831), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5635) );
  AND2_X1 U6330 ( .A1(n8641), .A2(n8636), .ZN(n6183) );
  INV_X1 U6331 ( .A(n8921), .ZN(n8923) );
  NAND2_X1 U6332 ( .A1(n5948), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5965) );
  INV_X1 U6333 ( .A(n8619), .ZN(n7881) );
  INV_X1 U6334 ( .A(n7714), .ZN(n6924) );
  AND2_X1 U6335 ( .A1(n4829), .A2(n6871), .ZN(n6846) );
  OR2_X1 U6336 ( .A1(n8372), .A2(n8371), .ZN(n8649) );
  OR2_X1 U6337 ( .A1(n8340), .A2(n9238), .ZN(n8355) );
  INV_X1 U6338 ( .A(n6800), .ZN(n8676) );
  OR2_X1 U6339 ( .A1(n8297), .A2(n8296), .ZN(n8309) );
  NAND2_X1 U6340 ( .A1(n9546), .A2(n9559), .ZN(n8692) );
  INV_X1 U6341 ( .A(n9418), .ZN(n7900) );
  NAND2_X1 U6342 ( .A1(n8244), .A2(n8243), .ZN(n8248) );
  NAND2_X1 U6343 ( .A1(n6086), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6121) );
  OR2_X1 U6344 ( .A1(n5945), .A2(n5613), .ZN(n5615) );
  OR2_X1 U6345 ( .A1(n6065), .A2(n8816), .ZN(n6087) );
  AND2_X1 U6346 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  NAND2_X1 U6347 ( .A1(n6076), .A2(n6075), .ZN(n6077) );
  INV_X1 U6348 ( .A(n6183), .ZN(n6761) );
  OR2_X1 U6349 ( .A1(n5988), .A2(n8839), .ZN(n6026) );
  INV_X1 U6350 ( .A(n9122), .ZN(n8989) );
  INV_X1 U6351 ( .A(n10638), .ZN(n10150) );
  NAND2_X1 U6352 ( .A1(n6924), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U6353 ( .A1(n6921), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7285) );
  AND2_X1 U6354 ( .A1(n7671), .A2(n7670), .ZN(n7672) );
  OR2_X1 U6355 ( .A1(n7285), .A2(n7284), .ZN(n7313) );
  OR2_X1 U6356 ( .A1(n7688), .A2(n7687), .ZN(n7714) );
  AND2_X1 U6358 ( .A1(n8649), .A2(n8373), .ZN(n9281) );
  INV_X1 U6359 ( .A(n9790), .ZN(n9587) );
  INV_X1 U6360 ( .A(n8401), .ZN(n8402) );
  OR2_X1 U6361 ( .A1(n6715), .A2(n6727), .ZN(n9745) );
  INV_X1 U6362 ( .A(n9697), .ZN(n10493) );
  XNOR2_X1 U6363 ( .A(n5540), .B(n5534), .ZN(n5837) );
  AND2_X1 U6364 ( .A1(n6748), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8820) );
  OAI22_X1 U6365 ( .A1(n7371), .A2(n7370), .B1(n5783), .B2(n5782), .ZN(n7390)
         );
  INV_X1 U6366 ( .A(n10397), .ZN(n8844) );
  OR2_X1 U6367 ( .A1(n6761), .A2(n6184), .ZN(n10439) );
  AND2_X1 U6368 ( .A1(n6051), .A2(n6050), .ZN(n8813) );
  AND4_X1 U6369 ( .A1(n5817), .A2(n5816), .A3(n5815), .A4(n5814), .ZN(n7776)
         );
  INV_X1 U6370 ( .A(n8896), .ZN(n10301) );
  INV_X1 U6371 ( .A(n8956), .ZN(n8948) );
  INV_X1 U6372 ( .A(n8918), .ZN(n9033) );
  INV_X1 U6373 ( .A(n10439), .ZN(n9080) );
  AND2_X1 U6374 ( .A1(n7154), .A2(n7153), .ZN(n10461) );
  NAND2_X1 U6375 ( .A1(n7450), .A2(n6764), .ZN(n10644) );
  AND2_X1 U6376 ( .A1(n5746), .A2(n5745), .ZN(n6459) );
  INV_X1 U6377 ( .A(n9274), .ZN(n9280) );
  AND2_X1 U6378 ( .A1(n8679), .A2(n8678), .ZN(n9578) );
  AND2_X1 U6379 ( .A1(n8184), .A2(n8183), .ZN(n9746) );
  INV_X1 U6380 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n6317) );
  INV_X1 U6381 ( .A(n8393), .ZN(n9617) );
  AND2_X1 U6382 ( .A1(n9411), .A2(n9412), .ZN(n9409) );
  AND2_X1 U6383 ( .A1(n10539), .A2(n7106), .ZN(n10534) );
  AND2_X1 U6384 ( .A1(n6632), .A2(n9903), .ZN(n7639) );
  OR2_X1 U6385 ( .A1(n9488), .A2(n9538), .ZN(n10552) );
  INV_X1 U6386 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6286) );
  INV_X1 U6387 ( .A(n7889), .ZN(n10630) );
  INV_X1 U6388 ( .A(n7771), .ZN(n10622) );
  INV_X1 U6389 ( .A(n8957), .ZN(n8920) );
  NAND2_X1 U6390 ( .A1(n4833), .A2(n7148), .ZN(n9089) );
  INV_X1 U6391 ( .A(n10646), .ZN(n10645) );
  INV_X1 U6392 ( .A(n10650), .ZN(n10647) );
  AND2_X1 U6393 ( .A1(n6366), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10274) );
  INV_X1 U6394 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6533) );
  INV_X1 U6395 ( .A(n9287), .ZN(n9224) );
  OR2_X1 U6396 ( .A1(n6819), .A2(n6719), .ZN(n9289) );
  INV_X1 U6397 ( .A(n8771), .ZN(n9576) );
  INV_X1 U6398 ( .A(n7535), .ZN(n9554) );
  NAND2_X1 U6399 ( .A1(n7263), .A2(n10488), .ZN(n10539) );
  INV_X1 U6400 ( .A(n10591), .ZN(n10589) );
  INV_X1 U6401 ( .A(n10595), .ZN(n10592) );
  AND2_X1 U6402 ( .A1(n6815), .A2(n6489), .ZN(n6728) );
  INV_X1 U6403 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6530) );
  NAND3_X1 U6404 ( .A1(n5479), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5481) );
  AND2_X1 U6405 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U6406 ( .A1(n5491), .A2(n5480), .ZN(n6636) );
  NAND2_X1 U6407 ( .A1(n5481), .A2(n6636), .ZN(n5483) );
  INV_X1 U6408 ( .A(SI_1_), .ZN(n5482) );
  XNOR2_X1 U6409 ( .A(n5483), .B(n5482), .ZN(n5612) );
  MUX2_X1 U6410 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5491), .Z(n5611) );
  NAND2_X1 U6411 ( .A1(n5612), .A2(n5611), .ZN(n5639) );
  NAND2_X1 U6412 ( .A1(n5483), .A2(SI_1_), .ZN(n5638) );
  NAND2_X1 U6413 ( .A1(n5486), .A2(SI_2_), .ZN(n5487) );
  AND2_X1 U6414 ( .A1(n5638), .A2(n5487), .ZN(n5484) );
  NAND2_X1 U6415 ( .A1(n5639), .A2(n5484), .ZN(n5490) );
  INV_X1 U6416 ( .A(SI_2_), .ZN(n5485) );
  INV_X1 U6417 ( .A(n5640), .ZN(n5488) );
  MUX2_X1 U6418 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5491), .Z(n5493) );
  INV_X1 U6419 ( .A(SI_3_), .ZN(n9988) );
  XNOR2_X1 U6420 ( .A(n5493), .B(n9988), .ZN(n5658) );
  MUX2_X1 U6421 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5491), .Z(n5492) );
  XNOR2_X1 U6422 ( .A(n5492), .B(SI_4_), .ZN(n5662) );
  NAND2_X1 U6423 ( .A1(n5492), .A2(SI_4_), .ZN(n5494) );
  NAND2_X1 U6424 ( .A1(n5493), .A2(SI_3_), .ZN(n5660) );
  MUX2_X1 U6425 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5491), .Z(n5496) );
  XNOR2_X1 U6426 ( .A(n5496), .B(SI_5_), .ZN(n5683) );
  INV_X1 U6427 ( .A(n5683), .ZN(n5495) );
  NAND2_X1 U6428 ( .A1(n5496), .A2(SI_5_), .ZN(n5497) );
  MUX2_X1 U6429 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8257), .Z(n5499) );
  NAND2_X1 U6430 ( .A1(n5499), .A2(SI_6_), .ZN(n5500) );
  MUX2_X1 U6431 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8257), .Z(n5502) );
  NAND2_X1 U6432 ( .A1(n5502), .A2(SI_7_), .ZN(n5503) );
  INV_X1 U6433 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5505) );
  MUX2_X1 U6434 ( .A(n6512), .B(n5505), .S(n8257), .Z(n5506) );
  INV_X1 U6435 ( .A(n5506), .ZN(n5507) );
  NAND2_X1 U6436 ( .A1(n5507), .A2(SI_8_), .ZN(n5508) );
  INV_X1 U6437 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6513) );
  INV_X1 U6438 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5510) );
  MUX2_X1 U6439 ( .A(n6513), .B(n5510), .S(n8257), .Z(n5511) );
  INV_X1 U6440 ( .A(SI_9_), .ZN(n10086) );
  INV_X1 U6441 ( .A(n5511), .ZN(n5512) );
  NAND2_X1 U6442 ( .A1(n5512), .A2(SI_9_), .ZN(n5513) );
  MUX2_X1 U6443 ( .A(n6533), .B(n6530), .S(n8257), .Z(n5514) );
  INV_X1 U6444 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U6445 ( .A1(n5515), .A2(SI_10_), .ZN(n5516) );
  NAND2_X1 U6446 ( .A1(n5767), .A2(n5517), .ZN(n5521) );
  INV_X1 U6447 ( .A(n5770), .ZN(n5518) );
  MUX2_X1 U6448 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n8257), .Z(n5522) );
  NAND2_X1 U6449 ( .A1(n5522), .A2(SI_11_), .ZN(n5523) );
  MUX2_X1 U6450 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n8257), .Z(n5525) );
  INV_X1 U6451 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6740) );
  INV_X1 U6452 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5529) );
  MUX2_X1 U6453 ( .A(n6740), .B(n5529), .S(n8257), .Z(n5530) );
  INV_X1 U6454 ( .A(SI_13_), .ZN(n9949) );
  NAND2_X1 U6455 ( .A1(n5530), .A2(n9949), .ZN(n5533) );
  INV_X1 U6456 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U6457 ( .A1(n5531), .A2(SI_13_), .ZN(n5532) );
  MUX2_X1 U6458 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n8257), .Z(n5540) );
  INV_X1 U6459 ( .A(SI_14_), .ZN(n5534) );
  INV_X1 U6460 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6939) );
  INV_X1 U6461 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5536) );
  MUX2_X1 U6462 ( .A(n6939), .B(n5536), .S(n8257), .Z(n5537) );
  INV_X1 U6463 ( .A(SI_15_), .ZN(n9968) );
  NAND2_X1 U6464 ( .A1(n5537), .A2(n9968), .ZN(n5543) );
  INV_X1 U6465 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U6466 ( .A1(n5538), .A2(SI_15_), .ZN(n5539) );
  NAND2_X1 U6467 ( .A1(n5543), .A2(n5539), .ZN(n5860) );
  INV_X1 U6468 ( .A(n5860), .ZN(n5541) );
  NAND2_X1 U6469 ( .A1(n5540), .A2(SI_14_), .ZN(n5858) );
  INV_X1 U6470 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6942) );
  INV_X1 U6471 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6941) );
  MUX2_X1 U6472 ( .A(n6942), .B(n6941), .S(n8257), .Z(n5545) );
  INV_X1 U6473 ( .A(SI_16_), .ZN(n10071) );
  NAND2_X1 U6474 ( .A1(n5545), .A2(n10071), .ZN(n5548) );
  INV_X1 U6475 ( .A(n5545), .ZN(n5546) );
  NAND2_X1 U6476 ( .A1(n5546), .A2(SI_16_), .ZN(n5547) );
  MUX2_X1 U6477 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n8257), .Z(n5550) );
  INV_X1 U6478 ( .A(SI_17_), .ZN(n10070) );
  XNOR2_X1 U6479 ( .A(n5550), .B(n10070), .ZN(n5898) );
  INV_X1 U6480 ( .A(n5898), .ZN(n5549) );
  NAND2_X1 U6481 ( .A1(n5550), .A2(SI_17_), .ZN(n5551) );
  MUX2_X1 U6482 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n8257), .Z(n5553) );
  XNOR2_X1 U6483 ( .A(n5553), .B(SI_18_), .ZN(n5914) );
  INV_X1 U6484 ( .A(n5914), .ZN(n5552) );
  INV_X1 U6485 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7141) );
  INV_X1 U6486 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5554) );
  MUX2_X1 U6487 ( .A(n7141), .B(n5554), .S(n8257), .Z(n5555) );
  INV_X1 U6488 ( .A(SI_19_), .ZN(n10048) );
  NAND2_X1 U6489 ( .A1(n5555), .A2(n10048), .ZN(n5939) );
  INV_X1 U6490 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U6491 ( .A1(n5556), .A2(SI_19_), .ZN(n5557) );
  NAND2_X1 U6492 ( .A1(n5939), .A2(n5557), .ZN(n5940) );
  XNOR2_X1 U6493 ( .A(n5941), .B(n5940), .ZN(n8279) );
  NAND2_X1 U6494 ( .A1(n5558), .A2(n5591), .ZN(n5665) );
  NAND4_X1 U6495 ( .A1(n5561), .A2(n5560), .A3(n5716), .A4(n5795), .ZN(n5565)
         );
  INV_X1 U6496 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5563) );
  NAND4_X1 U6497 ( .A1(n5563), .A2(n5842), .A3(n5743), .A4(n5562), .ZN(n5564)
         );
  NOR2_X1 U6498 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5568) );
  NOR2_X1 U6499 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5567) );
  NAND4_X1 U6500 ( .A1(n5568), .A2(n5567), .A3(n5587), .A4(n5582), .ZN(n5570)
         );
  NAND4_X1 U6501 ( .A1(n5589), .A2(n6143), .A3(n6169), .A4(n6147), .ZN(n5569)
         );
  NAND2_X1 U6502 ( .A1(n6136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5573) );
  MUX2_X1 U6503 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5573), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5575) );
  NAND2_X1 U6504 ( .A1(n6382), .A2(n4832), .ZN(n5648) );
  NAND2_X1 U6506 ( .A1(n8279), .A2(n5657), .ZN(n5581) );
  INV_X2 U6507 ( .A(n5945), .ZN(n5918) );
  INV_X1 U6508 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U6509 ( .A1(n5584), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5916) );
  INV_X1 U6510 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U6511 ( .A1(n5916), .A2(n5583), .ZN(n5577) );
  NAND2_X1 U6512 ( .A1(n5577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U6513 ( .A1(n5578), .A2(n5582), .ZN(n5586) );
  OR2_X1 U6514 ( .A1(n5578), .A2(n5582), .ZN(n5579) );
  AOI22_X1 U6515 ( .A1(n4859), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8973), .B2(
        n5917), .ZN(n5580) );
  INV_X1 U6516 ( .A(n9155), .ZN(n8914) );
  INV_X1 U6517 ( .A(n6133), .ZN(n5585) );
  INV_X1 U6518 ( .A(n8423), .ZN(n8636) );
  XNOR2_X1 U6519 ( .A(n8914), .B(n6127), .ZN(n5937) );
  XNOR2_X1 U6520 ( .A(n5659), .B(n5658), .ZN(n6781) );
  NAND2_X1 U6521 ( .A1(n4859), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5596) );
  NOR2_X1 U6522 ( .A1(n5591), .A2(n8262), .ZN(n5643) );
  INV_X1 U6523 ( .A(n5643), .ZN(n5593) );
  INV_X1 U6524 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U6525 ( .A1(n5593), .A2(n5592), .ZN(n5644) );
  NAND2_X1 U6526 ( .A1(n5644), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5594) );
  XNOR2_X1 U6527 ( .A(n5594), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6403) );
  NAND2_X1 U6528 ( .A1(n5917), .A2(n6403), .ZN(n5595) );
  OAI211_X1 U6529 ( .C1(n5648), .C2(n6781), .A(n5596), .B(n5595), .ZN(n7237)
         );
  INV_X1 U6530 ( .A(n7237), .ZN(n10420) );
  XNOR2_X1 U6531 ( .A(n6127), .B(n10420), .ZN(n5655) );
  NAND2_X1 U6532 ( .A1(n5598), .A2(n5602), .ZN(n8263) );
  INV_X1 U6533 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5599) );
  XNOR2_X2 U6534 ( .A(n5600), .B(n5599), .ZN(n5605) );
  NAND2_X1 U6535 ( .A1(n5601), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5603) );
  INV_X1 U6536 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5602) );
  INV_X1 U6537 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6362) );
  OR2_X1 U6538 ( .A1(n5633), .A2(n6362), .ZN(n5608) );
  NAND2_X2 U6539 ( .A1(n5605), .A2(n8227), .ZN(n5720) );
  INV_X1 U6540 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6374) );
  OR2_X1 U6541 ( .A1(n5720), .A2(n6374), .ZN(n5607) );
  NAND2_X1 U6542 ( .A1(n4830), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5606) );
  OR2_X1 U6543 ( .A1(n5620), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U6544 ( .A1(n7074), .A2(n4858), .ZN(n5656) );
  XNOR2_X1 U6545 ( .A(n5612), .B(n5611), .ZN(n8412) );
  INV_X1 U6546 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U6547 ( .A1(n5917), .A2(n10292), .ZN(n5614) );
  OAI211_X2 U6548 ( .C1(n5648), .C2(n8412), .A(n5615), .B(n5614), .ZN(n6768)
         );
  XNOR2_X1 U6549 ( .A(n6127), .B(n10378), .ZN(n5629) );
  NAND2_X1 U6550 ( .A1(n6584), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5619) );
  INV_X1 U6551 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10372) );
  OR2_X1 U6552 ( .A1(n5620), .A2(n10372), .ZN(n5618) );
  INV_X1 U6553 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6372) );
  OR2_X1 U6554 ( .A1(n5720), .A2(n6372), .ZN(n5617) );
  INV_X1 U6555 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6360) );
  OR2_X1 U6556 ( .A1(n5633), .A2(n6360), .ZN(n5616) );
  AND4_X2 U6557 ( .A1(n5619), .A2(n5618), .A3(n5617), .A4(n5616), .ZN(n10392)
         );
  NAND2_X1 U6558 ( .A1(n6760), .A2(n4857), .ZN(n5631) );
  XNOR2_X1 U6559 ( .A(n5629), .B(n5631), .ZN(n6751) );
  INV_X1 U6560 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10283) );
  OR2_X1 U6561 ( .A1(n5620), .A2(n10283), .ZN(n5625) );
  INV_X1 U6562 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10277) );
  OR2_X1 U6563 ( .A1(n5720), .A2(n10277), .ZN(n5624) );
  INV_X1 U6564 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5621) );
  OR2_X1 U6565 ( .A1(n5633), .A2(n5621), .ZN(n5623) );
  NAND2_X1 U6566 ( .A1(n4831), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5622) );
  NAND4_X1 U6567 ( .A1(n5625), .A2(n5624), .A3(n5623), .A4(n5622), .ZN(n8862)
         );
  NAND2_X1 U6568 ( .A1(n4832), .A2(SI_0_), .ZN(n5626) );
  XNOR2_X1 U6569 ( .A(n5626), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9189) );
  MUX2_X1 U6570 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9189), .S(n6382), .Z(n10339)
         );
  NAND2_X1 U6571 ( .A1(n8862), .A2(n10339), .ZN(n7066) );
  INV_X1 U6572 ( .A(n7066), .ZN(n5627) );
  NAND2_X1 U6573 ( .A1(n5627), .A2(n4858), .ZN(n6914) );
  INV_X1 U6574 ( .A(n10339), .ZN(n7144) );
  NAND2_X1 U6575 ( .A1(n6127), .A2(n7144), .ZN(n5628) );
  AND2_X1 U6576 ( .A1(n6914), .A2(n5628), .ZN(n6750) );
  NAND2_X1 U6577 ( .A1(n6751), .A2(n6750), .ZN(n6749) );
  INV_X1 U6578 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U6579 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  NAND2_X1 U6580 ( .A1(n6749), .A2(n5632), .ZN(n10396) );
  INV_X1 U6581 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10403) );
  OR2_X1 U6582 ( .A1(n5620), .A2(n10403), .ZN(n5637) );
  NAND2_X1 U6583 ( .A1(n6536), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5636) );
  INV_X1 U6584 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6361) );
  OR2_X1 U6585 ( .A1(n5633), .A2(n6361), .ZN(n5634) );
  NAND2_X1 U6586 ( .A1(n5639), .A2(n5638), .ZN(n5641) );
  XNOR2_X1 U6587 ( .A(n5641), .B(n5640), .ZN(n6693) );
  INV_X1 U6588 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U6589 ( .A1(n5643), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U6590 ( .A1(n5917), .A2(n10307), .ZN(n5646) );
  OAI211_X1 U6591 ( .C1(n5648), .C2(n6693), .A(n5647), .B(n5646), .ZN(n7366)
         );
  XNOR2_X1 U6592 ( .A(n6127), .B(n10405), .ZN(n5650) );
  NAND2_X1 U6593 ( .A1(n5649), .A2(n5650), .ZN(n5654) );
  INV_X1 U6594 ( .A(n5649), .ZN(n5652) );
  INV_X1 U6595 ( .A(n5650), .ZN(n5651) );
  NAND2_X1 U6596 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  NAND2_X1 U6597 ( .A1(n5654), .A2(n5653), .ZN(n10395) );
  OAI21_X1 U6598 ( .B1(n10396), .B2(n10395), .A(n5654), .ZN(n6883) );
  XNOR2_X1 U6599 ( .A(n5656), .B(n5655), .ZN(n6882) );
  NAND2_X1 U6600 ( .A1(n5659), .A2(n5658), .ZN(n5661) );
  NAND2_X1 U6601 ( .A1(n5661), .A2(n5660), .ZN(n5663) );
  XNOR2_X1 U6602 ( .A(n5663), .B(n5662), .ZN(n6807) );
  NAND2_X1 U6603 ( .A1(n5657), .A2(n6807), .ZN(n5669) );
  NAND2_X1 U6604 ( .A1(n5918), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U6605 ( .A1(n5665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5664) );
  MUX2_X1 U6606 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5664), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5666) );
  OR2_X1 U6607 ( .A1(n5665), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U6608 ( .A1(n5917), .A2(n6430), .ZN(n5667) );
  XNOR2_X1 U6609 ( .A(n6129), .B(n10451), .ZN(n5677) );
  INV_X1 U6610 ( .A(n5677), .ZN(n5675) );
  NAND2_X1 U6611 ( .A1(n4831), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5673) );
  XNOR2_X1 U6612 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7014) );
  OR2_X1 U6613 ( .A1(n5620), .A2(n7014), .ZN(n5672) );
  NAND2_X1 U6614 ( .A1(n6535), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U6615 ( .A1(n6536), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U6616 ( .A1(n8860), .A2(n4858), .ZN(n5676) );
  INV_X1 U6617 ( .A(n5676), .ZN(n5674) );
  AND2_X1 U6618 ( .A1(n5675), .A2(n5674), .ZN(n7011) );
  NAND2_X1 U6619 ( .A1(n5677), .A2(n5676), .ZN(n7010) );
  INV_X1 U6620 ( .A(n5678), .ZN(n5682) );
  NAND2_X1 U6621 ( .A1(n5679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5680) );
  MUX2_X1 U6622 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5680), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5681) );
  NAND2_X1 U6623 ( .A1(n5682), .A2(n5681), .ZN(n6485) );
  XNOR2_X1 U6624 ( .A(n5684), .B(n5683), .ZN(n6850) );
  NAND2_X1 U6625 ( .A1(n6850), .A2(n5657), .ZN(n5686) );
  NAND2_X1 U6626 ( .A1(n4859), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5685) );
  OAI211_X1 U6627 ( .C1(n6382), .C2(n6485), .A(n5686), .B(n5685), .ZN(n7185)
         );
  INV_X1 U6628 ( .A(n7185), .ZN(n10501) );
  XNOR2_X1 U6629 ( .A(n10501), .B(n6127), .ZN(n5695) );
  NAND2_X1 U6630 ( .A1(n6535), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5693) );
  NAND3_X1 U6631 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5704) );
  INV_X1 U6632 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U6633 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5687) );
  NAND2_X1 U6634 ( .A1(n5688), .A2(n5687), .ZN(n5689) );
  NAND2_X1 U6635 ( .A1(n5704), .A2(n5689), .ZN(n7183) );
  OR2_X1 U6636 ( .A1(n5620), .A2(n7183), .ZN(n5692) );
  NAND2_X1 U6637 ( .A1(n4830), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U6638 ( .A1(n6536), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5690) );
  NAND4_X1 U6639 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .ZN(n7086)
         );
  AND2_X1 U6640 ( .A1(n7086), .A2(n4858), .ZN(n5694) );
  NOR2_X1 U6641 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  AOI21_X1 U6642 ( .B1(n5695), .B2(n5694), .A(n5696), .ZN(n6995) );
  INV_X1 U6643 ( .A(n5696), .ZN(n5697) );
  XNOR2_X1 U6644 ( .A(n5699), .B(n5698), .ZN(n6945) );
  NAND2_X1 U6645 ( .A1(n6945), .A2(n5657), .ZN(n5702) );
  OR2_X1 U6646 ( .A1(n5678), .A2(n8262), .ZN(n5700) );
  XNOR2_X1 U6647 ( .A(n5700), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6418) );
  AOI22_X1 U6648 ( .A1(n5918), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5917), .B2(
        n6418), .ZN(n5701) );
  NAND2_X1 U6649 ( .A1(n5702), .A2(n5701), .ZN(n7205) );
  INV_X1 U6650 ( .A(n7205), .ZN(n7216) );
  XNOR2_X1 U6651 ( .A(n7216), .B(n6127), .ZN(n5711) );
  NAND2_X1 U6652 ( .A1(n6535), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5709) );
  INV_X1 U6653 ( .A(n5704), .ZN(n5703) );
  INV_X1 U6654 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10137) );
  NAND2_X1 U6655 ( .A1(n5704), .A2(n10137), .ZN(n5705) );
  NAND2_X1 U6656 ( .A1(n5723), .A2(n5705), .ZN(n7160) );
  OR2_X1 U6657 ( .A1(n6089), .A2(n7160), .ZN(n5708) );
  NAND2_X1 U6658 ( .A1(n4830), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6659 ( .A1(n6536), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5706) );
  NAND4_X1 U6660 ( .A1(n5709), .A2(n5708), .A3(n5707), .A4(n5706), .ZN(n7206)
         );
  INV_X1 U6661 ( .A(n7206), .ZN(n7215) );
  NOR2_X1 U6662 ( .A1(n7215), .A2(n6911), .ZN(n5710) );
  NOR2_X1 U6663 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  AOI21_X1 U6664 ( .B1(n5711), .B2(n5710), .A(n5712), .ZN(n6985) );
  NAND2_X1 U6665 ( .A1(n6984), .A2(n6985), .ZN(n6983) );
  INV_X1 U6666 ( .A(n5712), .ZN(n5713) );
  NAND2_X1 U6667 ( .A1(n6983), .A2(n5713), .ZN(n7003) );
  XNOR2_X1 U6668 ( .A(n5715), .B(n5714), .ZN(n7022) );
  NAND2_X1 U6669 ( .A1(n7022), .A2(n5657), .ZN(n5719) );
  NAND2_X1 U6670 ( .A1(n5678), .A2(n5716), .ZN(n5741) );
  NAND2_X1 U6671 ( .A1(n5741), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5717) );
  XNOR2_X1 U6672 ( .A(n5717), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6444) );
  AOI22_X1 U6673 ( .A1(n5918), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5917), .B2(
        n6444), .ZN(n5718) );
  NAND2_X1 U6674 ( .A1(n5719), .A2(n5718), .ZN(n7411) );
  XNOR2_X1 U6675 ( .A(n7411), .B(n6127), .ZN(n5731) );
  NAND2_X1 U6676 ( .A1(n6535), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5729) );
  INV_X1 U6677 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6419) );
  OR2_X1 U6678 ( .A1(n5720), .A2(n6419), .ZN(n5728) );
  INV_X1 U6679 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U6680 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  NAND2_X1 U6681 ( .A1(n5733), .A2(n5724), .ZN(n7220) );
  OR2_X1 U6682 ( .A1(n6089), .A2(n7220), .ZN(n5727) );
  INV_X1 U6683 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5725) );
  OR2_X1 U6684 ( .A1(n6190), .A2(n5725), .ZN(n5726) );
  INV_X1 U6685 ( .A(n7403), .ZN(n7412) );
  NAND2_X1 U6686 ( .A1(n7412), .A2(n8434), .ZN(n5730) );
  XNOR2_X1 U6687 ( .A(n5731), .B(n5730), .ZN(n7004) );
  NAND2_X1 U6688 ( .A1(n4831), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5738) );
  INV_X1 U6689 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7407) );
  OR2_X1 U6690 ( .A1(n5633), .A2(n7407), .ZN(n5737) );
  INV_X1 U6691 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U6692 ( .A1(n5733), .A2(n7048), .ZN(n5734) );
  NAND2_X1 U6693 ( .A1(n5757), .A2(n5734), .ZN(n7406) );
  OR2_X1 U6694 ( .A1(n6089), .A2(n7406), .ZN(n5736) );
  INV_X1 U6695 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6445) );
  OR2_X1 U6696 ( .A1(n5720), .A2(n6445), .ZN(n5735) );
  INV_X1 U6697 ( .A(n7397), .ZN(n7423) );
  NAND2_X1 U6698 ( .A1(n7423), .A2(n8434), .ZN(n5750) );
  XNOR2_X1 U6699 ( .A(n5740), .B(n5739), .ZN(n7277) );
  NAND2_X1 U6700 ( .A1(n7277), .A2(n5657), .ZN(n5748) );
  INV_X1 U6701 ( .A(n5773), .ZN(n5746) );
  NAND2_X1 U6702 ( .A1(n5742), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5744) );
  MUX2_X1 U6703 ( .A(n5744), .B(P2_IR_REG_31__SCAN_IN), .S(n5743), .Z(n5745)
         );
  AOI22_X1 U6704 ( .A1(n5918), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5917), .B2(
        n6459), .ZN(n5747) );
  NAND2_X1 U6705 ( .A1(n5748), .A2(n5747), .ZN(n7419) );
  XNOR2_X1 U6706 ( .A(n7419), .B(n6127), .ZN(n5749) );
  XOR2_X1 U6707 ( .A(n5750), .B(n5749), .Z(n7046) );
  INV_X1 U6708 ( .A(n5749), .ZN(n5752) );
  INV_X1 U6709 ( .A(n5750), .ZN(n5751) );
  OR2_X1 U6710 ( .A1(n5773), .A2(n8262), .ZN(n5753) );
  XNOR2_X1 U6711 ( .A(n5753), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6472) );
  AOI22_X1 U6712 ( .A1(n5918), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5917), .B2(
        n6472), .ZN(n5754) );
  XNOR2_X1 U6713 ( .A(n10596), .B(n6129), .ZN(n5764) );
  NAND2_X1 U6714 ( .A1(n6535), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5762) );
  INV_X1 U6715 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5755) );
  OR2_X1 U6716 ( .A1(n6190), .A2(n5755), .ZN(n5761) );
  NAND2_X1 U6717 ( .A1(n5757), .A2(n5756), .ZN(n5758) );
  NAND2_X1 U6718 ( .A1(n5776), .A2(n5758), .ZN(n7431) );
  OR2_X1 U6719 ( .A1(n5620), .A2(n7431), .ZN(n5760) );
  INV_X1 U6720 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6460) );
  OR2_X1 U6721 ( .A1(n5720), .A2(n6460), .ZN(n5759) );
  NOR2_X1 U6722 ( .A1(n7446), .A2(n6911), .ZN(n5763) );
  NOR2_X1 U6723 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  AOI21_X1 U6724 ( .B1(n5764), .B2(n5763), .A(n5765), .ZN(n7167) );
  INV_X1 U6725 ( .A(n5765), .ZN(n5766) );
  NAND2_X1 U6726 ( .A1(n5767), .A2(n5471), .ZN(n5769) );
  NAND2_X1 U6727 ( .A1(n5769), .A2(n5768), .ZN(n5771) );
  XNOR2_X1 U6728 ( .A(n5771), .B(n5770), .ZN(n7482) );
  NAND2_X1 U6729 ( .A1(n7482), .A2(n5657), .ZN(n5775) );
  INV_X1 U6730 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U6731 ( .A1(n5773), .A2(n5772), .ZN(n5806) );
  NAND2_X1 U6732 ( .A1(n5806), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5796) );
  XNOR2_X1 U6733 ( .A(n5796), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7195) );
  AOI22_X1 U6734 ( .A1(n5918), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5917), .B2(
        n7195), .ZN(n5774) );
  NAND2_X1 U6735 ( .A1(n5775), .A2(n5774), .ZN(n7575) );
  XNOR2_X1 U6736 ( .A(n7575), .B(n6127), .ZN(n5783) );
  NAND2_X1 U6737 ( .A1(n4831), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5781) );
  INV_X1 U6738 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7452) );
  OR2_X1 U6739 ( .A1(n5633), .A2(n7452), .ZN(n5780) );
  NAND2_X1 U6740 ( .A1(n5776), .A2(n10105), .ZN(n5777) );
  NAND2_X1 U6741 ( .A1(n5786), .A2(n5777), .ZN(n7451) );
  OR2_X1 U6742 ( .A1(n6089), .A2(n7451), .ZN(n5779) );
  INV_X1 U6743 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6473) );
  OR2_X1 U6744 ( .A1(n5720), .A2(n6473), .ZN(n5778) );
  INV_X1 U6745 ( .A(n7442), .ZN(n8859) );
  NAND2_X1 U6746 ( .A1(n8859), .A2(n8434), .ZN(n5782) );
  XNOR2_X1 U6747 ( .A(n5783), .B(n5782), .ZN(n7370) );
  NAND2_X1 U6748 ( .A1(n6536), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5792) );
  INV_X1 U6749 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7580) );
  OR2_X1 U6750 ( .A1(n5633), .A2(n7580), .ZN(n5791) );
  INV_X1 U6751 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U6752 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  NAND2_X1 U6753 ( .A1(n5812), .A2(n5787), .ZN(n7579) );
  OR2_X1 U6754 ( .A1(n6089), .A2(n7579), .ZN(n5790) );
  INV_X1 U6755 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5788) );
  OR2_X1 U6756 ( .A1(n6190), .A2(n5788), .ZN(n5789) );
  INV_X1 U6757 ( .A(n7627), .ZN(n8858) );
  NAND2_X1 U6758 ( .A1(n8858), .A2(n8434), .ZN(n5802) );
  XNOR2_X1 U6759 ( .A(n5794), .B(n5793), .ZN(n7521) );
  NAND2_X1 U6760 ( .A1(n7521), .A2(n5657), .ZN(n5800) );
  NAND2_X1 U6761 ( .A1(n5796), .A2(n5795), .ZN(n5797) );
  NAND2_X1 U6762 ( .A1(n5797), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5798) );
  XNOR2_X1 U6763 ( .A(n5798), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7546) );
  AOI22_X1 U6764 ( .A1(n5918), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7546), .B2(
        n5917), .ZN(n5799) );
  XNOR2_X1 U6765 ( .A(n10612), .B(n6127), .ZN(n5801) );
  XOR2_X1 U6766 ( .A(n5802), .B(n5801), .Z(n7389) );
  INV_X1 U6767 ( .A(n5801), .ZN(n5804) );
  INV_X1 U6768 ( .A(n5802), .ZN(n5803) );
  XNOR2_X1 U6769 ( .A(n5805), .B(SI_12_), .ZN(n7675) );
  NAND2_X1 U6770 ( .A1(n7675), .A2(n5657), .ZN(n5809) );
  NAND2_X1 U6771 ( .A1(n5823), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5807) );
  XNOR2_X1 U6772 ( .A(n5807), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7567) );
  AOI22_X1 U6773 ( .A1(n5918), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5917), .B2(
        n7567), .ZN(n5808) );
  XNOR2_X1 U6774 ( .A(n10149), .B(n6129), .ZN(n5819) );
  NAND2_X1 U6775 ( .A1(n4830), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5817) );
  INV_X1 U6776 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5810) );
  OR2_X1 U6777 ( .A1(n5633), .A2(n5810), .ZN(n5816) );
  INV_X1 U6778 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10117) );
  NAND2_X1 U6779 ( .A1(n5812), .A2(n10117), .ZN(n5813) );
  NAND2_X1 U6780 ( .A1(n5827), .A2(n5813), .ZN(n7626) );
  OR2_X1 U6781 ( .A1(n5620), .A2(n7626), .ZN(n5815) );
  INV_X1 U6782 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7547) );
  OR2_X1 U6783 ( .A1(n5720), .A2(n7547), .ZN(n5814) );
  NOR2_X1 U6784 ( .A1(n7776), .A2(n6911), .ZN(n5818) );
  NOR2_X1 U6785 ( .A1(n5819), .A2(n5818), .ZN(n5820) );
  AOI21_X1 U6786 ( .B1(n5819), .B2(n5818), .A(n5820), .ZN(n7622) );
  NAND2_X1 U6787 ( .A1(n7623), .A2(n7622), .ZN(n7621) );
  INV_X1 U6788 ( .A(n5820), .ZN(n5821) );
  NAND2_X1 U6789 ( .A1(n7621), .A2(n5821), .ZN(n7661) );
  XNOR2_X1 U6790 ( .A(n5822), .B(n5470), .ZN(n7707) );
  NAND2_X1 U6791 ( .A1(n7707), .A2(n5657), .ZN(n5825) );
  OAI21_X1 U6792 ( .B1(n5823), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U6793 ( .A(n5840), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7650) );
  AOI22_X1 U6794 ( .A1(n5918), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7650), .B2(
        n5917), .ZN(n5824) );
  XNOR2_X1 U6795 ( .A(n7771), .B(n6129), .ZN(n5834) );
  NAND2_X1 U6796 ( .A1(n4831), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5832) );
  INV_X1 U6797 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7780) );
  OR2_X1 U6798 ( .A1(n5633), .A2(n7780), .ZN(n5831) );
  INV_X1 U6799 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7544) );
  OR2_X1 U6800 ( .A1(n5720), .A2(n7544), .ZN(n5830) );
  INV_X1 U6801 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U6802 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  NAND2_X1 U6803 ( .A1(n5848), .A2(n5828), .ZN(n7770) );
  OR2_X1 U6804 ( .A1(n5620), .A2(n7770), .ZN(n5829) );
  NOR2_X1 U6805 ( .A1(n7882), .A2(n6911), .ZN(n5833) );
  NOR2_X1 U6806 ( .A1(n5834), .A2(n5833), .ZN(n5835) );
  AOI21_X1 U6807 ( .B1(n5834), .B2(n5833), .A(n5835), .ZN(n7662) );
  NAND2_X1 U6808 ( .A1(n7661), .A2(n7662), .ZN(n7660) );
  INV_X1 U6809 ( .A(n5835), .ZN(n5836) );
  NAND2_X1 U6810 ( .A1(n7660), .A2(n5836), .ZN(n7741) );
  XNOR2_X1 U6811 ( .A(n5838), .B(n5837), .ZN(n7806) );
  NAND2_X1 U6812 ( .A1(n7806), .A2(n5657), .ZN(n5846) );
  INV_X1 U6813 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U6814 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  NAND2_X1 U6815 ( .A1(n5841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U6816 ( .A1(n5843), .A2(n5842), .ZN(n5862) );
  OR2_X1 U6817 ( .A1(n5843), .A2(n5842), .ZN(n5844) );
  AOI22_X1 U6818 ( .A1(n7973), .A2(n5917), .B1(n5918), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5845) );
  XNOR2_X1 U6819 ( .A(n7889), .B(n6129), .ZN(n5855) );
  NAND2_X1 U6820 ( .A1(n4831), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5853) );
  INV_X1 U6821 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7887) );
  OR2_X1 U6822 ( .A1(n5633), .A2(n7887), .ZN(n5852) );
  INV_X1 U6823 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7651) );
  OR2_X1 U6824 ( .A1(n5720), .A2(n7651), .ZN(n5851) );
  INV_X1 U6825 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U6826 ( .A1(n5848), .A2(n10037), .ZN(n5849) );
  NAND2_X1 U6827 ( .A1(n5869), .A2(n5849), .ZN(n7886) );
  OR2_X1 U6828 ( .A1(n5620), .A2(n7886), .ZN(n5850) );
  NOR2_X1 U6829 ( .A1(n7956), .A2(n6911), .ZN(n5854) );
  NOR2_X1 U6830 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  AOI21_X1 U6831 ( .B1(n5855), .B2(n5854), .A(n5856), .ZN(n7742) );
  INV_X1 U6832 ( .A(n5856), .ZN(n5857) );
  NAND2_X1 U6833 ( .A1(n5859), .A2(n5858), .ZN(n5861) );
  NAND2_X1 U6834 ( .A1(n8057), .A2(n5657), .ZN(n5867) );
  NAND2_X1 U6835 ( .A1(n5862), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5864) );
  INV_X1 U6836 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5863) );
  XNOR2_X1 U6837 ( .A(n5864), .B(n5863), .ZN(n8015) );
  OAI22_X1 U6838 ( .A1(n8015), .A2(n6382), .B1(n5945), .B2(n6939), .ZN(n5865)
         );
  INV_X1 U6839 ( .A(n5865), .ZN(n5866) );
  XNOR2_X1 U6840 ( .A(n10637), .B(n6129), .ZN(n5877) );
  NAND2_X1 U6841 ( .A1(n4831), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5875) );
  INV_X1 U6842 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7958) );
  OR2_X1 U6843 ( .A1(n5633), .A2(n7958), .ZN(n5874) );
  INV_X1 U6844 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U6845 ( .A1(n5869), .A2(n5868), .ZN(n5870) );
  NAND2_X1 U6846 ( .A1(n5888), .A2(n5870), .ZN(n7957) );
  OR2_X1 U6847 ( .A1(n6089), .A2(n7957), .ZN(n5873) );
  INV_X1 U6848 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5871) );
  OR2_X1 U6849 ( .A1(n5720), .A2(n5871), .ZN(n5872) );
  NOR2_X1 U6850 ( .A1(n7952), .A2(n6911), .ZN(n5876) );
  NOR2_X1 U6851 ( .A1(n5877), .A2(n5876), .ZN(n7753) );
  NAND2_X1 U6852 ( .A1(n5877), .A2(n5876), .ZN(n7754) );
  XNOR2_X1 U6853 ( .A(n5879), .B(n5878), .ZN(n8062) );
  NAND2_X1 U6854 ( .A1(n8062), .A2(n5657), .ZN(n5886) );
  AND2_X1 U6855 ( .A1(n5678), .A2(n5880), .ZN(n5881) );
  NOR2_X1 U6856 ( .A1(n5881), .A2(n8262), .ZN(n5882) );
  MUX2_X1 U6857 ( .A(n8262), .B(n5882), .S(P2_IR_REG_16__SCAN_IN), .Z(n5884)
         );
  OR2_X1 U6858 ( .A1(n5884), .A2(n5883), .ZN(n7969) );
  INV_X1 U6859 ( .A(n7969), .ZN(n8195) );
  AOI22_X1 U6860 ( .A1(n5918), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5917), .B2(
        n8195), .ZN(n5885) );
  XNOR2_X1 U6861 ( .A(n9169), .B(n6127), .ZN(n5896) );
  NAND2_X1 U6862 ( .A1(n4830), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5894) );
  INV_X1 U6863 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U6864 ( .A1(n5888), .A2(n10014), .ZN(n5889) );
  NAND2_X1 U6865 ( .A1(n5905), .A2(n5889), .ZN(n8046) );
  OR2_X1 U6866 ( .A1(n8046), .A2(n6089), .ZN(n5893) );
  INV_X1 U6867 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5890) );
  OR2_X1 U6868 ( .A1(n5633), .A2(n5890), .ZN(n5892) );
  INV_X1 U6869 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7968) );
  OR2_X1 U6870 ( .A1(n5720), .A2(n7968), .ZN(n5891) );
  INV_X1 U6871 ( .A(n8032), .ZN(n8855) );
  NAND2_X1 U6872 ( .A1(n8855), .A2(n8434), .ZN(n5895) );
  XNOR2_X1 U6873 ( .A(n5896), .B(n5895), .ZN(n7831) );
  XNOR2_X1 U6874 ( .A(n5899), .B(n5898), .ZN(n8161) );
  NAND2_X1 U6875 ( .A1(n8161), .A2(n5657), .ZN(n5903) );
  INV_X1 U6876 ( .A(n5883), .ZN(n5900) );
  NAND2_X1 U6877 ( .A1(n5900), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5901) );
  XNOR2_X1 U6878 ( .A(n5901), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8875) );
  AOI22_X1 U6879 ( .A1(n4859), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5917), .B2(
        n8875), .ZN(n5902) );
  XNOR2_X1 U6880 ( .A(n9165), .B(n6127), .ZN(n5913) );
  INV_X1 U6881 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U6882 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  AND2_X1 U6883 ( .A1(n5922), .A2(n5906), .ZN(n8026) );
  NAND2_X1 U6884 ( .A1(n8026), .A2(n6192), .ZN(n5911) );
  NAND2_X1 U6885 ( .A1(n4831), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U6886 ( .A1(n6535), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5907) );
  AND2_X1 U6887 ( .A1(n5908), .A2(n5907), .ZN(n5910) );
  NAND2_X1 U6888 ( .A1(n6536), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5909) );
  OR2_X1 U6889 ( .A1(n8229), .A2(n6911), .ZN(n5912) );
  NAND2_X1 U6890 ( .A1(n5913), .A2(n5912), .ZN(n7932) );
  NOR2_X1 U6891 ( .A1(n5913), .A2(n5912), .ZN(n7934) );
  XNOR2_X1 U6892 ( .A(n5915), .B(n5914), .ZN(n8275) );
  NAND2_X1 U6893 ( .A1(n8275), .A2(n5657), .ZN(n5920) );
  XNOR2_X1 U6894 ( .A(n5916), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8886) );
  AOI22_X1 U6895 ( .A1(n5918), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5917), .B2(
        n8886), .ZN(n5919) );
  XNOR2_X1 U6896 ( .A(n9158), .B(n6127), .ZN(n5930) );
  INV_X1 U6897 ( .A(n5930), .ZN(n5928) );
  INV_X1 U6898 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U6899 ( .A1(n5922), .A2(n10134), .ZN(n5923) );
  NAND2_X1 U6900 ( .A1(n5932), .A2(n5923), .ZN(n9073) );
  OR2_X1 U6901 ( .A1(n9073), .A2(n5620), .ZN(n5926) );
  AOI22_X1 U6902 ( .A1(n4830), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n6535), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n5925) );
  INV_X1 U6903 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8863) );
  OR2_X1 U6904 ( .A1(n5720), .A2(n8863), .ZN(n5924) );
  OR2_X1 U6905 ( .A1(n8234), .A2(n6911), .ZN(n5929) );
  INV_X1 U6906 ( .A(n5929), .ZN(n5927) );
  NAND2_X1 U6907 ( .A1(n5928), .A2(n5927), .ZN(n8138) );
  AND2_X1 U6908 ( .A1(n5930), .A2(n5929), .ZN(n8139) );
  INV_X1 U6909 ( .A(n8131), .ZN(n5938) );
  INV_X1 U6910 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U6911 ( .A1(n5932), .A2(n5931), .ZN(n5933) );
  AND2_X1 U6912 ( .A1(n5950), .A2(n5933), .ZN(n8132) );
  INV_X1 U6913 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U6914 ( .A1(n4830), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U6915 ( .A1(n6536), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5934) );
  OAI211_X1 U6916 ( .C1(n5633), .C2(n8887), .A(n5935), .B(n5934), .ZN(n5936)
         );
  AOI21_X1 U6917 ( .B1(n8132), .B2(n6192), .A(n5936), .ZN(n8913) );
  NOR2_X1 U6918 ( .A1(n8913), .A2(n6911), .ZN(n8129) );
  INV_X1 U6919 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7396) );
  INV_X1 U6920 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8293) );
  MUX2_X1 U6921 ( .A(n7396), .B(n8293), .S(n8257), .Z(n5942) );
  INV_X1 U6922 ( .A(SI_20_), .ZN(n10042) );
  NAND2_X1 U6923 ( .A1(n5942), .A2(n10042), .ZN(n5962) );
  INV_X1 U6924 ( .A(n5942), .ZN(n5943) );
  NAND2_X1 U6925 ( .A1(n5943), .A2(SI_20_), .ZN(n5944) );
  XNOR2_X1 U6926 ( .A(n5961), .B(n5960), .ZN(n8292) );
  NAND2_X1 U6927 ( .A1(n8292), .A2(n5657), .ZN(n5947) );
  NAND2_X1 U6928 ( .A1(n5918), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5946) );
  XNOR2_X1 U6929 ( .A(n9148), .B(n6127), .ZN(n5959) );
  INV_X1 U6930 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U6931 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  NAND2_X1 U6932 ( .A1(n5965), .A2(n5951), .ZN(n9060) );
  OR2_X1 U6933 ( .A1(n9060), .A2(n6089), .ZN(n5957) );
  INV_X1 U6934 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U6935 ( .A1(n6536), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U6936 ( .A1(n6535), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5952) );
  OAI211_X1 U6937 ( .C1(n6190), .C2(n5954), .A(n5953), .B(n5952), .ZN(n5955)
         );
  INV_X1 U6938 ( .A(n5955), .ZN(n5956) );
  NAND2_X1 U6939 ( .A1(n5957), .A2(n5956), .ZN(n9050) );
  NAND2_X1 U6940 ( .A1(n9050), .A2(n8434), .ZN(n5958) );
  NOR2_X1 U6941 ( .A1(n5959), .A2(n5958), .ZN(n5975) );
  AOI21_X1 U6942 ( .B1(n5959), .B2(n5958), .A(n5975), .ZN(n8831) );
  MUX2_X1 U6943 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n8257), .Z(n5981) );
  INV_X1 U6944 ( .A(SI_21_), .ZN(n10043) );
  XNOR2_X1 U6945 ( .A(n5981), .B(n10043), .ZN(n5978) );
  XNOR2_X1 U6946 ( .A(n5980), .B(n5978), .ZN(n8305) );
  NAND2_X1 U6947 ( .A1(n8305), .A2(n5657), .ZN(n5964) );
  NAND2_X1 U6948 ( .A1(n5918), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U6949 ( .A(n9143), .B(n6127), .ZN(n5974) );
  INV_X1 U6950 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10112) );
  NAND2_X1 U6951 ( .A1(n5965), .A2(n10112), .ZN(n5966) );
  NAND2_X1 U6952 ( .A1(n5988), .A2(n5966), .ZN(n8803) );
  OR2_X1 U6953 ( .A1(n8803), .A2(n6089), .ZN(n5972) );
  INV_X1 U6954 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U6955 ( .A1(n6536), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U6956 ( .A1(n6535), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5967) );
  OAI211_X1 U6957 ( .C1(n6190), .C2(n5969), .A(n5968), .B(n5967), .ZN(n5970)
         );
  INV_X1 U6958 ( .A(n5970), .ZN(n5971) );
  NAND2_X1 U6959 ( .A1(n5972), .A2(n5971), .ZN(n9056) );
  NAND2_X1 U6960 ( .A1(n9056), .A2(n8434), .ZN(n5973) );
  AOI21_X1 U6961 ( .B1(n5974), .B2(n5973), .A(n6014), .ZN(n8801) );
  AND2_X1 U6962 ( .A1(n8831), .A2(n8801), .ZN(n5977) );
  INV_X1 U6963 ( .A(n8801), .ZN(n5976) );
  INV_X1 U6964 ( .A(n5975), .ZN(n8798) );
  INV_X1 U6965 ( .A(n6014), .ZN(n6012) );
  NAND2_X1 U6966 ( .A1(n8799), .A2(n6012), .ZN(n8837) );
  INV_X1 U6967 ( .A(n5978), .ZN(n5979) );
  NAND2_X1 U6968 ( .A1(n5981), .A2(SI_21_), .ZN(n5982) );
  INV_X1 U6969 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7620) );
  INV_X1 U6970 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8318) );
  MUX2_X1 U6971 ( .A(n7620), .B(n8318), .S(n8257), .Z(n5983) );
  INV_X1 U6972 ( .A(SI_22_), .ZN(n10049) );
  NAND2_X1 U6973 ( .A1(n5983), .A2(n10049), .ZN(n6036) );
  INV_X1 U6974 ( .A(n5983), .ZN(n5984) );
  NAND2_X1 U6975 ( .A1(n5984), .A2(SI_22_), .ZN(n5985) );
  NAND2_X1 U6976 ( .A1(n6036), .A2(n5985), .ZN(n5995) );
  XNOR2_X1 U6977 ( .A(n5996), .B(n5995), .ZN(n8317) );
  NAND2_X1 U6978 ( .A1(n8317), .A2(n5657), .ZN(n5987) );
  NAND2_X1 U6979 ( .A1(n5918), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5986) );
  XNOR2_X1 U6980 ( .A(n9138), .B(n6127), .ZN(n6010) );
  INV_X1 U6981 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U6982 ( .A1(n5988), .A2(n8839), .ZN(n5989) );
  NAND2_X1 U6983 ( .A1(n6026), .A2(n5989), .ZN(n9027) );
  INV_X1 U6984 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U6985 ( .A1(n6536), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U6986 ( .A1(n6535), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5990) );
  OAI211_X1 U6987 ( .C1(n6190), .C2(n5992), .A(n5991), .B(n5990), .ZN(n5993)
         );
  INV_X1 U6988 ( .A(n5993), .ZN(n5994) );
  OAI21_X1 U6989 ( .B1(n9027), .B2(n5620), .A(n5994), .ZN(n9049) );
  NAND2_X1 U6990 ( .A1(n9049), .A2(n8434), .ZN(n6011) );
  XNOR2_X1 U6991 ( .A(n6010), .B(n6011), .ZN(n8838) );
  INV_X1 U6992 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5997) );
  INV_X1 U6993 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8333) );
  MUX2_X1 U6994 ( .A(n5997), .B(n8333), .S(n8257), .Z(n5998) );
  INV_X1 U6995 ( .A(SI_23_), .ZN(n10046) );
  NAND2_X1 U6996 ( .A1(n5998), .A2(n10046), .ZN(n6035) );
  INV_X1 U6997 ( .A(n5998), .ZN(n5999) );
  NAND2_X1 U6998 ( .A1(n5999), .A2(SI_23_), .ZN(n6037) );
  NAND2_X1 U6999 ( .A1(n6035), .A2(n6037), .ZN(n6001) );
  NAND2_X1 U7000 ( .A1(n6000), .A2(n6001), .ZN(n6005) );
  INV_X1 U7001 ( .A(n6000), .ZN(n6003) );
  INV_X1 U7002 ( .A(n6001), .ZN(n6002) );
  NAND2_X1 U7003 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U7004 ( .A1(n4859), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6006) );
  XNOR2_X1 U7005 ( .A(n9132), .B(n6129), .ZN(n6009) );
  NAND2_X1 U7006 ( .A1(n6010), .A2(n6011), .ZN(n6017) );
  NAND2_X1 U7007 ( .A1(n6009), .A2(n6017), .ZN(n6034) );
  NOR2_X1 U7008 ( .A1(n8799), .A2(n6034), .ZN(n6023) );
  INV_X1 U7009 ( .A(n6011), .ZN(n6015) );
  INV_X1 U7010 ( .A(n6010), .ZN(n6007) );
  AOI211_X1 U7011 ( .C1(n6015), .C2(n6007), .A(n6014), .B(n6009), .ZN(n6008)
         );
  INV_X1 U7012 ( .A(n6009), .ZN(n6018) );
  AOI21_X1 U7013 ( .B1(n6012), .B2(n6011), .A(n6010), .ZN(n6013) );
  AOI211_X1 U7014 ( .C1(n6015), .C2(n6014), .A(n6018), .B(n6013), .ZN(n6016)
         );
  AOI21_X1 U7015 ( .B1(n6018), .B2(n6017), .A(n6016), .ZN(n6019) );
  INV_X1 U7016 ( .A(n6019), .ZN(n6020) );
  NAND2_X1 U7017 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  NOR2_X2 U7018 ( .A1(n6023), .A2(n6022), .ZN(n8790) );
  INV_X1 U7019 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U7020 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  NAND2_X1 U7021 ( .A1(n6044), .A2(n6027), .ZN(n8793) );
  OR2_X1 U7022 ( .A1(n8793), .A2(n5620), .ZN(n6033) );
  INV_X1 U7023 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7024 ( .A1(n6535), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7025 ( .A1(n6536), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6028) );
  OAI211_X1 U7026 ( .C1(n6030), .C2(n6190), .A(n6029), .B(n6028), .ZN(n6031)
         );
  INV_X1 U7027 ( .A(n6031), .ZN(n6032) );
  NOR2_X1 U7028 ( .A1(n9035), .A2(n6911), .ZN(n8792) );
  NAND2_X1 U7029 ( .A1(n8790), .A2(n8792), .ZN(n8791) );
  OAI21_X1 U7030 ( .B1(n8836), .B2(n6034), .A(n8791), .ZN(n6052) );
  AND2_X1 U7031 ( .A1(n6036), .A2(n6035), .ZN(n6039) );
  INV_X1 U7032 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7750) );
  INV_X1 U7033 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8337) );
  MUX2_X1 U7034 ( .A(n7750), .B(n8337), .S(n8257), .Z(n6057) );
  XNOR2_X1 U7035 ( .A(n6057), .B(SI_24_), .ZN(n6056) );
  XNOR2_X1 U7036 ( .A(n6055), .B(n6056), .ZN(n8336) );
  NAND2_X1 U7037 ( .A1(n8336), .A2(n5657), .ZN(n6042) );
  NAND2_X1 U7038 ( .A1(n4859), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6041) );
  XNOR2_X1 U7039 ( .A(n9005), .B(n6127), .ZN(n6053) );
  XNOR2_X1 U7040 ( .A(n6052), .B(n6053), .ZN(n8825) );
  INV_X1 U7041 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9943) );
  NAND2_X1 U7042 ( .A1(n6044), .A2(n9943), .ZN(n6045) );
  NAND2_X1 U7043 ( .A1(n6065), .A2(n6045), .ZN(n9003) );
  OR2_X1 U7044 ( .A1(n9003), .A2(n6089), .ZN(n6051) );
  INV_X1 U7045 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7046 ( .A1(n6536), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7047 ( .A1(n6535), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6046) );
  OAI211_X1 U7048 ( .C1(n6190), .C2(n6048), .A(n6047), .B(n6046), .ZN(n6049)
         );
  INV_X1 U7049 ( .A(n6049), .ZN(n6050) );
  NOR2_X1 U7050 ( .A1(n8813), .A2(n6911), .ZN(n8824) );
  NAND2_X1 U7051 ( .A1(n8825), .A2(n8824), .ZN(n8823) );
  INV_X1 U7052 ( .A(n6052), .ZN(n6054) );
  INV_X1 U7053 ( .A(n6057), .ZN(n6058) );
  NAND2_X1 U7054 ( .A1(n6058), .A2(SI_24_), .ZN(n6059) );
  INV_X1 U7055 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7828) );
  INV_X1 U7056 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8350) );
  MUX2_X1 U7057 ( .A(n7828), .B(n8350), .S(n8257), .Z(n6060) );
  INV_X1 U7058 ( .A(SI_25_), .ZN(n10064) );
  NAND2_X1 U7059 ( .A1(n6060), .A2(n10064), .ZN(n6078) );
  INV_X1 U7060 ( .A(n6060), .ZN(n6061) );
  NAND2_X1 U7061 ( .A1(n6061), .A2(SI_25_), .ZN(n6062) );
  NAND2_X1 U7062 ( .A1(n6078), .A2(n6062), .ZN(n6079) );
  XNOR2_X1 U7063 ( .A(n6080), .B(n6079), .ZN(n8349) );
  NAND2_X1 U7064 ( .A1(n8349), .A2(n5657), .ZN(n6064) );
  NAND2_X1 U7065 ( .A1(n4859), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6063) );
  XNOR2_X1 U7066 ( .A(n8989), .B(n6127), .ZN(n6073) );
  INV_X1 U7067 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U7068 ( .A1(n6065), .A2(n8816), .ZN(n6066) );
  NAND2_X1 U7069 ( .A1(n8986), .A2(n6192), .ZN(n6072) );
  INV_X1 U7070 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7071 ( .A1(n6535), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7072 ( .A1(n6536), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6067) );
  OAI211_X1 U7073 ( .C1(n6069), .C2(n6190), .A(n6068), .B(n6067), .ZN(n6070)
         );
  INV_X1 U7074 ( .A(n6070), .ZN(n6071) );
  NOR2_X1 U7075 ( .A1(n8997), .A2(n6911), .ZN(n6074) );
  XNOR2_X1 U7076 ( .A(n6073), .B(n6074), .ZN(n8812) );
  INV_X1 U7077 ( .A(n6074), .ZN(n6075) );
  INV_X1 U7078 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8002) );
  INV_X1 U7079 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8368) );
  MUX2_X1 U7080 ( .A(n8002), .B(n8368), .S(n8257), .Z(n6081) );
  INV_X1 U7081 ( .A(SI_26_), .ZN(n10063) );
  NAND2_X1 U7082 ( .A1(n6081), .A2(n10063), .ZN(n6101) );
  INV_X1 U7083 ( .A(n6081), .ZN(n6082) );
  NAND2_X1 U7084 ( .A1(n6082), .A2(SI_26_), .ZN(n6083) );
  AND2_X1 U7085 ( .A1(n6101), .A2(n6083), .ZN(n6099) );
  NAND2_X1 U7086 ( .A1(n8367), .A2(n5657), .ZN(n6085) );
  NAND2_X1 U7087 ( .A1(n5918), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7088 ( .A(n9117), .B(n6127), .ZN(n6097) );
  INV_X1 U7089 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10140) );
  NAND2_X1 U7090 ( .A1(n6087), .A2(n10140), .ZN(n6088) );
  NAND2_X1 U7091 ( .A1(n6121), .A2(n6088), .ZN(n8972) );
  INV_X1 U7092 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7093 ( .A1(n6536), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7094 ( .A1(n6535), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6090) );
  OAI211_X1 U7095 ( .C1(n6190), .C2(n6092), .A(n6091), .B(n6090), .ZN(n6093)
         );
  INV_X1 U7096 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U7097 ( .A1(n8920), .A2(n8434), .ZN(n6096) );
  NOR2_X1 U7098 ( .A1(n6097), .A2(n6096), .ZN(n6098) );
  AOI21_X1 U7099 ( .B1(n6097), .B2(n6096), .A(n6098), .ZN(n8846) );
  NAND2_X1 U7100 ( .A1(n6100), .A2(n6099), .ZN(n6102) );
  INV_X1 U7101 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8054) );
  INV_X1 U7102 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8665) );
  MUX2_X1 U7103 ( .A(n8054), .B(n8665), .S(n8257), .Z(n6103) );
  INV_X1 U7104 ( .A(SI_27_), .ZN(n9955) );
  NAND2_X1 U7105 ( .A1(n6103), .A2(n9955), .ZN(n6117) );
  INV_X1 U7106 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7107 ( .A1(n6104), .A2(SI_27_), .ZN(n6105) );
  AND2_X1 U7108 ( .A1(n6117), .A2(n6105), .ZN(n6115) );
  NAND2_X1 U7109 ( .A1(n8664), .A2(n5657), .ZN(n6107) );
  NAND2_X1 U7110 ( .A1(n5918), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6106) );
  XNOR2_X1 U7111 ( .A(n9110), .B(n6127), .ZN(n6113) );
  XNOR2_X1 U7112 ( .A(n6121), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8953) );
  INV_X1 U7113 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7114 ( .A1(n6535), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7115 ( .A1(n6536), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6108) );
  OAI211_X1 U7116 ( .C1(n6110), .C2(n6190), .A(n6109), .B(n6108), .ZN(n6111)
         );
  OR2_X1 U7117 ( .A1(n8970), .A2(n6911), .ZN(n6112) );
  NOR2_X1 U7118 ( .A1(n6113), .A2(n6112), .ZN(n6114) );
  AOI21_X1 U7119 ( .B1(n6113), .B2(n6112), .A(n6114), .ZN(n8783) );
  NAND2_X1 U7120 ( .A1(n8784), .A2(n8783), .ZN(n8782) );
  MUX2_X1 U7121 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n8257), .Z(n8225) );
  INV_X1 U7122 ( .A(SI_28_), .ZN(n10058) );
  XNOR2_X1 U7123 ( .A(n8225), .B(n10058), .ZN(n8223) );
  NAND2_X1 U7124 ( .A1(n8778), .A2(n5657), .ZN(n6119) );
  NAND2_X1 U7125 ( .A1(n5918), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6118) );
  INV_X1 U7126 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8785) );
  INV_X1 U7127 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10002) );
  OAI21_X1 U7128 ( .B1(n6121), .B2(n8785), .A(n10002), .ZN(n6122) );
  NAND2_X1 U7129 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6120) );
  INV_X1 U7130 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7131 ( .A1(n6536), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7132 ( .A1(n6535), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6123) );
  OAI211_X1 U7133 ( .C1(n6190), .C2(n6125), .A(n6124), .B(n6123), .ZN(n6126)
         );
  NAND2_X1 U7134 ( .A1(n6127), .A2(n8434), .ZN(n6128) );
  OR2_X1 U7135 ( .A1(n8958), .A2(n6128), .ZN(n6131) );
  NAND2_X1 U7136 ( .A1(n8958), .A2(n6129), .ZN(n6130) );
  NAND2_X1 U7137 ( .A1(n6131), .A2(n6130), .ZN(n6177) );
  AND3_X1 U7138 ( .A1(n6143), .A2(n6169), .A3(n6147), .ZN(n6132) );
  AND2_X1 U7139 ( .A1(n6133), .A2(n6132), .ZN(n6138) );
  INV_X1 U7140 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7141 ( .A1(n6138), .A2(n6134), .ZN(n6141) );
  NAND2_X1 U7142 ( .A1(n6141), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6135) );
  MUX2_X1 U7143 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6135), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6137) );
  NAND2_X1 U7144 ( .A1(n6137), .A2(n6136), .ZN(n8004) );
  NOR2_X1 U7145 ( .A1(n6138), .A2(n8262), .ZN(n6139) );
  MUX2_X1 U7146 ( .A(n8262), .B(n6139), .S(P2_IR_REG_25__SCAN_IN), .Z(n6140)
         );
  INV_X1 U7147 ( .A(n6140), .ZN(n6142) );
  NAND2_X1 U7148 ( .A1(n6142), .A2(n6141), .ZN(n7827) );
  NAND2_X1 U7149 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  NAND2_X1 U7150 ( .A1(n6145), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7151 ( .A1(n6170), .A2(n6169), .ZN(n6146) );
  NAND2_X1 U7152 ( .A1(n6146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6148) );
  XNOR2_X1 U7153 ( .A(n6148), .B(n6147), .ZN(n7752) );
  INV_X1 U7154 ( .A(P2_B_REG_SCAN_IN), .ZN(n8901) );
  INV_X1 U7155 ( .A(n7752), .ZN(n6149) );
  AOI221_X1 U7156 ( .B1(P2_B_REG_SCAN_IN), .B2(n7752), .C1(n8901), .C2(n6149), 
        .A(n8004), .ZN(n6150) );
  OR2_X1 U7157 ( .A1(n9937), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7158 ( .A1(n7752), .A2(n8004), .ZN(n10270) );
  NAND2_X1 U7159 ( .A1(n6151), .A2(n10270), .ZN(n6774) );
  NOR4_X1 U7160 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6155) );
  NOR4_X1 U7161 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6154) );
  NOR4_X1 U7162 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6153) );
  NOR4_X1 U7163 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6152) );
  NAND4_X1 U7164 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n6162)
         );
  NOR2_X1 U7165 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6159) );
  NOR4_X1 U7166 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6158) );
  NOR4_X1 U7167 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6157) );
  NOR4_X1 U7168 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6156) );
  NAND4_X1 U7169 ( .A1(n6159), .A2(n6158), .A3(n6157), .A4(n6156), .ZN(n6161)
         );
  INV_X1 U7170 ( .A(n9937), .ZN(n6160) );
  OAI21_X1 U7171 ( .B1(n6162), .B2(n6161), .A(n6160), .ZN(n6758) );
  INV_X1 U7172 ( .A(n6758), .ZN(n6163) );
  NOR2_X1 U7173 ( .A1(n6774), .A2(n6163), .ZN(n6166) );
  OR2_X1 U7174 ( .A1(n9937), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6165) );
  AND2_X1 U7175 ( .A1(n7827), .A2(n8004), .ZN(n9938) );
  INV_X1 U7176 ( .A(n9938), .ZN(n6164) );
  NAND2_X1 U7177 ( .A1(n6165), .A2(n6164), .ZN(n7152) );
  INV_X1 U7178 ( .A(n7152), .ZN(n7145) );
  INV_X1 U7179 ( .A(n6167), .ZN(n6168) );
  XNOR2_X1 U7180 ( .A(n6170), .B(n6169), .ZN(n6366) );
  NAND2_X1 U7181 ( .A1(n6367), .A2(n10274), .ZN(n6383) );
  OR2_X1 U7182 ( .A1(n6171), .A2(n5610), .ZN(n10377) );
  NOR2_X1 U7183 ( .A1(n6383), .A2(n10377), .ZN(n6172) );
  NAND2_X1 U7184 ( .A1(n6193), .A2(n6172), .ZN(n6174) );
  AND2_X1 U7185 ( .A1(n5610), .A2(n8973), .ZN(n7147) );
  NAND2_X1 U7186 ( .A1(n10609), .A2(n8423), .ZN(n6755) );
  NOR3_X1 U7187 ( .A1(n5148), .A2(n6177), .A3(n8851), .ZN(n6175) );
  AOI21_X1 U7188 ( .B1(n5148), .B2(n6177), .A(n6175), .ZN(n6181) );
  NAND3_X1 U7189 ( .A1(n9105), .A2(n10399), .A3(n6177), .ZN(n6176) );
  OAI21_X1 U7190 ( .B1(n9105), .B2(n6177), .A(n6176), .ZN(n6178) );
  INV_X1 U7191 ( .A(n6173), .ZN(n8641) );
  OR2_X1 U7192 ( .A1(n6383), .A2(n6183), .ZN(n6756) );
  NAND2_X1 U7193 ( .A1(n5610), .A2(n8890), .ZN(n6195) );
  NAND2_X1 U7194 ( .A1(n10340), .A2(n6195), .ZN(n10638) );
  NOR2_X1 U7195 ( .A1(n6756), .A2(n10150), .ZN(n6179) );
  NAND2_X1 U7196 ( .A1(n6193), .A2(n6179), .ZN(n10397) );
  OAI21_X1 U7197 ( .B1(n5148), .B2(n10399), .A(n10397), .ZN(n6180) );
  OR2_X1 U7198 ( .A1(n6383), .A2(n6195), .ZN(n8640) );
  INV_X1 U7199 ( .A(n8640), .ZN(n6182) );
  INV_X1 U7200 ( .A(n8970), .ZN(n8944) );
  AOI22_X1 U7201 ( .A1(n8804), .A2(n8944), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6201) );
  INV_X1 U7202 ( .A(n6184), .ZN(n6185) );
  INV_X1 U7203 ( .A(n6186), .ZN(n8930) );
  INV_X1 U7204 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7205 ( .A1(n6536), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7206 ( .A1(n6535), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6187) );
  OAI211_X1 U7207 ( .C1(n6190), .C2(n6189), .A(n6188), .B(n6187), .ZN(n6191)
         );
  AOI21_X1 U7208 ( .B1(n8930), .B2(n6192), .A(n6191), .ZN(n8419) );
  INV_X1 U7209 ( .A(n8419), .ZN(n8943) );
  INV_X1 U7210 ( .A(n6193), .ZN(n6194) );
  NAND2_X1 U7211 ( .A1(n6194), .A2(n6755), .ZN(n6199) );
  INV_X1 U7212 ( .A(n6195), .ZN(n6196) );
  OAI211_X1 U7213 ( .C1(n6196), .C2(n6761), .A(n6367), .B(n6366), .ZN(n6197)
         );
  INV_X1 U7214 ( .A(n6197), .ZN(n6198) );
  NAND2_X1 U7215 ( .A1(n6199), .A2(n6198), .ZN(n6748) );
  AOI22_X1 U7216 ( .A1(n8802), .A2(n8943), .B1(n8820), .B2(n8940), .ZN(n6200)
         );
  AND2_X1 U7217 ( .A1(n6201), .A2(n6200), .ZN(n6202) );
  INV_X1 U7218 ( .A(n6367), .ZN(n6203) );
  NOR2_X1 U7219 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6206) );
  INV_X1 U7220 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7221 ( .A1(n6236), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7222 ( .A1(n6214), .A2(n6238), .ZN(n6216) );
  NAND2_X1 U7223 ( .A1(n6216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6213) );
  OR2_X1 U7224 ( .A1(n6214), .A2(n6238), .ZN(n6215) );
  NAND2_X1 U7225 ( .A1(n6216), .A2(n6215), .ZN(n6490) );
  NAND2_X1 U7226 ( .A1(n6217), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7227 ( .A1(n5266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6222) );
  XNOR2_X1 U7228 ( .A(n6222), .B(n6221), .ZN(n7702) );
  AND2_X1 U7229 ( .A1(n7702), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6489) );
  INV_X1 U7230 ( .A(n6489), .ZN(n6223) );
  OR2_X2 U7231 ( .A1(n6815), .A2(n6223), .ZN(n9557) );
  INV_X1 U7232 ( .A(n9557), .ZN(P1_U4006) );
  NOR2_X1 U7233 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6224) );
  INV_X1 U7234 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6251) );
  AND2_X1 U7235 ( .A1(n6252), .A2(n6251), .ZN(n6245) );
  INV_X1 U7236 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6225) );
  AND3_X1 U7237 ( .A1(n6249), .A2(n6226), .A3(n6225), .ZN(n6227) );
  NAND2_X1 U7238 ( .A1(n6617), .A2(n6616), .ZN(n6229) );
  NAND2_X1 U7239 ( .A1(n6233), .A2(n6230), .ZN(n6231) );
  NAND2_X1 U7240 ( .A1(n6698), .A2(n6234), .ZN(n6715) );
  NAND2_X1 U7241 ( .A1(n6715), .A2(n6815), .ZN(n6235) );
  NAND2_X1 U7242 ( .A1(n6235), .A2(n7702), .ZN(n10221) );
  INV_X1 U7243 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7244 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n6240) );
  XNOR2_X2 U7245 ( .A(n6242), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6311) );
  NAND2_X2 U7246 ( .A1(n6313), .A2(n6311), .ZN(n6694) );
  NAND2_X1 U7247 ( .A1(n10221), .A2(n6694), .ZN(n6243) );
  NAND2_X1 U7248 ( .A1(n6243), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U7249 ( .A1(n6244), .A2(n6245), .ZN(n6246) );
  NAND2_X1 U7250 ( .A1(n6246), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7251 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n6247) );
  NAND2_X1 U7252 ( .A1(n6253), .A2(n6247), .ZN(n6250) );
  OAI21_X1 U7253 ( .B1(n6250), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6248) );
  XNOR2_X1 U7254 ( .A(n6248), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10250) );
  XNOR2_X1 U7255 ( .A(n6249), .B(n6250), .ZN(n8162) );
  XNOR2_X1 U7256 ( .A(n6253), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8063) );
  AND2_X1 U7257 ( .A1(n6244), .A2(n6251), .ZN(n6257) );
  NOR2_X1 U7258 ( .A1(n6257), .A2(n6277), .ZN(n6254) );
  MUX2_X1 U7259 ( .A(n6254), .B(n6253), .S(n6252), .Z(n7790) );
  NOR2_X1 U7260 ( .A1(n6244), .A2(n6277), .ZN(n6255) );
  MUX2_X1 U7261 ( .A(n6277), .B(n6255), .S(P1_IR_REG_14__SCAN_IN), .Z(n6256)
         );
  INV_X1 U7262 ( .A(n6256), .ZN(n6259) );
  INV_X1 U7263 ( .A(n6257), .ZN(n6258) );
  AND2_X1 U7264 ( .A1(n6259), .A2(n6258), .ZN(n7807) );
  INV_X1 U7265 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6260) );
  XNOR2_X1 U7266 ( .A(n7807), .B(n6260), .ZN(n7614) );
  OR2_X1 U7267 ( .A1(n6261), .A2(n6277), .ZN(n6266) );
  NAND2_X1 U7268 ( .A1(n6266), .A2(n6262), .ZN(n6263) );
  NAND2_X1 U7269 ( .A1(n6263), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6264) );
  XNOR2_X1 U7270 ( .A(n6264), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7708) );
  INV_X1 U7271 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6265) );
  XNOR2_X1 U7272 ( .A(n7708), .B(n6265), .ZN(n7384) );
  XNOR2_X1 U7273 ( .A(n6266), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7676) );
  XOR2_X1 U7274 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7676), .Z(n7055) );
  NOR2_X1 U7275 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6278) );
  NOR2_X1 U7276 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n6267) );
  NAND3_X1 U7277 ( .A1(n6268), .A2(n6278), .A3(n6267), .ZN(n6273) );
  NOR2_X1 U7278 ( .A1(n6275), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6297) );
  OR2_X1 U7279 ( .A1(n6297), .A2(n6277), .ZN(n6271) );
  INV_X1 U7280 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7281 ( .A1(n6271), .A2(n6296), .ZN(n6269) );
  NAND2_X1 U7282 ( .A1(n6269), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6270) );
  XNOR2_X1 U7283 ( .A(n6270), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7271) );
  INV_X1 U7284 ( .A(n7271), .ZN(n6610) );
  INV_X1 U7285 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10590) );
  INV_X1 U7286 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10570) );
  XNOR2_X1 U7287 ( .A(n6271), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7278) );
  INV_X1 U7288 ( .A(n7278), .ZN(n6594) );
  NAND2_X1 U7289 ( .A1(n6275), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6272) );
  XNOR2_X1 U7290 ( .A(n6272), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7023) );
  NOR2_X1 U7291 ( .A1(n7023), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7292 ( .A1(n6273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6274) );
  MUX2_X1 U7293 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6274), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6276) );
  AND2_X1 U7294 ( .A1(n6276), .A2(n6275), .ZN(n10207) );
  NAND2_X1 U7295 ( .A1(n10207), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6293) );
  OAI21_X1 U7296 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(P1_IR_REG_2__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6279) );
  OAI21_X1 U7297 ( .B1(n6282), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6280) );
  XNOR2_X1 U7298 ( .A(n6280), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U7299 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n10258), .ZN(n6291) );
  MUX2_X1 U7300 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10481), .S(n10258), .Z(
        n10264) );
  INV_X1 U7301 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6281) );
  XNOR2_X1 U7302 ( .A(n6282), .B(n6281), .ZN(n6670) );
  NOR2_X1 U7303 ( .A1(n6670), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6290) );
  INV_X1 U7304 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7305 ( .A1(n6287), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6284) );
  INV_X1 U7306 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6283) );
  XNOR2_X1 U7307 ( .A(n6284), .B(n6283), .ZN(n6780) );
  INV_X1 U7308 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6576) );
  INV_X1 U7309 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10361) );
  NAND2_X1 U7310 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6285) );
  XNOR2_X1 U7311 ( .A(n6286), .B(n6285), .ZN(n6702) );
  XNOR2_X1 U7312 ( .A(n6702), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n6557) );
  NAND3_X1 U7313 ( .A1(n6557), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6555) );
  OAI21_X1 U7314 ( .B1(n10361), .B2(n6702), .A(n6555), .ZN(n10326) );
  XNOR2_X1 U7315 ( .A(n10319), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10327) );
  INV_X1 U7316 ( .A(n10319), .ZN(n6328) );
  AOI22_X1 U7317 ( .A1(n10326), .A2(n10327), .B1(P1_REG1_REG_2__SCAN_IN), .B2(
        n6328), .ZN(n6577) );
  MUX2_X1 U7318 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6576), .S(n6780), .Z(n6289)
         );
  OR2_X1 U7319 ( .A1(n6577), .A2(n6289), .ZN(n6578) );
  OAI21_X1 U7320 ( .B1(n6780), .B2(n6576), .A(n6578), .ZN(n6665) );
  INV_X1 U7321 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10432) );
  INV_X1 U7322 ( .A(n6670), .ZN(n6811) );
  AOI22_X1 U7323 ( .A1(n6670), .A2(n10432), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n6811), .ZN(n6664) );
  NOR2_X1 U7324 ( .A1(n6665), .A2(n6664), .ZN(n6663) );
  NOR2_X1 U7325 ( .A1(n6290), .A2(n6663), .ZN(n10265) );
  NAND2_X1 U7326 ( .A1(n10264), .A2(n10265), .ZN(n10263) );
  NAND2_X1 U7327 ( .A1(n6291), .A2(n10263), .ZN(n10213) );
  INV_X1 U7328 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10529) );
  INV_X1 U7329 ( .A(n10207), .ZN(n6505) );
  INV_X1 U7330 ( .A(n6293), .ZN(n6292) );
  AOI21_X1 U7331 ( .B1(n10529), .B2(n6505), .A(n6292), .ZN(n10214) );
  NAND2_X1 U7332 ( .A1(n10213), .A2(n10214), .ZN(n10212) );
  NAND2_X1 U7333 ( .A1(n6293), .A2(n10212), .ZN(n6549) );
  INV_X1 U7334 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10555) );
  INV_X1 U7335 ( .A(n7023), .ZN(n6506) );
  AOI22_X1 U7336 ( .A1(n7023), .A2(n10555), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n6506), .ZN(n6548) );
  NOR2_X1 U7337 ( .A1(n6549), .A2(n6548), .ZN(n6547) );
  NOR2_X1 U7338 ( .A1(n6294), .A2(n6547), .ZN(n6597) );
  AOI22_X1 U7339 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6594), .B1(n7278), .B2(
        n10570), .ZN(n6596) );
  NOR2_X1 U7340 ( .A1(n6597), .A2(n6596), .ZN(n6595) );
  AOI21_X1 U7341 ( .B1(n10570), .B2(n6594), .A(n6595), .ZN(n6605) );
  AOI22_X1 U7342 ( .A1(n7271), .A2(n10590), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6610), .ZN(n6604) );
  NOR2_X1 U7343 ( .A1(n6605), .A2(n6604), .ZN(n6603) );
  AOI21_X1 U7344 ( .B1(n6610), .B2(n10590), .A(n6603), .ZN(n6679) );
  INV_X1 U7345 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6295) );
  NAND3_X1 U7346 ( .A1(n6297), .A2(n6296), .A3(n6295), .ZN(n6298) );
  NAND2_X1 U7347 ( .A1(n6298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6299) );
  XNOR2_X1 U7348 ( .A(n6299), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7483) );
  INV_X1 U7349 ( .A(n7483), .ZN(n6681) );
  INV_X1 U7350 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7643) );
  AOI22_X1 U7351 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6681), .B1(n7483), .B2(
        n7643), .ZN(n6678) );
  NOR2_X1 U7352 ( .A1(n6679), .A2(n6678), .ZN(n6677) );
  NOR2_X1 U7353 ( .A1(n7483), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6300) );
  INV_X1 U7354 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U7355 ( .A1(n10232), .A2(n10231), .ZN(n10235) );
  NAND2_X1 U7356 ( .A1(n6301), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6302) );
  XNOR2_X1 U7357 ( .A(n6302), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10238) );
  INV_X1 U7358 ( .A(n10232), .ZN(n6303) );
  OAI22_X1 U7359 ( .A1(n10235), .A2(n10238), .B1(P1_REG1_REG_11__SCAN_IN), 
        .B2(n6303), .ZN(n10234) );
  NAND2_X1 U7360 ( .A1(n7055), .A2(n10234), .ZN(n7054) );
  OAI21_X1 U7361 ( .B1(n7676), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7054), .ZN(
        n7383) );
  NAND2_X1 U7362 ( .A1(n7384), .A2(n7383), .ZN(n7382) );
  OAI21_X1 U7363 ( .B1(n7708), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7382), .ZN(
        n7613) );
  NAND2_X1 U7364 ( .A1(n7614), .A2(n7613), .ZN(n7612) );
  OAI21_X1 U7365 ( .B1(n7807), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7612), .ZN(
        n6304) );
  NOR2_X1 U7366 ( .A1(n7790), .A2(n6304), .ZN(n6305) );
  INV_X1 U7367 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7793) );
  XNOR2_X1 U7368 ( .A(n7790), .B(n6304), .ZN(n7792) );
  NOR2_X1 U7369 ( .A1(n7793), .A2(n7792), .ZN(n7791) );
  NOR2_X1 U7370 ( .A1(n6305), .A2(n7791), .ZN(n7946) );
  XNOR2_X1 U7371 ( .A(n8063), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7945) );
  NOR2_X1 U7372 ( .A1(n7946), .A2(n7945), .ZN(n7944) );
  AOI21_X1 U7373 ( .B1(n8063), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7944), .ZN(
        n8151) );
  XNOR2_X1 U7374 ( .A(n8162), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8152) );
  NOR2_X1 U7375 ( .A1(n8151), .A2(n8152), .ZN(n8150) );
  AOI21_X1 U7376 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n8162), .A(n8150), .ZN(
        n10253) );
  INV_X1 U7377 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8181) );
  INV_X1 U7378 ( .A(n10250), .ZN(n7093) );
  AOI22_X1 U7379 ( .A1(n10250), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8181), .B2(
        n7093), .ZN(n10252) );
  NAND2_X1 U7380 ( .A1(n10253), .A2(n10252), .ZN(n10251) );
  OAI21_X1 U7381 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n10250), .A(n10251), .ZN(
        n6310) );
  NAND2_X1 U7382 ( .A1(n6307), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6308) );
  XNOR2_X2 U7383 ( .A(n6306), .B(n6308), .ZN(n9697) );
  XNOR2_X1 U7384 ( .A(n10493), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n6309) );
  XNOR2_X1 U7385 ( .A(n6310), .B(n6309), .ZN(n6314) );
  OR2_X1 U7386 ( .A1(n6311), .A2(P1_U3084), .ZN(n8148) );
  INV_X1 U7387 ( .A(n8148), .ZN(n6312) );
  NAND2_X1 U7388 ( .A1(n10221), .A2(n6312), .ZN(n6318) );
  INV_X1 U7389 ( .A(n10220), .ZN(n10198) );
  OR2_X1 U7390 ( .A1(n6318), .A2(n10198), .ZN(n10236) );
  NOR2_X1 U7391 ( .A1(n6314), .A2(n10236), .ZN(n6359) );
  INV_X1 U7392 ( .A(n7702), .ZN(n6315) );
  NOR2_X1 U7393 ( .A1(n6815), .A2(n6315), .ZN(n6316) );
  OR2_X1 U7394 ( .A1(P1_U3083), .A2(n6316), .ZN(n10312) );
  NOR2_X1 U7395 ( .A1(n10312), .A2(n6317), .ZN(n6358) );
  OR2_X1 U7396 ( .A1(n6318), .A2(n10220), .ZN(n10321) );
  NAND2_X1 U7397 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7483), .ZN(n6342) );
  INV_X1 U7398 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6319) );
  MUX2_X1 U7399 ( .A(n6319), .B(P1_REG2_REG_10__SCAN_IN), .S(n7483), .Z(n6320)
         );
  INV_X1 U7400 ( .A(n6320), .ZN(n6684) );
  NAND2_X1 U7401 ( .A1(n7271), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6341) );
  INV_X1 U7402 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6321) );
  MUX2_X1 U7403 ( .A(n6321), .B(P1_REG2_REG_9__SCAN_IN), .S(n7271), .Z(n6322)
         );
  INV_X1 U7404 ( .A(n6322), .ZN(n6607) );
  NOR2_X1 U7405 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7278), .ZN(n6340) );
  NOR2_X1 U7406 ( .A1(n7023), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6337) );
  INV_X1 U7407 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6334) );
  NOR2_X1 U7408 ( .A1(n6670), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6331) );
  INV_X1 U7409 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6329) );
  INV_X1 U7410 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6323) );
  MUX2_X1 U7411 ( .A(n6323), .B(P1_REG2_REG_2__SCAN_IN), .S(n10319), .Z(n6327)
         );
  INV_X1 U7412 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6325) );
  MUX2_X1 U7413 ( .A(n6325), .B(P1_REG2_REG_1__SCAN_IN), .S(n6702), .Z(n6561)
         );
  AND2_X1 U7414 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6324) );
  NAND2_X1 U7415 ( .A1(n6561), .A2(n6324), .ZN(n10314) );
  OR2_X1 U7416 ( .A1(n6702), .A2(n6325), .ZN(n10313) );
  NAND2_X1 U7417 ( .A1(n10314), .A2(n10313), .ZN(n6326) );
  MUX2_X1 U7418 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6329), .S(n6780), .Z(n6572)
         );
  OAI21_X1 U7419 ( .B1(n6780), .B2(n6329), .A(n6570), .ZN(n6669) );
  INV_X1 U7420 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6330) );
  AOI22_X1 U7421 ( .A1(n6670), .A2(n6330), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n6811), .ZN(n6668) );
  INV_X1 U7422 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6332) );
  MUX2_X1 U7423 ( .A(n6332), .B(P1_REG2_REG_5__SCAN_IN), .S(n10258), .Z(n10260) );
  MUX2_X1 U7424 ( .A(n6334), .B(P1_REG2_REG_6__SCAN_IN), .S(n10207), .Z(n6333)
         );
  INV_X1 U7425 ( .A(n6333), .ZN(n10210) );
  NAND2_X1 U7426 ( .A1(n10211), .A2(n10210), .ZN(n10209) );
  OAI21_X1 U7427 ( .B1(n6334), .B2(n6505), .A(n10209), .ZN(n6546) );
  INV_X1 U7428 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6335) );
  MUX2_X1 U7429 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6335), .S(n7023), .Z(n6336)
         );
  INV_X1 U7430 ( .A(n6336), .ZN(n6545) );
  NOR2_X1 U7431 ( .A1(n6546), .A2(n6545), .ZN(n6544) );
  NOR2_X1 U7432 ( .A1(n6337), .A2(n6544), .ZN(n6592) );
  INV_X1 U7433 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6338) );
  MUX2_X1 U7434 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6338), .S(n7278), .Z(n6339)
         );
  INV_X1 U7435 ( .A(n6339), .ZN(n6591) );
  NAND2_X1 U7436 ( .A1(n6684), .A2(n6685), .ZN(n6683) );
  NAND2_X1 U7437 ( .A1(n6342), .A2(n6683), .ZN(n10229) );
  AND2_X1 U7438 ( .A1(n10229), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6343) );
  OAI22_X1 U7439 ( .A1(n6343), .A2(n10238), .B1(n10229), .B2(
        P1_REG2_REG_11__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U7440 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7676), .ZN(n6344) );
  OAI21_X1 U7441 ( .B1(n7676), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6344), .ZN(
        n7060) );
  NOR2_X1 U7442 ( .A1(n10227), .A2(n7060), .ZN(n7059) );
  AOI21_X1 U7443 ( .B1(n7676), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7059), .ZN(
        n7379) );
  NAND2_X1 U7444 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7708), .ZN(n6345) );
  OAI21_X1 U7445 ( .B1(n7708), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6345), .ZN(
        n7378) );
  INV_X1 U7446 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6347) );
  NOR2_X1 U7447 ( .A1(n7807), .A2(n6347), .ZN(n6346) );
  AOI21_X1 U7448 ( .B1(n7807), .B2(n6347), .A(n6346), .ZN(n7608) );
  NOR2_X1 U7449 ( .A1(n7790), .A2(n6348), .ZN(n6349) );
  INV_X1 U7450 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7798) );
  XNOR2_X1 U7451 ( .A(n7790), .B(n6348), .ZN(n7797) );
  NOR2_X1 U7452 ( .A1(n7798), .A2(n7797), .ZN(n7796) );
  NAND2_X1 U7453 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8063), .ZN(n6350) );
  OAI21_X1 U7454 ( .B1(n8063), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6350), .ZN(
        n7942) );
  NAND2_X1 U7455 ( .A1(n8162), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6351) );
  OAI21_X1 U7456 ( .B1(n8162), .B2(P1_REG2_REG_17__SCAN_IN), .A(n6351), .ZN(
        n8156) );
  AOI21_X1 U7457 ( .B1(n8162), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8155), .ZN(
        n10247) );
  INV_X1 U7458 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n6353) );
  NOR2_X1 U7459 ( .A1(n10250), .A2(n6353), .ZN(n6352) );
  AOI21_X1 U7460 ( .B1(n10250), .B2(n6353), .A(n6352), .ZN(n10246) );
  NOR2_X1 U7461 ( .A1(n10247), .A2(n10246), .ZN(n10245) );
  INV_X1 U7462 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6354) );
  MUX2_X1 U7463 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n6354), .S(n9697), .Z(n6355)
         );
  INV_X1 U7464 ( .A(n6311), .ZN(n6727) );
  OR2_X1 U7465 ( .A1(n10220), .A2(P1_U3084), .ZN(n8005) );
  NOR2_X1 U7466 ( .A1(n6727), .A2(n8005), .ZN(n6356) );
  NAND2_X1 U7467 ( .A1(n10221), .A2(n6356), .ZN(n10318) );
  NAND2_X1 U7468 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9209) );
  OAI21_X1 U7469 ( .B1(n10318), .B2(n9697), .A(n9209), .ZN(n6357) );
  INV_X1 U7470 ( .A(n6485), .ZN(n6376) );
  INV_X1 U7471 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10275) );
  MUX2_X1 U7472 ( .A(n6360), .B(P2_REG2_REG_1__SCAN_IN), .S(n10292), .Z(n10288) );
  NOR3_X1 U7473 ( .A1(n10275), .A2(n5621), .A3(n10288), .ZN(n10287) );
  AOI21_X1 U7474 ( .B1(n10292), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10287), .ZN(
        n10304) );
  MUX2_X1 U7475 ( .A(n6361), .B(P2_REG2_REG_2__SCAN_IN), .S(n10307), .Z(n10303) );
  NOR2_X1 U7476 ( .A1(n10304), .A2(n10303), .ZN(n10302) );
  AOI21_X1 U7477 ( .B1(n10307), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10302), .ZN(
        n6402) );
  MUX2_X1 U7478 ( .A(n6362), .B(P2_REG2_REG_3__SCAN_IN), .S(n6403), .Z(n6401)
         );
  NOR2_X1 U7479 ( .A1(n6402), .A2(n6401), .ZN(n6400) );
  AOI21_X1 U7480 ( .B1(n6403), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6400), .ZN(
        n6429) );
  XNOR2_X1 U7481 ( .A(n6430), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6428) );
  INV_X1 U7482 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6363) );
  MUX2_X1 U7483 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6363), .S(n6485), .Z(n6391)
         );
  INV_X1 U7484 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6364) );
  MUX2_X1 U7485 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6364), .S(n6418), .Z(n6365)
         );
  INV_X1 U7486 ( .A(n6365), .ZN(n6370) );
  NOR2_X1 U7487 ( .A1(n4886), .A2(n6370), .ZN(n6413) );
  OR2_X1 U7488 ( .A1(n6366), .A2(P2_U3152), .ZN(n8644) );
  OAI211_X1 U7489 ( .C1(n6367), .C2(P2_U3152), .A(n6756), .B(n8644), .ZN(n6379) );
  NAND2_X1 U7490 ( .A1(n6379), .A2(n6382), .ZN(n6368) );
  NAND2_X1 U7491 ( .A1(n6368), .A2(n8861), .ZN(n6371) );
  NOR2_X1 U7492 ( .A1(n6184), .A2(n8902), .ZN(n6369) );
  AOI211_X1 U7493 ( .C1(n4886), .C2(n6370), .A(n6413), .B(n10301), .ZN(n6389)
         );
  NAND2_X1 U7494 ( .A1(n6371), .A2(n6184), .ZN(n8891) );
  INV_X1 U7495 ( .A(n6418), .ZN(n6502) );
  NOR2_X1 U7496 ( .A1(n8891), .A2(n6502), .ZN(n6388) );
  MUX2_X1 U7497 ( .A(n6372), .B(P2_REG1_REG_1__SCAN_IN), .S(n10292), .Z(n10285) );
  NOR3_X1 U7498 ( .A1(n10275), .A2(n10277), .A3(n10285), .ZN(n10284) );
  AOI21_X1 U7499 ( .B1(n10292), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10284), .ZN(
        n10300) );
  INV_X1 U7500 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6373) );
  MUX2_X1 U7501 ( .A(n6373), .B(P2_REG1_REG_2__SCAN_IN), .S(n10307), .Z(n10299) );
  NOR2_X1 U7502 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  AOI21_X1 U7503 ( .B1(n10307), .B2(P2_REG1_REG_2__SCAN_IN), .A(n10298), .ZN(
        n6406) );
  MUX2_X1 U7504 ( .A(n6374), .B(P2_REG1_REG_3__SCAN_IN), .S(n6403), .Z(n6405)
         );
  NOR2_X1 U7505 ( .A1(n6406), .A2(n6405), .ZN(n6404) );
  AOI21_X1 U7506 ( .B1(n6403), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6404), .ZN(
        n6433) );
  XNOR2_X1 U7507 ( .A(n6430), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6432) );
  NOR2_X1 U7508 ( .A1(n6433), .A2(n6432), .ZN(n6431) );
  AOI21_X1 U7509 ( .B1(n6430), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6431), .ZN(
        n6395) );
  INV_X1 U7510 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6375) );
  MUX2_X1 U7511 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6375), .S(n6485), .Z(n6394)
         );
  NOR2_X1 U7512 ( .A1(n6395), .A2(n6394), .ZN(n6393) );
  AOI21_X1 U7513 ( .B1(n6376), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6393), .ZN(
        n6381) );
  INV_X1 U7514 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6377) );
  MUX2_X1 U7515 ( .A(n6377), .B(P2_REG1_REG_6__SCAN_IN), .S(n6418), .Z(n6380)
         );
  NOR2_X1 U7516 ( .A1(n6381), .A2(n6380), .ZN(n6417) );
  AND2_X1 U7517 ( .A1(n6382), .A2(n8902), .ZN(n6378) );
  NAND2_X1 U7518 ( .A1(n6379), .A2(n6378), .ZN(n10297) );
  AOI211_X1 U7519 ( .C1(n6381), .C2(n6380), .A(n6417), .B(n10297), .ZN(n6387)
         );
  OAI21_X1 U7520 ( .B1(n6383), .B2(n6761), .A(n6382), .ZN(n6385) );
  NAND2_X1 U7521 ( .A1(n6383), .A2(n8644), .ZN(n6384) );
  NAND2_X1 U7522 ( .A1(n6385), .A2(n6384), .ZN(n8893) );
  INV_X1 U7523 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U7524 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6987) );
  OAI21_X1 U7525 ( .B1(n8893), .B2(n10171), .A(n6987), .ZN(n6386) );
  OR4_X1 U7526 ( .A1(n6389), .A2(n6388), .A3(n6387), .A4(n6386), .ZN(P2_U3251)
         );
  AOI211_X1 U7527 ( .C1(n6392), .C2(n6391), .A(n6390), .B(n10301), .ZN(n6399)
         );
  NOR2_X1 U7528 ( .A1(n8891), .A2(n6485), .ZN(n6398) );
  AOI211_X1 U7529 ( .C1(n6395), .C2(n6394), .A(n6393), .B(n10297), .ZN(n6397)
         );
  INV_X1 U7530 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U7531 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n6997) );
  OAI21_X1 U7532 ( .B1(n8893), .B2(n10169), .A(n6997), .ZN(n6396) );
  OR4_X1 U7533 ( .A1(n6399), .A2(n6398), .A3(n6397), .A4(n6396), .ZN(P2_U3250)
         );
  AOI211_X1 U7534 ( .C1(n6402), .C2(n6401), .A(n6400), .B(n10301), .ZN(n6412)
         );
  INV_X1 U7535 ( .A(n6403), .ZN(n6483) );
  NOR2_X1 U7536 ( .A1(n8891), .A2(n6483), .ZN(n6411) );
  AOI211_X1 U7537 ( .C1(n6406), .C2(n6405), .A(n6404), .B(n10297), .ZN(n6410)
         );
  INV_X1 U7538 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U7539 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n6407) );
  OAI21_X1 U7540 ( .B1(n8893), .B2(n6408), .A(n6407), .ZN(n6409) );
  OR4_X1 U7541 ( .A1(n6412), .A2(n6411), .A3(n6410), .A4(n6409), .ZN(P2_U3248)
         );
  INV_X1 U7542 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6414) );
  MUX2_X1 U7543 ( .A(n6414), .B(P2_REG2_REG_7__SCAN_IN), .S(n6444), .Z(n6415)
         );
  AOI211_X1 U7544 ( .C1(n6416), .C2(n6415), .A(n6439), .B(n10301), .ZN(n6426)
         );
  INV_X1 U7545 ( .A(n6444), .ZN(n6507) );
  NOR2_X1 U7546 ( .A1(n8891), .A2(n6507), .ZN(n6425) );
  AOI21_X1 U7547 ( .B1(n6418), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6417), .ZN(
        n6421) );
  MUX2_X1 U7548 ( .A(n6419), .B(P2_REG1_REG_7__SCAN_IN), .S(n6444), .Z(n6420)
         );
  NOR2_X1 U7549 ( .A1(n6421), .A2(n6420), .ZN(n6443) );
  AOI211_X1 U7550 ( .C1(n6421), .C2(n6420), .A(n10297), .B(n6443), .ZN(n6424)
         );
  INV_X1 U7551 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10173) );
  NAND2_X1 U7552 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n6422) );
  OAI21_X1 U7553 ( .B1(n8893), .B2(n10173), .A(n6422), .ZN(n6423) );
  OR4_X1 U7554 ( .A1(n6426), .A2(n6425), .A3(n6424), .A4(n6423), .ZN(P2_U3252)
         );
  AOI211_X1 U7555 ( .C1(n6429), .C2(n6428), .A(n6427), .B(n10301), .ZN(n6438)
         );
  NOR2_X1 U7556 ( .A1(n8891), .A2(n5004), .ZN(n6437) );
  AOI211_X1 U7557 ( .C1(n6433), .C2(n6432), .A(n6431), .B(n10297), .ZN(n6436)
         );
  INV_X1 U7558 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U7559 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7015) );
  OAI21_X1 U7560 ( .B1(n8893), .B2(n6434), .A(n7015), .ZN(n6435) );
  OR4_X1 U7561 ( .A1(n6438), .A2(n6437), .A3(n6436), .A4(n6435), .ZN(P2_U3249)
         );
  MUX2_X1 U7562 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7407), .S(n6459), .Z(n6440)
         );
  INV_X1 U7563 ( .A(n6440), .ZN(n6441) );
  AOI211_X1 U7564 ( .C1(n6442), .C2(n6441), .A(n10301), .B(n6453), .ZN(n6452)
         );
  AOI21_X1 U7565 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n6444), .A(n6443), .ZN(
        n6447) );
  MUX2_X1 U7566 ( .A(n6445), .B(P2_REG1_REG_8__SCAN_IN), .S(n6459), .Z(n6446)
         );
  NOR2_X1 U7567 ( .A1(n6447), .A2(n6446), .ZN(n6458) );
  AOI211_X1 U7568 ( .C1(n6447), .C2(n6446), .A(n10297), .B(n6458), .ZN(n6451)
         );
  INV_X1 U7569 ( .A(n6459), .ZN(n6510) );
  NOR2_X1 U7570 ( .A1(n8891), .A2(n6510), .ZN(n6450) );
  INV_X1 U7571 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U7572 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6448) );
  OAI21_X1 U7573 ( .B1(n8893), .B2(n10175), .A(n6448), .ZN(n6449) );
  OR4_X1 U7574 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(P2_U3253)
         );
  AOI21_X1 U7575 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6459), .A(n6453), .ZN(
        n6457) );
  INV_X1 U7576 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6454) );
  MUX2_X1 U7577 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6454), .S(n6472), .Z(n6455)
         );
  INV_X1 U7578 ( .A(n6455), .ZN(n6456) );
  NOR2_X1 U7579 ( .A1(n6457), .A2(n6456), .ZN(n6467) );
  AOI211_X1 U7580 ( .C1(n6457), .C2(n6456), .A(n10301), .B(n6467), .ZN(n6466)
         );
  AOI21_X1 U7581 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n6459), .A(n6458), .ZN(
        n6462) );
  MUX2_X1 U7582 ( .A(n6460), .B(P2_REG1_REG_9__SCAN_IN), .S(n6472), .Z(n6461)
         );
  NOR2_X1 U7583 ( .A1(n6462), .A2(n6461), .ZN(n6471) );
  AOI211_X1 U7584 ( .C1(n6462), .C2(n6461), .A(n10297), .B(n6471), .ZN(n6465)
         );
  INV_X1 U7585 ( .A(n6472), .ZN(n6515) );
  NOR2_X1 U7586 ( .A1(n8891), .A2(n6515), .ZN(n6464) );
  INV_X1 U7587 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10177) );
  NAND2_X1 U7588 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7169) );
  OAI21_X1 U7589 ( .B1(n8893), .B2(n10177), .A(n7169), .ZN(n6463) );
  OR4_X1 U7590 ( .A1(n6466), .A2(n6465), .A3(n6464), .A4(n6463), .ZN(P2_U3254)
         );
  NAND2_X1 U7591 ( .A1(n7195), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6468) );
  OAI21_X1 U7592 ( .B1(n7195), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6468), .ZN(
        n6469) );
  AOI211_X1 U7593 ( .C1(n6470), .C2(n6469), .A(n7189), .B(n10301), .ZN(n6481)
         );
  AOI21_X1 U7594 ( .B1(n6472), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6471), .ZN(
        n6475) );
  MUX2_X1 U7595 ( .A(n6473), .B(P2_REG1_REG_10__SCAN_IN), .S(n7195), .Z(n6474)
         );
  NOR2_X1 U7596 ( .A1(n6475), .A2(n6474), .ZN(n7194) );
  AOI211_X1 U7597 ( .C1(n6475), .C2(n6474), .A(n7194), .B(n10297), .ZN(n6480)
         );
  INV_X1 U7598 ( .A(n7195), .ZN(n6531) );
  NOR2_X1 U7599 ( .A1(n8891), .A2(n6531), .ZN(n6479) );
  INV_X1 U7600 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U7601 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n6476) );
  OAI21_X1 U7602 ( .B1(n8893), .B2(n6477), .A(n6476), .ZN(n6478) );
  OR4_X1 U7603 ( .A1(n6481), .A2(n6480), .A3(n6479), .A4(n6478), .ZN(P2_U3255)
         );
  AND2_X1 U7604 ( .A1(n8257), .A2(P2_U3152), .ZN(n8410) );
  AOI22_X1 U7605 ( .A1(n10307), .A2(P2_STATE_REG_SCAN_IN), .B1(n8410), .B2(
        P1_DATAO_REG_2__SCAN_IN), .ZN(n6482) );
  OAI21_X1 U7606 ( .B1(n6693), .B2(n7619), .A(n6482), .ZN(P2_U3356) );
  AND2_X1 U7607 ( .A1(n4832), .A2(P1_U3084), .ZN(n6980) );
  INV_X2 U7608 ( .A(n6980), .ZN(n8775) );
  INV_X1 U7609 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6701) );
  AND2_X1 U7610 ( .A1(n8257), .A2(P1_U3084), .ZN(n8147) );
  INV_X2 U7611 ( .A(n8147), .ZN(n8777) );
  OAI222_X1 U7612 ( .A1(n8775), .A2(n6701), .B1(n8777), .B2(n8412), .C1(
        P1_U3084), .C2(n6702), .ZN(P1_U3352) );
  INV_X1 U7613 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6808) );
  INV_X1 U7614 ( .A(n6807), .ZN(n6487) );
  OAI222_X1 U7615 ( .A1(n8775), .A2(n6808), .B1(n8777), .B2(n6487), .C1(
        P1_U3084), .C2(n6811), .ZN(P1_U3349) );
  INV_X1 U7616 ( .A(n8410), .ZN(n8781) );
  INV_X1 U7617 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6484) );
  OAI222_X1 U7618 ( .A1(n8781), .A2(n6484), .B1(n7619), .B2(n6781), .C1(
        P2_U3152), .C2(n6483), .ZN(P2_U3355) );
  INV_X1 U7619 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6486) );
  INV_X1 U7620 ( .A(n6850), .ZN(n6500) );
  OAI222_X1 U7621 ( .A1(n8781), .A2(n6486), .B1(n7619), .B2(n6500), .C1(
        P2_U3152), .C2(n6485), .ZN(P2_U3353) );
  INV_X1 U7622 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6488) );
  OAI222_X1 U7623 ( .A1(n8781), .A2(n6488), .B1(n7619), .B2(n6487), .C1(
        P2_U3152), .C2(n5004), .ZN(P2_U3354) );
  INV_X1 U7624 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6499) );
  NAND3_X1 U7625 ( .A1(n6490), .A2(P1_B_REG_SCAN_IN), .A3(n7749), .ZN(n6493)
         );
  INV_X1 U7626 ( .A(n7749), .ZN(n6491) );
  INV_X1 U7627 ( .A(P1_B_REG_SCAN_IN), .ZN(n9545) );
  NAND2_X1 U7628 ( .A1(n6491), .A2(n9545), .ZN(n6492) );
  AND2_X1 U7629 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  NAND2_X1 U7630 ( .A1(n6495), .A2(n6494), .ZN(n6629) );
  INV_X1 U7631 ( .A(n6629), .ZN(n9901) );
  NAND2_X1 U7632 ( .A1(n9901), .A2(n6499), .ZN(n6497) );
  INV_X1 U7633 ( .A(n6495), .ZN(n7964) );
  NAND2_X1 U7634 ( .A1(n7964), .A2(n6490), .ZN(n6496) );
  NAND2_X1 U7635 ( .A1(n6497), .A2(n6496), .ZN(n7101) );
  INV_X1 U7636 ( .A(n7101), .ZN(n6718) );
  NAND2_X1 U7637 ( .A1(n6718), .A2(n6728), .ZN(n6498) );
  OAI21_X1 U7638 ( .B1(n6728), .B2(n6499), .A(n6498), .ZN(P1_U3441) );
  INV_X1 U7639 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6919) );
  OAI222_X1 U7640 ( .A1(n10319), .A2(P1_U3084), .B1(n8777), .B2(n6693), .C1(
        n8775), .C2(n6919), .ZN(P1_U3351) );
  INV_X1 U7641 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6900) );
  OAI222_X1 U7642 ( .A1(n6780), .A2(P1_U3084), .B1(n8777), .B2(n6781), .C1(
        n8775), .C2(n6900), .ZN(P1_U3350) );
  INV_X1 U7643 ( .A(n10258), .ZN(n6501) );
  INV_X1 U7644 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6909) );
  OAI222_X1 U7645 ( .A1(n6501), .A2(P1_U3084), .B1(n8777), .B2(n6500), .C1(
        n8775), .C2(n6909), .ZN(P1_U3348) );
  INV_X1 U7646 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6503) );
  INV_X1 U7647 ( .A(n6945), .ZN(n6504) );
  OAI222_X1 U7648 ( .A1(n8781), .A2(n6503), .B1(n7619), .B2(n6504), .C1(
        P2_U3152), .C2(n6502), .ZN(P2_U3352) );
  INV_X1 U7649 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6903) );
  OAI222_X1 U7650 ( .A1(n6505), .A2(P1_U3084), .B1(n8777), .B2(n6504), .C1(
        n8775), .C2(n6903), .ZN(P1_U3347) );
  INV_X1 U7651 ( .A(n7022), .ZN(n6508) );
  INV_X1 U7652 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6906) );
  OAI222_X1 U7653 ( .A1(n6506), .A2(P1_U3084), .B1(n8777), .B2(n6508), .C1(
        n8775), .C2(n6906), .ZN(P1_U3346) );
  INV_X1 U7654 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6509) );
  OAI222_X1 U7655 ( .A1(n8781), .A2(n6509), .B1(n7619), .B2(n6508), .C1(
        P2_U3152), .C2(n6507), .ZN(P2_U3351) );
  INV_X1 U7656 ( .A(n7277), .ZN(n6511) );
  OAI222_X1 U7657 ( .A1(n6594), .A2(P1_U3084), .B1(n8777), .B2(n6511), .C1(
        n8775), .C2(n5505), .ZN(P1_U3345) );
  OAI222_X1 U7658 ( .A1(n8781), .A2(n6512), .B1(n7619), .B2(n6511), .C1(
        P2_U3152), .C2(n6510), .ZN(P2_U3350) );
  INV_X1 U7659 ( .A(n7270), .ZN(n6514) );
  OAI222_X1 U7660 ( .A1(n8777), .A2(n6514), .B1(n8775), .B2(n5510), .C1(
        P1_U3084), .C2(n6610), .ZN(P1_U3344) );
  OAI222_X1 U7661 ( .A1(P2_U3152), .A2(n6515), .B1(n7619), .B2(n6514), .C1(
        n6513), .C2(n8781), .ZN(P2_U3349) );
  INV_X1 U7662 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6529) );
  INV_X1 U7663 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6517) );
  INV_X1 U7664 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U7665 ( .A1(n6519), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n6520) );
  AND2_X2 U7666 ( .A1(n6521), .A2(n6523), .ZN(n6823) );
  NAND2_X1 U7667 ( .A1(n6823), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U7668 ( .A1(n6801), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U7669 ( .A1(n4874), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U7670 ( .A1(n6800), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U7671 ( .A1(n10355), .A2(P1_U4006), .ZN(n6528) );
  OAI21_X1 U7672 ( .B1(P1_U4006), .B2(n6529), .A(n6528), .ZN(P1_U3555) );
  INV_X1 U7673 ( .A(n7482), .ZN(n6532) );
  OAI222_X1 U7674 ( .A1(n8777), .A2(n6532), .B1(n6681), .B2(P1_U3084), .C1(
        n6530), .C2(n8775), .ZN(P1_U3343) );
  OAI222_X1 U7675 ( .A1(n8781), .A2(n6533), .B1(n7619), .B2(n6532), .C1(n6531), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7676 ( .A(n7521), .ZN(n6541) );
  INV_X1 U7677 ( .A(n10238), .ZN(n10230) );
  INV_X1 U7678 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6534) );
  OAI222_X1 U7679 ( .A1(n8777), .A2(n6541), .B1(n10230), .B2(P1_U3084), .C1(
        n6534), .C2(n8775), .ZN(P1_U3342) );
  NAND2_X1 U7680 ( .A1(n4830), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U7681 ( .A1(n6535), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U7682 ( .A1(n6536), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6537) );
  AND3_X1 U7683 ( .A1(n6539), .A2(n6538), .A3(n6537), .ZN(n8926) );
  NAND2_X1 U7684 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n8861), .ZN(n6540) );
  OAI21_X1 U7685 ( .B1(n8926), .B2(n8861), .A(n6540), .ZN(P2_U3582) );
  INV_X1 U7686 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6542) );
  INV_X1 U7687 ( .A(n7546), .ZN(n7203) );
  OAI222_X1 U7688 ( .A1(n8781), .A2(n6542), .B1(n7619), .B2(n6541), .C1(n7203), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  NAND2_X1 U7689 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n8861), .ZN(n6543) );
  OAI21_X1 U7690 ( .B1(n8234), .B2(n8861), .A(n6543), .ZN(P2_U3570) );
  AOI21_X1 U7691 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(n6554) );
  INV_X1 U7692 ( .A(n10312), .ZN(n10259) );
  AOI21_X1 U7693 ( .B1(n6549), .B2(n6548), .A(n6547), .ZN(n6551) );
  INV_X1 U7694 ( .A(n10318), .ZN(n10257) );
  AND2_X1 U7695 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7041) );
  AOI21_X1 U7696 ( .B1(n10257), .B2(n7023), .A(n7041), .ZN(n6550) );
  OAI21_X1 U7697 ( .B1(n6551), .B2(n10236), .A(n6550), .ZN(n6552) );
  AOI21_X1 U7698 ( .B1(n10259), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6552), .ZN(
        n6553) );
  OAI21_X1 U7699 ( .B1(n6554), .B2(n10321), .A(n6553), .ZN(P1_U3248) );
  INV_X1 U7700 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6564) );
  INV_X1 U7701 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6652) );
  NOR2_X1 U7702 ( .A1(n10200), .A2(n6652), .ZN(n6556) );
  INV_X1 U7703 ( .A(n10236), .ZN(n10329) );
  OAI211_X1 U7704 ( .C1(n6557), .C2(n6556), .A(n10329), .B(n6555), .ZN(n6559)
         );
  NAND2_X1 U7705 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n6558) );
  OAI211_X1 U7706 ( .C1(n10318), .C2(n6702), .A(n6559), .B(n6558), .ZN(n6560)
         );
  INV_X1 U7707 ( .A(n6560), .ZN(n6563) );
  NAND2_X1 U7708 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6659) );
  INV_X1 U7709 ( .A(n10321), .ZN(n10226) );
  OAI211_X1 U7710 ( .C1(n6324), .C2(n6561), .A(n10226), .B(n10314), .ZN(n6562)
         );
  OAI211_X1 U7711 ( .C1(n10312), .C2(n6564), .A(n6563), .B(n6562), .ZN(
        P1_U3242) );
  INV_X1 U7712 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U7713 ( .A1(n6800), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U7714 ( .A1(n6801), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U7715 ( .A1(n4874), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6565) );
  AND3_X1 U7716 ( .A1(n6567), .A2(n6566), .A3(n6565), .ZN(n9351) );
  INV_X1 U7717 ( .A(n9351), .ZN(n9558) );
  NAND2_X1 U7718 ( .A1(n9558), .A2(P1_U4006), .ZN(n6568) );
  OAI21_X1 U7719 ( .B1(P1_U4006), .B2(n6569), .A(n6568), .ZN(P1_U3586) );
  INV_X1 U7720 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6583) );
  INV_X1 U7721 ( .A(n6780), .ZN(n6575) );
  AND2_X1 U7722 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6874) );
  INV_X1 U7723 ( .A(n6570), .ZN(n6571) );
  AOI211_X1 U7724 ( .C1(n6573), .C2(n6572), .A(n6571), .B(n10321), .ZN(n6574)
         );
  AOI211_X1 U7725 ( .C1(n10257), .C2(n6575), .A(n6874), .B(n6574), .ZN(n6582)
         );
  MUX2_X1 U7726 ( .A(n6576), .B(P1_REG1_REG_3__SCAN_IN), .S(n6780), .Z(n6580)
         );
  INV_X1 U7727 ( .A(n6577), .ZN(n6579) );
  OAI211_X1 U7728 ( .C1(n6580), .C2(n6579), .A(n10329), .B(n6578), .ZN(n6581)
         );
  OAI211_X1 U7729 ( .C1(n10312), .C2(n6583), .A(n6582), .B(n6581), .ZN(
        P1_U3244) );
  INV_X1 U7730 ( .A(n8893), .ZN(n10296) );
  NOR2_X1 U7731 ( .A1(n10296), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7732 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6589) );
  INV_X1 U7733 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U7734 ( .A1(n4831), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6587) );
  INV_X1 U7735 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6585) );
  OR2_X1 U7736 ( .A1(n5720), .A2(n6585), .ZN(n6586) );
  OAI211_X1 U7737 ( .C1(n5633), .C2(n8905), .A(n6587), .B(n6586), .ZN(n8588)
         );
  NAND2_X1 U7738 ( .A1(n8588), .A2(P2_U3966), .ZN(n6588) );
  OAI21_X1 U7739 ( .B1(n6589), .B2(P2_U3966), .A(n6588), .ZN(P2_U3583) );
  AOI21_X1 U7740 ( .B1(n6592), .B2(n6591), .A(n6590), .ZN(n6602) );
  INV_X1 U7741 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7034) );
  NOR2_X1 U7742 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7034), .ZN(n7329) );
  INV_X1 U7743 ( .A(n7329), .ZN(n6593) );
  OAI21_X1 U7744 ( .B1(n10318), .B2(n6594), .A(n6593), .ZN(n6600) );
  AOI21_X1 U7745 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(n6598) );
  NOR2_X1 U7746 ( .A1(n6598), .A2(n10236), .ZN(n6599) );
  AOI211_X1 U7747 ( .C1(n10259), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n6600), .B(
        n6599), .ZN(n6601) );
  OAI21_X1 U7748 ( .B1(n6602), .B2(n10321), .A(n6601), .ZN(P1_U3249) );
  AOI21_X1 U7749 ( .B1(n6605), .B2(n6604), .A(n6603), .ZN(n6614) );
  OAI211_X1 U7750 ( .C1(n6608), .C2(n6607), .A(n10226), .B(n6606), .ZN(n6613)
         );
  AND2_X1 U7751 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7319) );
  INV_X1 U7752 ( .A(n7319), .ZN(n6609) );
  OAI21_X1 U7753 ( .B1(n10318), .B2(n6610), .A(n6609), .ZN(n6611) );
  AOI21_X1 U7754 ( .B1(n10259), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n6611), .ZN(
        n6612) );
  OAI211_X1 U7755 ( .C1(n6614), .C2(n10236), .A(n6613), .B(n6612), .ZN(
        P1_U3250) );
  INV_X1 U7756 ( .A(n7675), .ZN(n6645) );
  AOI22_X1 U7757 ( .A1(n7567), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8410), .ZN(n6615) );
  OAI21_X1 U7758 ( .B1(n6645), .B2(n7619), .A(n6615), .ZN(P2_U3346) );
  XNOR2_X1 U7759 ( .A(n6617), .B(n6616), .ZN(n7388) );
  OR2_X1 U7760 ( .A1(n6715), .A2(n7105), .ZN(n6816) );
  NAND2_X1 U7761 ( .A1(n6816), .A2(n6728), .ZN(n6722) );
  NOR4_X1 U7762 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6621) );
  NOR4_X1 U7763 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6620) );
  NOR4_X1 U7764 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6619) );
  NOR4_X1 U7765 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6618) );
  NAND4_X1 U7766 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n6627)
         );
  NOR2_X1 U7767 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n6625) );
  NOR4_X1 U7768 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6624) );
  NOR4_X1 U7769 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6623) );
  NOR4_X1 U7770 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6622) );
  NAND4_X1 U7771 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6626)
         );
  NOR2_X1 U7772 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  NOR2_X1 U7773 ( .A1(n6629), .A2(n6628), .ZN(n6716) );
  INV_X1 U7774 ( .A(n7388), .ZN(n9538) );
  OAI21_X1 U7775 ( .B1(n10552), .B2(n6234), .A(n7101), .ZN(n6630) );
  NOR2_X1 U7776 ( .A1(n7100), .A2(n6630), .ZN(n7640) );
  INV_X1 U7777 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U7778 ( .A1(n9901), .A2(n6631), .ZN(n6632) );
  NAND2_X1 U7779 ( .A1(n7964), .A2(n7749), .ZN(n9903) );
  INV_X1 U7780 ( .A(n7639), .ZN(n6633) );
  AND2_X2 U7781 ( .A1(n7640), .A2(n6633), .ZN(n10595) );
  INV_X1 U7782 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U7783 ( .A1(n8257), .A2(SI_0_), .ZN(n6635) );
  INV_X1 U7784 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U7785 ( .A1(n6635), .A2(n6634), .ZN(n6637) );
  AND2_X1 U7786 ( .A1(n6637), .A2(n6636), .ZN(n9904) );
  MUX2_X1 U7787 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9904), .S(n6694), .Z(n7097) );
  INV_X1 U7788 ( .A(n6234), .ZN(n7462) );
  INV_X1 U7789 ( .A(n7261), .ZN(n6641) );
  INV_X1 U7790 ( .A(n9745), .ZN(n10514) );
  NAND2_X1 U7791 ( .A1(n6800), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U7792 ( .A1(n6823), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6638) );
  NOR2_X1 U7793 ( .A1(n10355), .A2(n10350), .ZN(n10352) );
  AND2_X1 U7794 ( .A1(n10355), .A2(n10350), .ZN(n9505) );
  NOR2_X1 U7795 ( .A1(n10352), .A2(n9505), .ZN(n9354) );
  INV_X1 U7796 ( .A(n7105), .ZN(n9540) );
  OR2_X1 U7797 ( .A1(n6715), .A2(n9540), .ZN(n7112) );
  INV_X1 U7798 ( .A(n7112), .ZN(n7489) );
  NOR3_X1 U7799 ( .A1(n9354), .A2(n7489), .A3(n7261), .ZN(n6640) );
  AOI21_X1 U7800 ( .B1(n10514), .B2(n9765), .A(n6640), .ZN(n10334) );
  OAI21_X1 U7801 ( .B1(n10350), .B2(n6641), .A(n10334), .ZN(n9881) );
  NAND2_X1 U7802 ( .A1(n9881), .A2(n10595), .ZN(n6642) );
  OAI21_X1 U7803 ( .B1(n10595), .B2(n6643), .A(n6642), .ZN(P1_U3454) );
  INV_X1 U7804 ( .A(n7676), .ZN(n7058) );
  INV_X1 U7805 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6644) );
  OAI222_X1 U7806 ( .A1(n8777), .A2(n6645), .B1(n7058), .B2(P1_U3084), .C1(
        n6644), .C2(n8775), .ZN(P1_U3341) );
  OAI22_X1 U7807 ( .A1(n8763), .A2(n10350), .B1(n6815), .B2(n10200), .ZN(n6648) );
  INV_X1 U7808 ( .A(n6648), .ZN(n6651) );
  OR2_X1 U7809 ( .A1(n6698), .A2(n9540), .ZN(n6649) );
  NAND2_X1 U7810 ( .A1(n6950), .A2(n10355), .ZN(n6650) );
  AND2_X1 U7811 ( .A1(n6651), .A2(n6650), .ZN(n6657) );
  NAND2_X1 U7812 ( .A1(n6951), .A2(n10355), .ZN(n6656) );
  OR2_X1 U7813 ( .A1(n10350), .A2(n8764), .ZN(n6654) );
  AND2_X1 U7814 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  NAND2_X1 U7815 ( .A1(n6656), .A2(n6655), .ZN(n6713) );
  NAND2_X1 U7816 ( .A1(n6657), .A2(n6713), .ZN(n6712) );
  OR2_X1 U7817 ( .A1(n6657), .A2(n6713), .ZN(n6658) );
  NAND2_X1 U7818 ( .A1(n6712), .A2(n6658), .ZN(n6742) );
  MUX2_X1 U7819 ( .A(n6742), .B(n6659), .S(n10198), .Z(n6662) );
  NOR2_X1 U7820 ( .A1(n10220), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6660) );
  OR2_X1 U7821 ( .A1(n6311), .A2(n6660), .ZN(n10201) );
  AOI21_X1 U7822 ( .B1(n10200), .B2(n10201), .A(n9557), .ZN(n6661) );
  OAI21_X1 U7823 ( .B1(n6662), .B2(n6311), .A(n6661), .ZN(n10325) );
  AOI21_X1 U7824 ( .B1(n6665), .B2(n6664), .A(n6663), .ZN(n6666) );
  NOR2_X1 U7825 ( .A1(n10236), .A2(n6666), .ZN(n6674) );
  AOI21_X1 U7826 ( .B1(n6669), .B2(n6668), .A(n6667), .ZN(n6672) );
  NAND2_X1 U7827 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n6831) );
  NAND2_X1 U7828 ( .A1(n10257), .A2(n6670), .ZN(n6671) );
  OAI211_X1 U7829 ( .C1(n10321), .C2(n6672), .A(n6831), .B(n6671), .ZN(n6673)
         );
  AOI211_X1 U7830 ( .C1(n10259), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n6674), .B(
        n6673), .ZN(n6675) );
  NAND2_X1 U7831 ( .A1(n10325), .A2(n6675), .ZN(P1_U3245) );
  INV_X1 U7832 ( .A(n7707), .ZN(n6741) );
  INV_X1 U7833 ( .A(n7708), .ZN(n6676) );
  OAI222_X1 U7834 ( .A1(n8777), .A2(n6741), .B1(n8775), .B2(n5529), .C1(
        P1_U3084), .C2(n6676), .ZN(P1_U3340) );
  AOI21_X1 U7835 ( .B1(n6679), .B2(n6678), .A(n6677), .ZN(n6688) );
  INV_X1 U7836 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7312) );
  NOR2_X1 U7837 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7312), .ZN(n7512) );
  INV_X1 U7838 ( .A(n7512), .ZN(n6680) );
  OAI21_X1 U7839 ( .B1(n10318), .B2(n6681), .A(n6680), .ZN(n6682) );
  AOI21_X1 U7840 ( .B1(n10259), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6682), .ZN(
        n6687) );
  OAI211_X1 U7841 ( .C1(n6685), .C2(n6684), .A(n10226), .B(n6683), .ZN(n6686)
         );
  OAI211_X1 U7842 ( .C1(n6688), .C2(n10236), .A(n6687), .B(n6686), .ZN(
        P1_U3251) );
  NAND2_X1 U7843 ( .A1(n6823), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U7844 ( .A1(n6800), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U7845 ( .A1(n4874), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U7846 ( .A1(n6801), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U7847 ( .A1(n6694), .A2(n8257), .ZN(n6806) );
  OR2_X1 U7848 ( .A1(n6806), .A2(n6693), .ZN(n6696) );
  NAND2_X4 U7849 ( .A1(n6694), .A2(n4832), .ZN(n9345) );
  NAND2_X1 U7850 ( .A1(n6698), .A2(n9697), .ZN(n6699) );
  NAND2_X4 U7851 ( .A1(n6699), .A2(n7110), .ZN(n8761) );
  XNOR2_X1 U7852 ( .A(n6700), .B(n4836), .ZN(n6797) );
  OAI22_X1 U7853 ( .A1(n8760), .A2(n7118), .B1(n10385), .B2(n8763), .ZN(n6795)
         );
  XNOR2_X1 U7854 ( .A(n6797), .B(n6795), .ZN(n6793) );
  OR2_X1 U7855 ( .A1(n6806), .A2(n8412), .ZN(n6706) );
  INV_X2 U7856 ( .A(n6694), .ZN(n6704) );
  INV_X1 U7857 ( .A(n6702), .ZN(n6703) );
  INV_X1 U7858 ( .A(n10351), .ZN(n6708) );
  NAND2_X1 U7859 ( .A1(n6708), .A2(n4856), .ZN(n6709) );
  NAND2_X1 U7860 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  OAI22_X1 U7861 ( .A1(n8760), .A2(n7113), .B1(n10351), .B2(n8763), .ZN(n6890)
         );
  NAND2_X1 U7862 ( .A1(n6892), .A2(n6890), .ZN(n6714) );
  OAI21_X1 U7863 ( .B1(n4854), .B2(n6713), .A(n6712), .ZN(n6889) );
  XOR2_X1 U7864 ( .A(n6793), .B(n6794), .Z(n6739) );
  INV_X1 U7865 ( .A(n6715), .ZN(n9498) );
  OR2_X1 U7866 ( .A1(n10549), .A2(n9498), .ZN(n6819) );
  INV_X1 U7867 ( .A(n6716), .ZN(n6717) );
  AND3_X1 U7868 ( .A1(n6718), .A2(n7639), .A3(n6717), .ZN(n6818) );
  INV_X1 U7869 ( .A(n6818), .ZN(n6729) );
  INV_X1 U7870 ( .A(n6728), .ZN(n9902) );
  NOR2_X1 U7871 ( .A1(n6729), .A2(n9902), .ZN(n6724) );
  INV_X1 U7872 ( .A(n6724), .ZN(n6719) );
  NAND2_X1 U7873 ( .A1(n7261), .A2(n9538), .ZN(n10485) );
  NAND2_X1 U7874 ( .A1(n10485), .A2(n7112), .ZN(n6721) );
  AND2_X1 U7875 ( .A1(n6729), .A2(n6728), .ZN(n6720) );
  NAND2_X1 U7876 ( .A1(n6721), .A2(n6720), .ZN(n6821) );
  INV_X1 U7877 ( .A(n6722), .ZN(n6723) );
  OAI211_X1 U7878 ( .C1(n10549), .C2(n6818), .A(n6821), .B(n6723), .ZN(n6895)
         );
  INV_X1 U7879 ( .A(n10485), .ZN(n10364) );
  NAND2_X1 U7880 ( .A1(n10364), .A2(n6724), .ZN(n6726) );
  OR2_X1 U7881 ( .A1(n6234), .A2(n9902), .ZN(n6725) );
  NAND2_X1 U7882 ( .A1(n6726), .A2(n10488), .ZN(n9287) );
  NAND2_X1 U7883 ( .A1(n7105), .A2(n6728), .ZN(n9291) );
  OR2_X1 U7884 ( .A1(n6729), .A2(n9291), .ZN(n6731) );
  INV_X1 U7885 ( .A(n6731), .ZN(n6730) );
  NAND2_X1 U7886 ( .A1(n10516), .A2(n6730), .ZN(n9284) );
  INV_X1 U7887 ( .A(n9284), .ZN(n9250) );
  NAND2_X1 U7888 ( .A1(n6800), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6735) );
  INV_X1 U7889 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U7890 ( .A1(n6801), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U7891 ( .A1(n4874), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6732) );
  AOI22_X1 U7892 ( .A1(n9250), .A2(n9765), .B1(n9262), .B2(n6779), .ZN(n6736)
         );
  OAI21_X1 U7893 ( .B1(n10385), .B2(n9224), .A(n6736), .ZN(n6737) );
  AOI21_X1 U7894 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6895), .A(n6737), .ZN(
        n6738) );
  OAI21_X1 U7895 ( .B1(n6739), .B2(n9289), .A(n6738), .ZN(P1_U3235) );
  INV_X1 U7896 ( .A(n7650), .ZN(n7555) );
  OAI222_X1 U7897 ( .A1(P2_U3152), .A2(n7555), .B1(n7619), .B2(n6741), .C1(
        n6740), .C2(n8781), .ZN(P2_U3345) );
  INV_X1 U7898 ( .A(n6742), .ZN(n6745) );
  INV_X1 U7899 ( .A(n9262), .ZN(n9242) );
  OAI22_X1 U7900 ( .A1(n9224), .A2(n10350), .B1(n9242), .B2(n7113), .ZN(n6743)
         );
  AOI21_X1 U7901 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6895), .A(n6743), .ZN(
        n6744) );
  OAI21_X1 U7902 ( .B1(n6745), .B2(n9289), .A(n6744), .ZN(P1_U3230) );
  INV_X1 U7903 ( .A(n7806), .ZN(n6838) );
  AOI22_X1 U7904 ( .A1(n7807), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n6980), .ZN(n6746) );
  OAI21_X1 U7905 ( .B1(n6838), .B2(n8777), .A(n6746), .ZN(P1_U3339) );
  INV_X1 U7906 ( .A(n8913), .ZN(n9083) );
  NAND2_X1 U7907 ( .A1(n9083), .A2(P2_U3966), .ZN(n6747) );
  OAI21_X1 U7908 ( .B1(n5554), .B2(P2_U3966), .A(n6747), .ZN(P2_U3571) );
  NOR2_X1 U7909 ( .A1(n6748), .A2(P2_U3152), .ZN(n10404) );
  OAI21_X1 U7910 ( .B1(n6751), .B2(n6750), .A(n6749), .ZN(n6752) );
  INV_X1 U7911 ( .A(n8862), .ZN(n6912) );
  OAI22_X1 U7912 ( .A1(n6912), .A2(n10439), .B1(n7071), .B2(n10441), .ZN(n6765) );
  AOI22_X1 U7913 ( .A1(n8844), .A2(n6752), .B1(n8815), .B2(n6765), .ZN(n6754)
         );
  NAND2_X1 U7914 ( .A1(n8851), .A2(n6768), .ZN(n6753) );
  OAI211_X1 U7915 ( .C1(n10404), .C2(n10372), .A(n6754), .B(n6753), .ZN(
        P2_U3224) );
  NAND2_X1 U7916 ( .A1(n6756), .A2(n8640), .ZN(n6757) );
  NAND2_X1 U7917 ( .A1(n6758), .A2(n6757), .ZN(n6773) );
  INV_X1 U7918 ( .A(n6773), .ZN(n6759) );
  AND2_X2 U7919 ( .A1(n6776), .A2(n7154), .ZN(n10650) );
  INV_X1 U7920 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U7921 ( .A1(n6760), .A2(n10378), .ZN(n7081) );
  NAND2_X1 U7922 ( .A1(n10392), .A2(n6768), .ZN(n8464) );
  NAND2_X1 U7923 ( .A1(n7081), .A2(n8464), .ZN(n7067) );
  XNOR2_X1 U7924 ( .A(n7067), .B(n7066), .ZN(n10380) );
  INV_X1 U7925 ( .A(n10380), .ZN(n6770) );
  NOR2_X1 U7926 ( .A1(n6761), .A2(n8598), .ZN(n6762) );
  OR2_X1 U7927 ( .A1(n6763), .A2(n6762), .ZN(n7450) );
  INV_X1 U7928 ( .A(n10609), .ZN(n6764) );
  XNOR2_X1 U7929 ( .A(n8599), .B(n7067), .ZN(n6766) );
  NAND2_X1 U7930 ( .A1(n8641), .A2(n8973), .ZN(n8593) );
  AOI21_X1 U7931 ( .B1(n6766), .B2(n9085), .A(n6765), .ZN(n10376) );
  AND2_X1 U7932 ( .A1(n6768), .A2(n10339), .ZN(n6767) );
  NOR2_X1 U7933 ( .A1(n7361), .A2(n6767), .ZN(n10375) );
  AOI22_X1 U7934 ( .A1(n10375), .A2(n10449), .B1(n10150), .B2(n6768), .ZN(
        n6769) );
  OAI211_X1 U7935 ( .C1(n6770), .C2(n10620), .A(n10376), .B(n6769), .ZN(n6777)
         );
  NAND2_X1 U7936 ( .A1(n10650), .A2(n6777), .ZN(n6771) );
  OAI21_X1 U7937 ( .B1(n10650), .B2(n6772), .A(n6771), .ZN(P2_U3454) );
  NOR2_X1 U7938 ( .A1(n6774), .A2(n6773), .ZN(n6775) );
  AND2_X2 U7939 ( .A1(n6776), .A2(n6775), .ZN(n10646) );
  NAND2_X1 U7940 ( .A1(n10646), .A2(n6777), .ZN(n6778) );
  OAI21_X1 U7941 ( .B1(n10646), .B2(n6372), .A(n6778), .ZN(P2_U3521) );
  NAND2_X1 U7942 ( .A1(n6779), .A2(n6951), .ZN(n6786) );
  OR2_X1 U7943 ( .A1(n6694), .A2(n6780), .ZN(n6784) );
  OR2_X1 U7944 ( .A1(n9345), .A2(n6900), .ZN(n6783) );
  OR2_X1 U7945 ( .A1(n6806), .A2(n6781), .ZN(n6782) );
  NAND2_X1 U7946 ( .A1(n7104), .A2(n4856), .ZN(n6785) );
  NAND2_X1 U7947 ( .A1(n6786), .A2(n6785), .ZN(n6787) );
  XNOR2_X1 U7948 ( .A(n6787), .B(n4836), .ZN(n6791) );
  INV_X1 U7949 ( .A(n7104), .ZN(n10413) );
  XNOR2_X1 U7950 ( .A(n6791), .B(n6789), .ZN(n6870) );
  INV_X1 U7951 ( .A(n6870), .ZN(n6792) );
  INV_X1 U7952 ( .A(n6789), .ZN(n6790) );
  NAND2_X1 U7953 ( .A1(n6792), .A2(n4829), .ZN(n6839) );
  INV_X1 U7954 ( .A(n6795), .ZN(n6796) );
  NAND2_X1 U7955 ( .A1(n6797), .A2(n6796), .ZN(n6871) );
  NAND2_X1 U7956 ( .A1(n6847), .A2(n6846), .ZN(n6798) );
  AND2_X1 U7957 ( .A1(n6839), .A2(n6798), .ZN(n6814) );
  NAND2_X1 U7958 ( .A1(n4874), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6805) );
  INV_X1 U7959 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6799) );
  XNOR2_X1 U7960 ( .A(n6799), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7127) );
  NAND2_X1 U7961 ( .A1(n6823), .A2(n7127), .ZN(n6804) );
  NAND2_X1 U7962 ( .A1(n6800), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U7963 ( .A1(n6801), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U7964 ( .A1(n6944), .A2(n6807), .ZN(n6810) );
  OR2_X1 U7965 ( .A1(n9345), .A2(n6808), .ZN(n6809) );
  OAI211_X1 U7966 ( .C1(n6811), .C2(n6694), .A(n6810), .B(n6809), .ZN(n7125)
         );
  OAI22_X1 U7967 ( .A1(n7240), .A2(n8763), .B1(n4835), .B2(n8764), .ZN(n6812)
         );
  XNOR2_X1 U7968 ( .A(n6812), .B(n8761), .ZN(n6841) );
  OAI22_X1 U7969 ( .A1(n8760), .A2(n7240), .B1(n4835), .B2(n8763), .ZN(n6840)
         );
  XNOR2_X1 U7970 ( .A(n6841), .B(n6840), .ZN(n6813) );
  XNOR2_X1 U7971 ( .A(n6814), .B(n6813), .ZN(n6836) );
  AND3_X1 U7972 ( .A1(n6816), .A2(n6815), .A3(n7702), .ZN(n6817) );
  OAI21_X1 U7973 ( .B1(n6819), .B2(n6818), .A(n6817), .ZN(n6820) );
  NAND2_X1 U7974 ( .A1(n6820), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6822) );
  NAND3_X1 U7975 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6858) );
  INV_X1 U7976 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U7977 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6824) );
  NAND2_X1 U7978 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  AND2_X1 U7979 ( .A1(n6858), .A2(n6826), .ZN(n10484) );
  NAND2_X1 U7980 ( .A1(n6823), .A2(n10484), .ZN(n6830) );
  NAND2_X1 U7981 ( .A1(n6800), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U7982 ( .A1(n4874), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U7983 ( .A1(n6801), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6827) );
  OAI21_X1 U7984 ( .B1(n9242), .B2(n7247), .A(n6831), .ZN(n6832) );
  AOI21_X1 U7985 ( .B1(n9250), .B2(n6779), .A(n6832), .ZN(n6833) );
  OAI21_X1 U7986 ( .B1(n4835), .B2(n9224), .A(n6833), .ZN(n6834) );
  AOI21_X1 U7987 ( .B1(n7127), .B2(n9280), .A(n6834), .ZN(n6835) );
  OAI21_X1 U7988 ( .B1(n6836), .B2(n9289), .A(n6835), .ZN(P1_U3228) );
  INV_X1 U7989 ( .A(n7973), .ZN(n7659) );
  INV_X1 U7990 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6837) );
  OAI222_X1 U7991 ( .A1(P2_U3152), .A2(n7659), .B1(n7619), .B2(n6838), .C1(
        n6837), .C2(n8781), .ZN(P2_U3344) );
  NOR2_X1 U7992 ( .A1(n6841), .A2(n6840), .ZN(n6844) );
  NOR2_X1 U7993 ( .A1(n6839), .A2(n6844), .ZN(n6843) );
  AND2_X1 U7994 ( .A1(n6841), .A2(n6840), .ZN(n6842) );
  NOR2_X1 U7995 ( .A1(n6843), .A2(n6842), .ZN(n6849) );
  INV_X1 U7996 ( .A(n6844), .ZN(n6845) );
  NAND2_X1 U7997 ( .A1(n6849), .A2(n6848), .ZN(n6961) );
  AOI22_X1 U7998 ( .A1(n8280), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6704), .B2(
        n10258), .ZN(n6852) );
  NAND2_X1 U7999 ( .A1(n6850), .A2(n6944), .ZN(n6851) );
  NAND2_X1 U8000 ( .A1(n6852), .A2(n6851), .ZN(n7259) );
  NAND2_X1 U8001 ( .A1(n8752), .A2(n7259), .ZN(n6853) );
  OAI21_X1 U8002 ( .B1(n8760), .B2(n7247), .A(n6853), .ZN(n6959) );
  NAND2_X1 U8003 ( .A1(n4856), .A2(n7259), .ZN(n6854) );
  OAI21_X1 U8004 ( .B1(n7247), .B2(n8763), .A(n6854), .ZN(n6855) );
  XNOR2_X1 U8005 ( .A(n6855), .B(n8761), .ZN(n6960) );
  XOR2_X1 U8006 ( .A(n6959), .B(n6960), .Z(n6856) );
  XNOR2_X1 U8007 ( .A(n6961), .B(n6856), .ZN(n6869) );
  INV_X1 U8008 ( .A(n7259), .ZN(n10486) );
  NAND2_X1 U8009 ( .A1(n6800), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6863) );
  INV_X1 U8010 ( .A(n6858), .ZN(n6857) );
  INV_X1 U8011 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U8012 ( .A1(n6858), .A2(n6973), .ZN(n6859) );
  AND2_X1 U8013 ( .A1(n6967), .A2(n6859), .ZN(n10543) );
  NAND2_X1 U8014 ( .A1(n6823), .A2(n10543), .ZN(n6862) );
  NAND2_X1 U8015 ( .A1(n4874), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6861) );
  NAND2_X1 U8016 ( .A1(n6801), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U8017 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10268) );
  INV_X1 U8018 ( .A(n10268), .ZN(n6865) );
  NOR2_X1 U8019 ( .A1(n9284), .A2(n7240), .ZN(n6864) );
  AOI211_X1 U8020 ( .C1(n9262), .C2(n10474), .A(n6865), .B(n6864), .ZN(n6866)
         );
  OAI21_X1 U8021 ( .B1(n10486), .B2(n9224), .A(n6866), .ZN(n6867) );
  AOI21_X1 U8022 ( .B1(n10484), .B2(n9280), .A(n6867), .ZN(n6868) );
  OAI21_X1 U8023 ( .B1(n6869), .B2(n9289), .A(n6868), .ZN(P1_U3225) );
  NAND2_X1 U8024 ( .A1(n6847), .A2(n6871), .ZN(n6872) );
  XOR2_X1 U8025 ( .A(n6870), .B(n6872), .Z(n6879) );
  INV_X1 U8026 ( .A(n7240), .ZN(n10475) );
  NOR2_X1 U8027 ( .A1(n9284), .A2(n7118), .ZN(n6873) );
  AOI211_X1 U8028 ( .C1(n9262), .C2(n10475), .A(n6874), .B(n6873), .ZN(n6875)
         );
  OAI21_X1 U8029 ( .B1(n10413), .B2(n9224), .A(n6875), .ZN(n6876) );
  AOI21_X1 U8030 ( .B1(n6877), .B2(n9280), .A(n6876), .ZN(n6878) );
  OAI21_X1 U8031 ( .B1(n6879), .B2(n9289), .A(n6878), .ZN(P1_U3216) );
  INV_X1 U8032 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6880) );
  OAI22_X1 U8033 ( .A1(n10399), .A2(n10420), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6880), .ZN(n6881) );
  AOI21_X1 U8034 ( .B1(n8804), .B2(n7070), .A(n6881), .ZN(n6888) );
  NOR2_X1 U8035 ( .A1(n6883), .A2(n6882), .ZN(n6884) );
  NOR2_X1 U8036 ( .A1(n10397), .A2(n6884), .ZN(n6886) );
  AOI22_X1 U8037 ( .A1(n8802), .A2(n8860), .B1(n6886), .B2(n6885), .ZN(n6887)
         );
  OAI211_X1 U8038 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8848), .A(n6888), .B(
        n6887), .ZN(P2_U3220) );
  XNOR2_X1 U8039 ( .A(n6889), .B(n6890), .ZN(n6891) );
  XNOR2_X1 U8040 ( .A(n6892), .B(n6891), .ZN(n6897) );
  INV_X1 U8041 ( .A(n7118), .ZN(n10356) );
  AOI22_X1 U8042 ( .A1(n9250), .A2(n10355), .B1(n9262), .B2(n10356), .ZN(n6893) );
  OAI21_X1 U8043 ( .B1(n10351), .B2(n9224), .A(n6893), .ZN(n6894) );
  AOI21_X1 U8044 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6895), .A(n6894), .ZN(
        n6896) );
  OAI21_X1 U8045 ( .B1(n6897), .B2(n9289), .A(n6896), .ZN(P1_U3220) );
  INV_X1 U8046 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U8047 ( .A1(n9056), .A2(P2_U3966), .ZN(n6898) );
  OAI21_X1 U8048 ( .B1(n7463), .B2(P2_U3966), .A(n6898), .ZN(P2_U3573) );
  NAND2_X1 U8049 ( .A1(n7074), .A2(P2_U3966), .ZN(n6899) );
  OAI21_X1 U8050 ( .B1(n6900), .B2(P2_U3966), .A(n6899), .ZN(P2_U3555) );
  INV_X1 U8051 ( .A(n7952), .ZN(n8020) );
  NAND2_X1 U8052 ( .A1(n8020), .A2(P2_U3966), .ZN(n6901) );
  OAI21_X1 U8053 ( .B1(n5536), .B2(P2_U3966), .A(n6901), .ZN(P2_U3567) );
  NAND2_X1 U8054 ( .A1(n7206), .A2(P2_U3966), .ZN(n6902) );
  OAI21_X1 U8055 ( .B1(n6903), .B2(P2_U3966), .A(n6902), .ZN(P2_U3558) );
  NAND2_X1 U8056 ( .A1(n7423), .A2(P2_U3966), .ZN(n6904) );
  OAI21_X1 U8057 ( .B1(n5505), .B2(P2_U3966), .A(n6904), .ZN(P2_U3560) );
  NAND2_X1 U8058 ( .A1(n7412), .A2(P2_U3966), .ZN(n6905) );
  OAI21_X1 U8059 ( .B1(n6906), .B2(P2_U3966), .A(n6905), .ZN(P2_U3559) );
  INV_X1 U8060 ( .A(n7446), .ZN(n7439) );
  NAND2_X1 U8061 ( .A1(n7439), .A2(P2_U3966), .ZN(n6907) );
  OAI21_X1 U8062 ( .B1(n5510), .B2(P2_U3966), .A(n6907), .ZN(P2_U3561) );
  NAND2_X1 U8063 ( .A1(n7086), .A2(P2_U3966), .ZN(n6908) );
  OAI21_X1 U8064 ( .B1(n6909), .B2(P2_U3966), .A(n6908), .ZN(P2_U3557) );
  INV_X1 U8065 ( .A(n7882), .ZN(n7630) );
  NAND2_X1 U8066 ( .A1(n7630), .A2(P2_U3966), .ZN(n6910) );
  OAI21_X1 U8067 ( .B1(n5529), .B2(P2_U3966), .A(n6910), .ZN(P2_U3565) );
  OAI21_X1 U8068 ( .B1(n6912), .B2(n6911), .A(n7144), .ZN(n6913) );
  NAND3_X1 U8069 ( .A1(n8844), .A2(n6914), .A3(n6913), .ZN(n6915) );
  OAI21_X1 U8070 ( .B1(n10399), .B2(n7144), .A(n6915), .ZN(n6916) );
  AOI21_X1 U8071 ( .B1(n8802), .B2(n6760), .A(n6916), .ZN(n6917) );
  OAI21_X1 U8072 ( .B1(n10404), .B2(n10283), .A(n6917), .ZN(P2_U3234) );
  INV_X1 U8073 ( .A(n7071), .ZN(n7070) );
  NAND2_X1 U8074 ( .A1(n7070), .A2(P2_U3966), .ZN(n6918) );
  OAI21_X1 U8075 ( .B1(n6919), .B2(P2_U3966), .A(n6918), .ZN(P2_U3554) );
  INV_X1 U8076 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7687) );
  INV_X1 U8077 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7814) );
  INV_X1 U8078 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8077) );
  INV_X1 U8079 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8296) );
  INV_X1 U8080 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8308) );
  INV_X1 U8081 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U8082 ( .A1(n8323), .A2(n6930), .ZN(n6931) );
  NAND2_X1 U8083 ( .A1(n8340), .A2(n6931), .ZN(n9645) );
  OR2_X1 U8084 ( .A1(n9645), .A2(n8672), .ZN(n6937) );
  INV_X1 U8085 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U8086 ( .A1(n4874), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U8087 ( .A1(n6801), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6932) );
  OAI211_X1 U8088 ( .C1(n6934), .C2(n8676), .A(n6933), .B(n6932), .ZN(n6935)
         );
  INV_X1 U8089 ( .A(n6935), .ZN(n6936) );
  INV_X1 U8090 ( .A(n9239), .ZN(n9670) );
  NAND2_X1 U8091 ( .A1(n9670), .A2(P1_U4006), .ZN(n6938) );
  OAI21_X1 U8092 ( .B1(P1_U4006), .B2(n5997), .A(n6938), .ZN(P1_U3578) );
  INV_X1 U8093 ( .A(n8057), .ZN(n6940) );
  OAI222_X1 U8094 ( .A1(n8781), .A2(n6939), .B1(n7619), .B2(n6940), .C1(
        P2_U3152), .C2(n8015), .ZN(P2_U3343) );
  OAI222_X1 U8095 ( .A1(n8775), .A2(n5536), .B1(n8777), .B2(n6940), .C1(
        P1_U3084), .C2(n7790), .ZN(P1_U3338) );
  INV_X1 U8096 ( .A(n8062), .ZN(n6943) );
  INV_X1 U8097 ( .A(n8063), .ZN(n7948) );
  OAI222_X1 U8098 ( .A1(n8777), .A2(n6943), .B1(n7948), .B2(P1_U3084), .C1(
        n6941), .C2(n8775), .ZN(P1_U3337) );
  OAI222_X1 U8099 ( .A1(P2_U3152), .A2(n7969), .B1(n7619), .B2(n6943), .C1(
        n6942), .C2(n8781), .ZN(P2_U3342) );
  NAND2_X1 U8100 ( .A1(n6945), .A2(n6944), .ZN(n6947) );
  AOI22_X1 U8101 ( .A1(n8280), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6704), .B2(
        n10207), .ZN(n6946) );
  NAND2_X1 U8102 ( .A1(n6947), .A2(n6946), .ZN(n7260) );
  NAND2_X1 U8103 ( .A1(n7260), .A2(n4856), .ZN(n6948) );
  XNOR2_X1 U8104 ( .A(n6949), .B(n4854), .ZN(n6957) );
  INV_X1 U8105 ( .A(n6957), .ZN(n6955) );
  NAND2_X1 U8106 ( .A1(n10474), .A2(n8744), .ZN(n6953) );
  NAND2_X1 U8107 ( .A1(n7260), .A2(n8752), .ZN(n6952) );
  AND2_X1 U8108 ( .A1(n6953), .A2(n6952), .ZN(n6956) );
  INV_X1 U8109 ( .A(n6956), .ZN(n6954) );
  NAND2_X1 U8110 ( .A1(n6955), .A2(n6954), .ZN(n6958) );
  NAND2_X1 U8111 ( .A1(n6957), .A2(n6956), .ZN(n7029) );
  INV_X1 U8112 ( .A(n7030), .ZN(n6963) );
  AOI21_X1 U8113 ( .B1(n6965), .B2(n6964), .A(n6963), .ZN(n6978) );
  NAND2_X1 U8114 ( .A1(n6800), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6972) );
  INV_X1 U8115 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U8116 ( .A1(n6967), .A2(n6966), .ZN(n6968) );
  AND2_X1 U8117 ( .A1(n7035), .A2(n6968), .ZN(n7264) );
  NAND2_X1 U8118 ( .A1(n6823), .A2(n7264), .ZN(n6971) );
  NAND2_X1 U8119 ( .A1(n4874), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6970) );
  NAND2_X1 U8120 ( .A1(n6801), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U8121 ( .A1(n9280), .A2(n10543), .ZN(n6975) );
  NOR2_X1 U8122 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6973), .ZN(n10208) );
  AOI21_X1 U8123 ( .B1(n9250), .B2(n10515), .A(n10208), .ZN(n6974) );
  OAI211_X1 U8124 ( .C1(n7342), .C2(n9242), .A(n6975), .B(n6974), .ZN(n6976)
         );
  AOI21_X1 U8125 ( .B1(n7260), .B2(n9287), .A(n6976), .ZN(n6977) );
  OAI21_X1 U8126 ( .B1(n6978), .B2(n9289), .A(n6977), .ZN(P1_U3237) );
  INV_X1 U8127 ( .A(n8161), .ZN(n6982) );
  AOI22_X1 U8128 ( .A1(n8875), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8410), .ZN(n6979) );
  OAI21_X1 U8129 ( .B1(n6982), .B2(n7619), .A(n6979), .ZN(P2_U3341) );
  AOI22_X1 U8130 ( .A1(n8162), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6980), .ZN(n6981) );
  OAI21_X1 U8131 ( .B1(n6982), .B2(n8777), .A(n6981), .ZN(P1_U3336) );
  OAI21_X1 U8132 ( .B1(n6985), .B2(n6984), .A(n6983), .ZN(n6991) );
  INV_X1 U8133 ( .A(n7160), .ZN(n6986) );
  NAND2_X1 U8134 ( .A1(n8820), .A2(n6986), .ZN(n6988) );
  OAI211_X1 U8135 ( .C1(n7216), .C2(n10399), .A(n6988), .B(n6987), .ZN(n6990)
         );
  INV_X1 U8136 ( .A(n7086), .ZN(n10442) );
  OAI22_X1 U8137 ( .A1(n10442), .A2(n10393), .B1(n10394), .B2(n7403), .ZN(
        n6989) );
  AOI211_X1 U8138 ( .C1(n8844), .C2(n6991), .A(n6990), .B(n6989), .ZN(n6992)
         );
  INV_X1 U8139 ( .A(n6992), .ZN(P2_U3241) );
  OAI21_X1 U8140 ( .B1(n6995), .B2(n6994), .A(n6993), .ZN(n7001) );
  INV_X1 U8141 ( .A(n7183), .ZN(n6996) );
  NAND2_X1 U8142 ( .A1(n8820), .A2(n6996), .ZN(n6998) );
  OAI211_X1 U8143 ( .C1(n10501), .C2(n10399), .A(n6998), .B(n6997), .ZN(n7000)
         );
  INV_X1 U8144 ( .A(n8860), .ZN(n8477) );
  OAI22_X1 U8145 ( .A1(n8477), .A2(n10393), .B1(n10394), .B2(n7215), .ZN(n6999) );
  AOI211_X1 U8146 ( .C1(n8844), .C2(n7001), .A(n7000), .B(n6999), .ZN(n7002)
         );
  INV_X1 U8147 ( .A(n7002), .ZN(P2_U3229) );
  XNOR2_X1 U8148 ( .A(n7003), .B(n7004), .ZN(n7009) );
  AOI22_X1 U8149 ( .A1(n8804), .A2(n7206), .B1(n8802), .B2(n7423), .ZN(n7008)
         );
  INV_X1 U8150 ( .A(n7220), .ZN(n7006) );
  INV_X1 U8151 ( .A(n7411), .ZN(n10558) );
  OAI22_X1 U8152 ( .A1(n10399), .A2(n10558), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5722), .ZN(n7005) );
  AOI21_X1 U8153 ( .B1(n7006), .B2(n8820), .A(n7005), .ZN(n7007) );
  OAI211_X1 U8154 ( .C1(n7009), .C2(n10397), .A(n7008), .B(n7007), .ZN(
        P2_U3215) );
  NOR2_X1 U8155 ( .A1(n5321), .A2(n7011), .ZN(n7012) );
  XNOR2_X1 U8156 ( .A(n7013), .B(n7012), .ZN(n7019) );
  INV_X1 U8157 ( .A(n7014), .ZN(n10459) );
  OAI21_X1 U8158 ( .B1(n10399), .B2(n10451), .A(n7015), .ZN(n7017) );
  OAI22_X1 U8159 ( .A1(n10440), .A2(n10393), .B1(n10394), .B2(n10442), .ZN(
        n7016) );
  AOI211_X1 U8160 ( .C1(n10459), .C2(n8820), .A(n7017), .B(n7016), .ZN(n7018)
         );
  OAI21_X1 U8161 ( .B1(n7019), .B2(n10397), .A(n7018), .ZN(P2_U3232) );
  INV_X1 U8162 ( .A(n8997), .ZN(n7020) );
  NAND2_X1 U8163 ( .A1(n7020), .A2(P2_U3966), .ZN(n7021) );
  OAI21_X1 U8164 ( .B1(n8350), .B2(P2_U3966), .A(n7021), .ZN(P2_U3577) );
  NAND2_X1 U8165 ( .A1(n7022), .A2(n6944), .ZN(n7025) );
  AOI22_X1 U8166 ( .A1(n8280), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6704), .B2(
        n7023), .ZN(n7024) );
  NAND2_X1 U8167 ( .A1(n7025), .A2(n7024), .ZN(n10548) );
  INV_X1 U8168 ( .A(n10548), .ZN(n7266) );
  NAND2_X1 U8169 ( .A1(n10548), .A2(n4856), .ZN(n7027) );
  NAND2_X1 U8170 ( .A1(n10513), .A2(n8752), .ZN(n7026) );
  NAND2_X1 U8171 ( .A1(n7027), .A2(n7026), .ZN(n7028) );
  XNOR2_X1 U8172 ( .A(n7028), .B(n8761), .ZN(n7274) );
  AOI22_X1 U8173 ( .A1(n10548), .A2(n8752), .B1(n8744), .B2(n10513), .ZN(n7275) );
  XNOR2_X1 U8174 ( .A(n7274), .B(n7275), .ZN(n7032) );
  NAND2_X1 U8175 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  OAI21_X1 U8176 ( .B1(n7032), .B2(n7031), .A(n7301), .ZN(n7033) );
  NAND2_X1 U8177 ( .A1(n7033), .A2(n4834), .ZN(n7045) );
  NAND2_X1 U8178 ( .A1(n7035), .A2(n7034), .ZN(n7036) );
  AND2_X1 U8179 ( .A1(n7285), .A2(n7036), .ZN(n7349) );
  NAND2_X1 U8180 ( .A1(n6823), .A2(n7349), .ZN(n7040) );
  NAND2_X1 U8181 ( .A1(n6800), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7039) );
  NAND2_X1 U8182 ( .A1(n4874), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7038) );
  NAND2_X1 U8183 ( .A1(n6801), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7037) );
  AOI21_X1 U8184 ( .B1(n9262), .B2(n9556), .A(n7041), .ZN(n7042) );
  OAI21_X1 U8185 ( .B1(n7249), .B2(n9284), .A(n7042), .ZN(n7043) );
  AOI21_X1 U8186 ( .B1(n9280), .B2(n7264), .A(n7043), .ZN(n7044) );
  OAI211_X1 U8187 ( .C1(n7266), .C2(n9224), .A(n7045), .B(n7044), .ZN(P1_U3211) );
  XNOR2_X1 U8188 ( .A(n7047), .B(n7046), .ZN(n7053) );
  INV_X1 U8189 ( .A(n7406), .ZN(n7051) );
  OAI22_X1 U8190 ( .A1(n10399), .A2(n5131), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7048), .ZN(n7050) );
  OAI22_X1 U8191 ( .A1(n7403), .A2(n10393), .B1(n10394), .B2(n7446), .ZN(n7049) );
  AOI211_X1 U8192 ( .C1(n7051), .C2(n8820), .A(n7050), .B(n7049), .ZN(n7052)
         );
  OAI21_X1 U8193 ( .B1(n7053), .B2(n10397), .A(n7052), .ZN(P2_U3223) );
  OAI21_X1 U8194 ( .B1(n10234), .B2(n7055), .A(n7054), .ZN(n7063) );
  NAND2_X1 U8195 ( .A1(n10259), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7057) );
  INV_X1 U8196 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7526) );
  NOR2_X1 U8197 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7526), .ZN(n7694) );
  INV_X1 U8198 ( .A(n7694), .ZN(n7056) );
  OAI211_X1 U8199 ( .C1(n10318), .C2(n7058), .A(n7057), .B(n7056), .ZN(n7062)
         );
  AOI211_X1 U8200 ( .C1(n10227), .C2(n7060), .A(n7059), .B(n10321), .ZN(n7061)
         );
  AOI211_X1 U8201 ( .C1(n7063), .C2(n10329), .A(n7062), .B(n7061), .ZN(n7064)
         );
  INV_X1 U8202 ( .A(n7064), .ZN(P1_U3253) );
  INV_X1 U8203 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7090) );
  NAND2_X1 U8204 ( .A1(n7216), .A2(n7206), .ZN(n8487) );
  INV_X1 U8205 ( .A(n8487), .ZN(n7065) );
  AND2_X1 U8206 ( .A1(n7215), .A2(n7205), .ZN(n8486) );
  NOR2_X1 U8207 ( .A1(n7065), .A2(n8486), .ZN(n8606) );
  NAND2_X1 U8208 ( .A1(n7067), .A2(n7066), .ZN(n7069) );
  NAND2_X1 U8209 ( .A1(n10392), .A2(n10378), .ZN(n7068) );
  NAND2_X1 U8210 ( .A1(n7069), .A2(n7068), .ZN(n7355) );
  NAND2_X1 U8211 ( .A1(n7071), .A2(n7366), .ZN(n7084) );
  NAND2_X1 U8212 ( .A1(n7355), .A2(n7356), .ZN(n7073) );
  NAND2_X1 U8213 ( .A1(n7071), .A2(n10405), .ZN(n7072) );
  NAND2_X1 U8214 ( .A1(n7073), .A2(n7072), .ZN(n7226) );
  NAND2_X1 U8215 ( .A1(n8472), .A2(n8471), .ZN(n8475) );
  NAND2_X1 U8216 ( .A1(n7226), .A2(n8475), .ZN(n7076) );
  NAND2_X1 U8217 ( .A1(n10440), .A2(n10420), .ZN(n7075) );
  NAND2_X1 U8218 ( .A1(n7076), .A2(n7075), .ZN(n10435) );
  NAND2_X1 U8219 ( .A1(n10435), .A2(n10438), .ZN(n7078) );
  NAND2_X1 U8220 ( .A1(n8477), .A2(n10451), .ZN(n7077) );
  NAND2_X1 U8221 ( .A1(n7078), .A2(n7077), .ZN(n7181) );
  INV_X1 U8222 ( .A(n7181), .ZN(n7079) );
  NAND2_X1 U8223 ( .A1(n7086), .A2(n7185), .ZN(n7080) );
  XOR2_X1 U8224 ( .A(n8606), .B(n7204), .Z(n7165) );
  NAND2_X1 U8225 ( .A1(n8599), .A2(n8464), .ZN(n7082) );
  NAND2_X1 U8226 ( .A1(n7357), .A2(n7084), .ZN(n7227) );
  NAND2_X1 U8227 ( .A1(n7227), .A2(n8602), .ZN(n7228) );
  NAND2_X1 U8228 ( .A1(n7228), .A2(n8472), .ZN(n10436) );
  NAND2_X1 U8229 ( .A1(n8860), .A2(n10451), .ZN(n7085) );
  AND2_X1 U8230 ( .A1(n7086), .A2(n10501), .ZN(n7175) );
  NAND2_X1 U8231 ( .A1(n10442), .A2(n7185), .ZN(n8482) );
  XNOR2_X1 U8232 ( .A(n7209), .B(n8606), .ZN(n7087) );
  AOI222_X1 U8233 ( .A1(n9085), .A2(n7087), .B1(n7412), .B2(n9082), .C1(n7086), 
        .C2(n9080), .ZN(n7158) );
  NAND2_X1 U8234 ( .A1(n7361), .A2(n10405), .ZN(n7363) );
  OR2_X1 U8235 ( .A1(n7363), .A2(n7237), .ZN(n10446) );
  INV_X1 U8236 ( .A(n10451), .ZN(n10465) );
  XNOR2_X1 U8237 ( .A(n7217), .B(n7205), .ZN(n7159) );
  AOI22_X1 U8238 ( .A1(n7159), .A2(n10449), .B1(n10150), .B2(n7205), .ZN(n7088) );
  OAI211_X1 U8239 ( .C1(n10620), .C2(n7165), .A(n7158), .B(n7088), .ZN(n7091)
         );
  NAND2_X1 U8240 ( .A1(n7091), .A2(n10650), .ZN(n7089) );
  OAI21_X1 U8241 ( .B1(n10650), .B2(n7090), .A(n7089), .ZN(P2_U3469) );
  NAND2_X1 U8242 ( .A1(n7091), .A2(n10646), .ZN(n7092) );
  OAI21_X1 U8243 ( .B1(n10646), .B2(n6377), .A(n7092), .ZN(P2_U3526) );
  INV_X1 U8244 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7094) );
  INV_X1 U8245 ( .A(n8275), .ZN(n7095) );
  OAI222_X1 U8246 ( .A1(n8775), .A2(n7094), .B1(n8777), .B2(n7095), .C1(
        P1_U3084), .C2(n7093), .ZN(P1_U3335) );
  INV_X1 U8247 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7096) );
  INV_X1 U8248 ( .A(n8886), .ZN(n8872) );
  OAI222_X1 U8249 ( .A1(n8781), .A2(n7096), .B1(n7619), .B2(n7095), .C1(
        P2_U3152), .C2(n8872), .ZN(P2_U3340) );
  AND2_X1 U8250 ( .A1(n10355), .A2(n7097), .ZN(n10347) );
  NAND2_X1 U8251 ( .A1(n9765), .A2(n6708), .ZN(n7098) );
  NAND2_X1 U8252 ( .A1(n7118), .A2(n6697), .ZN(n9509) );
  NAND2_X1 U8253 ( .A1(n7118), .A2(n10385), .ZN(n7099) );
  XNOR2_X1 U8254 ( .A(n6779), .B(n10413), .ZN(n9356) );
  INV_X1 U8255 ( .A(n9356), .ZN(n7133) );
  XNOR2_X1 U8256 ( .A(n7124), .B(n7133), .ZN(n10412) );
  INV_X1 U8257 ( .A(n7100), .ZN(n7103) );
  NOR2_X1 U8258 ( .A1(n7639), .A2(n7101), .ZN(n7102) );
  NAND2_X1 U8259 ( .A1(n7103), .A2(n7102), .ZN(n7263) );
  NOR2_X1 U8260 ( .A1(n7110), .A2(n9697), .ZN(n10370) );
  NAND2_X1 U8261 ( .A1(n10539), .A2(n10370), .ZN(n9757) );
  NAND2_X1 U8262 ( .A1(n10539), .A2(n10364), .ZN(n10538) );
  INV_X1 U8263 ( .A(n10538), .ZN(n9702) );
  OAI22_X1 U8264 ( .A1(n10539), .A2(n6329), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10488), .ZN(n7109) );
  AND2_X1 U8265 ( .A1(n7261), .A2(n7105), .ZN(n7106) );
  INV_X1 U8266 ( .A(n10534), .ZN(n10333) );
  NAND2_X1 U8267 ( .A1(n10351), .A2(n10350), .ZN(n10349) );
  AND2_X1 U8268 ( .A1(n9771), .A2(n7104), .ZN(n7107) );
  OR2_X1 U8269 ( .A1(n7107), .A2(n7129), .ZN(n10414) );
  NOR2_X1 U8270 ( .A1(n10333), .A2(n10414), .ZN(n7108) );
  AOI211_X1 U8271 ( .C1(n9702), .C2(n7104), .A(n7109), .B(n7108), .ZN(n7123)
         );
  AOI21_X1 U8272 ( .B1(n9502), .B2(n7110), .A(n10493), .ZN(n7111) );
  NAND2_X1 U8273 ( .A1(n7112), .A2(n7111), .ZN(n10526) );
  NAND2_X1 U8274 ( .A1(n7113), .A2(n6708), .ZN(n7114) );
  NAND2_X1 U8275 ( .A1(n7115), .A2(n9509), .ZN(n7134) );
  XNOR2_X1 U8276 ( .A(n7134), .B(n7133), .ZN(n7120) );
  NAND2_X1 U8277 ( .A1(n6698), .A2(n10493), .ZN(n7117) );
  NAND2_X1 U8278 ( .A1(n6234), .A2(n9538), .ZN(n7116) );
  NAND2_X1 U8279 ( .A1(n7117), .A2(n7116), .ZN(n10473) );
  INV_X1 U8280 ( .A(n10516), .ZN(n9743) );
  OAI22_X1 U8281 ( .A1(n9743), .A2(n7118), .B1(n7240), .B2(n9745), .ZN(n7119)
         );
  AOI21_X1 U8282 ( .B1(n7120), .B2(n10473), .A(n7119), .ZN(n7121) );
  OAI21_X1 U8283 ( .B1(n10412), .B2(n10526), .A(n7121), .ZN(n10415) );
  NAND2_X1 U8284 ( .A1(n10415), .A2(n10539), .ZN(n7122) );
  OAI211_X1 U8285 ( .C1(n10412), .C2(n9757), .A(n7123), .B(n7122), .ZN(
        P1_U3288) );
  NAND2_X1 U8286 ( .A1(n6788), .A2(n10413), .ZN(n7241) );
  NAND2_X1 U8287 ( .A1(n7243), .A2(n7241), .ZN(n7126) );
  NAND2_X1 U8288 ( .A1(n7240), .A2(n7125), .ZN(n9516) );
  NAND2_X1 U8289 ( .A1(n10475), .A2(n4835), .ZN(n9514) );
  NAND2_X1 U8290 ( .A1(n9516), .A2(n9514), .ZN(n7245) );
  INV_X1 U8291 ( .A(n7245), .ZN(n9355) );
  XNOR2_X1 U8292 ( .A(n7126), .B(n9355), .ZN(n10427) );
  INV_X1 U8293 ( .A(n7127), .ZN(n7128) );
  OAI22_X1 U8294 ( .A1(n10539), .A2(n6330), .B1(n7128), .B2(n10488), .ZN(n7132) );
  OR2_X1 U8295 ( .A1(n7129), .A2(n4835), .ZN(n7130) );
  NAND2_X1 U8296 ( .A1(n10476), .A2(n7130), .ZN(n10428) );
  NOR2_X1 U8297 ( .A1(n10333), .A2(n10428), .ZN(n7131) );
  AOI211_X1 U8298 ( .C1(n9702), .C2(n7125), .A(n7132), .B(n7131), .ZN(n7140)
         );
  NAND2_X1 U8299 ( .A1(n7134), .A2(n7133), .ZN(n7135) );
  NAND2_X1 U8300 ( .A1(n6788), .A2(n7104), .ZN(n9512) );
  NAND2_X1 U8301 ( .A1(n7135), .A2(n9512), .ZN(n7251) );
  XNOR2_X1 U8302 ( .A(n7251), .B(n9355), .ZN(n7137) );
  OAI22_X1 U8303 ( .A1(n9743), .A2(n6788), .B1(n7247), .B2(n9745), .ZN(n7136)
         );
  AOI21_X1 U8304 ( .B1(n7137), .B2(n10473), .A(n7136), .ZN(n7138) );
  OAI21_X1 U8305 ( .B1(n10427), .B2(n10526), .A(n7138), .ZN(n10429) );
  NAND2_X1 U8306 ( .A1(n10429), .A2(n10539), .ZN(n7139) );
  OAI211_X1 U8307 ( .C1(n10427), .C2(n9757), .A(n7140), .B(n7139), .ZN(
        P1_U3287) );
  INV_X1 U8308 ( .A(n8279), .ZN(n7142) );
  OAI222_X1 U8309 ( .A1(n8781), .A2(n7141), .B1(n7619), .B2(n7142), .C1(
        P2_U3152), .C2(n8890), .ZN(P2_U3339) );
  OAI222_X1 U8310 ( .A1(n9697), .A2(P1_U3084), .B1(n8777), .B2(n7142), .C1(
        n8775), .C2(n5554), .ZN(P1_U3334) );
  NAND2_X1 U8311 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8861), .ZN(n7143) );
  OAI21_X1 U8312 ( .B1(n8958), .B2(n8861), .A(n7143), .ZN(P2_U3580) );
  NAND2_X1 U8313 ( .A1(n8862), .A2(n7144), .ZN(n8597) );
  NAND2_X1 U8314 ( .A1(n8599), .A2(n8597), .ZN(n10341) );
  INV_X1 U8315 ( .A(n10341), .ZN(n7157) );
  NAND2_X1 U8316 ( .A1(n7154), .A2(n7145), .ZN(n7146) );
  AND2_X2 U8317 ( .A1(n7146), .A2(n10373), .ZN(n10469) );
  NAND2_X1 U8318 ( .A1(n7147), .A2(n8636), .ZN(n7234) );
  NAND2_X1 U8319 ( .A1(n7450), .A2(n7234), .ZN(n7148) );
  AOI22_X1 U8320 ( .A1(n10341), .A2(n9085), .B1(n9082), .B2(n6760), .ZN(n10343) );
  OAI21_X1 U8321 ( .B1(n10283), .B2(n10373), .A(n10343), .ZN(n7150) );
  NOR2_X1 U8322 ( .A1(n4833), .A2(n5621), .ZN(n7149) );
  AOI21_X1 U8323 ( .B1(n4833), .B2(n7150), .A(n7149), .ZN(n7156) );
  INV_X1 U8324 ( .A(n10377), .ZN(n7151) );
  NAND2_X1 U8325 ( .A1(n4833), .A2(n7151), .ZN(n9076) );
  NOR2_X1 U8326 ( .A1(n7152), .A2(n8434), .ZN(n7153) );
  OAI21_X1 U8327 ( .B1(n10466), .B2(n10461), .A(n10339), .ZN(n7155) );
  OAI211_X1 U8328 ( .C1(n7157), .C2(n9089), .A(n7156), .B(n7155), .ZN(P2_U3296) );
  MUX2_X1 U8329 ( .A(n6364), .B(n7158), .S(n4833), .Z(n7164) );
  INV_X1 U8330 ( .A(n10461), .ZN(n9008) );
  INV_X1 U8331 ( .A(n7159), .ZN(n7161) );
  OAI22_X1 U8332 ( .A1(n9008), .A2(n7161), .B1(n7160), .B2(n10373), .ZN(n7162)
         );
  AOI21_X1 U8333 ( .B1(n10466), .B2(n7205), .A(n7162), .ZN(n7163) );
  OAI211_X1 U8334 ( .C1(n9089), .C2(n7165), .A(n7164), .B(n7163), .ZN(P2_U3290) );
  OAI21_X1 U8335 ( .B1(n7168), .B2(n7167), .A(n7166), .ZN(n7173) );
  OAI22_X1 U8336 ( .A1(n7397), .A2(n10393), .B1(n10394), .B2(n7442), .ZN(n7172) );
  NAND2_X1 U8337 ( .A1(n8851), .A2(n10596), .ZN(n7170) );
  OAI211_X1 U8338 ( .C1(n8848), .C2(n7431), .A(n7170), .B(n7169), .ZN(n7171)
         );
  AOI211_X1 U8339 ( .C1(n7173), .C2(n8844), .A(n7172), .B(n7171), .ZN(n7174)
         );
  INV_X1 U8340 ( .A(n7174), .ZN(P2_U3233) );
  INV_X1 U8341 ( .A(n7175), .ZN(n8483) );
  AND2_X1 U8342 ( .A1(n8483), .A2(n8482), .ZN(n8601) );
  INV_X1 U8343 ( .A(n8601), .ZN(n7176) );
  XNOR2_X1 U8344 ( .A(n7177), .B(n7176), .ZN(n7178) );
  NAND2_X1 U8345 ( .A1(n7178), .A2(n9085), .ZN(n7180) );
  AOI22_X1 U8346 ( .A1(n9080), .A2(n8860), .B1(n7206), .B2(n9082), .ZN(n7179)
         );
  AND2_X1 U8347 ( .A1(n7180), .A2(n7179), .ZN(n10502) );
  INV_X1 U8348 ( .A(n9089), .ZN(n10457) );
  XOR2_X1 U8349 ( .A(n7181), .B(n8601), .Z(n10505) );
  AND2_X1 U8350 ( .A1(n4833), .A2(n8890), .ZN(n8985) );
  INV_X1 U8351 ( .A(n10448), .ZN(n7182) );
  INV_X1 U8352 ( .A(n10449), .ZN(n10639) );
  AOI211_X1 U8353 ( .C1(n7185), .C2(n7182), .A(n10639), .B(n7217), .ZN(n10499)
         );
  AOI22_X1 U8354 ( .A1(n10457), .A2(n10505), .B1(n8985), .B2(n10499), .ZN(
        n7187) );
  OAI22_X1 U8355 ( .A1(n4833), .A2(n6363), .B1(n7183), .B2(n10373), .ZN(n7184)
         );
  AOI21_X1 U8356 ( .B1(n10466), .B2(n7185), .A(n7184), .ZN(n7186) );
  OAI211_X1 U8357 ( .C1(n10469), .C2(n10502), .A(n7187), .B(n7186), .ZN(
        P2_U3291) );
  NOR2_X1 U8358 ( .A1(n7546), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7188) );
  AOI21_X1 U8359 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7546), .A(n7188), .ZN(
        n7191) );
  OAI21_X1 U8360 ( .B1(n7191), .B2(n7190), .A(n7539), .ZN(n7192) );
  NAND2_X1 U8361 ( .A1(n7192), .A2(n8896), .ZN(n7202) );
  INV_X1 U8362 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7193) );
  NOR2_X1 U8363 ( .A1(n8893), .A2(n7193), .ZN(n7200) );
  AOI21_X1 U8364 ( .B1(n7195), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7194), .ZN(
        n7198) );
  INV_X1 U8365 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7196) );
  MUX2_X1 U8366 ( .A(n7196), .B(P2_REG1_REG_11__SCAN_IN), .S(n7546), .Z(n7197)
         );
  NOR2_X1 U8367 ( .A1(n7198), .A2(n7197), .ZN(n7545) );
  AOI211_X1 U8368 ( .C1(n7198), .C2(n7197), .A(n7545), .B(n10297), .ZN(n7199)
         );
  AOI211_X1 U8369 ( .C1(P2_REG3_REG_11__SCAN_IN), .C2(P2_U3152), .A(n7200), 
        .B(n7199), .ZN(n7201) );
  OAI211_X1 U8370 ( .C1(n8891), .C2(n7203), .A(n7202), .B(n7201), .ZN(P2_U3256) );
  NAND2_X1 U8371 ( .A1(n7215), .A2(n7216), .ZN(n7207) );
  NAND2_X1 U8372 ( .A1(n7208), .A2(n7207), .ZN(n7410) );
  OR2_X1 U8373 ( .A1(n7403), .A2(n7411), .ZN(n8492) );
  NAND2_X1 U8374 ( .A1(n7411), .A2(n7403), .ZN(n8491) );
  NAND2_X1 U8375 ( .A1(n8492), .A2(n8491), .ZN(n7409) );
  XNOR2_X1 U8376 ( .A(n7410), .B(n7409), .ZN(n10562) );
  INV_X1 U8377 ( .A(n10562), .ZN(n7225) );
  INV_X1 U8378 ( .A(n7211), .ZN(n7213) );
  INV_X1 U8379 ( .A(n7409), .ZN(n8605) );
  NAND2_X1 U8380 ( .A1(n7211), .A2(n8605), .ZN(n7399) );
  INV_X1 U8381 ( .A(n7399), .ZN(n7212) );
  AOI21_X1 U8382 ( .B1(n7409), .B2(n7213), .A(n7212), .ZN(n7214) );
  OAI222_X1 U8383 ( .A1(n10441), .A2(n7397), .B1(n10439), .B2(n7215), .C1(
        n10437), .C2(n7214), .ZN(n10560) );
  NAND2_X1 U8384 ( .A1(n10560), .A2(n4833), .ZN(n7224) );
  NOR2_X1 U8385 ( .A1(n4833), .A2(n6414), .ZN(n7222) );
  NAND2_X1 U8386 ( .A1(n7217), .A2(n7216), .ZN(n7218) );
  INV_X1 U8387 ( .A(n7218), .ZN(n7219) );
  OAI21_X1 U8388 ( .B1(n7219), .B2(n10558), .A(n7404), .ZN(n10559) );
  OAI22_X1 U8389 ( .A1(n9008), .A2(n10559), .B1(n7220), .B2(n10373), .ZN(n7221) );
  AOI211_X1 U8390 ( .C1(n10466), .C2(n7411), .A(n7222), .B(n7221), .ZN(n7223)
         );
  OAI211_X1 U8391 ( .C1(n7225), .C2(n9089), .A(n7224), .B(n7223), .ZN(P2_U3289) );
  XNOR2_X1 U8392 ( .A(n7226), .B(n8602), .ZN(n7236) );
  OAI21_X1 U8393 ( .B1(n8602), .B2(n7227), .A(n7228), .ZN(n7230) );
  OAI22_X1 U8394 ( .A1(n8477), .A2(n10441), .B1(n7071), .B2(n10439), .ZN(n7229) );
  AOI21_X1 U8395 ( .B1(n7230), .B2(n9085), .A(n7229), .ZN(n7231) );
  OAI21_X1 U8396 ( .B1(n7236), .B2(n7450), .A(n7231), .ZN(n10422) );
  NAND2_X1 U8397 ( .A1(n7363), .A2(n7237), .ZN(n7232) );
  NAND2_X1 U8398 ( .A1(n10446), .A2(n7232), .ZN(n10421) );
  OAI22_X1 U8399 ( .A1(n9008), .A2(n10421), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10373), .ZN(n7233) );
  AOI21_X1 U8400 ( .B1(n4833), .B2(n10422), .A(n7233), .ZN(n7239) );
  INV_X1 U8401 ( .A(n7234), .ZN(n7235) );
  NAND2_X1 U8402 ( .A1(n4833), .A2(n7235), .ZN(n7459) );
  INV_X1 U8403 ( .A(n7459), .ZN(n7367) );
  INV_X1 U8404 ( .A(n7236), .ZN(n10424) );
  AOI22_X1 U8405 ( .A1(n7367), .A2(n10424), .B1(n10466), .B2(n7237), .ZN(n7238) );
  OAI211_X1 U8406 ( .C1(n6362), .C2(n4833), .A(n7239), .B(n7238), .ZN(P2_U3293) );
  NAND2_X1 U8407 ( .A1(n7240), .A2(n4835), .ZN(n7244) );
  AND2_X1 U8408 ( .A1(n7241), .A2(n7244), .ZN(n7242) );
  INV_X1 U8409 ( .A(n7244), .ZN(n7246) );
  NAND2_X1 U8410 ( .A1(n7247), .A2(n7259), .ZN(n9517) );
  OR2_X1 U8411 ( .A1(n7249), .A2(n7260), .ZN(n10517) );
  NAND2_X1 U8412 ( .A1(n7260), .A2(n7249), .ZN(n9522) );
  NAND2_X1 U8413 ( .A1(n10517), .A2(n9522), .ZN(n10519) );
  NAND2_X1 U8414 ( .A1(n10509), .A2(n10519), .ZN(n10508) );
  INV_X1 U8415 ( .A(n7260), .ZN(n10537) );
  NAND2_X1 U8416 ( .A1(n10537), .A2(n7249), .ZN(n7250) );
  NAND2_X1 U8417 ( .A1(n10508), .A2(n7250), .ZN(n7335) );
  OR2_X1 U8418 ( .A1(n10548), .A2(n7342), .ZN(n9397) );
  NAND2_X1 U8419 ( .A1(n10548), .A2(n7342), .ZN(n9395) );
  NAND2_X1 U8420 ( .A1(n9397), .A2(n9395), .ZN(n7334) );
  XNOR2_X1 U8421 ( .A(n7335), .B(n7334), .ZN(n7258) );
  INV_X1 U8422 ( .A(n7258), .ZN(n10553) );
  INV_X1 U8423 ( .A(n10526), .ZN(n9764) );
  NAND2_X1 U8424 ( .A1(n7251), .A2(n9355), .ZN(n7252) );
  NAND2_X1 U8425 ( .A1(n7252), .A2(n9516), .ZN(n9391) );
  INV_X1 U8426 ( .A(n9522), .ZN(n7253) );
  NAND2_X1 U8427 ( .A1(n10523), .A2(n10517), .ZN(n7254) );
  INV_X1 U8428 ( .A(n7334), .ZN(n9358) );
  XNOR2_X1 U8429 ( .A(n7254), .B(n9358), .ZN(n7256) );
  INV_X1 U8430 ( .A(n10473), .ZN(n10518) );
  AOI22_X1 U8431 ( .A1(n10516), .A2(n10474), .B1(n10514), .B2(n9556), .ZN(
        n7255) );
  OAI21_X1 U8432 ( .B1(n7256), .B2(n10518), .A(n7255), .ZN(n7257) );
  AOI21_X1 U8433 ( .B1(n7258), .B2(n9764), .A(n7257), .ZN(n10551) );
  MUX2_X1 U8434 ( .A(n6335), .B(n10551), .S(n10539), .Z(n7269) );
  NOR2_X1 U8435 ( .A1(n10510), .A2(n7260), .ZN(n7262) );
  INV_X1 U8436 ( .A(n7262), .ZN(n10511) );
  AND2_X1 U8437 ( .A1(n7261), .A2(n7388), .ZN(n10477) );
  AOI211_X1 U8438 ( .C1(n10548), .C2(n10511), .A(n10565), .B(n7347), .ZN(
        n10547) );
  NOR2_X1 U8439 ( .A1(n7263), .A2(n10493), .ZN(n8076) );
  INV_X1 U8440 ( .A(n7264), .ZN(n7265) );
  OAI22_X1 U8441 ( .A1(n10538), .A2(n7266), .B1(n10488), .B2(n7265), .ZN(n7267) );
  AOI21_X1 U8442 ( .B1(n10547), .B2(n8076), .A(n7267), .ZN(n7268) );
  OAI211_X1 U8443 ( .C1(n10553), .C2(n9757), .A(n7269), .B(n7268), .ZN(
        P1_U3284) );
  NAND2_X1 U8444 ( .A1(n7270), .A2(n6944), .ZN(n7273) );
  AOI22_X1 U8445 ( .A1(n8280), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6704), .B2(
        n7271), .ZN(n7272) );
  NAND2_X1 U8446 ( .A1(n7273), .A2(n7272), .ZN(n7486) );
  INV_X1 U8447 ( .A(n7486), .ZN(n10583) );
  INV_X1 U8448 ( .A(n7274), .ZN(n7276) );
  NAND2_X1 U8449 ( .A1(n7276), .A2(n7275), .ZN(n7300) );
  NAND2_X1 U8450 ( .A1(n7277), .A2(n6944), .ZN(n7280) );
  AOI22_X1 U8451 ( .A1(n8280), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6704), .B2(
        n7278), .ZN(n7279) );
  NAND2_X1 U8452 ( .A1(n7280), .A2(n7279), .ZN(n7464) );
  NOR2_X1 U8453 ( .A1(n8760), .A2(n7337), .ZN(n7281) );
  AOI21_X1 U8454 ( .B1(n7464), .B2(n8752), .A(n7281), .ZN(n7302) );
  INV_X1 U8455 ( .A(n7302), .ZN(n7282) );
  AND2_X1 U8456 ( .A1(n7300), .A2(n7282), .ZN(n7283) );
  NAND2_X1 U8457 ( .A1(n7301), .A2(n7283), .ZN(n7308) );
  NAND2_X1 U8458 ( .A1(n7486), .A2(n4856), .ZN(n7292) );
  NAND2_X1 U8459 ( .A1(n6800), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7290) );
  NAND2_X1 U8460 ( .A1(n7285), .A2(n7284), .ZN(n7286) );
  AND2_X1 U8461 ( .A1(n7313), .A2(n7286), .ZN(n7474) );
  NAND2_X1 U8462 ( .A1(n6823), .A2(n7474), .ZN(n7289) );
  NAND2_X1 U8463 ( .A1(n4874), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7288) );
  NAND2_X1 U8464 ( .A1(n6801), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7287) );
  NAND4_X1 U8465 ( .A1(n7290), .A2(n7289), .A3(n7288), .A4(n7287), .ZN(n9555)
         );
  NAND2_X1 U8466 ( .A1(n8752), .A2(n9555), .ZN(n7291) );
  NAND2_X1 U8467 ( .A1(n7292), .A2(n7291), .ZN(n7293) );
  XNOR2_X1 U8468 ( .A(n7293), .B(n4854), .ZN(n7295) );
  INV_X1 U8469 ( .A(n9555), .ZN(n7515) );
  NOR2_X1 U8470 ( .A1(n8760), .A2(n7515), .ZN(n7294) );
  AOI21_X1 U8471 ( .B1(n7486), .B2(n8752), .A(n7294), .ZN(n7296) );
  NAND2_X1 U8472 ( .A1(n7295), .A2(n7296), .ZN(n7506) );
  INV_X1 U8473 ( .A(n7295), .ZN(n7298) );
  INV_X1 U8474 ( .A(n7296), .ZN(n7297) );
  NAND2_X1 U8475 ( .A1(n7298), .A2(n7297), .ZN(n7299) );
  AND2_X1 U8476 ( .A1(n7506), .A2(n7299), .ZN(n7309) );
  AND2_X1 U8477 ( .A1(n7308), .A2(n7309), .ZN(n7306) );
  NAND2_X1 U8478 ( .A1(n7464), .A2(n4855), .ZN(n7304) );
  NAND2_X1 U8479 ( .A1(n9556), .A2(n8752), .ZN(n7303) );
  NAND2_X1 U8480 ( .A1(n7304), .A2(n7303), .ZN(n7305) );
  XNOR2_X1 U8481 ( .A(n7305), .B(n8761), .ZN(n7324) );
  INV_X1 U8482 ( .A(n7507), .ZN(n7311) );
  AOI21_X1 U8483 ( .B1(n7307), .B2(n7308), .A(n7309), .ZN(n7310) );
  OAI21_X1 U8484 ( .B1(n7311), .B2(n7310), .A(n4834), .ZN(n7323) );
  NAND2_X1 U8485 ( .A1(n4874), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7318) );
  NAND2_X1 U8486 ( .A1(n6800), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7317) );
  NAND2_X1 U8487 ( .A1(n7313), .A2(n7312), .ZN(n7314) );
  AND2_X1 U8488 ( .A1(n7491), .A2(n7314), .ZN(n7511) );
  NAND2_X1 U8489 ( .A1(n6823), .A2(n7511), .ZN(n7316) );
  NAND2_X1 U8490 ( .A1(n6801), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7315) );
  AOI21_X1 U8491 ( .B1(n9262), .B2(n9554), .A(n7319), .ZN(n7320) );
  OAI21_X1 U8492 ( .B1(n7337), .B2(n9284), .A(n7320), .ZN(n7321) );
  AOI21_X1 U8493 ( .B1(n9280), .B2(n7474), .A(n7321), .ZN(n7322) );
  OAI211_X1 U8494 ( .C1(n10583), .C2(n9224), .A(n7323), .B(n7322), .ZN(
        P1_U3229) );
  INV_X1 U8495 ( .A(n7464), .ZN(n10564) );
  INV_X1 U8496 ( .A(n7308), .ZN(n7328) );
  AOI21_X1 U8497 ( .B1(n7325), .B2(n7308), .A(n7324), .ZN(n7326) );
  NOR2_X1 U8498 ( .A1(n7326), .A2(n9289), .ZN(n7327) );
  OAI21_X1 U8499 ( .B1(n7328), .B2(n7307), .A(n7327), .ZN(n7333) );
  AOI21_X1 U8500 ( .B1(n9262), .B2(n9555), .A(n7329), .ZN(n7330) );
  OAI21_X1 U8501 ( .B1(n7342), .B2(n9284), .A(n7330), .ZN(n7331) );
  AOI21_X1 U8502 ( .B1(n9280), .B2(n7349), .A(n7331), .ZN(n7332) );
  OAI211_X1 U8503 ( .C1(n10564), .C2(n9224), .A(n7333), .B(n7332), .ZN(
        P1_U3219) );
  OR2_X1 U8504 ( .A1(n10548), .A2(n10513), .ZN(n7336) );
  OR2_X1 U8505 ( .A1(n7464), .A2(n7337), .ZN(n9402) );
  NAND2_X1 U8506 ( .A1(n7464), .A2(n7337), .ZN(n9403) );
  NAND2_X1 U8507 ( .A1(n7339), .A2(n9401), .ZN(n7340) );
  NAND2_X1 U8508 ( .A1(n7466), .A2(n7340), .ZN(n7346) );
  AND2_X1 U8509 ( .A1(n9397), .A2(n10517), .ZN(n9521) );
  NAND2_X1 U8510 ( .A1(n9328), .A2(n9395), .ZN(n7341) );
  XNOR2_X1 U8511 ( .A(n7341), .B(n9401), .ZN(n7344) );
  OAI22_X1 U8512 ( .A1(n9743), .A2(n7342), .B1(n7515), .B2(n9745), .ZN(n7343)
         );
  AOI21_X1 U8513 ( .B1(n7344), .B2(n10473), .A(n7343), .ZN(n7345) );
  OAI21_X1 U8514 ( .B1(n7346), .B2(n10526), .A(n7345), .ZN(n10567) );
  INV_X1 U8515 ( .A(n10567), .ZN(n7354) );
  INV_X1 U8516 ( .A(n7346), .ZN(n10569) );
  INV_X1 U8517 ( .A(n9757), .ZN(n10535) );
  OR2_X1 U8518 ( .A1(n7347), .A2(n10564), .ZN(n7348) );
  NAND2_X1 U8519 ( .A1(n7467), .A2(n7348), .ZN(n10566) );
  INV_X1 U8520 ( .A(n10488), .ZN(n10544) );
  AOI22_X1 U8521 ( .A1(n10498), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7349), .B2(
        n10544), .ZN(n7351) );
  NAND2_X1 U8522 ( .A1(n9702), .A2(n7464), .ZN(n7350) );
  OAI211_X1 U8523 ( .C1(n10566), .C2(n10333), .A(n7351), .B(n7350), .ZN(n7352)
         );
  AOI21_X1 U8524 ( .B1(n10569), .B2(n10535), .A(n7352), .ZN(n7353) );
  OAI21_X1 U8525 ( .B1(n7354), .B2(n10498), .A(n7353), .ZN(P1_U3283) );
  XOR2_X1 U8526 ( .A(n7355), .B(n7356), .Z(n7365) );
  OAI21_X1 U8527 ( .B1(n5475), .B2(n7083), .A(n7357), .ZN(n7359) );
  OAI22_X1 U8528 ( .A1(n10440), .A2(n10441), .B1(n10392), .B2(n10439), .ZN(
        n7358) );
  AOI21_X1 U8529 ( .B1(n7359), .B2(n9085), .A(n7358), .ZN(n7360) );
  OAI21_X1 U8530 ( .B1(n7365), .B2(n7450), .A(n7360), .ZN(n10407) );
  OR2_X1 U8531 ( .A1(n7361), .A2(n10405), .ZN(n7362) );
  NAND2_X1 U8532 ( .A1(n7363), .A2(n7362), .ZN(n10406) );
  OAI22_X1 U8533 ( .A1(n9008), .A2(n10406), .B1(n10403), .B2(n10373), .ZN(
        n7364) );
  AOI21_X1 U8534 ( .B1(n4833), .B2(n10407), .A(n7364), .ZN(n7369) );
  INV_X1 U8535 ( .A(n7365), .ZN(n10409) );
  AOI22_X1 U8536 ( .A1(n7367), .A2(n10409), .B1(n10466), .B2(n7366), .ZN(n7368) );
  OAI211_X1 U8537 ( .C1(n6361), .C2(n4833), .A(n7369), .B(n7368), .ZN(P2_U3294) );
  XNOR2_X1 U8538 ( .A(n7371), .B(n7370), .ZN(n7376) );
  INV_X1 U8539 ( .A(n7451), .ZN(n7374) );
  INV_X1 U8540 ( .A(n7575), .ZN(n10604) );
  OAI22_X1 U8541 ( .A1(n10399), .A2(n10604), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10105), .ZN(n7373) );
  OAI22_X1 U8542 ( .A1(n7446), .A2(n10393), .B1(n10394), .B2(n7627), .ZN(n7372) );
  AOI211_X1 U8543 ( .C1(n7374), .C2(n8820), .A(n7373), .B(n7372), .ZN(n7375)
         );
  OAI21_X1 U8544 ( .B1(n7376), .B2(n10397), .A(n7375), .ZN(P2_U3219) );
  NAND2_X1 U8545 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7720) );
  INV_X1 U8546 ( .A(n7720), .ZN(n7381) );
  AOI211_X1 U8547 ( .C1(n7379), .C2(n7378), .A(n7377), .B(n10321), .ZN(n7380)
         );
  AOI211_X1 U8548 ( .C1(n10257), .C2(n7708), .A(n7381), .B(n7380), .ZN(n7387)
         );
  OAI21_X1 U8549 ( .B1(n7384), .B2(n7383), .A(n7382), .ZN(n7385) );
  AOI22_X1 U8550 ( .A1(n10259), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(n10329), 
        .B2(n7385), .ZN(n7386) );
  NAND2_X1 U8551 ( .A1(n7387), .A2(n7386), .ZN(P1_U3254) );
  INV_X1 U8552 ( .A(n8292), .ZN(n7395) );
  OAI222_X1 U8553 ( .A1(n8777), .A2(n7395), .B1(n7388), .B2(P1_U3084), .C1(
        n8293), .C2(n8775), .ZN(P1_U3333) );
  XNOR2_X1 U8554 ( .A(n7390), .B(n7389), .ZN(n7394) );
  OAI22_X1 U8555 ( .A1(n10394), .A2(n7776), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5785), .ZN(n7392) );
  OAI22_X1 U8556 ( .A1(n10393), .A2(n7442), .B1(n8848), .B2(n7579), .ZN(n7391)
         );
  AOI211_X1 U8557 ( .C1(n10612), .C2(n8851), .A(n7392), .B(n7391), .ZN(n7393)
         );
  OAI21_X1 U8558 ( .B1(n7394), .B2(n10397), .A(n7393), .ZN(P2_U3238) );
  OAI222_X1 U8559 ( .A1(n8781), .A2(n7396), .B1(n7619), .B2(n7395), .C1(n5610), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OR2_X1 U8560 ( .A1(n7419), .A2(n7397), .ZN(n8497) );
  NAND2_X1 U8561 ( .A1(n7419), .A2(n7397), .ZN(n8495) );
  INV_X1 U8562 ( .A(n8491), .ZN(n7398) );
  NOR2_X1 U8563 ( .A1(n8607), .A2(n7398), .ZN(n7401) );
  NAND2_X1 U8564 ( .A1(n7399), .A2(n8491), .ZN(n7400) );
  NAND2_X1 U8565 ( .A1(n7400), .A2(n8607), .ZN(n7427) );
  INV_X1 U8566 ( .A(n7427), .ZN(n7424) );
  AOI21_X1 U8567 ( .B1(n7401), .B2(n7399), .A(n7424), .ZN(n7402) );
  OAI222_X1 U8568 ( .A1(n10441), .A2(n7446), .B1(n10439), .B2(n7403), .C1(
        n10437), .C2(n7402), .ZN(n10578) );
  INV_X1 U8569 ( .A(n8985), .ZN(n7584) );
  AOI21_X1 U8570 ( .B1(n7404), .B2(n7419), .A(n10639), .ZN(n7405) );
  NAND2_X1 U8571 ( .A1(n7405), .A2(n7432), .ZN(n10575) );
  OAI22_X1 U8572 ( .A1(n4833), .A2(n7407), .B1(n7406), .B2(n10373), .ZN(n7408)
         );
  AOI21_X1 U8573 ( .B1(n10466), .B2(n7419), .A(n7408), .ZN(n7416) );
  OR2_X1 U8574 ( .A1(n7412), .A2(n7411), .ZN(n7413) );
  NAND2_X1 U8575 ( .A1(n7414), .A2(n8607), .ZN(n10573) );
  NAND3_X1 U8576 ( .A1(n10574), .A2(n10573), .A3(n10457), .ZN(n7415) );
  OAI211_X1 U8577 ( .C1(n7584), .C2(n10575), .A(n7416), .B(n7415), .ZN(n7417)
         );
  AOI21_X1 U8578 ( .B1(n10578), .B2(n4833), .A(n7417), .ZN(n7418) );
  INV_X1 U8579 ( .A(n7418), .ZN(P2_U3288) );
  NAND2_X1 U8580 ( .A1(n7419), .A2(n7423), .ZN(n7420) );
  AND2_X1 U8581 ( .A1(n10574), .A2(n7420), .ZN(n7422) );
  NAND2_X1 U8582 ( .A1(n10596), .A2(n7446), .ZN(n8500) );
  NAND2_X1 U8583 ( .A1(n8502), .A2(n8500), .ZN(n8609) );
  AND2_X1 U8584 ( .A1(n7420), .A2(n8609), .ZN(n7421) );
  NAND2_X1 U8585 ( .A1(n10574), .A2(n7421), .ZN(n7441) );
  OAI21_X1 U8586 ( .B1(n7422), .B2(n8609), .A(n7441), .ZN(n10601) );
  INV_X1 U8587 ( .A(n10601), .ZN(n7438) );
  AOI22_X1 U8588 ( .A1(n9080), .A2(n7423), .B1(n8859), .B2(n9082), .ZN(n7430)
         );
  INV_X1 U8589 ( .A(n8495), .ZN(n7425) );
  OAI21_X1 U8590 ( .B1(n7424), .B2(n7425), .A(n8609), .ZN(n7428) );
  NAND3_X1 U8591 ( .A1(n7428), .A2(n7445), .A3(n9085), .ZN(n7429) );
  OAI211_X1 U8592 ( .C1(n7438), .C2(n7450), .A(n7430), .B(n7429), .ZN(n10599)
         );
  NAND2_X1 U8593 ( .A1(n10599), .A2(n4833), .ZN(n7437) );
  OAI22_X1 U8594 ( .A1(n4833), .A2(n6454), .B1(n7431), .B2(n10373), .ZN(n7435)
         );
  AND2_X1 U8595 ( .A1(n7432), .A2(n10596), .ZN(n7433) );
  OR2_X1 U8596 ( .A1(n7433), .A2(n7454), .ZN(n10598) );
  NOR2_X1 U8597 ( .A1(n9008), .A2(n10598), .ZN(n7434) );
  AOI211_X1 U8598 ( .C1(n10466), .C2(n10596), .A(n7435), .B(n7434), .ZN(n7436)
         );
  OAI211_X1 U8599 ( .C1(n7438), .C2(n7459), .A(n7437), .B(n7436), .ZN(P2_U3287) );
  OR2_X1 U8600 ( .A1(n10596), .A2(n7439), .ZN(n7440) );
  NAND2_X1 U8601 ( .A1(n7441), .A2(n7440), .ZN(n7443) );
  OR2_X1 U8602 ( .A1(n7575), .A2(n7442), .ZN(n8507) );
  NAND2_X1 U8603 ( .A1(n7575), .A2(n7442), .ZN(n8505) );
  OR2_X2 U8604 ( .A1(n7443), .A2(n8613), .ZN(n7598) );
  NAND2_X1 U8605 ( .A1(n7443), .A2(n8613), .ZN(n7444) );
  NAND2_X1 U8606 ( .A1(n7598), .A2(n7444), .ZN(n10603) );
  OAI21_X1 U8607 ( .B1(n4934), .B2(n8613), .A(n7570), .ZN(n7448) );
  OAI22_X1 U8608 ( .A1(n7446), .A2(n10439), .B1(n7627), .B2(n10441), .ZN(n7447) );
  AOI21_X1 U8609 ( .B1(n7448), .B2(n9085), .A(n7447), .ZN(n7449) );
  OAI21_X1 U8610 ( .B1(n7450), .B2(n10603), .A(n7449), .ZN(n10606) );
  OAI22_X1 U8611 ( .A1(n4833), .A2(n7452), .B1(n7451), .B2(n10373), .ZN(n7453)
         );
  AOI21_X1 U8612 ( .B1(n10466), .B2(n7575), .A(n7453), .ZN(n7458) );
  OR2_X1 U8613 ( .A1(n7454), .A2(n10604), .ZN(n7455) );
  NAND2_X1 U8614 ( .A1(n7573), .A2(n7455), .ZN(n10605) );
  INV_X1 U8615 ( .A(n10605), .ZN(n7456) );
  NAND2_X1 U8616 ( .A1(n7456), .A2(n10461), .ZN(n7457) );
  OAI211_X1 U8617 ( .C1(n10603), .C2(n7459), .A(n7458), .B(n7457), .ZN(n7460)
         );
  AOI21_X1 U8618 ( .B1(n10606), .B2(n4833), .A(n7460), .ZN(n7461) );
  INV_X1 U8619 ( .A(n7461), .ZN(P2_U3286) );
  INV_X1 U8620 ( .A(n8305), .ZN(n7480) );
  OAI222_X1 U8621 ( .A1(n8777), .A2(n7480), .B1(n8775), .B2(n7463), .C1(n7462), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  NAND2_X1 U8622 ( .A1(n7464), .A2(n9556), .ZN(n7465) );
  OR2_X1 U8623 ( .A1(n7486), .A2(n7515), .ZN(n9406) );
  NAND2_X1 U8624 ( .A1(n7486), .A2(n7515), .ZN(n9407) );
  NAND2_X1 U8625 ( .A1(n9406), .A2(n9407), .ZN(n9361) );
  INV_X1 U8626 ( .A(n9361), .ZN(n9405) );
  XNOR2_X1 U8627 ( .A(n7487), .B(n9405), .ZN(n10586) );
  INV_X1 U8628 ( .A(n10586), .ZN(n7479) );
  AOI21_X1 U8629 ( .B1(n7467), .B2(n7486), .A(n10565), .ZN(n7468) );
  NAND2_X1 U8630 ( .A1(n7468), .A2(n7500), .ZN(n10581) );
  AND2_X1 U8631 ( .A1(n9403), .A2(n9395), .ZN(n9324) );
  NAND2_X1 U8632 ( .A1(n9328), .A2(n9324), .ZN(n7497) );
  NAND2_X1 U8633 ( .A1(n7497), .A2(n9402), .ZN(n7469) );
  XNOR2_X1 U8634 ( .A(n7469), .B(n9405), .ZN(n7471) );
  AOI22_X1 U8635 ( .A1(n10516), .A2(n9556), .B1(n10514), .B2(n9554), .ZN(n7470) );
  OAI21_X1 U8636 ( .B1(n7471), .B2(n10518), .A(n7470), .ZN(n7472) );
  AOI21_X1 U8637 ( .B1(n10586), .B2(n9764), .A(n7472), .ZN(n10588) );
  OAI21_X1 U8638 ( .B1(n10493), .B2(n10581), .A(n10588), .ZN(n7473) );
  NAND2_X1 U8639 ( .A1(n7473), .A2(n10539), .ZN(n7478) );
  INV_X1 U8640 ( .A(n7474), .ZN(n7475) );
  OAI22_X1 U8641 ( .A1(n10539), .A2(n6321), .B1(n7475), .B2(n10488), .ZN(n7476) );
  AOI21_X1 U8642 ( .B1(n9702), .B2(n7486), .A(n7476), .ZN(n7477) );
  OAI211_X1 U8643 ( .C1(n7479), .C2(n9757), .A(n7478), .B(n7477), .ZN(P1_U3282) );
  INV_X1 U8644 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7481) );
  OAI222_X1 U8645 ( .A1(n8781), .A2(n7481), .B1(n7619), .B2(n7480), .C1(n8423), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U8646 ( .A1(n7482), .A2(n6944), .ZN(n7485) );
  AOI22_X1 U8647 ( .A1(n8280), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6704), .B2(
        n7483), .ZN(n7484) );
  OR2_X1 U8648 ( .A1(n7728), .A2(n7535), .ZN(n9411) );
  NAND2_X1 U8649 ( .A1(n7728), .A2(n7535), .ZN(n9412) );
  AOI21_X1 U8650 ( .B1(n9409), .B2(n7488), .A(n4931), .ZN(n7636) );
  NOR2_X1 U8651 ( .A1(n7489), .A2(n4854), .ZN(n10496) );
  NAND2_X1 U8652 ( .A1(n10539), .A2(n10496), .ZN(n9718) );
  NAND2_X1 U8653 ( .A1(n4874), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7496) );
  INV_X1 U8654 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7490) );
  NAND2_X1 U8655 ( .A1(n7491), .A2(n7490), .ZN(n7492) );
  AND2_X1 U8656 ( .A1(n7527), .A2(n7492), .ZN(n7734) );
  NAND2_X1 U8657 ( .A1(n6823), .A2(n7734), .ZN(n7495) );
  NAND2_X1 U8658 ( .A1(n6800), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U8659 ( .A1(n6801), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7493) );
  AND2_X1 U8660 ( .A1(n9406), .A2(n9402), .ZN(n9313) );
  NAND2_X1 U8661 ( .A1(n7497), .A2(n9313), .ZN(n7498) );
  NAND2_X1 U8662 ( .A1(n7498), .A2(n9407), .ZN(n7726) );
  INV_X1 U8663 ( .A(n9409), .ZN(n9362) );
  XNOR2_X1 U8664 ( .A(n7726), .B(n9362), .ZN(n7499) );
  OAI222_X1 U8665 ( .A1(n9745), .A2(n7896), .B1(n7499), .B2(n10518), .C1(n9743), .C2(n7515), .ZN(n7633) );
  INV_X1 U8666 ( .A(n7728), .ZN(n7503) );
  AOI211_X1 U8667 ( .C1(n7728), .C2(n7500), .A(n10565), .B(n7733), .ZN(n7634)
         );
  NAND2_X1 U8668 ( .A1(n7634), .A2(n8076), .ZN(n7502) );
  AOI22_X1 U8669 ( .A1(n10498), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7511), .B2(
        n10544), .ZN(n7501) );
  OAI211_X1 U8670 ( .C1(n7503), .C2(n10538), .A(n7502), .B(n7501), .ZN(n7504)
         );
  AOI21_X1 U8671 ( .B1(n7633), .B2(n10539), .A(n7504), .ZN(n7505) );
  OAI21_X1 U8672 ( .B1(n7636), .B2(n9718), .A(n7505), .ZN(P1_U3281) );
  AOI22_X1 U8673 ( .A1(n7728), .A2(n4856), .B1(n8752), .B2(n9554), .ZN(n7508)
         );
  XOR2_X1 U8674 ( .A(n8761), .B(n7508), .Z(n7509) );
  NAND2_X1 U8675 ( .A1(n4933), .A2(n7519), .ZN(n7510) );
  AOI22_X1 U8676 ( .A1(n7728), .A2(n8752), .B1(n8744), .B2(n9554), .ZN(n7520)
         );
  XNOR2_X1 U8677 ( .A(n7510), .B(n7520), .ZN(n7518) );
  NAND2_X1 U8678 ( .A1(n9280), .A2(n7511), .ZN(n7514) );
  INV_X1 U8679 ( .A(n7896), .ZN(n9553) );
  AOI21_X1 U8680 ( .B1(n9262), .B2(n9553), .A(n7512), .ZN(n7513) );
  OAI211_X1 U8681 ( .C1(n7515), .C2(n9284), .A(n7514), .B(n7513), .ZN(n7516)
         );
  AOI21_X1 U8682 ( .B1(n7728), .B2(n9287), .A(n7516), .ZN(n7517) );
  OAI21_X1 U8683 ( .B1(n7518), .B2(n9289), .A(n7517), .ZN(P1_U3215) );
  NAND2_X1 U8684 ( .A1(n7521), .A2(n6944), .ZN(n7523) );
  AOI22_X1 U8685 ( .A1(n8280), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6704), .B2(
        n10238), .ZN(n7522) );
  NAND2_X1 U8686 ( .A1(n7523), .A2(n7522), .ZN(n7897) );
  INV_X1 U8687 ( .A(n7897), .ZN(n7762) );
  OAI22_X1 U8688 ( .A1(n7762), .A2(n8764), .B1(n7896), .B2(n8763), .ZN(n7524)
         );
  XNOR2_X1 U8689 ( .A(n7524), .B(n8761), .ZN(n7671) );
  NOR2_X1 U8690 ( .A1(n8760), .A2(n7896), .ZN(n7525) );
  AOI21_X1 U8691 ( .B1(n7897), .B2(n8752), .A(n7525), .ZN(n7669) );
  XNOR2_X1 U8692 ( .A(n7671), .B(n7669), .ZN(n7673) );
  XNOR2_X1 U8693 ( .A(n7674), .B(n7673), .ZN(n7538) );
  NAND2_X1 U8694 ( .A1(n9280), .A2(n7734), .ZN(n7534) );
  NAND2_X1 U8695 ( .A1(n6800), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U8696 ( .A1(n7527), .A2(n7526), .ZN(n7528) );
  AND2_X1 U8697 ( .A1(n7688), .A2(n7528), .ZN(n7910) );
  NAND2_X1 U8698 ( .A1(n6823), .A2(n7910), .ZN(n7531) );
  NAND2_X1 U8699 ( .A1(n4874), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7530) );
  NAND2_X1 U8700 ( .A1(n6801), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7529) );
  INV_X1 U8701 ( .A(n7985), .ZN(n9552) );
  AND2_X1 U8702 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10224) );
  AOI21_X1 U8703 ( .B1(n9262), .B2(n9552), .A(n10224), .ZN(n7533) );
  OAI211_X1 U8704 ( .C1(n7535), .C2(n9284), .A(n7534), .B(n7533), .ZN(n7536)
         );
  AOI21_X1 U8705 ( .B1(n7897), .B2(n9287), .A(n7536), .ZN(n7537) );
  OAI21_X1 U8706 ( .B1(n7538), .B2(n9289), .A(n7537), .ZN(P1_U3234) );
  OAI21_X1 U8707 ( .B1(n7546), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7539), .ZN(
        n7564) );
  XNOR2_X1 U8708 ( .A(n7567), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7563) );
  NOR2_X1 U8709 ( .A1(n7564), .A2(n7563), .ZN(n7562) );
  MUX2_X1 U8710 ( .A(n7780), .B(P2_REG2_REG_13__SCAN_IN), .S(n7650), .Z(n7540)
         );
  INV_X1 U8711 ( .A(n7540), .ZN(n7541) );
  OAI21_X1 U8712 ( .B1(n7542), .B2(n7541), .A(n7644), .ZN(n7543) );
  NAND2_X1 U8713 ( .A1(n7543), .A2(n8896), .ZN(n7554) );
  INV_X1 U8714 ( .A(n10297), .ZN(n10278) );
  MUX2_X1 U8715 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n7544), .S(n7650), .Z(n7549)
         );
  AOI21_X1 U8716 ( .B1(n7546), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7545), .ZN(
        n7557) );
  XNOR2_X1 U8717 ( .A(n7567), .B(n7547), .ZN(n7558) );
  NAND2_X1 U8718 ( .A1(n7557), .A2(n7558), .ZN(n7556) );
  OAI21_X1 U8719 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7567), .A(n7556), .ZN(
        n7548) );
  NAND2_X1 U8720 ( .A1(n7548), .A2(n7549), .ZN(n7649) );
  OAI21_X1 U8721 ( .B1(n7549), .B2(n7548), .A(n7649), .ZN(n7552) );
  INV_X1 U8722 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7550) );
  NAND2_X1 U8723 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n7664) );
  OAI21_X1 U8724 ( .B1(n8893), .B2(n7550), .A(n7664), .ZN(n7551) );
  AOI21_X1 U8725 ( .B1(n10278), .B2(n7552), .A(n7551), .ZN(n7553) );
  OAI211_X1 U8726 ( .C1(n8891), .C2(n7555), .A(n7554), .B(n7553), .ZN(P2_U3258) );
  INV_X1 U8727 ( .A(n8891), .ZN(n10308) );
  INV_X1 U8728 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7561) );
  OAI21_X1 U8729 ( .B1(n7558), .B2(n7557), .A(n7556), .ZN(n7559) );
  NAND2_X1 U8730 ( .A1(n10278), .A2(n7559), .ZN(n7560) );
  NAND2_X1 U8731 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7625) );
  OAI211_X1 U8732 ( .C1(n7561), .C2(n8893), .A(n7560), .B(n7625), .ZN(n7566)
         );
  AOI211_X1 U8733 ( .C1(n7564), .C2(n7563), .A(n10301), .B(n7562), .ZN(n7565)
         );
  AOI211_X1 U8734 ( .C1(n10308), .C2(n7567), .A(n7566), .B(n7565), .ZN(n7568)
         );
  INV_X1 U8735 ( .A(n7568), .ZN(P2_U3257) );
  OR2_X1 U8736 ( .A1(n10612), .A2(n7627), .ZN(n8508) );
  NAND2_X1 U8737 ( .A1(n10612), .A2(n7627), .ZN(n8506) );
  NAND2_X1 U8738 ( .A1(n8508), .A2(n8506), .ZN(n7592) );
  INV_X1 U8739 ( .A(n7592), .ZN(n8612) );
  NAND2_X1 U8740 ( .A1(n7569), .A2(n8612), .ZN(n7587) );
  NAND3_X1 U8741 ( .A1(n7570), .A2(n8505), .A3(n7592), .ZN(n7571) );
  NAND2_X1 U8742 ( .A1(n7587), .A2(n7571), .ZN(n7572) );
  INV_X1 U8743 ( .A(n7776), .ZN(n8857) );
  AOI222_X1 U8744 ( .A1(n9085), .A2(n7572), .B1(n8857), .B2(n9082), .C1(n8859), 
        .C2(n9080), .ZN(n10614) );
  AOI21_X1 U8745 ( .B1(n7573), .B2(n10612), .A(n10639), .ZN(n7574) );
  NAND2_X1 U8746 ( .A1(n7574), .A2(n7601), .ZN(n10613) );
  NAND2_X1 U8747 ( .A1(n7575), .A2(n8859), .ZN(n7590) );
  NAND2_X1 U8748 ( .A1(n7598), .A2(n7590), .ZN(n7577) );
  NAND2_X1 U8749 ( .A1(n7577), .A2(n7592), .ZN(n7576) );
  OAI21_X1 U8750 ( .B1(n7577), .B2(n7592), .A(n7576), .ZN(n7578) );
  INV_X1 U8751 ( .A(n7578), .ZN(n10617) );
  NAND2_X1 U8752 ( .A1(n10617), .A2(n10457), .ZN(n7583) );
  OAI22_X1 U8753 ( .A1(n4833), .A2(n7580), .B1(n7579), .B2(n10373), .ZN(n7581)
         );
  AOI21_X1 U8754 ( .B1(n10466), .B2(n10612), .A(n7581), .ZN(n7582) );
  OAI211_X1 U8755 ( .C1(n10613), .C2(n7584), .A(n7583), .B(n7582), .ZN(n7585)
         );
  INV_X1 U8756 ( .A(n7585), .ZN(n7586) );
  OAI21_X1 U8757 ( .B1(n10614), .B2(n10469), .A(n7586), .ZN(P2_U3285) );
  NAND2_X1 U8758 ( .A1(n10149), .A2(n7776), .ZN(n8456) );
  XNOR2_X1 U8759 ( .A(n7772), .B(n7599), .ZN(n7589) );
  OAI22_X1 U8760 ( .A1(n7627), .A2(n10439), .B1(n7882), .B2(n10441), .ZN(n7588) );
  AOI21_X1 U8761 ( .B1(n7589), .B2(n9085), .A(n7588), .ZN(n10153) );
  NAND2_X1 U8762 ( .A1(n10612), .A2(n8858), .ZN(n7591) );
  AND2_X1 U8763 ( .A1(n7590), .A2(n7591), .ZN(n7595) );
  NAND2_X1 U8764 ( .A1(n7598), .A2(n7595), .ZN(n7594) );
  INV_X1 U8765 ( .A(n7591), .ZN(n7593) );
  OR2_X1 U8766 ( .A1(n7593), .A2(n7592), .ZN(n7596) );
  NAND2_X1 U8767 ( .A1(n7594), .A2(n7596), .ZN(n7600) );
  AND2_X1 U8768 ( .A1(n7595), .A2(n7599), .ZN(n7597) );
  AOI21_X1 U8769 ( .B1(n7598), .B2(n7597), .A(n4871), .ZN(n7782) );
  OAI21_X1 U8770 ( .B1(n7600), .B2(n7599), .A(n7782), .ZN(n10148) );
  AOI21_X1 U8771 ( .B1(n10149), .B2(n7601), .A(n7778), .ZN(n10151) );
  NAND2_X1 U8772 ( .A1(n10151), .A2(n10461), .ZN(n7604) );
  INV_X1 U8773 ( .A(n7626), .ZN(n7602) );
  INV_X1 U8774 ( .A(n10373), .ZN(n10458) );
  AOI22_X1 U8775 ( .A1(n10469), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7602), .B2(
        n10458), .ZN(n7603) );
  OAI211_X1 U8776 ( .C1(n5139), .C2(n9076), .A(n7604), .B(n7603), .ZN(n7605)
         );
  AOI21_X1 U8777 ( .B1(n10148), .B2(n10457), .A(n7605), .ZN(n7606) );
  OAI21_X1 U8778 ( .B1(n10153), .B2(n10469), .A(n7606), .ZN(P2_U3284) );
  NAND2_X1 U8779 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7821) );
  INV_X1 U8780 ( .A(n7821), .ZN(n7611) );
  AOI211_X1 U8781 ( .C1(n7609), .C2(n7608), .A(n7607), .B(n10321), .ZN(n7610)
         );
  AOI211_X1 U8782 ( .C1(n7807), .C2(n10257), .A(n7611), .B(n7610), .ZN(n7617)
         );
  OAI21_X1 U8783 ( .B1(n7614), .B2(n7613), .A(n7612), .ZN(n7615) );
  AOI22_X1 U8784 ( .A1(n10259), .A2(P1_ADDR_REG_14__SCAN_IN), .B1(n10329), 
        .B2(n7615), .ZN(n7616) );
  NAND2_X1 U8785 ( .A1(n7617), .A2(n7616), .ZN(P1_U3255) );
  INV_X1 U8786 ( .A(n8317), .ZN(n7618) );
  OAI222_X1 U8787 ( .A1(n8775), .A2(n8318), .B1(n8777), .B2(n7618), .C1(n9502), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  OAI222_X1 U8788 ( .A1(n8781), .A2(n7620), .B1(n7619), .B2(n7618), .C1(
        P2_U3152), .C2(n6173), .ZN(P2_U3336) );
  OAI21_X1 U8789 ( .B1(n7623), .B2(n7622), .A(n7621), .ZN(n7624) );
  NAND2_X1 U8790 ( .A1(n7624), .A2(n8844), .ZN(n7632) );
  INV_X1 U8791 ( .A(n7625), .ZN(n7629) );
  OAI22_X1 U8792 ( .A1(n10393), .A2(n7627), .B1(n8848), .B2(n7626), .ZN(n7628)
         );
  AOI211_X1 U8793 ( .C1(n8802), .C2(n7630), .A(n7629), .B(n7628), .ZN(n7631)
         );
  OAI211_X1 U8794 ( .C1(n5139), .C2(n10399), .A(n7632), .B(n7631), .ZN(
        P2_U3226) );
  INV_X1 U8795 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7638) );
  AND2_X1 U8796 ( .A1(n10526), .A2(n10552), .ZN(n9863) );
  AOI211_X1 U8797 ( .C1(n10549), .C2(n7728), .A(n7634), .B(n7633), .ZN(n7635)
         );
  OAI21_X1 U8798 ( .B1(n7636), .B2(n9863), .A(n7635), .ZN(n7641) );
  NAND2_X1 U8799 ( .A1(n7641), .A2(n10595), .ZN(n7637) );
  OAI21_X1 U8800 ( .B1(n10595), .B2(n7638), .A(n7637), .ZN(P1_U3484) );
  AND2_X2 U8801 ( .A1(n7640), .A2(n7639), .ZN(n10591) );
  NAND2_X1 U8802 ( .A1(n7641), .A2(n10591), .ZN(n7642) );
  OAI21_X1 U8803 ( .B1(n10591), .B2(n7643), .A(n7642), .ZN(P1_U3533) );
  MUX2_X1 U8804 ( .A(n7887), .B(P2_REG2_REG_14__SCAN_IN), .S(n7973), .Z(n7645)
         );
  INV_X1 U8805 ( .A(n7645), .ZN(n7646) );
  OAI21_X1 U8806 ( .B1(n7647), .B2(n7646), .A(n7972), .ZN(n7648) );
  NAND2_X1 U8807 ( .A1(n7648), .A2(n8896), .ZN(n7658) );
  OAI21_X1 U8808 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7650), .A(n7649), .ZN(
        n7653) );
  MUX2_X1 U8809 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7651), .S(n7973), .Z(n7652)
         );
  NAND2_X1 U8810 ( .A1(n7652), .A2(n7653), .ZN(n7965) );
  OAI21_X1 U8811 ( .B1(n7653), .B2(n7652), .A(n7965), .ZN(n7656) );
  INV_X1 U8812 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7654) );
  NAND2_X1 U8813 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7744) );
  OAI21_X1 U8814 ( .B1(n8893), .B2(n7654), .A(n7744), .ZN(n7655) );
  AOI21_X1 U8815 ( .B1(n10278), .B2(n7656), .A(n7655), .ZN(n7657) );
  OAI211_X1 U8816 ( .C1(n8891), .C2(n7659), .A(n7658), .B(n7657), .ZN(P2_U3259) );
  OAI21_X1 U8817 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n7663) );
  NAND2_X1 U8818 ( .A1(n7663), .A2(n8844), .ZN(n7668) );
  INV_X1 U8819 ( .A(n7956), .ZN(n8856) );
  INV_X1 U8820 ( .A(n7664), .ZN(n7666) );
  OAI22_X1 U8821 ( .A1(n10393), .A2(n7776), .B1(n8848), .B2(n7770), .ZN(n7665)
         );
  AOI211_X1 U8822 ( .C1(n8802), .C2(n8856), .A(n7666), .B(n7665), .ZN(n7667)
         );
  OAI211_X1 U8823 ( .C1(n10622), .C2(n10399), .A(n7668), .B(n7667), .ZN(
        P2_U3236) );
  INV_X1 U8824 ( .A(n7669), .ZN(n7670) );
  NAND2_X1 U8825 ( .A1(n7675), .A2(n6944), .ZN(n7678) );
  AOI22_X1 U8826 ( .A1(n8280), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6704), .B2(
        n7676), .ZN(n7677) );
  NAND2_X1 U8827 ( .A1(n9877), .A2(n4855), .ZN(n7680) );
  NAND2_X1 U8828 ( .A1(n9552), .A2(n8752), .ZN(n7679) );
  NAND2_X1 U8829 ( .A1(n7680), .A2(n7679), .ZN(n7681) );
  XNOR2_X1 U8830 ( .A(n7681), .B(n4854), .ZN(n7684) );
  NOR2_X1 U8831 ( .A1(n8760), .A2(n7985), .ZN(n7682) );
  AOI21_X1 U8832 ( .B1(n9877), .B2(n8752), .A(n7682), .ZN(n7683) );
  AND2_X1 U8833 ( .A1(n7684), .A2(n7683), .ZN(n7705) );
  INV_X1 U8834 ( .A(n7705), .ZN(n7685) );
  OR2_X1 U8835 ( .A1(n7684), .A2(n7683), .ZN(n7704) );
  NAND2_X1 U8836 ( .A1(n7685), .A2(n7704), .ZN(n7686) );
  XNOR2_X1 U8837 ( .A(n7706), .B(n7686), .ZN(n7699) );
  NAND2_X1 U8838 ( .A1(n4874), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U8839 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  AND2_X1 U8840 ( .A1(n7714), .A2(n7689), .ZN(n7996) );
  NAND2_X1 U8841 ( .A1(n6823), .A2(n7996), .ZN(n7692) );
  NAND2_X1 U8842 ( .A1(n6800), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U8843 ( .A1(n6801), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7690) );
  NAND2_X1 U8844 ( .A1(n9280), .A2(n7910), .ZN(n7696) );
  AOI21_X1 U8845 ( .B1(n9250), .B2(n9553), .A(n7694), .ZN(n7695) );
  OAI211_X1 U8846 ( .C1(n9428), .C2(n9242), .A(n7696), .B(n7695), .ZN(n7697)
         );
  AOI21_X1 U8847 ( .B1(n9877), .B2(n9287), .A(n7697), .ZN(n7698) );
  OAI21_X1 U8848 ( .B1(n7699), .B2(n9289), .A(n7698), .ZN(P1_U3222) );
  INV_X1 U8849 ( .A(n8332), .ZN(n7701) );
  NAND2_X1 U8850 ( .A1(n8410), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7700) );
  OAI211_X1 U8851 ( .C1(n7701), .C2(n7619), .A(n7700), .B(n8644), .ZN(P2_U3335) );
  NAND2_X1 U8852 ( .A1(n8332), .A2(n8147), .ZN(n7703) );
  OR2_X1 U8853 ( .A1(n7702), .A2(P1_U3084), .ZN(n9542) );
  OAI211_X1 U8854 ( .C1(n8333), .C2(n8775), .A(n7703), .B(n9542), .ZN(P1_U3330) );
  NAND2_X1 U8855 ( .A1(n7707), .A2(n6944), .ZN(n7710) );
  AOI22_X1 U8856 ( .A1(n8280), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6704), .B2(
        n7708), .ZN(n7709) );
  INV_X1 U8857 ( .A(n9428), .ZN(n9551) );
  AOI22_X1 U8858 ( .A1(n9871), .A2(n4856), .B1(n8752), .B2(n9551), .ZN(n7711)
         );
  XOR2_X1 U8859 ( .A(n8761), .B(n7711), .Z(n7804) );
  AOI22_X1 U8860 ( .A1(n9871), .A2(n8752), .B1(n8744), .B2(n9551), .ZN(n7802)
         );
  XNOR2_X1 U8861 ( .A(n7804), .B(n7802), .ZN(n7712) );
  XNOR2_X1 U8862 ( .A(n7805), .B(n7712), .ZN(n7725) );
  NAND2_X1 U8863 ( .A1(n6800), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7719) );
  NAND2_X1 U8864 ( .A1(n4874), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7718) );
  INV_X1 U8865 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U8866 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  AND2_X1 U8867 ( .A1(n7815), .A2(n7715), .ZN(n7925) );
  NAND2_X1 U8868 ( .A1(n6823), .A2(n7925), .ZN(n7717) );
  NAND2_X1 U8869 ( .A1(n6801), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7716) );
  INV_X1 U8870 ( .A(n9430), .ZN(n9550) );
  NAND2_X1 U8871 ( .A1(n9262), .A2(n9550), .ZN(n7721) );
  OAI211_X1 U8872 ( .C1(n7985), .C2(n9284), .A(n7721), .B(n7720), .ZN(n7723)
         );
  INV_X1 U8873 ( .A(n9871), .ZN(n7998) );
  NOR2_X1 U8874 ( .A1(n7998), .A2(n9224), .ZN(n7722) );
  AOI211_X1 U8875 ( .C1(n7996), .C2(n9280), .A(n7723), .B(n7722), .ZN(n7724)
         );
  OAI21_X1 U8876 ( .B1(n7725), .B2(n9289), .A(n7724), .ZN(P1_U3232) );
  NAND2_X1 U8877 ( .A1(n7726), .A2(n9409), .ZN(n7727) );
  NAND2_X1 U8878 ( .A1(n7727), .A2(n9412), .ZN(n7893) );
  OR2_X1 U8879 ( .A1(n7897), .A2(n7896), .ZN(n9415) );
  NAND2_X1 U8880 ( .A1(n7897), .A2(n7896), .ZN(n9416) );
  NAND2_X1 U8881 ( .A1(n9415), .A2(n9416), .ZN(n9410) );
  XNOR2_X1 U8882 ( .A(n7893), .B(n9410), .ZN(n7732) );
  NAND2_X1 U8883 ( .A1(n7729), .A2(n9410), .ZN(n7899) );
  OAI21_X1 U8884 ( .B1(n7729), .B2(n9410), .A(n7899), .ZN(n7766) );
  NAND2_X1 U8885 ( .A1(n7766), .A2(n9764), .ZN(n7731) );
  AOI22_X1 U8886 ( .A1(n10516), .A2(n9554), .B1(n10514), .B2(n9552), .ZN(n7730) );
  OAI211_X1 U8887 ( .C1(n10518), .C2(n7732), .A(n7731), .B(n7730), .ZN(n7764)
         );
  INV_X1 U8888 ( .A(n7764), .ZN(n7739) );
  AND2_X1 U8889 ( .A1(n7733), .A2(n7762), .ZN(n7907) );
  INV_X1 U8890 ( .A(n7907), .ZN(n7909) );
  OAI21_X1 U8891 ( .B1(n7762), .B2(n7733), .A(n7909), .ZN(n7763) );
  AOI22_X1 U8892 ( .A1(n10498), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7734), .B2(
        n10544), .ZN(n7736) );
  NAND2_X1 U8893 ( .A1(n7897), .A2(n9702), .ZN(n7735) );
  OAI211_X1 U8894 ( .C1(n7763), .C2(n10333), .A(n7736), .B(n7735), .ZN(n7737)
         );
  AOI21_X1 U8895 ( .B1(n7766), .B2(n10535), .A(n7737), .ZN(n7738) );
  OAI21_X1 U8896 ( .B1(n7739), .B2(n10498), .A(n7738), .ZN(P1_U3280) );
  OAI21_X1 U8897 ( .B1(n7742), .B2(n7741), .A(n7740), .ZN(n7743) );
  NAND2_X1 U8898 ( .A1(n7743), .A2(n8844), .ZN(n7748) );
  INV_X1 U8899 ( .A(n7744), .ZN(n7746) );
  OAI22_X1 U8900 ( .A1(n10393), .A2(n7882), .B1(n8848), .B2(n7886), .ZN(n7745)
         );
  AOI211_X1 U8901 ( .C1(n8802), .C2(n8020), .A(n7746), .B(n7745), .ZN(n7747)
         );
  OAI211_X1 U8902 ( .C1(n10630), .C2(n10399), .A(n7748), .B(n7747), .ZN(
        P2_U3217) );
  INV_X1 U8903 ( .A(n8336), .ZN(n7751) );
  OAI222_X1 U8904 ( .A1(n8777), .A2(n7751), .B1(P1_U3084), .B2(n7749), .C1(
        n8337), .C2(n8775), .ZN(P1_U3329) );
  OAI222_X1 U8905 ( .A1(P2_U3152), .A2(n7752), .B1(n7619), .B2(n7751), .C1(
        n7750), .C2(n8781), .ZN(P2_U3334) );
  INV_X1 U8906 ( .A(n7753), .ZN(n7755) );
  NAND2_X1 U8907 ( .A1(n7755), .A2(n7754), .ZN(n7756) );
  XNOR2_X1 U8908 ( .A(n7757), .B(n7756), .ZN(n7761) );
  NAND2_X1 U8909 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8012) );
  OAI21_X1 U8910 ( .B1(n10394), .B2(n8032), .A(n8012), .ZN(n7759) );
  OAI22_X1 U8911 ( .A1(n10393), .A2(n7956), .B1(n8848), .B2(n7957), .ZN(n7758)
         );
  AOI211_X1 U8912 ( .C1(n10637), .C2(n8851), .A(n7759), .B(n7758), .ZN(n7760)
         );
  OAI21_X1 U8913 ( .B1(n7761), .B2(n10397), .A(n7760), .ZN(P2_U3243) );
  INV_X1 U8914 ( .A(n10552), .ZN(n10585) );
  INV_X1 U8915 ( .A(n10549), .ZN(n10582) );
  OAI22_X1 U8916 ( .A1(n7763), .A2(n10565), .B1(n7762), .B2(n10582), .ZN(n7765) );
  AOI211_X1 U8917 ( .C1(n10585), .C2(n7766), .A(n7765), .B(n7764), .ZN(n7769)
         );
  NAND2_X1 U8918 ( .A1(n10592), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7767) );
  OAI21_X1 U8919 ( .B1(n7769), .B2(n10592), .A(n7767), .ZN(P1_U3487) );
  NAND2_X1 U8920 ( .A1(n10589), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7768) );
  OAI21_X1 U8921 ( .B1(n7769), .B2(n10589), .A(n7768), .ZN(P1_U3534) );
  INV_X1 U8922 ( .A(n7770), .ZN(n7777) );
  OR2_X1 U8923 ( .A1(n7771), .A2(n7882), .ZN(n8516) );
  NAND2_X1 U8924 ( .A1(n7771), .A2(n7882), .ZN(n8517) );
  NAND2_X1 U8925 ( .A1(n8516), .A2(n8517), .ZN(n8616) );
  INV_X1 U8926 ( .A(n8616), .ZN(n8515) );
  OAI21_X1 U8927 ( .B1(n8515), .B2(n7773), .A(n7879), .ZN(n7774) );
  INV_X1 U8928 ( .A(n7774), .ZN(n7775) );
  OAI222_X1 U8929 ( .A1(n10441), .A2(n7956), .B1(n10439), .B2(n7776), .C1(
        n10437), .C2(n7775), .ZN(n10624) );
  AOI21_X1 U8930 ( .B1(n7777), .B2(n10458), .A(n10624), .ZN(n7789) );
  NOR2_X1 U8931 ( .A1(n7778), .A2(n10622), .ZN(n7779) );
  OR2_X1 U8932 ( .A1(n7885), .A2(n7779), .ZN(n10623) );
  INV_X1 U8933 ( .A(n10623), .ZN(n7787) );
  OAI22_X1 U8934 ( .A1(n10622), .A2(n9076), .B1(n7780), .B2(n4833), .ZN(n7786)
         );
  OR2_X1 U8935 ( .A1(n10149), .A2(n8857), .ZN(n7781) );
  NOR2_X1 U8936 ( .A1(n7783), .A2(n8616), .ZN(n10621) );
  INV_X1 U8937 ( .A(n7877), .ZN(n7784) );
  NOR3_X1 U8938 ( .A1(n10621), .A2(n7784), .A3(n9089), .ZN(n7785) );
  AOI211_X1 U8939 ( .C1(n10461), .C2(n7787), .A(n7786), .B(n7785), .ZN(n7788)
         );
  OAI21_X1 U8940 ( .B1(n10469), .B2(n7789), .A(n7788), .ZN(P2_U3283) );
  INV_X1 U8941 ( .A(n7790), .ZN(n8058) );
  NAND2_X1 U8942 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8123) );
  INV_X1 U8943 ( .A(n8123), .ZN(n7795) );
  AOI211_X1 U8944 ( .C1(n7793), .C2(n7792), .A(n7791), .B(n10236), .ZN(n7794)
         );
  AOI211_X1 U8945 ( .C1(n10257), .C2(n8058), .A(n7795), .B(n7794), .ZN(n7801)
         );
  AOI211_X1 U8946 ( .C1(n7798), .C2(n7797), .A(n7796), .B(n10321), .ZN(n7799)
         );
  AOI21_X1 U8947 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n10259), .A(n7799), .ZN(
        n7800) );
  NAND2_X1 U8948 ( .A1(n7801), .A2(n7800), .ZN(P1_U3256) );
  INV_X1 U8949 ( .A(n7802), .ZN(n7803) );
  NAND2_X1 U8950 ( .A1(n7806), .A2(n6944), .ZN(n7809) );
  AOI22_X1 U8951 ( .A1(n8280), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6704), .B2(
        n7807), .ZN(n7808) );
  NAND2_X1 U8952 ( .A1(n9434), .A2(n4855), .ZN(n7811) );
  NAND2_X1 U8953 ( .A1(n9550), .A2(n8752), .ZN(n7810) );
  NAND2_X1 U8954 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  XNOR2_X1 U8955 ( .A(n7812), .B(n4854), .ZN(n8105) );
  INV_X1 U8956 ( .A(n9434), .ZN(n9866) );
  OAI22_X1 U8957 ( .A1(n9866), .A2(n8763), .B1(n9430), .B2(n8760), .ZN(n8092)
         );
  XNOR2_X1 U8958 ( .A(n8105), .B(n8092), .ZN(n7813) );
  XNOR2_X1 U8959 ( .A(n8093), .B(n7813), .ZN(n7826) );
  NAND2_X1 U8960 ( .A1(n7815), .A2(n7814), .ZN(n7816) );
  AND2_X1 U8961 ( .A1(n8067), .A2(n7816), .ZN(n8216) );
  NAND2_X1 U8962 ( .A1(n8216), .A2(n6823), .ZN(n7820) );
  NAND2_X1 U8963 ( .A1(n4874), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U8964 ( .A1(n6800), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U8965 ( .A1(n6801), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7817) );
  INV_X1 U8966 ( .A(n8094), .ZN(n9549) );
  NAND2_X1 U8967 ( .A1(n9262), .A2(n9549), .ZN(n7822) );
  OAI211_X1 U8968 ( .C1(n9428), .C2(n9284), .A(n7822), .B(n7821), .ZN(n7824)
         );
  NOR2_X1 U8969 ( .A1(n9866), .A2(n9224), .ZN(n7823) );
  AOI211_X1 U8970 ( .C1(n7925), .C2(n9280), .A(n7824), .B(n7823), .ZN(n7825)
         );
  OAI21_X1 U8971 ( .B1(n7826), .B2(n9289), .A(n7825), .ZN(P1_U3213) );
  INV_X1 U8972 ( .A(n8349), .ZN(n7829) );
  OAI222_X1 U8973 ( .A1(n8781), .A2(n7828), .B1(n7619), .B2(n7829), .C1(n7827), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U8974 ( .A1(P1_U3084), .A2(n6490), .B1(n8777), .B2(n7829), .C1(
        n8775), .C2(n8350), .ZN(P1_U3328) );
  AOI21_X1 U8975 ( .B1(n7831), .B2(n7830), .A(n4926), .ZN(n7835) );
  OAI22_X1 U8976 ( .A1(n8229), .A2(n10441), .B1(n7952), .B2(n10439), .ZN(n8038) );
  AOI22_X1 U8977 ( .A1(n8815), .A2(n8038), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n7832) );
  OAI21_X1 U8978 ( .B1(n8848), .B2(n8046), .A(n7832), .ZN(n7833) );
  AOI21_X1 U8979 ( .B1(n9169), .B2(n8851), .A(n7833), .ZN(n7834) );
  OAI21_X1 U8980 ( .B1(n7835), .B2(n10397), .A(n7834), .ZN(P2_U3228) );
  NOR2_X1 U8981 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7872) );
  NOR2_X1 U8982 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7870) );
  NOR2_X1 U8983 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7868) );
  NOR2_X1 U8984 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7866) );
  NOR2_X1 U8985 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7864) );
  NOR2_X1 U8986 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7862) );
  NAND2_X1 U8987 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7860) );
  XOR2_X1 U8988 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10182) );
  NAND2_X1 U8989 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7858) );
  XOR2_X1 U8990 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10180) );
  NOR2_X1 U8991 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7842) );
  XNOR2_X1 U8992 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10166) );
  NAND2_X1 U8993 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7840) );
  XOR2_X1 U8994 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10164) );
  NAND2_X1 U8995 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7838) );
  XOR2_X1 U8996 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10162) );
  AOI21_X1 U8997 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10157) );
  INV_X1 U8998 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7836) );
  NAND3_X1 U8999 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10159) );
  OAI21_X1 U9000 ( .B1(n10157), .B2(n7836), .A(n10159), .ZN(n10161) );
  NAND2_X1 U9001 ( .A1(n10162), .A2(n10161), .ZN(n7837) );
  NAND2_X1 U9002 ( .A1(n7838), .A2(n7837), .ZN(n10163) );
  NAND2_X1 U9003 ( .A1(n10164), .A2(n10163), .ZN(n7839) );
  NAND2_X1 U9004 ( .A1(n7840), .A2(n7839), .ZN(n10165) );
  NOR2_X1 U9005 ( .A1(n10166), .A2(n10165), .ZN(n7841) );
  NOR2_X1 U9006 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  NOR2_X1 U9007 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7843), .ZN(n10167) );
  AND2_X1 U9008 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7843), .ZN(n10168) );
  NOR2_X1 U9009 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10168), .ZN(n7844) );
  NOR2_X1 U9010 ( .A1(n10167), .A2(n7844), .ZN(n7845) );
  NAND2_X1 U9011 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7845), .ZN(n7847) );
  XOR2_X1 U9012 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7845), .Z(n10172) );
  NAND2_X1 U9013 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10172), .ZN(n7846) );
  NAND2_X1 U9014 ( .A1(n7847), .A2(n7846), .ZN(n7848) );
  NAND2_X1 U9015 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7848), .ZN(n7850) );
  XOR2_X1 U9016 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7848), .Z(n10174) );
  NAND2_X1 U9017 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10174), .ZN(n7849) );
  NAND2_X1 U9018 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  NAND2_X1 U9019 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7851), .ZN(n7853) );
  XOR2_X1 U9020 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7851), .Z(n10176) );
  NAND2_X1 U9021 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10176), .ZN(n7852) );
  NAND2_X1 U9022 ( .A1(n7853), .A2(n7852), .ZN(n7854) );
  NAND2_X1 U9023 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7854), .ZN(n7856) );
  XOR2_X1 U9024 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7854), .Z(n10178) );
  NAND2_X1 U9025 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10178), .ZN(n7855) );
  NAND2_X1 U9026 ( .A1(n7856), .A2(n7855), .ZN(n10179) );
  NAND2_X1 U9027 ( .A1(n10180), .A2(n10179), .ZN(n7857) );
  NAND2_X1 U9028 ( .A1(n7858), .A2(n7857), .ZN(n10181) );
  NAND2_X1 U9029 ( .A1(n10182), .A2(n10181), .ZN(n7859) );
  NAND2_X1 U9030 ( .A1(n7860), .A2(n7859), .ZN(n10184) );
  XNOR2_X1 U9031 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10183) );
  NOR2_X1 U9032 ( .A1(n10184), .A2(n10183), .ZN(n7861) );
  NOR2_X1 U9033 ( .A1(n7862), .A2(n7861), .ZN(n10186) );
  XNOR2_X1 U9034 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10185) );
  NOR2_X1 U9035 ( .A1(n10186), .A2(n10185), .ZN(n7863) );
  NOR2_X1 U9036 ( .A1(n7864), .A2(n7863), .ZN(n10188) );
  XNOR2_X1 U9037 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10187) );
  NOR2_X1 U9038 ( .A1(n10188), .A2(n10187), .ZN(n7865) );
  NOR2_X1 U9039 ( .A1(n7866), .A2(n7865), .ZN(n10190) );
  XNOR2_X1 U9040 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10189) );
  NOR2_X1 U9041 ( .A1(n10190), .A2(n10189), .ZN(n7867) );
  NOR2_X1 U9042 ( .A1(n7868), .A2(n7867), .ZN(n10192) );
  XNOR2_X1 U9043 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10191) );
  NOR2_X1 U9044 ( .A1(n10192), .A2(n10191), .ZN(n7869) );
  NOR2_X1 U9045 ( .A1(n7870), .A2(n7869), .ZN(n10194) );
  XNOR2_X1 U9046 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10193) );
  NOR2_X1 U9047 ( .A1(n10194), .A2(n10193), .ZN(n7871) );
  NOR2_X1 U9048 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  AND2_X1 U9049 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7873), .ZN(n10195) );
  NOR2_X1 U9050 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10195), .ZN(n7874) );
  NOR2_X1 U9051 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7873), .ZN(n10196) );
  NOR2_X1 U9052 ( .A1(n7874), .A2(n10196), .ZN(n7876) );
  XNOR2_X1 U9053 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7875) );
  XNOR2_X1 U9054 ( .A(n7876), .B(n7875), .ZN(ADD_1071_U4) );
  NAND2_X1 U9055 ( .A1(n7889), .A2(n7956), .ZN(n8454) );
  AOI21_X1 U9056 ( .B1(n8619), .B2(n7878), .A(n4927), .ZN(n10629) );
  AOI211_X1 U9057 ( .C1(n7881), .C2(n7880), .A(n10437), .B(n7954), .ZN(n7884)
         );
  OAI22_X1 U9058 ( .A1(n7882), .A2(n10439), .B1(n7952), .B2(n10441), .ZN(n7883) );
  OR2_X1 U9059 ( .A1(n7884), .A2(n7883), .ZN(n10632) );
  OAI21_X1 U9060 ( .B1(n7885), .B2(n10630), .A(n8024), .ZN(n10631) );
  OAI22_X1 U9061 ( .A1(n4833), .A2(n7887), .B1(n7886), .B2(n10373), .ZN(n7888)
         );
  AOI21_X1 U9062 ( .B1(n7889), .B2(n10466), .A(n7888), .ZN(n7890) );
  OAI21_X1 U9063 ( .B1(n10631), .B2(n9008), .A(n7890), .ZN(n7891) );
  AOI21_X1 U9064 ( .B1(n10632), .B2(n4833), .A(n7891), .ZN(n7892) );
  OAI21_X1 U9065 ( .B1(n10629), .B2(n9089), .A(n7892), .ZN(P2_U3282) );
  OR2_X1 U9066 ( .A1(n9877), .A2(n7985), .ZN(n9423) );
  NAND2_X1 U9067 ( .A1(n9877), .A2(n7985), .ZN(n9421) );
  NAND2_X1 U9068 ( .A1(n7893), .A2(n9415), .ZN(n7894) );
  NAND2_X1 U9069 ( .A1(n7894), .A2(n9416), .ZN(n7895) );
  NAND2_X1 U9070 ( .A1(n7895), .A2(n9418), .ZN(n7920) );
  OAI21_X1 U9071 ( .B1(n9418), .B2(n7895), .A(n7920), .ZN(n7906) );
  OAI22_X1 U9072 ( .A1(n9743), .A2(n7896), .B1(n9428), .B2(n9745), .ZN(n7905)
         );
  OR2_X1 U9073 ( .A1(n7897), .A2(n9553), .ZN(n7898) );
  NAND2_X1 U9074 ( .A1(n7899), .A2(n7898), .ZN(n7902) );
  INV_X1 U9075 ( .A(n7902), .ZN(n7901) );
  NAND2_X1 U9076 ( .A1(n7902), .A2(n9418), .ZN(n7903) );
  NAND2_X1 U9077 ( .A1(n7917), .A2(n7903), .ZN(n9880) );
  NOR2_X1 U9078 ( .A1(n9880), .A2(n10526), .ZN(n7904) );
  AOI211_X1 U9079 ( .C1(n10473), .C2(n7906), .A(n7905), .B(n7904), .ZN(n9879)
         );
  INV_X1 U9080 ( .A(n9877), .ZN(n7912) );
  INV_X1 U9081 ( .A(n7995), .ZN(n7908) );
  AOI211_X1 U9082 ( .C1(n9877), .C2(n7909), .A(n10565), .B(n7908), .ZN(n9876)
         );
  AOI22_X1 U9083 ( .A1(n10498), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7910), .B2(
        n10544), .ZN(n7911) );
  OAI21_X1 U9084 ( .B1(n7912), .B2(n10538), .A(n7911), .ZN(n7914) );
  NOR2_X1 U9085 ( .A1(n9880), .A2(n9757), .ZN(n7913) );
  AOI211_X1 U9086 ( .C1(n9876), .C2(n8076), .A(n7914), .B(n7913), .ZN(n7915)
         );
  OAI21_X1 U9087 ( .B1(n9879), .B2(n10498), .A(n7915), .ZN(P1_U3279) );
  NAND2_X1 U9088 ( .A1(n9877), .A2(n9552), .ZN(n7916) );
  OR2_X1 U9089 ( .A1(n9871), .A2(n9428), .ZN(n9438) );
  NAND2_X1 U9090 ( .A1(n9871), .A2(n9428), .ZN(n9425) );
  NAND2_X1 U9091 ( .A1(n9438), .A2(n9425), .ZN(n7987) );
  NAND2_X1 U9092 ( .A1(n9434), .A2(n9430), .ZN(n9426) );
  NAND2_X1 U9093 ( .A1(n9422), .A2(n9426), .ZN(n8083) );
  NAND2_X1 U9094 ( .A1(n7918), .A2(n8083), .ZN(n8056) );
  OR2_X1 U9095 ( .A1(n7918), .A2(n8083), .ZN(n7919) );
  NAND2_X1 U9096 ( .A1(n8056), .A2(n7919), .ZN(n9864) );
  INV_X1 U9097 ( .A(n9864), .ZN(n7931) );
  NAND2_X1 U9098 ( .A1(n7920), .A2(n9421), .ZN(n7984) );
  INV_X1 U9099 ( .A(n7987), .ZN(n9364) );
  NAND2_X1 U9100 ( .A1(n7984), .A2(n9364), .ZN(n7983) );
  NAND2_X1 U9101 ( .A1(n7983), .A2(n9425), .ZN(n8084) );
  INV_X1 U9102 ( .A(n8083), .ZN(n9365) );
  XNOR2_X1 U9103 ( .A(n8084), .B(n9365), .ZN(n7921) );
  NAND2_X1 U9104 ( .A1(n7921), .A2(n10473), .ZN(n7923) );
  AOI22_X1 U9105 ( .A1(n10516), .A2(n9551), .B1(n10514), .B2(n9549), .ZN(n7922) );
  NAND2_X1 U9106 ( .A1(n7923), .A2(n7922), .ZN(n9868) );
  AOI21_X1 U9107 ( .B1(n9434), .B2(n7993), .A(n10565), .ZN(n7924) );
  NAND2_X1 U9108 ( .A1(n7924), .A2(n8215), .ZN(n9865) );
  INV_X1 U9109 ( .A(n8076), .ZN(n7928) );
  AOI22_X1 U9110 ( .A1(n10498), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7925), .B2(
        n10544), .ZN(n7927) );
  NAND2_X1 U9111 ( .A1(n9434), .A2(n9702), .ZN(n7926) );
  OAI211_X1 U9112 ( .C1(n9865), .C2(n7928), .A(n7927), .B(n7926), .ZN(n7929)
         );
  AOI21_X1 U9113 ( .B1(n9868), .B2(n10539), .A(n7929), .ZN(n7930) );
  OAI21_X1 U9114 ( .B1(n7931), .B2(n9718), .A(n7930), .ZN(P1_U3277) );
  INV_X1 U9115 ( .A(n7932), .ZN(n7933) );
  NOR2_X1 U9116 ( .A1(n7934), .A2(n7933), .ZN(n7935) );
  XNOR2_X1 U9117 ( .A(n7936), .B(n7935), .ZN(n7940) );
  AOI22_X1 U9118 ( .A1(n8804), .A2(n8855), .B1(n8820), .B2(n8026), .ZN(n7937)
         );
  NAND2_X1 U9119 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n8200) );
  OAI211_X1 U9120 ( .C1(n8234), .C2(n10394), .A(n7937), .B(n8200), .ZN(n7938)
         );
  AOI21_X1 U9121 ( .B1(n9165), .B2(n8851), .A(n7938), .ZN(n7939) );
  OAI21_X1 U9122 ( .B1(n7940), .B2(n10397), .A(n7939), .ZN(P2_U3230) );
  AOI211_X1 U9123 ( .C1(n7943), .C2(n7942), .A(n7941), .B(n10321), .ZN(n7951)
         );
  AOI211_X1 U9124 ( .C1(n7946), .C2(n7945), .A(n7944), .B(n10236), .ZN(n7950)
         );
  NAND2_X1 U9125 ( .A1(n10259), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7947) );
  NAND2_X1 U9126 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8113) );
  OAI211_X1 U9127 ( .C1(n7948), .C2(n10318), .A(n7947), .B(n8113), .ZN(n7949)
         );
  OR3_X1 U9128 ( .A1(n7951), .A2(n7950), .A3(n7949), .ZN(P1_U3257) );
  NAND2_X1 U9129 ( .A1(n10637), .A2(n7952), .ZN(n8452) );
  XNOR2_X1 U9130 ( .A(n8021), .B(n8618), .ZN(n10643) );
  INV_X1 U9131 ( .A(n10643), .ZN(n7963) );
  INV_X1 U9132 ( .A(n8453), .ZN(n7953) );
  XOR2_X1 U9133 ( .A(n8618), .B(n8036), .Z(n7955) );
  OAI222_X1 U9134 ( .A1(n10441), .A2(n8032), .B1(n10439), .B2(n7956), .C1(
        n10437), .C2(n7955), .ZN(n10641) );
  XNOR2_X1 U9135 ( .A(n8024), .B(n10637), .ZN(n10640) );
  OAI22_X1 U9136 ( .A1(n4833), .A2(n7958), .B1(n7957), .B2(n10373), .ZN(n7959)
         );
  AOI21_X1 U9137 ( .B1(n10637), .B2(n10466), .A(n7959), .ZN(n7960) );
  OAI21_X1 U9138 ( .B1(n10640), .B2(n9008), .A(n7960), .ZN(n7961) );
  AOI21_X1 U9139 ( .B1(n10641), .B2(n4833), .A(n7961), .ZN(n7962) );
  OAI21_X1 U9140 ( .B1(n7963), .B2(n9089), .A(n7962), .ZN(P2_U3281) );
  INV_X1 U9141 ( .A(n8367), .ZN(n8003) );
  OAI222_X1 U9142 ( .A1(n8777), .A2(n8003), .B1(P1_U3084), .B2(n7964), .C1(
        n8368), .C2(n8775), .ZN(P1_U3327) );
  OAI21_X1 U9143 ( .B1(n7973), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7965), .ZN(
        n7966) );
  NOR2_X1 U9144 ( .A1(n8015), .A2(n7966), .ZN(n7967) );
  XNOR2_X1 U9145 ( .A(n8015), .B(n7966), .ZN(n8009) );
  NOR2_X1 U9146 ( .A1(n5871), .A2(n8009), .ZN(n8010) );
  NOR2_X1 U9147 ( .A1(n7967), .A2(n8010), .ZN(n8194) );
  XNOR2_X1 U9148 ( .A(n7969), .B(n7968), .ZN(n8196) );
  XNOR2_X1 U9149 ( .A(n8194), .B(n8196), .ZN(n7982) );
  INV_X1 U9150 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U9151 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n7970) );
  OAI21_X1 U9152 ( .B1(n8893), .B2(n7971), .A(n7970), .ZN(n7980) );
  OAI21_X1 U9153 ( .B1(n7973), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7972), .ZN(
        n7974) );
  NAND2_X1 U9154 ( .A1(n8015), .A2(n7974), .ZN(n7976) );
  INV_X1 U9155 ( .A(n7974), .ZN(n7975) );
  XNOR2_X1 U9156 ( .A(n8015), .B(n7975), .ZN(n8008) );
  NAND2_X1 U9157 ( .A1(n8008), .A2(n7958), .ZN(n8007) );
  NAND2_X1 U9158 ( .A1(n7976), .A2(n8007), .ZN(n7978) );
  XNOR2_X1 U9159 ( .A(n8195), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n7977) );
  NOR2_X1 U9160 ( .A1(n7978), .A2(n7977), .ZN(n8190) );
  AOI211_X1 U9161 ( .C1(n7978), .C2(n7977), .A(n10301), .B(n8190), .ZN(n7979)
         );
  AOI211_X1 U9162 ( .C1(n10308), .C2(n8195), .A(n7980), .B(n7979), .ZN(n7981)
         );
  OAI21_X1 U9163 ( .B1(n7982), .B2(n10297), .A(n7981), .ZN(P2_U3261) );
  OAI21_X1 U9164 ( .B1(n9364), .B2(n7984), .A(n7983), .ZN(n7992) );
  OAI22_X1 U9165 ( .A1(n9743), .A2(n7985), .B1(n9430), .B2(n9745), .ZN(n7991)
         );
  OAI21_X1 U9166 ( .B1(n7988), .B2(n7987), .A(n7986), .ZN(n7989) );
  INV_X1 U9167 ( .A(n7989), .ZN(n9875) );
  NOR2_X1 U9168 ( .A1(n9875), .A2(n10526), .ZN(n7990) );
  AOI211_X1 U9169 ( .C1(n10473), .C2(n7992), .A(n7991), .B(n7990), .ZN(n9874)
         );
  INV_X1 U9170 ( .A(n7993), .ZN(n7994) );
  AOI21_X1 U9171 ( .B1(n9871), .B2(n7995), .A(n7994), .ZN(n9872) );
  AOI22_X1 U9172 ( .A1(n10498), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7996), .B2(
        n10544), .ZN(n7997) );
  OAI21_X1 U9173 ( .B1(n7998), .B2(n10538), .A(n7997), .ZN(n8000) );
  NOR2_X1 U9174 ( .A1(n9875), .A2(n9757), .ZN(n7999) );
  AOI211_X1 U9175 ( .C1(n9872), .C2(n10534), .A(n8000), .B(n7999), .ZN(n8001)
         );
  OAI21_X1 U9176 ( .B1(n9874), .B2(n10498), .A(n8001), .ZN(P1_U3278) );
  OAI222_X1 U9177 ( .A1(n8004), .A2(P2_U3152), .B1(n7619), .B2(n8003), .C1(
        n8002), .C2(n8781), .ZN(P2_U3332) );
  NAND2_X1 U9178 ( .A1(n8664), .A2(n8147), .ZN(n8006) );
  OAI211_X1 U9179 ( .C1(n8775), .C2(n8665), .A(n8006), .B(n8005), .ZN(P1_U3326) );
  OAI21_X1 U9180 ( .B1(n8008), .B2(n7958), .A(n8007), .ZN(n8018) );
  INV_X1 U9181 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8014) );
  AND2_X1 U9182 ( .A1(n8009), .A2(n5871), .ZN(n8011) );
  OR3_X1 U9183 ( .A1(n10297), .A2(n8011), .A3(n8010), .ZN(n8013) );
  OAI211_X1 U9184 ( .C1(n8014), .C2(n8893), .A(n8013), .B(n8012), .ZN(n8017)
         );
  NOR2_X1 U9185 ( .A1(n8891), .A2(n8015), .ZN(n8016) );
  AOI211_X1 U9186 ( .C1(n8896), .C2(n8018), .A(n8017), .B(n8016), .ZN(n8019)
         );
  INV_X1 U9187 ( .A(n8019), .ZN(P2_U3260) );
  NAND2_X1 U9188 ( .A1(n9169), .A2(n8032), .ZN(n8449) );
  AOI21_X1 U9189 ( .B1(n8855), .B2(n9169), .A(n8047), .ZN(n8022) );
  NAND2_X1 U9190 ( .A1(n9165), .A2(n8229), .ZN(n8527) );
  NAND2_X1 U9191 ( .A1(n8528), .A2(n8527), .ZN(n8621) );
  NAND2_X1 U9192 ( .A1(n8022), .A2(n8621), .ZN(n8230) );
  OAI21_X1 U9193 ( .B1(n8022), .B2(n8621), .A(n8230), .ZN(n8023) );
  INV_X1 U9194 ( .A(n8023), .ZN(n9167) );
  NOR2_X2 U9195 ( .A1(n9169), .A2(n8040), .ZN(n8043) );
  INV_X1 U9196 ( .A(n8043), .ZN(n8025) );
  INV_X1 U9197 ( .A(n9165), .ZN(n8028) );
  AOI211_X1 U9198 ( .C1(n9165), .C2(n8025), .A(n10639), .B(n9069), .ZN(n9164)
         );
  AOI22_X1 U9199 ( .A1(n10469), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8026), .B2(
        n10458), .ZN(n8027) );
  OAI21_X1 U9200 ( .B1(n8028), .B2(n9076), .A(n8027), .ZN(n8029) );
  AOI21_X1 U9201 ( .B1(n9164), .B2(n8985), .A(n8029), .ZN(n8034) );
  INV_X1 U9202 ( .A(n8449), .ZN(n8030) );
  INV_X1 U9203 ( .A(n8452), .ZN(n8035) );
  XNOR2_X1 U9204 ( .A(n8232), .B(n8621), .ZN(n8031) );
  OAI222_X1 U9205 ( .A1(n10441), .A2(n8234), .B1(n10439), .B2(n8032), .C1(
        n10437), .C2(n8031), .ZN(n9163) );
  NAND2_X1 U9206 ( .A1(n9163), .A2(n4833), .ZN(n8033) );
  OAI211_X1 U9207 ( .C1(n9167), .C2(n9089), .A(n8034), .B(n8033), .ZN(P2_U3279) );
  OAI21_X1 U9208 ( .B1(n8036), .B2(n8035), .A(n8451), .ZN(n8037) );
  XOR2_X1 U9209 ( .A(n8620), .B(n8037), .Z(n8039) );
  AOI21_X1 U9210 ( .B1(n8039), .B2(n9085), .A(n8038), .ZN(n9171) );
  NAND2_X1 U9211 ( .A1(n9169), .A2(n8040), .ZN(n8041) );
  NAND2_X1 U9212 ( .A1(n8041), .A2(n10449), .ZN(n8042) );
  NOR2_X1 U9213 ( .A1(n8043), .A2(n8042), .ZN(n9168) );
  NAND2_X1 U9214 ( .A1(n9169), .A2(n10466), .ZN(n8045) );
  NAND2_X1 U9215 ( .A1(n10469), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8044) );
  OAI211_X1 U9216 ( .C1(n10373), .C2(n8046), .A(n8045), .B(n8044), .ZN(n8051)
         );
  AOI21_X1 U9217 ( .B1(n8620), .B2(n8048), .A(n8047), .ZN(n8049) );
  INV_X1 U9218 ( .A(n8049), .ZN(n9172) );
  NOR2_X1 U9219 ( .A1(n9172), .A2(n9089), .ZN(n8050) );
  AOI211_X1 U9220 ( .C1(n9168), .C2(n8985), .A(n8051), .B(n8050), .ZN(n8052)
         );
  OAI21_X1 U9221 ( .B1(n10469), .B2(n9171), .A(n8052), .ZN(P2_U3280) );
  INV_X1 U9222 ( .A(n8664), .ZN(n8053) );
  OAI222_X1 U9223 ( .A1(n8781), .A2(n8054), .B1(n7619), .B2(n8053), .C1(n8902), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  OR2_X1 U9224 ( .A1(n9434), .A2(n9550), .ZN(n8055) );
  NAND2_X1 U9225 ( .A1(n8057), .A2(n6944), .ZN(n8060) );
  AOI22_X1 U9226 ( .A1(n8280), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6704), .B2(
        n8058), .ZN(n8059) );
  OR2_X1 U9227 ( .A1(n9858), .A2(n8094), .ZN(n9445) );
  NAND2_X1 U9228 ( .A1(n9858), .A2(n8094), .ZN(n9444) );
  NAND2_X1 U9229 ( .A1(n9858), .A2(n9549), .ZN(n8061) );
  NAND2_X1 U9230 ( .A1(n8062), .A2(n6944), .ZN(n8065) );
  AOI22_X1 U9231 ( .A1(n8280), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6704), .B2(
        n8063), .ZN(n8064) );
  AOI22_X1 U9232 ( .A1(n6800), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n4874), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n8071) );
  INV_X1 U9233 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8066) );
  NAND2_X1 U9234 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U9235 ( .A1(n8078), .A2(n8068), .ZN(n8114) );
  OR2_X1 U9236 ( .A1(n8672), .A2(n8114), .ZN(n8070) );
  NAND2_X1 U9237 ( .A1(n6801), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U9238 ( .A1(n9855), .A2(n9744), .ZN(n9388) );
  NAND2_X1 U9239 ( .A1(n9389), .A2(n9388), .ZN(n9390) );
  XNOR2_X1 U9240 ( .A(n8272), .B(n9390), .ZN(n9857) );
  INV_X1 U9241 ( .A(n8214), .ZN(n8072) );
  INV_X1 U9242 ( .A(n9855), .ZN(n8119) );
  AOI211_X1 U9243 ( .C1(n9855), .C2(n8072), .A(n10565), .B(n9749), .ZN(n9854)
         );
  NOR2_X1 U9244 ( .A1(n8119), .A2(n10538), .ZN(n8075) );
  INV_X1 U9245 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8073) );
  OAI22_X1 U9246 ( .A1(n10539), .A2(n8073), .B1(n8114), .B2(n10488), .ZN(n8074) );
  AOI211_X1 U9247 ( .C1(n9854), .C2(n8076), .A(n8075), .B(n8074), .ZN(n8088)
         );
  NAND2_X1 U9248 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  AND2_X1 U9249 ( .A1(n8177), .A2(n8079), .ZN(n9753) );
  NAND2_X1 U9250 ( .A1(n9753), .A2(n6823), .ZN(n8082) );
  AOI22_X1 U9251 ( .A1(n6801), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n4874), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U9252 ( .A1(n6800), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8080) );
  INV_X1 U9253 ( .A(n9443), .ZN(n9367) );
  XNOR2_X1 U9254 ( .A(n8381), .B(n9390), .ZN(n8086) );
  OAI222_X1 U9255 ( .A1(n9745), .A2(n9271), .B1(n8086), .B2(n10518), .C1(n9743), .C2(n8094), .ZN(n9853) );
  NAND2_X1 U9256 ( .A1(n9853), .A2(n10539), .ZN(n8087) );
  OAI211_X1 U9257 ( .C1(n9857), .C2(n9718), .A(n8088), .B(n8087), .ZN(P1_U3275) );
  NAND2_X1 U9258 ( .A1(n9858), .A2(n4856), .ZN(n8090) );
  NAND2_X1 U9259 ( .A1(n9549), .A2(n8752), .ZN(n8089) );
  NAND2_X1 U9260 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  XNOR2_X1 U9261 ( .A(n8091), .B(n4854), .ZN(n8106) );
  INV_X1 U9262 ( .A(n9858), .ZN(n8218) );
  OAI22_X1 U9263 ( .A1(n8218), .A2(n8763), .B1(n8094), .B2(n8760), .ZN(n8122)
         );
  NAND2_X1 U9264 ( .A1(n8120), .A2(n8122), .ZN(n8109) );
  NAND2_X1 U9265 ( .A1(n9855), .A2(n4856), .ZN(n8096) );
  INV_X1 U9266 ( .A(n9744), .ZN(n9548) );
  NAND2_X1 U9267 ( .A1(n9548), .A2(n8752), .ZN(n8095) );
  NAND2_X1 U9268 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  XNOR2_X1 U9269 ( .A(n8097), .B(n4854), .ZN(n8099) );
  NOR2_X1 U9270 ( .A1(n9744), .A2(n8760), .ZN(n8098) );
  AOI21_X1 U9271 ( .B1(n9855), .B2(n8752), .A(n8098), .ZN(n8100) );
  NAND2_X1 U9272 ( .A1(n8099), .A2(n8100), .ZN(n8174) );
  INV_X1 U9273 ( .A(n8099), .ZN(n8102) );
  INV_X1 U9274 ( .A(n8100), .ZN(n8101) );
  NAND2_X1 U9275 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  AND2_X1 U9276 ( .A1(n8174), .A2(n8103), .ZN(n8110) );
  INV_X1 U9277 ( .A(n8104), .ZN(n8108) );
  INV_X1 U9278 ( .A(n8106), .ZN(n8107) );
  INV_X1 U9279 ( .A(n8172), .ZN(n8112) );
  OAI21_X1 U9280 ( .B1(n8112), .B2(n8111), .A(n4834), .ZN(n8118) );
  OAI21_X1 U9281 ( .B1(n9242), .B2(n9271), .A(n8113), .ZN(n8116) );
  NOR2_X1 U9282 ( .A1(n9274), .A2(n8114), .ZN(n8115) );
  AOI211_X1 U9283 ( .C1(n9250), .C2(n9549), .A(n8116), .B(n8115), .ZN(n8117)
         );
  OAI211_X1 U9284 ( .C1(n8119), .C2(n9224), .A(n8118), .B(n8117), .ZN(P1_U3224) );
  XOR2_X1 U9285 ( .A(n8122), .B(n8121), .Z(n8128) );
  NAND2_X1 U9286 ( .A1(n9262), .A2(n9548), .ZN(n8124) );
  OAI211_X1 U9287 ( .C1(n9430), .C2(n9284), .A(n8124), .B(n8123), .ZN(n8126)
         );
  NOR2_X1 U9288 ( .A1(n8218), .A2(n9224), .ZN(n8125) );
  AOI211_X1 U9289 ( .C1(n8216), .C2(n9280), .A(n8126), .B(n8125), .ZN(n8127)
         );
  OAI21_X1 U9290 ( .B1(n8128), .B2(n9289), .A(n8127), .ZN(P1_U3239) );
  XNOR2_X1 U9291 ( .A(n5310), .B(n8129), .ZN(n8130) );
  XNOR2_X1 U9292 ( .A(n8131), .B(n8130), .ZN(n8136) );
  INV_X1 U9293 ( .A(n9050), .ZN(n8235) );
  NAND2_X1 U9294 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8892) );
  OAI21_X1 U9295 ( .B1(n10394), .B2(n8235), .A(n8892), .ZN(n8134) );
  INV_X1 U9296 ( .A(n8132), .ZN(n8236) );
  OAI22_X1 U9297 ( .A1(n10393), .A2(n8234), .B1(n8848), .B2(n8236), .ZN(n8133)
         );
  AOI211_X1 U9298 ( .C1(n9155), .C2(n8851), .A(n8134), .B(n8133), .ZN(n8135)
         );
  OAI21_X1 U9299 ( .B1(n8136), .B2(n10397), .A(n8135), .ZN(P2_U3221) );
  INV_X1 U9300 ( .A(n9158), .ZN(n9077) );
  INV_X1 U9301 ( .A(n8137), .ZN(n8143) );
  INV_X1 U9302 ( .A(n8138), .ZN(n8140) );
  NOR2_X1 U9303 ( .A1(n8140), .A2(n8139), .ZN(n8142) );
  NAND2_X1 U9304 ( .A1(n8143), .A2(n8142), .ZN(n8141) );
  OAI211_X1 U9305 ( .C1(n8143), .C2(n8142), .A(n8141), .B(n8844), .ZN(n8146)
         );
  NOR2_X1 U9306 ( .A1(n10134), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8870) );
  OAI22_X1 U9307 ( .A1(n10393), .A2(n8229), .B1(n8848), .B2(n9073), .ZN(n8144)
         );
  AOI211_X1 U9308 ( .C1(n8802), .C2(n9083), .A(n8870), .B(n8144), .ZN(n8145)
         );
  OAI211_X1 U9309 ( .C1(n9077), .C2(n10399), .A(n8146), .B(n8145), .ZN(
        P2_U3240) );
  INV_X1 U9310 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U9311 ( .A1(n8778), .A2(n8147), .ZN(n8149) );
  OAI211_X1 U9312 ( .C1(n8775), .C2(n8645), .A(n8149), .B(n8148), .ZN(P1_U3325) );
  NAND2_X1 U9313 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8185) );
  INV_X1 U9314 ( .A(n8185), .ZN(n8154) );
  AOI211_X1 U9315 ( .C1(n8152), .C2(n8151), .A(n8150), .B(n10236), .ZN(n8153)
         );
  AOI211_X1 U9316 ( .C1(n10257), .C2(n8162), .A(n8154), .B(n8153), .ZN(n8160)
         );
  AOI211_X1 U9317 ( .C1(n8157), .C2(n8156), .A(n8155), .B(n10321), .ZN(n8158)
         );
  AOI21_X1 U9318 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n10259), .A(n8158), .ZN(
        n8159) );
  NAND2_X1 U9319 ( .A1(n8160), .A2(n8159), .ZN(P1_U3258) );
  NAND2_X1 U9320 ( .A1(n8161), .A2(n6944), .ZN(n8164) );
  AOI22_X1 U9321 ( .A1(n8280), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6704), .B2(
        n8162), .ZN(n8163) );
  INV_X1 U9322 ( .A(n9848), .ZN(n9755) );
  NAND2_X1 U9323 ( .A1(n9848), .A2(n4856), .ZN(n8166) );
  OR2_X1 U9324 ( .A1(n9271), .A2(n8763), .ZN(n8165) );
  NAND2_X1 U9325 ( .A1(n8166), .A2(n8165), .ZN(n8167) );
  XNOR2_X1 U9326 ( .A(n8167), .B(n4854), .ZN(n8170) );
  NOR2_X1 U9327 ( .A1(n9271), .A2(n8760), .ZN(n8168) );
  AOI21_X1 U9328 ( .B1(n9848), .B2(n8752), .A(n8168), .ZN(n8169) );
  NAND2_X1 U9329 ( .A1(n8170), .A2(n8169), .ZN(n8702) );
  OR2_X1 U9330 ( .A1(n8170), .A2(n8169), .ZN(n8171) );
  NAND2_X1 U9331 ( .A1(n8702), .A2(n8171), .ZN(n8173) );
  AND3_X1 U9332 ( .A1(n8172), .A2(n8174), .A3(n8173), .ZN(n8175) );
  OAI21_X1 U9333 ( .B1(n8704), .B2(n8175), .A(n4834), .ZN(n8189) );
  INV_X1 U9334 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8176) );
  NAND2_X1 U9335 ( .A1(n8177), .A2(n8176), .ZN(n8178) );
  NAND2_X1 U9336 ( .A1(n8284), .A2(n8178), .ZN(n9733) );
  OR2_X1 U9337 ( .A1(n9733), .A2(n8672), .ZN(n8184) );
  NAND2_X1 U9338 ( .A1(n4874), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U9339 ( .A1(n6801), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8179) );
  OAI211_X1 U9340 ( .C1(n8181), .C2(n8676), .A(n8180), .B(n8179), .ZN(n8182)
         );
  INV_X1 U9341 ( .A(n8182), .ZN(n8183) );
  NAND2_X1 U9342 ( .A1(n9250), .A2(n9548), .ZN(n8186) );
  OAI211_X1 U9343 ( .C1(n9242), .C2(n9746), .A(n8186), .B(n8185), .ZN(n8187)
         );
  AOI21_X1 U9344 ( .B1(n9280), .B2(n9753), .A(n8187), .ZN(n8188) );
  OAI211_X1 U9345 ( .C1(n9755), .C2(n9224), .A(n8189), .B(n8188), .ZN(P1_U3226) );
  AOI21_X1 U9346 ( .B1(n8195), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8190), .ZN(
        n8193) );
  NAND2_X1 U9347 ( .A1(n8875), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8191) );
  OAI21_X1 U9348 ( .B1(n8875), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8191), .ZN(
        n8192) );
  NOR2_X1 U9349 ( .A1(n8193), .A2(n8192), .ZN(n8874) );
  AOI211_X1 U9350 ( .C1(n8193), .C2(n8192), .A(n10301), .B(n8874), .ZN(n8205)
         );
  INV_X1 U9351 ( .A(n8194), .ZN(n8197) );
  OAI22_X1 U9352 ( .A1(n8197), .A2(n8196), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n8195), .ZN(n8199) );
  XNOR2_X1 U9353 ( .A(n8875), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8198) );
  NOR2_X1 U9354 ( .A1(n8199), .A2(n8198), .ZN(n8864) );
  AOI211_X1 U9355 ( .C1(n8199), .C2(n8198), .A(n10297), .B(n8864), .ZN(n8204)
         );
  INV_X1 U9356 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U9357 ( .A1(n10308), .A2(n8875), .ZN(n8201) );
  OAI211_X1 U9358 ( .C1(n8202), .C2(n8893), .A(n8201), .B(n8200), .ZN(n8203)
         );
  OR3_X1 U9359 ( .A1(n8205), .A2(n8204), .A3(n8203), .ZN(P2_U3262) );
  INV_X1 U9360 ( .A(n8206), .ZN(n8207) );
  AOI21_X1 U9361 ( .B1(n9443), .B2(n8208), .A(n8207), .ZN(n8219) );
  NAND2_X1 U9362 ( .A1(n8209), .A2(n9367), .ZN(n8210) );
  AOI21_X1 U9363 ( .B1(n8211), .B2(n8210), .A(n10518), .ZN(n8213) );
  OAI22_X1 U9364 ( .A1(n9743), .A2(n9430), .B1(n9744), .B2(n9745), .ZN(n8212)
         );
  AOI211_X1 U9365 ( .C1(n8219), .C2(n9764), .A(n8213), .B(n8212), .ZN(n9861)
         );
  AOI21_X1 U9366 ( .B1(n9858), .B2(n8215), .A(n8214), .ZN(n9859) );
  AOI22_X1 U9367 ( .A1(n10498), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8216), .B2(
        n10544), .ZN(n8217) );
  OAI21_X1 U9368 ( .B1(n8218), .B2(n10538), .A(n8217), .ZN(n8221) );
  INV_X1 U9369 ( .A(n8219), .ZN(n9862) );
  NOR2_X1 U9370 ( .A1(n9862), .A2(n9757), .ZN(n8220) );
  AOI211_X1 U9371 ( .C1(n9859), .C2(n10534), .A(n8221), .B(n8220), .ZN(n8222)
         );
  OAI21_X1 U9372 ( .B1(n10498), .B2(n9861), .A(n8222), .ZN(P1_U3276) );
  INV_X1 U9373 ( .A(n8225), .ZN(n8226) );
  MUX2_X1 U9374 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n8257), .Z(n8245) );
  INV_X1 U9375 ( .A(SI_29_), .ZN(n10055) );
  XNOR2_X1 U9376 ( .A(n8245), .B(n10055), .ZN(n8243) );
  INV_X1 U9377 ( .A(n8668), .ZN(n8242) );
  AOI22_X1 U9378 ( .A1(n8227), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8410), .ZN(n8228) );
  OAI21_X1 U9379 ( .B1(n8242), .B2(n7619), .A(n8228), .ZN(P2_U3329) );
  INV_X1 U9380 ( .A(n8229), .ZN(n9081) );
  NAND2_X1 U9381 ( .A1(n9158), .A2(n8234), .ZN(n8448) );
  NAND2_X1 U9382 ( .A1(n8447), .A2(n8448), .ZN(n9078) );
  NAND2_X1 U9383 ( .A1(n9155), .A2(n8913), .ZN(n8536) );
  NAND2_X1 U9384 ( .A1(n8535), .A2(n8536), .ZN(n8624) );
  OAI21_X1 U9385 ( .B1(n8231), .B2(n8624), .A(n8915), .ZN(n9157) );
  AOI22_X1 U9386 ( .A1(n9155), .A2(n10466), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n10469), .ZN(n8240) );
  INV_X1 U9387 ( .A(n9078), .ZN(n9067) );
  XNOR2_X1 U9388 ( .A(n8413), .B(n8624), .ZN(n8233) );
  OAI222_X1 U9389 ( .A1(n10441), .A2(n8235), .B1(n10439), .B2(n8234), .C1(
        n10437), .C2(n8233), .ZN(n9153) );
  AOI211_X1 U9390 ( .C1(n9155), .C2(n9070), .A(n10639), .B(n4921), .ZN(n9154)
         );
  INV_X1 U9391 ( .A(n9154), .ZN(n8237) );
  OAI22_X1 U9392 ( .A1(n8237), .A2(n8973), .B1(n10373), .B2(n8236), .ZN(n8238)
         );
  OAI21_X1 U9393 ( .B1(n9153), .B2(n8238), .A(n4833), .ZN(n8239) );
  OAI211_X1 U9394 ( .C1(n9157), .C2(n9089), .A(n8240), .B(n8239), .ZN(P2_U3277) );
  INV_X1 U9395 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8669) );
  OAI222_X1 U9396 ( .A1(n8777), .A2(n8242), .B1(P1_U3084), .B2(n8241), .C1(
        n8669), .C2(n8775), .ZN(P1_U3324) );
  INV_X1 U9397 ( .A(n8245), .ZN(n8246) );
  NAND2_X1 U9398 ( .A1(n8246), .A2(n10055), .ZN(n8247) );
  MUX2_X1 U9399 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n8257), .Z(n8253) );
  INV_X1 U9400 ( .A(SI_30_), .ZN(n10056) );
  XNOR2_X1 U9401 ( .A(n8253), .B(n10056), .ZN(n8251) );
  INV_X1 U9402 ( .A(n9339), .ZN(n8776) );
  AOI22_X1 U9403 ( .A1(n8249), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8410), .ZN(n8250) );
  OAI21_X1 U9404 ( .B1(n8776), .B2(n7619), .A(n8250), .ZN(P2_U3328) );
  NAND2_X1 U9405 ( .A1(n8252), .A2(n8251), .ZN(n8256) );
  INV_X1 U9406 ( .A(n8253), .ZN(n8254) );
  NAND2_X1 U9407 ( .A1(n8254), .A2(n10056), .ZN(n8255) );
  MUX2_X1 U9408 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n8257), .Z(n8259) );
  INV_X1 U9409 ( .A(SI_31_), .ZN(n8258) );
  XNOR2_X1 U9410 ( .A(n8259), .B(n8258), .ZN(n8260) );
  INV_X1 U9411 ( .A(n9344), .ZN(n8271) );
  NOR4_X1 U9412 ( .A1(n8263), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8262), .A4(
        P2_U3152), .ZN(n8264) );
  AOI21_X1 U9413 ( .B1(n8410), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8264), .ZN(
        n8265) );
  OAI21_X1 U9414 ( .B1(n8271), .B2(n7619), .A(n8265), .ZN(P2_U3327) );
  NAND3_X1 U9415 ( .A1(n8266), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n8267) );
  OAI22_X1 U9416 ( .A1(n8268), .A2(n8267), .B1(n6589), .B2(n8775), .ZN(n8269)
         );
  INV_X1 U9417 ( .A(n8269), .ZN(n8270) );
  OAI21_X1 U9418 ( .B1(n8271), .B2(n8777), .A(n8270), .ZN(P1_U3322) );
  NAND2_X1 U9419 ( .A1(n9855), .A2(n9548), .ZN(n8273) );
  NAND2_X1 U9420 ( .A1(n9848), .A2(n9271), .ZN(n9451) );
  INV_X1 U9421 ( .A(n9271), .ZN(n9722) );
  OR2_X1 U9422 ( .A1(n9848), .A2(n9722), .ZN(n8274) );
  NAND2_X1 U9423 ( .A1(n8275), .A2(n6944), .ZN(n8277) );
  AOI22_X1 U9424 ( .A1(n8280), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10250), 
        .B2(n6704), .ZN(n8276) );
  OR2_X1 U9425 ( .A1(n9843), .A2(n9746), .ZN(n9386) );
  NAND2_X1 U9426 ( .A1(n9843), .A2(n9746), .ZN(n9387) );
  NAND2_X1 U9427 ( .A1(n9386), .A2(n9387), .ZN(n9720) );
  NAND2_X1 U9428 ( .A1(n9721), .A2(n9720), .ZN(n9719) );
  INV_X1 U9429 ( .A(n9746), .ZN(n9712) );
  NAND2_X1 U9430 ( .A1(n9843), .A2(n9712), .ZN(n8278) );
  NAND2_X1 U9431 ( .A1(n8279), .A2(n6944), .ZN(n8282) );
  AOI22_X1 U9432 ( .A1(n8280), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10493), 
        .B2(n6704), .ZN(n8281) );
  INV_X1 U9433 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U9434 ( .A1(n8284), .A2(n8283), .ZN(n8285) );
  NAND2_X1 U9435 ( .A1(n8297), .A2(n8285), .ZN(n9708) );
  OR2_X1 U9436 ( .A1(n9708), .A2(n8672), .ZN(n8290) );
  NAND2_X1 U9437 ( .A1(n6800), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U9438 ( .A1(n4874), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8286) );
  OAI211_X1 U9439 ( .C1(n5173), .C2(n6354), .A(n8287), .B(n8286), .ZN(n8288)
         );
  INV_X1 U9440 ( .A(n8288), .ZN(n8289) );
  NAND2_X1 U9441 ( .A1(n8290), .A2(n8289), .ZN(n9723) );
  AND2_X1 U9442 ( .A1(n9837), .A2(n9723), .ZN(n8291) );
  NAND2_X1 U9443 ( .A1(n8292), .A2(n6944), .ZN(n8295) );
  OR2_X1 U9444 ( .A1(n9345), .A2(n8293), .ZN(n8294) );
  NAND2_X1 U9445 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U9446 ( .A1(n8309), .A2(n8298), .ZN(n9698) );
  OR2_X1 U9447 ( .A1(n9698), .A2(n8672), .ZN(n8304) );
  INV_X1 U9448 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U9449 ( .A1(n4874), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U9450 ( .A1(n6801), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8299) );
  OAI211_X1 U9451 ( .C1(n8676), .C2(n8301), .A(n8300), .B(n8299), .ZN(n8302)
         );
  INV_X1 U9452 ( .A(n8302), .ZN(n8303) );
  NAND2_X1 U9453 ( .A1(n8304), .A2(n8303), .ZN(n9713) );
  NAND2_X1 U9454 ( .A1(n8305), .A2(n6944), .ZN(n8307) );
  OR2_X1 U9455 ( .A1(n9345), .A2(n7463), .ZN(n8306) );
  NAND2_X1 U9456 ( .A1(n8309), .A2(n8308), .ZN(n8310) );
  AND2_X1 U9457 ( .A1(n8321), .A2(n8310), .ZN(n9684) );
  INV_X1 U9458 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U9459 ( .A1(n6801), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U9460 ( .A1(n4874), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8311) );
  OAI211_X1 U9461 ( .C1(n8676), .C2(n8313), .A(n8312), .B(n8311), .ZN(n8314)
         );
  AOI21_X1 U9462 ( .B1(n9684), .B2(n6823), .A(n8314), .ZN(n9260) );
  OR2_X1 U9463 ( .A1(n9828), .A2(n9260), .ZN(n9297) );
  NAND2_X1 U9464 ( .A1(n9828), .A2(n9260), .ZN(n9381) );
  NAND2_X1 U9465 ( .A1(n9297), .A2(n9381), .ZN(n9678) );
  INV_X1 U9466 ( .A(n9260), .ZN(n9693) );
  NAND2_X1 U9467 ( .A1(n9828), .A2(n9693), .ZN(n8315) );
  NAND2_X1 U9468 ( .A1(n8316), .A2(n8315), .ZN(n9661) );
  NAND2_X1 U9469 ( .A1(n8317), .A2(n6944), .ZN(n8320) );
  OR2_X1 U9470 ( .A1(n9345), .A2(n8318), .ZN(n8319) );
  INV_X1 U9471 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U9472 ( .A1(n8321), .A2(n9259), .ZN(n8322) );
  NAND2_X1 U9473 ( .A1(n8323), .A2(n8322), .ZN(n9663) );
  OR2_X1 U9474 ( .A1(n9663), .A2(n8672), .ZN(n8329) );
  INV_X1 U9475 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U9476 ( .A1(n4874), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U9477 ( .A1(n6801), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8324) );
  OAI211_X1 U9478 ( .C1(n8326), .C2(n8676), .A(n8325), .B(n8324), .ZN(n8327)
         );
  INV_X1 U9479 ( .A(n8327), .ZN(n8328) );
  NAND2_X1 U9480 ( .A1(n8329), .A2(n8328), .ZN(n9653) );
  OR2_X1 U9481 ( .A1(n9821), .A2(n9653), .ZN(n8330) );
  NAND2_X1 U9482 ( .A1(n9821), .A2(n9653), .ZN(n8331) );
  NAND2_X1 U9483 ( .A1(n8332), .A2(n6944), .ZN(n8335) );
  OR2_X1 U9484 ( .A1(n9345), .A2(n8333), .ZN(n8334) );
  NAND2_X1 U9485 ( .A1(n9816), .A2(n9239), .ZN(n9378) );
  NAND2_X1 U9486 ( .A1(n9648), .A2(n9239), .ZN(n9623) );
  NAND2_X1 U9487 ( .A1(n8336), .A2(n6944), .ZN(n8339) );
  OR2_X1 U9488 ( .A1(n9345), .A2(n8337), .ZN(n8338) );
  INV_X1 U9489 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U9490 ( .A1(n8340), .A2(n9238), .ZN(n8341) );
  AND2_X1 U9491 ( .A1(n8355), .A2(n8341), .ZN(n9634) );
  NAND2_X1 U9492 ( .A1(n9634), .A2(n6823), .ZN(n8347) );
  INV_X1 U9493 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8344) );
  NAND2_X1 U9494 ( .A1(n4874), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U9495 ( .A1(n6801), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8342) );
  OAI211_X1 U9496 ( .C1(n8676), .C2(n8344), .A(n8343), .B(n8342), .ZN(n8345)
         );
  INV_X1 U9497 ( .A(n8345), .ZN(n8346) );
  NAND2_X1 U9498 ( .A1(n8347), .A2(n8346), .ZN(n9654) );
  OR2_X1 U9499 ( .A1(n9812), .A2(n9654), .ZN(n8348) );
  AND2_X1 U9500 ( .A1(n9623), .A2(n8348), .ZN(n9605) );
  NAND2_X1 U9501 ( .A1(n8349), .A2(n6944), .ZN(n8352) );
  OR2_X1 U9502 ( .A1(n9345), .A2(n8350), .ZN(n8351) );
  INV_X1 U9503 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U9504 ( .A1(n8355), .A2(n8354), .ZN(n8356) );
  NAND2_X1 U9505 ( .A1(n8372), .A2(n8356), .ZN(n9230) );
  INV_X1 U9506 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U9507 ( .A1(n4874), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U9508 ( .A1(n6801), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8357) );
  OAI211_X1 U9509 ( .C1(n8676), .C2(n8359), .A(n8358), .B(n8357), .ZN(n8360)
         );
  INV_X1 U9510 ( .A(n8360), .ZN(n8361) );
  OR2_X1 U9511 ( .A1(n9806), .A2(n9631), .ZN(n8363) );
  AND2_X1 U9512 ( .A1(n9605), .A2(n8363), .ZN(n8660) );
  INV_X1 U9513 ( .A(n8363), .ZN(n8365) );
  OR2_X1 U9514 ( .A1(n9806), .A2(n9285), .ZN(n9472) );
  NAND2_X1 U9515 ( .A1(n9806), .A2(n9285), .ZN(n9471) );
  NAND2_X1 U9516 ( .A1(n9472), .A2(n9471), .ZN(n8393) );
  NAND2_X1 U9517 ( .A1(n9812), .A2(n9654), .ZN(n9606) );
  AND2_X1 U9518 ( .A1(n8393), .A2(n9606), .ZN(n8364) );
  INV_X1 U9519 ( .A(n8662), .ZN(n8366) );
  OR2_X1 U9520 ( .A1(n9345), .A2(n8368), .ZN(n8369) );
  INV_X1 U9521 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U9522 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  NAND2_X1 U9523 ( .A1(n9281), .A2(n6823), .ZN(n8379) );
  INV_X1 U9524 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U9525 ( .A1(n6801), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U9526 ( .A1(n4874), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8374) );
  OAI211_X1 U9527 ( .C1(n8676), .C2(n8376), .A(n8375), .B(n8374), .ZN(n8377)
         );
  INV_X1 U9528 ( .A(n8377), .ZN(n8378) );
  INV_X1 U9529 ( .A(n9618), .ZN(n9597) );
  NAND2_X1 U9530 ( .A1(n9801), .A2(n9597), .ZN(n9376) );
  NAND2_X1 U9531 ( .A1(n8382), .A2(n9388), .ZN(n9741) );
  OR2_X1 U9532 ( .A1(n9742), .A2(n9720), .ZN(n8383) );
  OR2_X1 U9533 ( .A1(n9720), .A2(n9724), .ZN(n8384) );
  AND2_X2 U9534 ( .A1(n8385), .A2(n8384), .ZN(n9725) );
  INV_X1 U9535 ( .A(n9724), .ZN(n8386) );
  NAND2_X1 U9536 ( .A1(n9387), .A2(n8386), .ZN(n8387) );
  AND2_X1 U9537 ( .A1(n8387), .A2(n9386), .ZN(n9300) );
  INV_X1 U9538 ( .A(n9723), .ZN(n8388) );
  OR2_X1 U9539 ( .A1(n9837), .A2(n8388), .ZN(n9457) );
  NAND2_X1 U9540 ( .A1(n9837), .A2(n8388), .ZN(n9458) );
  NAND2_X1 U9541 ( .A1(n9457), .A2(n9458), .ZN(n9705) );
  INV_X1 U9542 ( .A(n9713), .ZN(n9680) );
  OR2_X1 U9543 ( .A1(n9833), .A2(n9680), .ZN(n9676) );
  NAND2_X1 U9544 ( .A1(n9833), .A2(n9680), .ZN(n9295) );
  AND2_X1 U9545 ( .A1(n9297), .A2(n9676), .ZN(n9383) );
  NAND2_X1 U9546 ( .A1(n9675), .A2(n9383), .ZN(n8389) );
  NAND2_X1 U9547 ( .A1(n8389), .A2(n9381), .ZN(n9668) );
  INV_X1 U9548 ( .A(n9653), .ZN(n9681) );
  OR2_X1 U9549 ( .A1(n9821), .A2(n9681), .ZN(n9462) );
  NAND2_X1 U9550 ( .A1(n9821), .A2(n9681), .ZN(n9463) );
  INV_X1 U9551 ( .A(n9651), .ZN(n9625) );
  INV_X1 U9552 ( .A(n9654), .ZN(n9305) );
  NAND2_X1 U9553 ( .A1(n9812), .A2(n9305), .ZN(n9467) );
  INV_X1 U9554 ( .A(n9467), .ZN(n8391) );
  OR2_X1 U9555 ( .A1(n9625), .A2(n8391), .ZN(n8390) );
  XNOR2_X1 U9556 ( .A(n9812), .B(n9654), .ZN(n9629) );
  AND2_X1 U9557 ( .A1(n9629), .A2(n9626), .ZN(n9627) );
  OR2_X1 U9558 ( .A1(n8391), .A2(n9627), .ZN(n8392) );
  NAND2_X1 U9559 ( .A1(n9616), .A2(n9617), .ZN(n9615) );
  NAND2_X1 U9560 ( .A1(n9615), .A2(n9471), .ZN(n8684) );
  XNOR2_X1 U9561 ( .A(n8684), .B(n9475), .ZN(n8394) );
  XNOR2_X1 U9562 ( .A(n8649), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9592) );
  NAND2_X1 U9563 ( .A1(n9592), .A2(n6823), .ZN(n8400) );
  INV_X1 U9564 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U9565 ( .A1(n6801), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U9566 ( .A1(n4874), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8395) );
  OAI211_X1 U9567 ( .C1(n8676), .C2(n8397), .A(n8396), .B(n8395), .ZN(n8398)
         );
  INV_X1 U9568 ( .A(n8398), .ZN(n8399) );
  OAI22_X1 U9569 ( .A1(n8771), .A2(n9745), .B1(n9285), .B2(n9743), .ZN(n8401)
         );
  INV_X1 U9570 ( .A(n9806), .ZN(n9614) );
  OR2_X2 U9571 ( .A1(n9828), .A2(n9690), .ZN(n9682) );
  NAND2_X1 U9572 ( .A1(n9648), .A2(n9662), .ZN(n9642) );
  NOR2_X2 U9573 ( .A1(n9812), .A2(n9642), .ZN(n9633) );
  AOI21_X1 U9574 ( .B1(n9801), .B2(n9609), .A(n5158), .ZN(n9802) );
  AOI22_X1 U9575 ( .A1(n9281), .A2(n10544), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n10498), .ZN(n8406) );
  OAI21_X1 U9576 ( .B1(n5161), .B2(n10538), .A(n8406), .ZN(n8408) );
  NOR2_X1 U9577 ( .A1(n9805), .A2(n9757), .ZN(n8407) );
  AOI211_X1 U9578 ( .C1(n9802), .C2(n10534), .A(n8408), .B(n8407), .ZN(n8409)
         );
  OAI21_X1 U9579 ( .B1(n9804), .B2(n10498), .A(n8409), .ZN(P1_U3265) );
  AOI22_X1 U9580 ( .A1(n8410), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n10292), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n8411) );
  OAI21_X1 U9581 ( .B1(n8412), .B2(n7619), .A(n8411), .ZN(P2_U3357) );
  OR2_X1 U9582 ( .A1(n9148), .A2(n9050), .ZN(n8541) );
  NAND2_X1 U9583 ( .A1(n9148), .A2(n9050), .ZN(n8916) );
  INV_X1 U9584 ( .A(n9062), .ZN(n8627) );
  AOI22_X1 U9585 ( .A1(n9055), .A2(n8627), .B1(n5141), .B2(n9050), .ZN(n9048)
         );
  INV_X1 U9586 ( .A(n9056), .ZN(n9034) );
  NAND2_X1 U9587 ( .A1(n9048), .A2(n8415), .ZN(n8416) );
  XNOR2_X1 U9588 ( .A(n9138), .B(n9049), .ZN(n8918) );
  INV_X1 U9589 ( .A(n9049), .ZN(n8551) );
  NAND2_X1 U9590 ( .A1(n9132), .A2(n9035), .ZN(n8442) );
  INV_X1 U9591 ( .A(n8442), .ZN(n8555) );
  NAND2_X1 U9592 ( .A1(n9005), .A2(n8813), .ZN(n8443) );
  NAND2_X1 U9593 ( .A1(n8563), .A2(n8443), .ZN(n8999) );
  INV_X1 U9594 ( .A(n8999), .ZN(n8993) );
  NAND2_X1 U9595 ( .A1(n9122), .A2(n8997), .ZN(n8561) );
  AND2_X1 U9596 ( .A1(n8596), .A2(n8966), .ZN(n8440) );
  NAND2_X1 U9597 ( .A1(n9117), .A2(n8957), .ZN(n8595) );
  INV_X1 U9598 ( .A(n8595), .ZN(n8567) );
  NAND2_X1 U9599 ( .A1(n9110), .A2(n8970), .ZN(n8572) );
  NAND2_X1 U9600 ( .A1(n9105), .A2(n8958), .ZN(n8577) );
  NAND2_X1 U9601 ( .A1(n8668), .A2(n5657), .ZN(n8418) );
  NAND2_X1 U9602 ( .A1(n4859), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8417) );
  NAND2_X1 U9603 ( .A1(n8929), .A2(n8419), .ZN(n8582) );
  INV_X1 U9604 ( .A(n8582), .ZN(n8420) );
  OAI21_X1 U9605 ( .B1(n8924), .B2(n8420), .A(n8581), .ZN(n8424) );
  INV_X1 U9606 ( .A(n8424), .ZN(n8426) );
  NAND2_X1 U9607 ( .A1(n9339), .A2(n5657), .ZN(n8422) );
  NAND2_X1 U9608 ( .A1(n4859), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8421) );
  NOR2_X1 U9609 ( .A1(n9094), .A2(n8926), .ZN(n8437) );
  OAI22_X1 U9610 ( .A1(n8424), .A2(n8437), .B1(n8423), .B2(n8588), .ZN(n8425)
         );
  OAI21_X1 U9611 ( .B1(n8426), .B2(n9094), .A(n8425), .ZN(n8431) );
  NAND2_X1 U9612 ( .A1(n9344), .A2(n5657), .ZN(n8429) );
  NAND2_X1 U9613 ( .A1(n5918), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8428) );
  INV_X1 U9614 ( .A(n8588), .ZN(n8904) );
  OR2_X1 U9615 ( .A1(n9090), .A2(n8904), .ZN(n8430) );
  NAND2_X1 U9616 ( .A1(n9094), .A2(n8926), .ZN(n8584) );
  AND2_X1 U9617 ( .A1(n9090), .A2(n8904), .ZN(n8436) );
  INV_X1 U9618 ( .A(n8435), .ZN(n8632) );
  INV_X1 U9619 ( .A(n8436), .ZN(n8438) );
  INV_X1 U9620 ( .A(n8437), .ZN(n8585) );
  NAND2_X1 U9621 ( .A1(n8438), .A2(n8585), .ZN(n8633) );
  AND2_X1 U9622 ( .A1(n8636), .A2(n8973), .ZN(n8439) );
  MUX2_X1 U9623 ( .A(n8632), .B(n8633), .S(n8587), .Z(n8592) );
  AND2_X1 U9624 ( .A1(n8595), .A2(n8561), .ZN(n8441) );
  MUX2_X1 U9625 ( .A(n8441), .B(n8440), .S(n8587), .Z(n8571) );
  NAND2_X1 U9626 ( .A1(n8563), .A2(n8552), .ZN(n8445) );
  NAND2_X1 U9627 ( .A1(n8443), .A2(n8442), .ZN(n8444) );
  MUX2_X1 U9628 ( .A(n8445), .B(n8444), .S(n8587), .Z(n8446) );
  INV_X1 U9629 ( .A(n8446), .ZN(n8560) );
  INV_X1 U9630 ( .A(n8624), .ZN(n8534) );
  MUX2_X1 U9631 ( .A(n8448), .B(n8447), .S(n8587), .Z(n8533) );
  INV_X1 U9632 ( .A(n8621), .ZN(n8526) );
  MUX2_X1 U9633 ( .A(n8450), .B(n8449), .S(n8587), .Z(n8525) );
  MUX2_X1 U9634 ( .A(n8452), .B(n8451), .S(n8587), .Z(n8523) );
  MUX2_X1 U9635 ( .A(n8454), .B(n8453), .S(n8580), .Z(n8521) );
  NAND2_X1 U9636 ( .A1(n8457), .A2(n8508), .ZN(n8455) );
  NAND2_X1 U9637 ( .A1(n8455), .A2(n8456), .ZN(n8460) );
  NAND2_X1 U9638 ( .A1(n8456), .A2(n8506), .ZN(n8458) );
  NAND2_X1 U9639 ( .A1(n8458), .A2(n8457), .ZN(n8459) );
  MUX2_X1 U9640 ( .A(n8460), .B(n8459), .S(n8587), .Z(n8514) );
  AND2_X1 U9641 ( .A1(n7081), .A2(n8597), .ZN(n8463) );
  NAND2_X1 U9642 ( .A1(n8463), .A2(n8636), .ZN(n8461) );
  NOR2_X1 U9643 ( .A1(n8461), .A2(n7356), .ZN(n8462) );
  NOR2_X1 U9644 ( .A1(n7227), .A2(n8462), .ZN(n8470) );
  INV_X1 U9645 ( .A(n8463), .ZN(n8465) );
  NAND2_X1 U9646 ( .A1(n8465), .A2(n8464), .ZN(n8467) );
  OAI21_X1 U9647 ( .B1(n8467), .B2(n7356), .A(n8466), .ZN(n8468) );
  INV_X1 U9648 ( .A(n8468), .ZN(n8469) );
  MUX2_X1 U9649 ( .A(n8470), .B(n8469), .S(n8580), .Z(n8476) );
  INV_X1 U9650 ( .A(n10438), .ZN(n8474) );
  MUX2_X1 U9651 ( .A(n8472), .B(n8471), .S(n8580), .Z(n8473) );
  OAI211_X1 U9652 ( .C1(n8476), .C2(n8475), .A(n8474), .B(n8473), .ZN(n8481)
         );
  NAND2_X1 U9653 ( .A1(n8477), .A2(n8580), .ZN(n8479) );
  NAND2_X1 U9654 ( .A1(n8860), .A2(n8587), .ZN(n8478) );
  MUX2_X1 U9655 ( .A(n8479), .B(n8478), .S(n10451), .Z(n8480) );
  NAND3_X1 U9656 ( .A1(n8481), .A2(n8601), .A3(n8480), .ZN(n8485) );
  MUX2_X1 U9657 ( .A(n8483), .B(n8482), .S(n8587), .Z(n8484) );
  NAND3_X1 U9658 ( .A1(n8485), .A2(n8606), .A3(n8484), .ZN(n8490) );
  INV_X1 U9659 ( .A(n8486), .ZN(n8488) );
  MUX2_X1 U9660 ( .A(n8488), .B(n8487), .S(n8587), .Z(n8489) );
  NAND3_X1 U9661 ( .A1(n8490), .A2(n8605), .A3(n8489), .ZN(n8494) );
  MUX2_X1 U9662 ( .A(n8492), .B(n8491), .S(n8587), .Z(n8493) );
  NAND3_X1 U9663 ( .A1(n8494), .A2(n8607), .A3(n8493), .ZN(n8499) );
  AND2_X1 U9664 ( .A1(n8500), .A2(n8495), .ZN(n8496) );
  MUX2_X1 U9665 ( .A(n8497), .B(n8496), .S(n8580), .Z(n8498) );
  NAND3_X1 U9666 ( .A1(n8499), .A2(n8502), .A3(n8498), .ZN(n8504) );
  AND2_X1 U9667 ( .A1(n8505), .A2(n8500), .ZN(n8501) );
  MUX2_X1 U9668 ( .A(n8502), .B(n8501), .S(n8587), .Z(n8503) );
  NAND3_X1 U9669 ( .A1(n8504), .A2(n8503), .A3(n8507), .ZN(n8512) );
  AND2_X1 U9670 ( .A1(n8506), .A2(n8505), .ZN(n8510) );
  AND2_X1 U9671 ( .A1(n8508), .A2(n8507), .ZN(n8509) );
  MUX2_X1 U9672 ( .A(n8510), .B(n8509), .S(n8587), .Z(n8511) );
  NAND3_X1 U9673 ( .A1(n8614), .A2(n8512), .A3(n8511), .ZN(n8513) );
  NAND3_X1 U9674 ( .A1(n8515), .A2(n8514), .A3(n8513), .ZN(n8519) );
  MUX2_X1 U9675 ( .A(n8517), .B(n8516), .S(n8587), .Z(n8518) );
  NAND3_X1 U9676 ( .A1(n8619), .A2(n8519), .A3(n8518), .ZN(n8520) );
  NAND3_X1 U9677 ( .A1(n8618), .A2(n8521), .A3(n8520), .ZN(n8522) );
  NAND3_X1 U9678 ( .A1(n8620), .A2(n8523), .A3(n8522), .ZN(n8524) );
  NAND3_X1 U9679 ( .A1(n8526), .A2(n8525), .A3(n8524), .ZN(n8530) );
  MUX2_X1 U9680 ( .A(n8528), .B(n8527), .S(n8580), .Z(n8529) );
  NAND2_X1 U9681 ( .A1(n8530), .A2(n8529), .ZN(n8531) );
  NAND2_X1 U9682 ( .A1(n9067), .A2(n8531), .ZN(n8532) );
  NAND3_X1 U9683 ( .A1(n8534), .A2(n8533), .A3(n8532), .ZN(n8538) );
  MUX2_X1 U9684 ( .A(n8536), .B(n8535), .S(n8580), .Z(n8537) );
  NAND2_X1 U9685 ( .A1(n8538), .A2(n8537), .ZN(n8543) );
  MUX2_X1 U9686 ( .A(n9050), .B(n9148), .S(n8580), .Z(n8539) );
  INV_X1 U9687 ( .A(n8539), .ZN(n8540) );
  OAI21_X1 U9688 ( .B1(n8543), .B2(n8541), .A(n8540), .ZN(n8545) );
  INV_X1 U9689 ( .A(n8916), .ZN(n8542) );
  NAND2_X1 U9690 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  NAND2_X1 U9691 ( .A1(n8545), .A2(n8544), .ZN(n8547) );
  NAND2_X1 U9692 ( .A1(n9143), .A2(n9056), .ZN(n8625) );
  INV_X1 U9693 ( .A(n8625), .ZN(n8546) );
  NAND2_X1 U9694 ( .A1(n8547), .A2(n8546), .ZN(n8550) );
  MUX2_X1 U9695 ( .A(n9056), .B(n9143), .S(n8580), .Z(n8549) );
  INV_X1 U9696 ( .A(n8547), .ZN(n8548) );
  INV_X1 U9697 ( .A(n8626), .ZN(n8917) );
  AOI22_X1 U9698 ( .A1(n8550), .A2(n8549), .B1(n8548), .B2(n8917), .ZN(n8558)
         );
  AND2_X1 U9699 ( .A1(n9138), .A2(n8551), .ZN(n8554) );
  MUX2_X1 U9700 ( .A(n8554), .B(n8553), .S(n8587), .Z(n8556) );
  NOR2_X1 U9701 ( .A1(n8556), .A2(n8555), .ZN(n8557) );
  OAI21_X1 U9702 ( .B1(n9033), .B2(n8558), .A(n8557), .ZN(n8559) );
  NAND2_X1 U9703 ( .A1(n8560), .A2(n8559), .ZN(n8562) );
  INV_X1 U9704 ( .A(n9005), .ZN(n9125) );
  AOI21_X1 U9705 ( .B1(n8562), .B2(n9125), .A(n8919), .ZN(n8566) );
  AND2_X1 U9706 ( .A1(n8561), .A2(n8587), .ZN(n8565) );
  OAI211_X1 U9707 ( .C1(n8587), .C2(n9013), .A(n8563), .B(n8562), .ZN(n8564)
         );
  OAI21_X1 U9708 ( .B1(n8566), .B2(n8565), .A(n8564), .ZN(n8570) );
  INV_X1 U9709 ( .A(n8596), .ZN(n8568) );
  MUX2_X1 U9710 ( .A(n8568), .B(n8567), .S(n8587), .Z(n8569) );
  AOI21_X1 U9711 ( .B1(n8571), .B2(n8570), .A(n8569), .ZN(n8575) );
  MUX2_X1 U9712 ( .A(n8573), .B(n8572), .S(n8587), .Z(n8574) );
  OAI211_X1 U9713 ( .C1(n8575), .C2(n8956), .A(n8936), .B(n8574), .ZN(n8579)
         );
  MUX2_X1 U9714 ( .A(n8577), .B(n8576), .S(n8587), .Z(n8578) );
  NAND3_X1 U9715 ( .A1(n8579), .A2(n8921), .A3(n8578), .ZN(n8586) );
  MUX2_X1 U9716 ( .A(n8582), .B(n8581), .S(n8580), .Z(n8583) );
  INV_X1 U9717 ( .A(n9090), .ZN(n8590) );
  MUX2_X1 U9718 ( .A(n9090), .B(n8588), .S(n8587), .Z(n8589) );
  OAI21_X1 U9719 ( .B1(n8590), .B2(n8904), .A(n8589), .ZN(n8591) );
  NOR3_X1 U9720 ( .A1(n8594), .A2(n8598), .A3(n10340), .ZN(n8639) );
  NOR2_X1 U9721 ( .A1(n7067), .A2(n7356), .ZN(n8603) );
  AND3_X1 U9722 ( .A1(n8599), .A2(n8598), .A3(n8597), .ZN(n8600) );
  NAND4_X1 U9723 ( .A1(n8603), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n8604)
         );
  NOR2_X1 U9724 ( .A1(n8604), .A2(n10438), .ZN(n8608) );
  NAND4_X1 U9725 ( .A1(n8608), .A2(n8607), .A3(n8606), .A4(n8605), .ZN(n8610)
         );
  NOR2_X1 U9726 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  NAND4_X1 U9727 ( .A1(n8614), .A2(n8613), .A3(n8612), .A4(n8611), .ZN(n8615)
         );
  NOR2_X1 U9728 ( .A1(n8616), .A2(n8615), .ZN(n8617) );
  NAND4_X1 U9729 ( .A1(n8620), .A2(n8619), .A3(n8618), .A4(n8617), .ZN(n8622)
         );
  OR3_X1 U9730 ( .A1(n8622), .A2(n9078), .A3(n8621), .ZN(n8623) );
  NOR2_X1 U9731 ( .A1(n8624), .A2(n8623), .ZN(n8628) );
  NAND2_X1 U9732 ( .A1(n8626), .A2(n8625), .ZN(n9047) );
  NAND4_X1 U9733 ( .A1(n9015), .A2(n8628), .A3(n9047), .A4(n8627), .ZN(n8629)
         );
  NOR4_X1 U9734 ( .A1(n8919), .A2(n8999), .A3(n9033), .A4(n8629), .ZN(n8630)
         );
  NAND4_X1 U9735 ( .A1(n8936), .A2(n8948), .A3(n8967), .A4(n8630), .ZN(n8631)
         );
  NOR4_X1 U9736 ( .A1(n8633), .A2(n8632), .A3(n8923), .A4(n8631), .ZN(n8634)
         );
  XNOR2_X1 U9737 ( .A(n8634), .B(n8973), .ZN(n8635) );
  AOI211_X1 U9738 ( .C1(n5610), .C2(n8637), .A(n8636), .B(n8635), .ZN(n8638)
         );
  NOR3_X1 U9739 ( .A1(n8640), .A2(n8902), .A3(n10439), .ZN(n8643) );
  OAI21_X1 U9740 ( .B1(n8644), .B2(n8641), .A(P2_B_REG_SCAN_IN), .ZN(n8642) );
  NAND2_X1 U9741 ( .A1(n8778), .A2(n6944), .ZN(n8647) );
  OR2_X1 U9742 ( .A1(n9345), .A2(n8645), .ZN(n8646) );
  INV_X1 U9743 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8648) );
  INV_X1 U9744 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8768) );
  OAI21_X1 U9745 ( .B1(n8649), .B2(n8648), .A(n8768), .ZN(n8652) );
  INV_X1 U9746 ( .A(n8649), .ZN(n8651) );
  AND2_X1 U9747 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n8650) );
  NAND2_X1 U9748 ( .A1(n8651), .A2(n8650), .ZN(n8680) );
  NAND2_X1 U9749 ( .A1(n8652), .A2(n8680), .ZN(n9584) );
  INV_X1 U9750 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U9751 ( .A1(n6801), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U9752 ( .A1(n4874), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8653) );
  OAI211_X1 U9753 ( .C1(n8676), .C2(n8655), .A(n8654), .B(n8653), .ZN(n8656)
         );
  INV_X1 U9754 ( .A(n8656), .ZN(n8657) );
  NOR2_X1 U9755 ( .A1(n9801), .A2(n9618), .ZN(n8663) );
  INV_X1 U9756 ( .A(n8663), .ZN(n8659) );
  AND2_X1 U9757 ( .A1(n8660), .A2(n8659), .ZN(n8661) );
  NAND2_X1 U9758 ( .A1(n8664), .A2(n6944), .ZN(n8667) );
  OR2_X1 U9759 ( .A1(n9345), .A2(n8665), .ZN(n8666) );
  NAND2_X1 U9760 ( .A1(n9796), .A2(n8771), .ZN(n9374) );
  NAND2_X1 U9761 ( .A1(n9790), .A2(n9598), .ZN(n9481) );
  NAND2_X1 U9762 ( .A1(n8668), .A2(n6944), .ZN(n8671) );
  OR2_X1 U9763 ( .A1(n9345), .A2(n8669), .ZN(n8670) );
  OR2_X1 U9764 ( .A1(n8680), .A2(n8672), .ZN(n8679) );
  INV_X1 U9765 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U9766 ( .A1(n4874), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U9767 ( .A1(n6801), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8673) );
  OAI211_X1 U9768 ( .C1(n8676), .C2(n8675), .A(n8674), .B(n8673), .ZN(n8677)
         );
  INV_X1 U9769 ( .A(n8677), .ZN(n8678) );
  NAND2_X1 U9770 ( .A1(n9785), .A2(n9578), .ZN(n9489) );
  INV_X1 U9771 ( .A(n9796), .ZN(n9594) );
  NOR2_X2 U9772 ( .A1(n9785), .A2(n9583), .ZN(n9563) );
  AOI21_X1 U9773 ( .B1(n9785), .B2(n9583), .A(n9563), .ZN(n9786) );
  INV_X1 U9774 ( .A(n9785), .ZN(n8683) );
  INV_X1 U9775 ( .A(n8680), .ZN(n8681) );
  AOI22_X1 U9776 ( .A1(n8681), .A2(n10544), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10498), .ZN(n8682) );
  OAI21_X1 U9777 ( .B1(n8683), .B2(n10538), .A(n8682), .ZN(n8695) );
  NAND2_X1 U9778 ( .A1(n8684), .A2(n9475), .ZN(n8685) );
  NAND2_X1 U9779 ( .A1(n8685), .A2(n9376), .ZN(n9596) );
  XOR2_X1 U9780 ( .A(n9352), .B(n8687), .Z(n8694) );
  NAND2_X1 U9781 ( .A1(n6800), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U9782 ( .A1(n6801), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U9783 ( .A1(n4874), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8688) );
  NAND3_X1 U9784 ( .A1(n8690), .A2(n8689), .A3(n8688), .ZN(n9546) );
  NOR2_X1 U9785 ( .A1(n10220), .A2(n9545), .ZN(n8691) );
  NOR2_X1 U9786 ( .A1(n9745), .A2(n8691), .ZN(n9559) );
  AOI22_X1 U9787 ( .A1(n9801), .A2(n8752), .B1(n8744), .B2(n9618), .ZN(n8751)
         );
  NAND2_X1 U9788 ( .A1(n9801), .A2(n4855), .ZN(n8697) );
  NAND2_X1 U9789 ( .A1(n9618), .A2(n8752), .ZN(n8696) );
  NAND2_X1 U9790 ( .A1(n8697), .A2(n8696), .ZN(n8698) );
  XNOR2_X1 U9791 ( .A(n8698), .B(n8761), .ZN(n8750) );
  AOI22_X1 U9792 ( .A1(n9821), .A2(n8752), .B1(n8744), .B2(n9653), .ZN(n8729)
         );
  NAND2_X1 U9793 ( .A1(n9821), .A2(n4855), .ZN(n8700) );
  NAND2_X1 U9794 ( .A1(n9653), .A2(n8752), .ZN(n8699) );
  NAND2_X1 U9795 ( .A1(n8700), .A2(n8699), .ZN(n8701) );
  XNOR2_X1 U9796 ( .A(n8701), .B(n8761), .ZN(n8727) );
  INV_X1 U9797 ( .A(n8727), .ZN(n8728) );
  INV_X1 U9798 ( .A(n8702), .ZN(n8703) );
  AOI22_X1 U9799 ( .A1(n9843), .A2(n4856), .B1(n8752), .B2(n9712), .ZN(n8705)
         );
  XOR2_X1 U9800 ( .A(n8761), .B(n8705), .Z(n8706) );
  AOI22_X1 U9801 ( .A1(n9843), .A2(n8752), .B1(n8744), .B2(n9712), .ZN(n9269)
         );
  NAND2_X1 U9802 ( .A1(n9837), .A2(n4855), .ZN(n8708) );
  NAND2_X1 U9803 ( .A1(n9723), .A2(n8752), .ZN(n8707) );
  NAND2_X1 U9804 ( .A1(n8708), .A2(n8707), .ZN(n8709) );
  XNOR2_X1 U9805 ( .A(n8709), .B(n4854), .ZN(n8712) );
  AND2_X1 U9806 ( .A1(n9723), .A2(n8744), .ZN(n8710) );
  AOI21_X1 U9807 ( .B1(n9837), .B2(n8752), .A(n8710), .ZN(n8711) );
  NOR2_X1 U9808 ( .A1(n8712), .A2(n8711), .ZN(n9206) );
  NAND2_X1 U9809 ( .A1(n8712), .A2(n8711), .ZN(n9205) );
  NAND2_X1 U9810 ( .A1(n9833), .A2(n4856), .ZN(n8714) );
  NAND2_X1 U9811 ( .A1(n9713), .A2(n8752), .ZN(n8713) );
  NAND2_X1 U9812 ( .A1(n8714), .A2(n8713), .ZN(n8715) );
  XNOR2_X1 U9813 ( .A(n8715), .B(n8761), .ZN(n9247) );
  NAND2_X1 U9814 ( .A1(n9833), .A2(n8752), .ZN(n8717) );
  NAND2_X1 U9815 ( .A1(n9713), .A2(n8744), .ZN(n8716) );
  NAND2_X1 U9816 ( .A1(n8717), .A2(n8716), .ZN(n9246) );
  NOR2_X1 U9817 ( .A1(n9247), .A2(n9246), .ZN(n8720) );
  INV_X1 U9818 ( .A(n9247), .ZN(n8719) );
  INV_X1 U9819 ( .A(n9246), .ZN(n8718) );
  NAND2_X1 U9820 ( .A1(n9828), .A2(n4856), .ZN(n8722) );
  OR2_X1 U9821 ( .A1(n9260), .A2(n8763), .ZN(n8721) );
  NAND2_X1 U9822 ( .A1(n8722), .A2(n8721), .ZN(n8723) );
  XNOR2_X1 U9823 ( .A(n8723), .B(n4854), .ZN(n8726) );
  NOR2_X1 U9824 ( .A1(n9260), .A2(n8760), .ZN(n8724) );
  AOI21_X1 U9825 ( .B1(n9828), .B2(n8752), .A(n8724), .ZN(n8725) );
  NOR2_X1 U9826 ( .A1(n8726), .A2(n8725), .ZN(n9216) );
  XOR2_X1 U9827 ( .A(n8729), .B(n8727), .Z(n9257) );
  OAI22_X1 U9828 ( .A1(n9648), .A2(n8764), .B1(n9239), .B2(n8763), .ZN(n8730)
         );
  NOR2_X1 U9829 ( .A1(n9239), .A2(n8760), .ZN(n8731) );
  AOI21_X1 U9830 ( .B1(n9816), .B2(n8752), .A(n8731), .ZN(n9197) );
  NAND2_X1 U9831 ( .A1(n9812), .A2(n4856), .ZN(n8735) );
  NAND2_X1 U9832 ( .A1(n9654), .A2(n8752), .ZN(n8734) );
  NAND2_X1 U9833 ( .A1(n8735), .A2(n8734), .ZN(n8736) );
  XNOR2_X1 U9834 ( .A(n8736), .B(n8761), .ZN(n8739) );
  AOI22_X1 U9835 ( .A1(n9812), .A2(n8752), .B1(n8744), .B2(n9654), .ZN(n8737)
         );
  INV_X1 U9836 ( .A(n8737), .ZN(n8738) );
  NAND2_X1 U9837 ( .A1(n9806), .A2(n4856), .ZN(n8742) );
  NAND2_X1 U9838 ( .A1(n9631), .A2(n8752), .ZN(n8741) );
  NAND2_X1 U9839 ( .A1(n8742), .A2(n8741), .ZN(n8743) );
  XNOR2_X1 U9840 ( .A(n8743), .B(n8761), .ZN(n9227) );
  NAND2_X1 U9841 ( .A1(n9806), .A2(n8752), .ZN(n8746) );
  NAND2_X1 U9842 ( .A1(n9631), .A2(n8744), .ZN(n8745) );
  NAND2_X1 U9843 ( .A1(n8746), .A2(n8745), .ZN(n9226) );
  NOR2_X1 U9844 ( .A1(n9227), .A2(n9226), .ZN(n8749) );
  INV_X1 U9845 ( .A(n9227), .ZN(n8748) );
  INV_X1 U9846 ( .A(n9226), .ZN(n8747) );
  XNOR2_X1 U9847 ( .A(n8750), .B(n8751), .ZN(n9278) );
  NAND2_X1 U9848 ( .A1(n9796), .A2(n4856), .ZN(n8754) );
  NAND2_X1 U9849 ( .A1(n9576), .A2(n8752), .ZN(n8753) );
  NAND2_X1 U9850 ( .A1(n8754), .A2(n8753), .ZN(n8755) );
  XNOR2_X1 U9851 ( .A(n8755), .B(n4854), .ZN(n8758) );
  NOR2_X1 U9852 ( .A1(n8771), .A2(n8760), .ZN(n8756) );
  AOI21_X1 U9853 ( .B1(n9796), .B2(n8752), .A(n8756), .ZN(n8757) );
  NAND2_X1 U9854 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  OAI21_X1 U9855 ( .B1(n8758), .B2(n8757), .A(n8759), .ZN(n9190) );
  OAI22_X1 U9856 ( .A1(n9587), .A2(n8763), .B1(n9598), .B2(n8760), .ZN(n8762)
         );
  XNOR2_X1 U9857 ( .A(n8762), .B(n8761), .ZN(n8766) );
  OAI22_X1 U9858 ( .A1(n9587), .A2(n8764), .B1(n9598), .B2(n8763), .ZN(n8765)
         );
  XNOR2_X1 U9859 ( .A(n8766), .B(n8765), .ZN(n8767) );
  INV_X1 U9860 ( .A(n9578), .ZN(n9547) );
  OAI22_X1 U9861 ( .A1(n9584), .A2(n9274), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8768), .ZN(n8769) );
  AOI21_X1 U9862 ( .B1(n9547), .B2(n9262), .A(n8769), .ZN(n8770) );
  OAI21_X1 U9863 ( .B1(n8771), .B2(n9284), .A(n8770), .ZN(n8772) );
  AOI21_X1 U9864 ( .B1(n9790), .B2(n9287), .A(n8772), .ZN(n8773) );
  OAI21_X1 U9865 ( .B1(n8774), .B2(n9289), .A(n8773), .ZN(P1_U3218) );
  INV_X1 U9866 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9337) );
  OAI222_X1 U9867 ( .A1(n8777), .A2(n8776), .B1(n6522), .B2(P1_U3084), .C1(
        n9337), .C2(n8775), .ZN(P1_U3323) );
  INV_X1 U9868 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8780) );
  INV_X1 U9869 ( .A(n8778), .ZN(n8779) );
  OAI222_X1 U9870 ( .A1(n8781), .A2(n8780), .B1(n7619), .B2(n8779), .C1(n6184), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  INV_X1 U9871 ( .A(n9110), .ZN(n8955) );
  OAI211_X1 U9872 ( .C1(n8784), .C2(n8783), .A(n8782), .B(n8844), .ZN(n8789)
         );
  NOR2_X1 U9873 ( .A1(n10393), .A2(n8957), .ZN(n8787) );
  OAI22_X1 U9874 ( .A1(n10394), .A2(n8958), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8785), .ZN(n8786) );
  AOI211_X1 U9875 ( .C1(n8820), .C2(n8953), .A(n8787), .B(n8786), .ZN(n8788)
         );
  OAI211_X1 U9876 ( .C1(n8955), .C2(n10399), .A(n8789), .B(n8788), .ZN(
        P2_U3216) );
  OAI211_X1 U9877 ( .C1(n8790), .C2(n8792), .A(n8791), .B(n8844), .ZN(n8797)
         );
  AOI22_X1 U9878 ( .A1(n8802), .A2(n9013), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8796) );
  INV_X1 U9879 ( .A(n8793), .ZN(n9018) );
  AOI22_X1 U9880 ( .A1(n8804), .A2(n9049), .B1(n8820), .B2(n9018), .ZN(n8795)
         );
  NAND2_X1 U9881 ( .A1(n9132), .A2(n8851), .ZN(n8794) );
  NAND4_X1 U9882 ( .A1(n8797), .A2(n8796), .A3(n8795), .A4(n8794), .ZN(
        P2_U3218) );
  NAND2_X1 U9883 ( .A1(n4891), .A2(n8831), .ZN(n8830) );
  NAND2_X1 U9884 ( .A1(n8830), .A2(n8798), .ZN(n8800) );
  OAI211_X1 U9885 ( .C1(n8801), .C2(n8800), .A(n8799), .B(n8844), .ZN(n8808)
         );
  AOI22_X1 U9886 ( .A1(n8802), .A2(n9049), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8807) );
  INV_X1 U9887 ( .A(n8803), .ZN(n9045) );
  AOI22_X1 U9888 ( .A1(n8804), .A2(n9050), .B1(n8820), .B2(n9045), .ZN(n8806)
         );
  NAND2_X1 U9889 ( .A1(n9143), .A2(n8851), .ZN(n8805) );
  NAND4_X1 U9890 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), .ZN(
        P2_U3225) );
  INV_X1 U9891 ( .A(n8810), .ZN(n8811) );
  AOI21_X1 U9892 ( .B1(n8812), .B2(n8809), .A(n8811), .ZN(n8822) );
  NOR2_X1 U9893 ( .A1(n8813), .A2(n10439), .ZN(n8814) );
  AOI21_X1 U9894 ( .B1(n8920), .B2(n9082), .A(n8814), .ZN(n8981) );
  INV_X1 U9895 ( .A(n8815), .ZN(n8817) );
  OAI22_X1 U9896 ( .A1(n8981), .A2(n8817), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8816), .ZN(n8819) );
  NOR2_X1 U9897 ( .A1(n8989), .A2(n10399), .ZN(n8818) );
  AOI211_X1 U9898 ( .C1(n8820), .C2(n8986), .A(n8819), .B(n8818), .ZN(n8821)
         );
  OAI21_X1 U9899 ( .B1(n8822), .B2(n10397), .A(n8821), .ZN(P2_U3227) );
  OAI211_X1 U9900 ( .C1(n8825), .C2(n8824), .A(n8823), .B(n8844), .ZN(n8829)
         );
  OAI22_X1 U9901 ( .A1(n10394), .A2(n8997), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9943), .ZN(n8827) );
  OAI22_X1 U9902 ( .A1(n10393), .A2(n9035), .B1(n8848), .B2(n9003), .ZN(n8826)
         );
  AOI211_X1 U9903 ( .C1(n9005), .C2(n8851), .A(n8827), .B(n8826), .ZN(n8828)
         );
  NAND2_X1 U9904 ( .A1(n8829), .A2(n8828), .ZN(P2_U3231) );
  OAI211_X1 U9905 ( .C1(n4891), .C2(n8831), .A(n8830), .B(n8844), .ZN(n8835)
         );
  NOR2_X1 U9906 ( .A1(n10394), .A2(n9034), .ZN(n8833) );
  OAI22_X1 U9907 ( .A1(n10393), .A2(n8913), .B1(n8848), .B2(n9060), .ZN(n8832)
         );
  AOI211_X1 U9908 ( .C1(P2_REG3_REG_20__SCAN_IN), .C2(P2_U3152), .A(n8833), 
        .B(n8832), .ZN(n8834) );
  OAI211_X1 U9909 ( .C1(n5141), .C2(n10399), .A(n8835), .B(n8834), .ZN(
        P2_U3235) );
  AOI21_X1 U9910 ( .B1(n8838), .B2(n8837), .A(n8836), .ZN(n8843) );
  OAI22_X1 U9911 ( .A1(n10394), .A2(n9035), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8839), .ZN(n8841) );
  OAI22_X1 U9912 ( .A1(n10393), .A2(n9034), .B1(n8848), .B2(n9027), .ZN(n8840)
         );
  AOI211_X1 U9913 ( .C1(n9138), .C2(n8851), .A(n8841), .B(n8840), .ZN(n8842)
         );
  OAI21_X1 U9914 ( .B1(n8843), .B2(n10397), .A(n8842), .ZN(P2_U3237) );
  OAI211_X1 U9915 ( .C1(n8847), .C2(n8846), .A(n8845), .B(n8844), .ZN(n8853)
         );
  OAI22_X1 U9916 ( .A1(n10394), .A2(n8970), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10140), .ZN(n8850) );
  OAI22_X1 U9917 ( .A1(n10393), .A2(n8997), .B1(n8848), .B2(n8972), .ZN(n8849)
         );
  AOI211_X1 U9918 ( .C1(n9117), .C2(n8851), .A(n8850), .B(n8849), .ZN(n8852)
         );
  NAND2_X1 U9919 ( .A1(n8853), .A2(n8852), .ZN(P2_U3242) );
  MUX2_X1 U9920 ( .A(n8943), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8861), .Z(
        P2_U3581) );
  MUX2_X1 U9921 ( .A(n8944), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8861), .Z(
        P2_U3579) );
  MUX2_X1 U9922 ( .A(n8920), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8861), .Z(
        P2_U3578) );
  MUX2_X1 U9923 ( .A(n9013), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8861), .Z(
        P2_U3576) );
  MUX2_X1 U9924 ( .A(n5113), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8861), .Z(
        P2_U3575) );
  MUX2_X1 U9925 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9049), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9926 ( .A(n9050), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8861), .Z(
        P2_U3572) );
  MUX2_X1 U9927 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9081), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9928 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8855), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9929 ( .A(n8856), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8861), .Z(
        P2_U3566) );
  MUX2_X1 U9930 ( .A(n8857), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8861), .Z(
        P2_U3564) );
  MUX2_X1 U9931 ( .A(n8858), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8861), .Z(
        P2_U3563) );
  MUX2_X1 U9932 ( .A(n8859), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8861), .Z(
        P2_U3562) );
  MUX2_X1 U9933 ( .A(n8860), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8861), .Z(
        P2_U3556) );
  MUX2_X1 U9934 ( .A(n6760), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8861), .Z(
        P2_U3553) );
  MUX2_X1 U9935 ( .A(n8862), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8861), .Z(
        P2_U3552) );
  XNOR2_X1 U9936 ( .A(n8886), .B(n8863), .ZN(n8866) );
  AOI21_X1 U9937 ( .B1(n8875), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8864), .ZN(
        n8865) );
  NAND2_X1 U9938 ( .A1(n8865), .A2(n8866), .ZN(n8882) );
  OAI21_X1 U9939 ( .B1(n8866), .B2(n8865), .A(n8882), .ZN(n8867) );
  INV_X1 U9940 ( .A(n8867), .ZN(n8881) );
  INV_X1 U9941 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8868) );
  NOR2_X1 U9942 ( .A1(n8893), .A2(n8868), .ZN(n8869) );
  AOI211_X1 U9943 ( .C1(n10308), .C2(n8886), .A(n8870), .B(n8869), .ZN(n8880)
         );
  INV_X1 U9944 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8873) );
  NOR2_X1 U9945 ( .A1(n8872), .A2(n8873), .ZN(n8871) );
  AOI21_X1 U9946 ( .B1(n8873), .B2(n8872), .A(n8871), .ZN(n8877) );
  AOI21_X1 U9947 ( .B1(n8875), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8874), .ZN(
        n8876) );
  NAND2_X1 U9948 ( .A1(n8876), .A2(n8877), .ZN(n8885) );
  OAI21_X1 U9949 ( .B1(n8877), .B2(n8876), .A(n8885), .ZN(n8878) );
  NAND2_X1 U9950 ( .A1(n8878), .A2(n8896), .ZN(n8879) );
  OAI211_X1 U9951 ( .C1(n8881), .C2(n10297), .A(n8880), .B(n8879), .ZN(
        P2_U3263) );
  OAI21_X1 U9952 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n8886), .A(n8882), .ZN(
        n8884) );
  XNOR2_X1 U9953 ( .A(n8973), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8883) );
  XNOR2_X1 U9954 ( .A(n8884), .B(n8883), .ZN(n8899) );
  OAI21_X1 U9955 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8886), .A(n8885), .ZN(
        n8889) );
  XNOR2_X1 U9956 ( .A(n8973), .B(n8887), .ZN(n8888) );
  XNOR2_X1 U9957 ( .A(n8889), .B(n8888), .ZN(n8897) );
  NOR2_X1 U9958 ( .A1(n8891), .A2(n8890), .ZN(n8895) );
  OAI21_X1 U9959 ( .B1(n8893), .B2(n5278), .A(n8892), .ZN(n8894) );
  AOI211_X1 U9960 ( .C1(n8897), .C2(n8896), .A(n8895), .B(n8894), .ZN(n8898)
         );
  OAI21_X1 U9961 ( .B1(n10297), .B2(n8899), .A(n8898), .ZN(P2_U3264) );
  INV_X1 U9962 ( .A(n9094), .ZN(n8908) );
  NAND2_X1 U9963 ( .A1(n9125), .A2(n9002), .ZN(n9001) );
  OR2_X2 U9964 ( .A1(n9122), .A2(n9001), .ZN(n8983) );
  NOR2_X2 U9965 ( .A1(n9117), .A2(n8983), .ZN(n8971) );
  NOR2_X1 U9966 ( .A1(n8902), .A2(n8901), .ZN(n8903) );
  OR2_X1 U9967 ( .A1(n10441), .A2(n8903), .ZN(n8927) );
  NOR2_X1 U9968 ( .A1(n8904), .A2(n8927), .ZN(n9093) );
  NAND2_X1 U9969 ( .A1(n4833), .A2(n9093), .ZN(n8909) );
  OAI21_X1 U9970 ( .B1(n4833), .B2(n8905), .A(n8909), .ZN(n8906) );
  AOI21_X1 U9971 ( .B1(n9090), .B2(n10466), .A(n8906), .ZN(n8907) );
  OAI21_X1 U9972 ( .B1(n9092), .B2(n9008), .A(n8907), .ZN(P2_U3265) );
  XNOR2_X1 U9973 ( .A(n8908), .B(n8928), .ZN(n9096) );
  INV_X1 U9974 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8910) );
  OAI21_X1 U9975 ( .B1(n4833), .B2(n8910), .A(n8909), .ZN(n8911) );
  AOI21_X1 U9976 ( .B1(n9094), .B2(n10466), .A(n8911), .ZN(n8912) );
  OAI21_X1 U9977 ( .B1(n9096), .B2(n9008), .A(n8912), .ZN(P2_U3266) );
  NAND2_X1 U9978 ( .A1(n9063), .A2(n9062), .ZN(n9061) );
  NAND2_X1 U9979 ( .A1(n9061), .A2(n8916), .ZN(n9042) );
  NOR2_X1 U9980 ( .A1(n9042), .A2(n9047), .ZN(n9041) );
  AOI21_X1 U9981 ( .B1(n8937), .B2(n8942), .A(n5466), .ZN(n8922) );
  XNOR2_X1 U9982 ( .A(n8922), .B(n8921), .ZN(n9097) );
  INV_X1 U9983 ( .A(n9097), .ZN(n8935) );
  XNOR2_X1 U9984 ( .A(n8924), .B(n8923), .ZN(n8925) );
  OAI222_X1 U9985 ( .A1(n10439), .A2(n8958), .B1(n8927), .B2(n8926), .C1(n8925), .C2(n10437), .ZN(n9099) );
  AOI21_X1 U9986 ( .B1(n8929), .B2(n8938), .A(n8928), .ZN(n9098) );
  NAND2_X1 U9987 ( .A1(n9098), .A2(n10461), .ZN(n8932) );
  AOI22_X1 U9988 ( .A1(n10469), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8930), .B2(
        n10458), .ZN(n8931) );
  OAI211_X1 U9989 ( .C1(n5147), .C2(n9076), .A(n8932), .B(n8931), .ZN(n8933)
         );
  AOI21_X1 U9990 ( .B1(n9099), .B2(n4833), .A(n8933), .ZN(n8934) );
  OAI21_X1 U9991 ( .B1(n8935), .B2(n9089), .A(n8934), .ZN(P2_U3267) );
  XNOR2_X1 U9992 ( .A(n8937), .B(n8936), .ZN(n9109) );
  INV_X1 U9993 ( .A(n8938), .ZN(n8939) );
  AOI21_X1 U9994 ( .B1(n9105), .B2(n8950), .A(n8939), .ZN(n9106) );
  AOI22_X1 U9995 ( .A1(n10469), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8940), .B2(
        n10458), .ZN(n8941) );
  OAI21_X1 U9996 ( .B1(n5148), .B2(n9076), .A(n8941), .ZN(n8946) );
  NOR2_X1 U9997 ( .A1(n9108), .A2(n10469), .ZN(n8945) );
  AOI211_X1 U9998 ( .C1(n10461), .C2(n9106), .A(n8946), .B(n8945), .ZN(n8947)
         );
  OAI21_X1 U9999 ( .B1(n9109), .B2(n9089), .A(n8947), .ZN(P2_U3268) );
  XNOR2_X1 U10000 ( .A(n8949), .B(n8948), .ZN(n9114) );
  INV_X1 U10001 ( .A(n8971), .ZN(n8952) );
  INV_X1 U10002 ( .A(n8950), .ZN(n8951) );
  AOI21_X1 U10003 ( .B1(n9110), .B2(n8952), .A(n8951), .ZN(n9111) );
  AOI22_X1 U10004 ( .A1(n10469), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8953), 
        .B2(n10458), .ZN(n8954) );
  OAI21_X1 U10005 ( .B1(n8955), .B2(n9076), .A(n8954), .ZN(n8963) );
  AOI21_X1 U10006 ( .B1(n4895), .B2(n8956), .A(n10437), .ZN(n8961) );
  OAI22_X1 U10007 ( .A1(n8958), .A2(n10441), .B1(n8957), .B2(n10439), .ZN(
        n8959) );
  AOI21_X1 U10008 ( .B1(n8961), .B2(n8960), .A(n8959), .ZN(n9113) );
  NOR2_X1 U10009 ( .A1(n9113), .A2(n10469), .ZN(n8962) );
  AOI211_X1 U10010 ( .C1(n10461), .C2(n9111), .A(n8963), .B(n8962), .ZN(n8964)
         );
  OAI21_X1 U10011 ( .B1(n9114), .B2(n9089), .A(n8964), .ZN(P2_U3269) );
  XOR2_X1 U10012 ( .A(n8967), .B(n8965), .Z(n9119) );
  AOI22_X1 U10013 ( .A1(n9117), .A2(n10466), .B1(n10469), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U10014 ( .A1(n8979), .A2(n8966), .ZN(n8968) );
  XNOR2_X1 U10015 ( .A(n8968), .B(n8967), .ZN(n8969) );
  OAI222_X1 U10016 ( .A1(n10441), .A2(n8970), .B1(n10439), .B2(n8997), .C1(
        n10437), .C2(n8969), .ZN(n9115) );
  AOI211_X1 U10017 ( .C1(n9117), .C2(n8983), .A(n10639), .B(n8971), .ZN(n9116)
         );
  INV_X1 U10018 ( .A(n9116), .ZN(n8974) );
  OAI22_X1 U10019 ( .A1(n8974), .A2(n8973), .B1(n10373), .B2(n8972), .ZN(n8975) );
  OAI21_X1 U10020 ( .B1(n9115), .B2(n8975), .A(n4833), .ZN(n8976) );
  OAI211_X1 U10021 ( .C1(n9119), .C2(n9089), .A(n8977), .B(n8976), .ZN(
        P2_U3270) );
  XNOR2_X1 U10022 ( .A(n8978), .B(n5384), .ZN(n9124) );
  OAI211_X1 U10023 ( .C1(n5384), .C2(n8980), .A(n8979), .B(n9085), .ZN(n8982)
         );
  NAND2_X1 U10024 ( .A1(n8982), .A2(n8981), .ZN(n9120) );
  INV_X1 U10025 ( .A(n8983), .ZN(n8984) );
  AOI211_X1 U10026 ( .C1(n9122), .C2(n9001), .A(n10639), .B(n8984), .ZN(n9121)
         );
  NAND2_X1 U10027 ( .A1(n9121), .A2(n8985), .ZN(n8988) );
  AOI22_X1 U10028 ( .A1(n10469), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8986), 
        .B2(n10458), .ZN(n8987) );
  OAI211_X1 U10029 ( .C1(n8989), .C2(n9076), .A(n8988), .B(n8987), .ZN(n8990)
         );
  AOI21_X1 U10030 ( .B1(n9120), .B2(n4833), .A(n8990), .ZN(n8991) );
  OAI21_X1 U10031 ( .B1(n9124), .B2(n9089), .A(n8991), .ZN(P2_U3271) );
  OAI211_X1 U10032 ( .C1(n8994), .C2(n8993), .A(n8992), .B(n9085), .ZN(n8996)
         );
  NAND2_X1 U10033 ( .A1(n5113), .A2(n9080), .ZN(n8995) );
  OAI211_X1 U10034 ( .C1(n8997), .C2(n10441), .A(n8996), .B(n8995), .ZN(n9128)
         );
  INV_X1 U10035 ( .A(n9128), .ZN(n9011) );
  OAI21_X1 U10036 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(n9129) );
  OAI21_X1 U10037 ( .B1(n9125), .B2(n9002), .A(n9001), .ZN(n9126) );
  INV_X1 U10038 ( .A(n9003), .ZN(n9004) );
  AOI22_X1 U10039 ( .A1(n10469), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9004), 
        .B2(n10458), .ZN(n9007) );
  NAND2_X1 U10040 ( .A1(n9005), .A2(n10466), .ZN(n9006) );
  OAI211_X1 U10041 ( .C1(n9126), .C2(n9008), .A(n9007), .B(n9006), .ZN(n9009)
         );
  AOI21_X1 U10042 ( .B1(n9129), .B2(n10457), .A(n9009), .ZN(n9010) );
  OAI21_X1 U10043 ( .B1(n10469), .B2(n9011), .A(n9010), .ZN(P2_U3272) );
  XNOR2_X1 U10044 ( .A(n9012), .B(n9015), .ZN(n9014) );
  AOI222_X1 U10045 ( .A1(n9085), .A2(n9014), .B1(n9049), .B2(n9080), .C1(n9013), .C2(n9082), .ZN(n9135) );
  INV_X1 U10046 ( .A(n9137), .ZN(n9017) );
  NAND2_X1 U10047 ( .A1(n9016), .A2(n9015), .ZN(n9131) );
  NAND3_X1 U10048 ( .A1(n9017), .A2(n10457), .A3(n9131), .ZN(n9023) );
  XOR2_X1 U10049 ( .A(n9025), .B(n9132), .Z(n9133) );
  INV_X1 U10050 ( .A(n9132), .ZN(n9020) );
  AOI22_X1 U10051 ( .A1(n10469), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9018), 
        .B2(n10458), .ZN(n9019) );
  OAI21_X1 U10052 ( .B1(n9020), .B2(n9076), .A(n9019), .ZN(n9021) );
  AOI21_X1 U10053 ( .B1(n9133), .B2(n10461), .A(n9021), .ZN(n9022) );
  OAI211_X1 U10054 ( .C1(n10469), .C2(n9135), .A(n9023), .B(n9022), .ZN(
        P2_U3273) );
  XNOR2_X1 U10055 ( .A(n9024), .B(n9033), .ZN(n9142) );
  INV_X1 U10056 ( .A(n9025), .ZN(n9026) );
  AOI21_X1 U10057 ( .B1(n9138), .B2(n9043), .A(n9026), .ZN(n9139) );
  INV_X1 U10058 ( .A(n9138), .ZN(n9030) );
  INV_X1 U10059 ( .A(n9027), .ZN(n9028) );
  AOI22_X1 U10060 ( .A1(n10469), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9028), 
        .B2(n10458), .ZN(n9029) );
  OAI21_X1 U10061 ( .B1(n9030), .B2(n9076), .A(n9029), .ZN(n9039) );
  AOI211_X1 U10062 ( .C1(n9033), .C2(n9031), .A(n10437), .B(n9032), .ZN(n9037)
         );
  OAI22_X1 U10063 ( .A1(n9035), .A2(n10441), .B1(n9034), .B2(n10439), .ZN(
        n9036) );
  NOR2_X1 U10064 ( .A1(n9037), .A2(n9036), .ZN(n9141) );
  NOR2_X1 U10065 ( .A1(n9141), .A2(n10469), .ZN(n9038) );
  AOI211_X1 U10066 ( .C1(n9139), .C2(n10461), .A(n9039), .B(n9038), .ZN(n9040)
         );
  OAI21_X1 U10067 ( .B1(n9089), .B2(n9142), .A(n9040), .ZN(P2_U3274) );
  AOI21_X1 U10068 ( .B1(n9047), .B2(n9042), .A(n9041), .ZN(n9147) );
  INV_X1 U10069 ( .A(n9043), .ZN(n9044) );
  AOI21_X1 U10070 ( .B1(n9143), .B2(n4924), .A(n9044), .ZN(n9144) );
  AOI22_X1 U10071 ( .A1(n10469), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9045), 
        .B2(n10458), .ZN(n9046) );
  OAI21_X1 U10072 ( .B1(n8414), .B2(n9076), .A(n9046), .ZN(n9053) );
  XNOR2_X1 U10073 ( .A(n9048), .B(n9047), .ZN(n9051) );
  AOI222_X1 U10074 ( .A1(n9085), .A2(n9051), .B1(n9050), .B2(n9080), .C1(n9049), .C2(n9082), .ZN(n9146) );
  NOR2_X1 U10075 ( .A1(n9146), .A2(n10469), .ZN(n9052) );
  AOI211_X1 U10076 ( .C1(n9144), .C2(n10461), .A(n9053), .B(n9052), .ZN(n9054)
         );
  OAI21_X1 U10077 ( .B1(n9147), .B2(n9089), .A(n9054), .ZN(P2_U3275) );
  XNOR2_X1 U10078 ( .A(n9055), .B(n9062), .ZN(n9057) );
  AOI222_X1 U10079 ( .A1(n9085), .A2(n9057), .B1(n9083), .B2(n9080), .C1(n9056), .C2(n9082), .ZN(n9151) );
  XNOR2_X1 U10080 ( .A(n4921), .B(n9148), .ZN(n9149) );
  NAND2_X1 U10081 ( .A1(n9148), .A2(n10466), .ZN(n9059) );
  NAND2_X1 U10082 ( .A1(n10469), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9058) );
  OAI211_X1 U10083 ( .C1(n10373), .C2(n9060), .A(n9059), .B(n9058), .ZN(n9065)
         );
  OAI21_X1 U10084 ( .B1(n9063), .B2(n9062), .A(n9061), .ZN(n9152) );
  NOR2_X1 U10085 ( .A1(n9152), .A2(n9089), .ZN(n9064) );
  AOI211_X1 U10086 ( .C1(n9149), .C2(n10461), .A(n9065), .B(n9064), .ZN(n9066)
         );
  OAI21_X1 U10087 ( .B1(n10469), .B2(n9151), .A(n9066), .ZN(P2_U3276) );
  XNOR2_X1 U10088 ( .A(n9068), .B(n9067), .ZN(n9162) );
  INV_X1 U10089 ( .A(n9069), .ZN(n9072) );
  INV_X1 U10090 ( .A(n9070), .ZN(n9071) );
  AOI21_X1 U10091 ( .B1(n9158), .B2(n9072), .A(n9071), .ZN(n9159) );
  INV_X1 U10092 ( .A(n9073), .ZN(n9074) );
  AOI22_X1 U10093 ( .A1(n10469), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9074), 
        .B2(n10458), .ZN(n9075) );
  OAI21_X1 U10094 ( .B1(n9077), .B2(n9076), .A(n9075), .ZN(n9087) );
  XNOR2_X1 U10095 ( .A(n9079), .B(n9078), .ZN(n9084) );
  AOI222_X1 U10096 ( .A1(n9085), .A2(n9084), .B1(n9083), .B2(n9082), .C1(n9081), .C2(n9080), .ZN(n9161) );
  NOR2_X1 U10097 ( .A1(n9161), .A2(n10469), .ZN(n9086) );
  AOI211_X1 U10098 ( .C1(n9159), .C2(n10461), .A(n9087), .B(n9086), .ZN(n9088)
         );
  OAI21_X1 U10099 ( .B1(n9162), .B2(n9089), .A(n9088), .ZN(P2_U3278) );
  AOI21_X1 U10100 ( .B1(n9090), .B2(n10150), .A(n9093), .ZN(n9091) );
  OAI21_X1 U10101 ( .B1(n9092), .B2(n10639), .A(n9091), .ZN(n9173) );
  MUX2_X1 U10102 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9173), .S(n10646), .Z(
        P2_U3551) );
  AOI21_X1 U10103 ( .B1(n9094), .B2(n10150), .A(n9093), .ZN(n9095) );
  OAI21_X1 U10104 ( .B1(n9096), .B2(n10639), .A(n9095), .ZN(n9174) );
  MUX2_X1 U10105 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9174), .S(n10646), .Z(
        P2_U3550) );
  NAND2_X1 U10106 ( .A1(n9097), .A2(n10644), .ZN(n9104) );
  INV_X1 U10107 ( .A(n9098), .ZN(n9101) );
  INV_X1 U10108 ( .A(n9099), .ZN(n9100) );
  OAI211_X1 U10109 ( .C1(n10639), .C2(n9101), .A(n5467), .B(n9100), .ZN(n9102)
         );
  INV_X1 U10110 ( .A(n9102), .ZN(n9103) );
  NAND2_X1 U10111 ( .A1(n9104), .A2(n9103), .ZN(n9175) );
  MUX2_X1 U10112 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9175), .S(n10646), .Z(
        P2_U3549) );
  AOI22_X1 U10113 ( .A1(n9106), .A2(n10449), .B1(n10150), .B2(n9105), .ZN(
        n9107) );
  OAI211_X1 U10114 ( .C1(n9109), .C2(n10620), .A(n9108), .B(n9107), .ZN(n9176)
         );
  MUX2_X1 U10115 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9176), .S(n10646), .Z(
        P2_U3548) );
  AOI22_X1 U10116 ( .A1(n9111), .A2(n10449), .B1(n10150), .B2(n9110), .ZN(
        n9112) );
  OAI211_X1 U10117 ( .C1(n9114), .C2(n10620), .A(n9113), .B(n9112), .ZN(n9177)
         );
  MUX2_X1 U10118 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9177), .S(n10646), .Z(
        P2_U3547) );
  AOI211_X1 U10119 ( .C1(n10150), .C2(n9117), .A(n9116), .B(n9115), .ZN(n9118)
         );
  OAI21_X1 U10120 ( .B1(n9119), .B2(n10620), .A(n9118), .ZN(n9178) );
  MUX2_X1 U10121 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9178), .S(n10646), .Z(
        P2_U3546) );
  AOI211_X1 U10122 ( .C1(n10150), .C2(n9122), .A(n9121), .B(n9120), .ZN(n9123)
         );
  OAI21_X1 U10123 ( .B1(n9124), .B2(n10620), .A(n9123), .ZN(n9179) );
  MUX2_X1 U10124 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9179), .S(n10646), .Z(
        P2_U3545) );
  OAI22_X1 U10125 ( .A1(n9126), .A2(n10639), .B1(n9125), .B2(n10638), .ZN(
        n9127) );
  AOI211_X1 U10126 ( .C1(n9129), .C2(n10644), .A(n9128), .B(n9127), .ZN(n9130)
         );
  INV_X1 U10127 ( .A(n9130), .ZN(n9180) );
  MUX2_X1 U10128 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9180), .S(n10646), .Z(
        P2_U3544) );
  NAND2_X1 U10129 ( .A1(n9131), .A2(n10644), .ZN(n9136) );
  AOI22_X1 U10130 ( .A1(n9133), .A2(n10449), .B1(n10150), .B2(n9132), .ZN(
        n9134) );
  OAI211_X1 U10131 ( .C1(n9137), .C2(n9136), .A(n9135), .B(n9134), .ZN(n9181)
         );
  MUX2_X1 U10132 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9181), .S(n10646), .Z(
        P2_U3543) );
  AOI22_X1 U10133 ( .A1(n9139), .A2(n10449), .B1(n10150), .B2(n9138), .ZN(
        n9140) );
  OAI211_X1 U10134 ( .C1(n9142), .C2(n10620), .A(n9141), .B(n9140), .ZN(n9182)
         );
  MUX2_X1 U10135 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9182), .S(n10646), .Z(
        P2_U3542) );
  AOI22_X1 U10136 ( .A1(n9144), .A2(n10449), .B1(n10150), .B2(n9143), .ZN(
        n9145) );
  OAI211_X1 U10137 ( .C1(n9147), .C2(n10620), .A(n9146), .B(n9145), .ZN(n9183)
         );
  MUX2_X1 U10138 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9183), .S(n10646), .Z(
        P2_U3541) );
  AOI22_X1 U10139 ( .A1(n9149), .A2(n10449), .B1(n10150), .B2(n9148), .ZN(
        n9150) );
  OAI211_X1 U10140 ( .C1(n9152), .C2(n10620), .A(n9151), .B(n9150), .ZN(n9184)
         );
  MUX2_X1 U10141 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9184), .S(n10646), .Z(
        P2_U3540) );
  AOI211_X1 U10142 ( .C1(n10150), .C2(n9155), .A(n9154), .B(n9153), .ZN(n9156)
         );
  OAI21_X1 U10143 ( .B1(n10620), .B2(n9157), .A(n9156), .ZN(n9185) );
  MUX2_X1 U10144 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9185), .S(n10646), .Z(
        P2_U3539) );
  AOI22_X1 U10145 ( .A1(n9159), .A2(n10449), .B1(n10150), .B2(n9158), .ZN(
        n9160) );
  OAI211_X1 U10146 ( .C1(n9162), .C2(n10620), .A(n9161), .B(n9160), .ZN(n9186)
         );
  MUX2_X1 U10147 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9186), .S(n10646), .Z(
        P2_U3538) );
  AOI211_X1 U10148 ( .C1(n10150), .C2(n9165), .A(n9164), .B(n9163), .ZN(n9166)
         );
  OAI21_X1 U10149 ( .B1(n10620), .B2(n9167), .A(n9166), .ZN(n9187) );
  MUX2_X1 U10150 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9187), .S(n10646), .Z(
        P2_U3537) );
  AOI21_X1 U10151 ( .B1(n10150), .B2(n9169), .A(n9168), .ZN(n9170) );
  OAI211_X1 U10152 ( .C1(n9172), .C2(n10620), .A(n9171), .B(n9170), .ZN(n9188)
         );
  MUX2_X1 U10153 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9188), .S(n10646), .Z(
        P2_U3536) );
  MUX2_X1 U10154 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9173), .S(n10650), .Z(
        P2_U3519) );
  MUX2_X1 U10155 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9174), .S(n10650), .Z(
        P2_U3518) );
  MUX2_X1 U10156 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9175), .S(n10650), .Z(
        P2_U3517) );
  MUX2_X1 U10157 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9176), .S(n10650), .Z(
        P2_U3516) );
  MUX2_X1 U10158 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9177), .S(n10650), .Z(
        P2_U3515) );
  MUX2_X1 U10159 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9178), .S(n10650), .Z(
        P2_U3514) );
  MUX2_X1 U10160 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9179), .S(n10650), .Z(
        P2_U3513) );
  MUX2_X1 U10161 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9180), .S(n10650), .Z(
        P2_U3512) );
  MUX2_X1 U10162 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9181), .S(n10650), .Z(
        P2_U3511) );
  MUX2_X1 U10163 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9182), .S(n10650), .Z(
        P2_U3510) );
  MUX2_X1 U10164 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9183), .S(n10650), .Z(
        P2_U3509) );
  MUX2_X1 U10165 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9184), .S(n10650), .Z(
        P2_U3508) );
  MUX2_X1 U10166 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9185), .S(n10650), .Z(
        P2_U3507) );
  MUX2_X1 U10167 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9186), .S(n10650), .Z(
        P2_U3505) );
  MUX2_X1 U10168 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9187), .S(n10650), .Z(
        P2_U3502) );
  MUX2_X1 U10169 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9188), .S(n10650), .Z(
        P2_U3499) );
  MUX2_X1 U10170 ( .A(n9189), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10171 ( .A(n9592), .ZN(n9193) );
  AOI22_X1 U10172 ( .A1(n9618), .A2(n9250), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9192) );
  OAI21_X1 U10173 ( .B1(n9274), .B2(n9193), .A(n9192), .ZN(n9194) );
  AOI21_X1 U10174 ( .B1(n9262), .B2(n5187), .A(n9194), .ZN(n9195) );
  OAI211_X1 U10175 ( .C1(n9594), .C2(n9224), .A(n9196), .B(n9195), .ZN(
        P1_U3212) );
  XNOR2_X1 U10176 ( .A(n5462), .B(n9197), .ZN(n9198) );
  XNOR2_X1 U10177 ( .A(n9199), .B(n9198), .ZN(n9204) );
  NAND2_X1 U10178 ( .A1(n9654), .A2(n9262), .ZN(n9201) );
  AOI22_X1 U10179 ( .A1(n9653), .A2(n9250), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9200) );
  OAI211_X1 U10180 ( .C1(n9274), .C2(n9645), .A(n9201), .B(n9200), .ZN(n9202)
         );
  AOI21_X1 U10181 ( .B1(n9816), .B2(n9287), .A(n9202), .ZN(n9203) );
  OAI21_X1 U10182 ( .B1(n9204), .B2(n9289), .A(n9203), .ZN(P1_U3214) );
  NOR2_X1 U10183 ( .A1(n9206), .A2(n5246), .ZN(n9207) );
  XNOR2_X1 U10184 ( .A(n9208), .B(n9207), .ZN(n9214) );
  OAI21_X1 U10185 ( .B1(n9680), .B2(n9242), .A(n9209), .ZN(n9210) );
  AOI21_X1 U10186 ( .B1(n9250), .B2(n9712), .A(n9210), .ZN(n9211) );
  OAI21_X1 U10187 ( .B1(n9274), .B2(n9708), .A(n9211), .ZN(n9212) );
  AOI21_X1 U10188 ( .B1(n9837), .B2(n9287), .A(n9212), .ZN(n9213) );
  OAI21_X1 U10189 ( .B1(n9214), .B2(n9289), .A(n9213), .ZN(P1_U3217) );
  INV_X1 U10190 ( .A(n9828), .ZN(n9225) );
  OAI21_X1 U10191 ( .B1(n9216), .B2(n9218), .A(n9215), .ZN(n9217) );
  OAI21_X1 U10192 ( .B1(n4892), .B2(n9218), .A(n9217), .ZN(n9219) );
  NAND2_X1 U10193 ( .A1(n9219), .A2(n4834), .ZN(n9223) );
  AOI22_X1 U10194 ( .A1(n9713), .A2(n9250), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9220) );
  OAI21_X1 U10195 ( .B1(n9681), .B2(n9242), .A(n9220), .ZN(n9221) );
  AOI21_X1 U10196 ( .B1(n9684), .B2(n9280), .A(n9221), .ZN(n9222) );
  OAI211_X1 U10197 ( .C1(n9225), .C2(n9224), .A(n9223), .B(n9222), .ZN(
        P1_U3221) );
  XNOR2_X1 U10198 ( .A(n9227), .B(n9226), .ZN(n9228) );
  XNOR2_X1 U10199 ( .A(n9229), .B(n9228), .ZN(n9235) );
  NAND2_X1 U10200 ( .A1(n9618), .A2(n9262), .ZN(n9232) );
  INV_X1 U10201 ( .A(n9230), .ZN(n9612) );
  AOI22_X1 U10202 ( .A1(n9612), .A2(n9280), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9231) );
  OAI211_X1 U10203 ( .C1(n9305), .C2(n9284), .A(n9232), .B(n9231), .ZN(n9233)
         );
  AOI21_X1 U10204 ( .B1(n9806), .B2(n9287), .A(n9233), .ZN(n9234) );
  OAI21_X1 U10205 ( .B1(n9235), .B2(n9289), .A(n9234), .ZN(P1_U3223) );
  XOR2_X1 U10206 ( .A(n9237), .B(n9236), .Z(n9245) );
  OAI22_X1 U10207 ( .A1(n9239), .A2(n9284), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9238), .ZN(n9240) );
  AOI21_X1 U10208 ( .B1(n9634), .B2(n9280), .A(n9240), .ZN(n9241) );
  OAI21_X1 U10209 ( .B1(n9285), .B2(n9242), .A(n9241), .ZN(n9243) );
  AOI21_X1 U10210 ( .B1(n9812), .B2(n9287), .A(n9243), .ZN(n9244) );
  OAI21_X1 U10211 ( .B1(n9245), .B2(n9289), .A(n9244), .ZN(P1_U3227) );
  XNOR2_X1 U10212 ( .A(n9247), .B(n9246), .ZN(n9248) );
  XNOR2_X1 U10213 ( .A(n9249), .B(n9248), .ZN(n9255) );
  NAND2_X1 U10214 ( .A1(n9693), .A2(n9262), .ZN(n9252) );
  AOI22_X1 U10215 ( .A1(n9723), .A2(n9250), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9251) );
  OAI211_X1 U10216 ( .C1(n9274), .C2(n9698), .A(n9252), .B(n9251), .ZN(n9253)
         );
  AOI21_X1 U10217 ( .B1(n9833), .B2(n9287), .A(n9253), .ZN(n9254) );
  OAI21_X1 U10218 ( .B1(n9255), .B2(n9289), .A(n9254), .ZN(P1_U3231) );
  AOI21_X1 U10219 ( .B1(n9258), .B2(n9257), .A(n9256), .ZN(n9266) );
  OAI22_X1 U10220 ( .A1(n9260), .A2(n9284), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9259), .ZN(n9261) );
  AOI21_X1 U10221 ( .B1(n9670), .B2(n9262), .A(n9261), .ZN(n9263) );
  OAI21_X1 U10222 ( .B1(n9274), .B2(n9663), .A(n9263), .ZN(n9264) );
  AOI21_X1 U10223 ( .B1(n9821), .B2(n9287), .A(n9264), .ZN(n9265) );
  OAI21_X1 U10224 ( .B1(n9266), .B2(n9289), .A(n9265), .ZN(P1_U3233) );
  NAND2_X1 U10225 ( .A1(n9267), .A2(n9268), .ZN(n9270) );
  XNOR2_X1 U10226 ( .A(n9270), .B(n9269), .ZN(n9277) );
  NAND2_X1 U10227 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10244)
         );
  OAI21_X1 U10228 ( .B1(n9284), .B2(n9271), .A(n10244), .ZN(n9272) );
  AOI21_X1 U10229 ( .B1(n9262), .B2(n9723), .A(n9272), .ZN(n9273) );
  OAI21_X1 U10230 ( .B1(n9274), .B2(n9733), .A(n9273), .ZN(n9275) );
  AOI21_X1 U10231 ( .B1(n9843), .B2(n9287), .A(n9275), .ZN(n9276) );
  OAI21_X1 U10232 ( .B1(n9277), .B2(n9289), .A(n9276), .ZN(P1_U3236) );
  XNOR2_X1 U10233 ( .A(n9279), .B(n9278), .ZN(n9290) );
  NAND2_X1 U10234 ( .A1(n9576), .A2(n9262), .ZN(n9283) );
  AOI22_X1 U10235 ( .A1(n9281), .A2(n9280), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9282) );
  OAI211_X1 U10236 ( .C1(n9285), .C2(n9284), .A(n9283), .B(n9282), .ZN(n9286)
         );
  AOI21_X1 U10237 ( .B1(n9801), .B2(n9287), .A(n9286), .ZN(n9288) );
  OAI21_X1 U10238 ( .B1(n9290), .B2(n9289), .A(n9288), .ZN(P1_U3238) );
  NOR3_X1 U10239 ( .A1(n9743), .A2(n9291), .A3(n10220), .ZN(n9544) );
  INV_X1 U10240 ( .A(n9376), .ZN(n9294) );
  INV_X1 U10241 ( .A(n9374), .ZN(n9293) );
  INV_X1 U10242 ( .A(n9481), .ZN(n9292) );
  AOI211_X1 U10243 ( .C1(n9294), .C2(n9375), .A(n9293), .B(n9292), .ZN(n9330)
         );
  INV_X1 U10244 ( .A(n9295), .ZN(n9296) );
  NAND2_X1 U10245 ( .A1(n9297), .A2(n9296), .ZN(n9298) );
  NAND2_X1 U10246 ( .A1(n9298), .A2(n9381), .ZN(n9385) );
  INV_X1 U10247 ( .A(n9385), .ZN(n9299) );
  NAND2_X1 U10248 ( .A1(n9299), .A2(n9463), .ZN(n9331) );
  NAND2_X1 U10249 ( .A1(n9300), .A2(n9457), .ZN(n9301) );
  NAND2_X1 U10250 ( .A1(n9301), .A2(n9458), .ZN(n9302) );
  AND2_X1 U10251 ( .A1(n9383), .A2(n9302), .ZN(n9303) );
  OAI21_X1 U10252 ( .B1(n9331), .B2(n9303), .A(n9462), .ZN(n9304) );
  AND2_X1 U10253 ( .A1(n9304), .A2(n9378), .ZN(n9306) );
  OR2_X1 U10254 ( .A1(n9812), .A2(n9305), .ZN(n9466) );
  NAND2_X1 U10255 ( .A1(n9466), .A2(n9626), .ZN(n9380) );
  OAI211_X1 U10256 ( .C1(n9306), .C2(n9380), .A(n9471), .B(n9467), .ZN(n9307)
         );
  NAND4_X1 U10257 ( .A1(n9375), .A2(n9377), .A3(n9472), .A4(n9307), .ZN(n9310)
         );
  AND2_X1 U10258 ( .A1(n9482), .A2(n9308), .ZN(n9487) );
  INV_X1 U10259 ( .A(n9487), .ZN(n9309) );
  AOI21_X1 U10260 ( .B1(n9330), .B2(n9310), .A(n9309), .ZN(n9532) );
  AND2_X1 U10261 ( .A1(n9451), .A2(n9388), .ZN(n9311) );
  NAND2_X1 U10262 ( .A1(n9387), .A2(n9311), .ZN(n9327) );
  INV_X1 U10263 ( .A(n9327), .ZN(n9323) );
  INV_X1 U10264 ( .A(n9407), .ZN(n9312) );
  OAI21_X1 U10265 ( .B1(n9313), .B2(n9312), .A(n9411), .ZN(n9314) );
  NAND3_X1 U10266 ( .A1(n9416), .A2(n9314), .A3(n9412), .ZN(n9315) );
  NAND3_X1 U10267 ( .A1(n9423), .A2(n9415), .A3(n9315), .ZN(n9316) );
  NAND2_X1 U10268 ( .A1(n9316), .A2(n9421), .ZN(n9317) );
  NAND2_X1 U10269 ( .A1(n9438), .A2(n9317), .ZN(n9318) );
  NAND2_X1 U10270 ( .A1(n9318), .A2(n9425), .ZN(n9319) );
  NAND2_X1 U10271 ( .A1(n9422), .A2(n9319), .ZN(n9320) );
  NAND3_X1 U10272 ( .A1(n9444), .A2(n9426), .A3(n9320), .ZN(n9321) );
  NAND3_X1 U10273 ( .A1(n9389), .A2(n9445), .A3(n9321), .ZN(n9322) );
  AND2_X1 U10274 ( .A1(n9323), .A2(n9322), .ZN(n9527) );
  AND4_X1 U10275 ( .A1(n9416), .A2(n9324), .A3(n9412), .A4(n9407), .ZN(n9325)
         );
  NAND4_X1 U10276 ( .A1(n9426), .A2(n9325), .A3(n9425), .A4(n9421), .ZN(n9326)
         );
  OR3_X1 U10277 ( .A1(n9327), .A2(n5412), .A3(n9326), .ZN(n9525) );
  INV_X1 U10278 ( .A(n9328), .ZN(n9329) );
  NOR2_X1 U10279 ( .A1(n9525), .A2(n9329), .ZN(n9336) );
  INV_X1 U10280 ( .A(n9330), .ZN(n9335) );
  INV_X1 U10281 ( .A(n9471), .ZN(n9334) );
  INV_X1 U10282 ( .A(n9331), .ZN(n9332) );
  NAND4_X1 U10283 ( .A1(n9467), .A2(n9332), .A3(n9378), .A4(n9458), .ZN(n9333)
         );
  NOR3_X1 U10284 ( .A1(n9335), .A2(n9334), .A3(n9333), .ZN(n9526) );
  OAI21_X1 U10285 ( .B1(n9527), .B2(n9336), .A(n9526), .ZN(n9342) );
  NOR2_X1 U10286 ( .A1(n9345), .A2(n9337), .ZN(n9338) );
  INV_X1 U10287 ( .A(n9564), .ZN(n9781) );
  NAND2_X1 U10288 ( .A1(n9558), .A2(n9546), .ZN(n9340) );
  NAND2_X1 U10289 ( .A1(n9781), .A2(n9340), .ZN(n9491) );
  INV_X1 U10290 ( .A(n9491), .ZN(n9341) );
  INV_X1 U10291 ( .A(n9489), .ZN(n9529) );
  AOI211_X1 U10292 ( .C1(n9532), .C2(n9342), .A(n9341), .B(n9529), .ZN(n9350)
         );
  AND2_X1 U10293 ( .A1(n9564), .A2(n9546), .ZN(n9534) );
  INV_X1 U10294 ( .A(n9534), .ZN(n9343) );
  NAND2_X1 U10295 ( .A1(n9343), .A2(n9558), .ZN(n9348) );
  NAND2_X1 U10296 ( .A1(n9344), .A2(n6944), .ZN(n9347) );
  OR2_X1 U10297 ( .A1(n9345), .A2(n6589), .ZN(n9346) );
  NAND2_X1 U10298 ( .A1(n9348), .A2(n9778), .ZN(n9485) );
  INV_X1 U10299 ( .A(n9485), .ZN(n9349) );
  OAI211_X1 U10300 ( .C1(n9350), .C2(n9349), .A(n6234), .B(n9533), .ZN(n9373)
         );
  NOR2_X1 U10301 ( .A1(n9564), .A2(n9546), .ZN(n9530) );
  INV_X1 U10302 ( .A(n9667), .ZN(n9660) );
  INV_X1 U10303 ( .A(n9720), .ZN(n9727) );
  NAND4_X1 U10304 ( .A1(n9355), .A2(n9354), .A3(n9353), .A4(n10353), .ZN(n9357) );
  NOR4_X1 U10305 ( .A1(n9357), .A2(n7248), .A3(n10519), .A4(n9356), .ZN(n9359)
         );
  NAND3_X1 U10306 ( .A1(n9359), .A2(n9401), .A3(n9358), .ZN(n9360) );
  NOR4_X1 U10307 ( .A1(n9410), .A2(n9362), .A3(n9361), .A4(n9360), .ZN(n9363)
         );
  NAND4_X1 U10308 ( .A1(n9365), .A2(n9418), .A3(n9364), .A4(n9363), .ZN(n9366)
         );
  NOR4_X1 U10309 ( .A1(n9742), .A2(n9367), .A3(n9390), .A4(n9366), .ZN(n9368)
         );
  NAND4_X1 U10310 ( .A1(n9694), .A2(n5415), .A3(n9727), .A4(n9368), .ZN(n9369)
         );
  NOR4_X1 U10311 ( .A1(n9625), .A2(n9660), .A3(n9678), .A4(n9369), .ZN(n9370)
         );
  AOI21_X1 U10312 ( .B1(n9371), .B2(n9533), .A(n6234), .ZN(n9497) );
  INV_X1 U10313 ( .A(n9497), .ZN(n9372) );
  NAND2_X1 U10314 ( .A1(n9373), .A2(n9372), .ZN(n9500) );
  MUX2_X1 U10315 ( .A(n9375), .B(n9374), .S(n9488), .Z(n9480) );
  INV_X1 U10316 ( .A(n9488), .ZN(n9492) );
  MUX2_X1 U10317 ( .A(n9377), .B(n9376), .S(n9492), .Z(n9477) );
  NAND2_X1 U10318 ( .A1(n9467), .A2(n9378), .ZN(n9379) );
  MUX2_X1 U10319 ( .A(n9380), .B(n9379), .S(n9488), .Z(n9470) );
  INV_X1 U10320 ( .A(n9381), .ZN(n9382) );
  NOR2_X1 U10321 ( .A1(n9383), .A2(n9382), .ZN(n9384) );
  MUX2_X1 U10322 ( .A(n9385), .B(n9384), .S(n9492), .Z(n9465) );
  MUX2_X1 U10323 ( .A(n9387), .B(n9386), .S(n9488), .Z(n9456) );
  MUX2_X1 U10324 ( .A(n9389), .B(n9388), .S(n9488), .Z(n9450) );
  INV_X1 U10325 ( .A(n9390), .ZN(n9447) );
  NOR2_X1 U10326 ( .A1(n9391), .A2(n7248), .ZN(n9392) );
  NAND2_X1 U10327 ( .A1(n9393), .A2(n9395), .ZN(n9400) );
  INV_X1 U10328 ( .A(n10519), .ZN(n9394) );
  NAND2_X1 U10329 ( .A1(n9394), .A2(n9519), .ZN(n9396) );
  NAND2_X1 U10330 ( .A1(n9398), .A2(n9397), .ZN(n9399) );
  MUX2_X1 U10331 ( .A(n9403), .B(n9402), .S(n9492), .Z(n9404) );
  MUX2_X1 U10332 ( .A(n9407), .B(n9406), .S(n9488), .Z(n9408) );
  INV_X1 U10333 ( .A(n9410), .ZN(n9414) );
  MUX2_X1 U10334 ( .A(n9412), .B(n9411), .S(n9492), .Z(n9413) );
  MUX2_X1 U10335 ( .A(n9416), .B(n9415), .S(n9488), .Z(n9417) );
  AND2_X1 U10336 ( .A1(n9418), .A2(n9417), .ZN(n9419) );
  NAND2_X1 U10337 ( .A1(n9420), .A2(n9419), .ZN(n9424) );
  NAND3_X1 U10338 ( .A1(n9871), .A2(n9428), .A3(n9488), .ZN(n9427) );
  OAI21_X1 U10339 ( .B1(n9492), .B2(n9550), .A(n9427), .ZN(n9435) );
  NAND3_X1 U10340 ( .A1(n9428), .A2(n9430), .A3(n9488), .ZN(n9429) );
  NAND2_X1 U10341 ( .A1(n9871), .A2(n9429), .ZN(n9433) );
  NOR2_X1 U10342 ( .A1(n9430), .A2(n9488), .ZN(n9436) );
  AND2_X1 U10343 ( .A1(n9436), .A2(n9551), .ZN(n9431) );
  OR2_X1 U10344 ( .A1(n9871), .A2(n9431), .ZN(n9432) );
  AOI22_X1 U10345 ( .A1(n9435), .A2(n9434), .B1(n9433), .B2(n9432), .ZN(n9441)
         );
  INV_X1 U10346 ( .A(n9436), .ZN(n9437) );
  OAI21_X1 U10347 ( .B1(n9438), .B2(n9488), .A(n9437), .ZN(n9439) );
  NAND2_X1 U10348 ( .A1(n9439), .A2(n9866), .ZN(n9440) );
  AND2_X1 U10349 ( .A1(n9441), .A2(n9440), .ZN(n9442) );
  MUX2_X1 U10350 ( .A(n9445), .B(n9444), .S(n9492), .Z(n9446) );
  NAND3_X1 U10351 ( .A1(n9450), .A2(n9449), .A3(n9448), .ZN(n9453) );
  MUX2_X1 U10352 ( .A(n9451), .B(n9724), .S(n9488), .Z(n9452) );
  NAND2_X1 U10353 ( .A1(n9453), .A2(n9452), .ZN(n9454) );
  NAND2_X1 U10354 ( .A1(n9727), .A2(n9454), .ZN(n9455) );
  NAND3_X1 U10355 ( .A1(n5415), .A2(n9456), .A3(n9455), .ZN(n9460) );
  MUX2_X1 U10356 ( .A(n9458), .B(n9457), .S(n9492), .Z(n9459) );
  NAND2_X1 U10357 ( .A1(n9460), .A2(n9459), .ZN(n9461) );
  MUX2_X1 U10358 ( .A(n9463), .B(n9462), .S(n9488), .Z(n9464) );
  MUX2_X1 U10359 ( .A(n9467), .B(n9466), .S(n9488), .Z(n9468) );
  OAI211_X1 U10360 ( .C1(n9470), .C2(n9469), .A(n9617), .B(n9468), .ZN(n9474)
         );
  MUX2_X1 U10361 ( .A(n9472), .B(n9471), .S(n9488), .Z(n9473) );
  NAND3_X1 U10362 ( .A1(n9475), .A2(n9474), .A3(n9473), .ZN(n9476) );
  NAND3_X1 U10363 ( .A1(n9478), .A2(n9477), .A3(n9476), .ZN(n9479) );
  NAND3_X1 U10364 ( .A1(n9568), .A2(n9480), .A3(n9479), .ZN(n9486) );
  NAND3_X1 U10365 ( .A1(n9486), .A2(n9481), .A3(n9489), .ZN(n9483) );
  NAND3_X1 U10366 ( .A1(n9483), .A2(n9492), .A3(n9482), .ZN(n9484) );
  NAND2_X1 U10367 ( .A1(n9487), .A2(n9486), .ZN(n9490) );
  NAND3_X1 U10368 ( .A1(n9490), .A2(n9489), .A3(n9488), .ZN(n9496) );
  OAI21_X1 U10369 ( .B1(n9492), .B2(n9491), .A(n9533), .ZN(n9494) );
  AND2_X1 U10370 ( .A1(n9494), .A2(n9536), .ZN(n9495) );
  AOI21_X1 U10371 ( .B1(n9501), .B2(n9498), .A(n9497), .ZN(n9499) );
  INV_X1 U10372 ( .A(n9501), .ZN(n9503) );
  INV_X1 U10373 ( .A(n9505), .ZN(n9507) );
  NAND2_X1 U10374 ( .A1(n9765), .A2(n10351), .ZN(n9506) );
  NAND3_X1 U10375 ( .A1(n9507), .A2(n6234), .A3(n9506), .ZN(n9508) );
  NAND2_X1 U10376 ( .A1(n9509), .A2(n9508), .ZN(n9511) );
  OAI21_X1 U10377 ( .B1(n9504), .B2(n9511), .A(n9510), .ZN(n9513) );
  NAND2_X1 U10378 ( .A1(n9513), .A2(n9512), .ZN(n9515) );
  OAI211_X1 U10379 ( .C1(n6788), .C2(n7104), .A(n9515), .B(n9514), .ZN(n9518)
         );
  NAND3_X1 U10380 ( .A1(n9518), .A2(n9517), .A3(n9516), .ZN(n9520) );
  NAND2_X1 U10381 ( .A1(n9520), .A2(n9519), .ZN(n9523) );
  AOI21_X1 U10382 ( .B1(n9523), .B2(n9522), .A(n5425), .ZN(n9524) );
  NOR2_X1 U10383 ( .A1(n9525), .A2(n9524), .ZN(n9528) );
  OAI21_X1 U10384 ( .B1(n9528), .B2(n9527), .A(n9526), .ZN(n9531) );
  AOI211_X1 U10385 ( .C1(n9532), .C2(n9531), .A(n9530), .B(n9529), .ZN(n9535)
         );
  OAI21_X1 U10386 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9537) );
  NAND2_X1 U10387 ( .A1(n9537), .A2(n9536), .ZN(n9539) );
  INV_X1 U10388 ( .A(n9539), .ZN(n9541) );
  NOR2_X1 U10389 ( .A1(n9541), .A2(n9540), .ZN(n9543) );
  MUX2_X1 U10390 ( .A(n9546), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9557), .Z(
        P1_U3585) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9547), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10392 ( .A(n5187), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9557), .Z(
        P1_U3583) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9576), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10394 ( .A(n9618), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9557), .Z(
        P1_U3581) );
  MUX2_X1 U10395 ( .A(n9631), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9557), .Z(
        P1_U3580) );
  MUX2_X1 U10396 ( .A(n9654), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9557), .Z(
        P1_U3579) );
  MUX2_X1 U10397 ( .A(n9653), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9557), .Z(
        P1_U3577) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9693), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10399 ( .A(n9713), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9557), .Z(
        P1_U3575) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9723), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9712), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9722), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10403 ( .A(n9548), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9557), .Z(
        P1_U3571) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9549), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9550), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10406 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9551), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10407 ( .A(n9552), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9557), .Z(
        P1_U3567) );
  MUX2_X1 U10408 ( .A(n9553), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9557), .Z(
        P1_U3566) );
  MUX2_X1 U10409 ( .A(n9554), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9557), .Z(
        P1_U3565) );
  MUX2_X1 U10410 ( .A(n9555), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9557), .Z(
        P1_U3564) );
  MUX2_X1 U10411 ( .A(n9556), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9557), .Z(
        P1_U3563) );
  MUX2_X1 U10412 ( .A(n10513), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9557), .Z(
        P1_U3562) );
  MUX2_X1 U10413 ( .A(n10474), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9557), .Z(
        P1_U3561) );
  MUX2_X1 U10414 ( .A(n10515), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9557), .Z(
        P1_U3560) );
  MUX2_X1 U10415 ( .A(n10475), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9557), .Z(
        P1_U3559) );
  MUX2_X1 U10416 ( .A(n6779), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9557), .Z(
        P1_U3558) );
  MUX2_X1 U10417 ( .A(n10356), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9557), .Z(
        P1_U3557) );
  MUX2_X1 U10418 ( .A(n9765), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9557), .Z(
        P1_U3556) );
  NAND2_X1 U10419 ( .A1(n9563), .A2(n9564), .ZN(n9562) );
  XNOR2_X1 U10420 ( .A(n9562), .B(n9778), .ZN(n9780) );
  NAND2_X1 U10421 ( .A1(n9559), .A2(n9558), .ZN(n9783) );
  NOR2_X1 U10422 ( .A1(n10498), .A2(n9783), .ZN(n9566) );
  AOI21_X1 U10423 ( .B1(n10498), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9566), .ZN(
        n9561) );
  NAND2_X1 U10424 ( .A1(n9778), .A2(n9702), .ZN(n9560) );
  OAI211_X1 U10425 ( .C1(n9780), .C2(n10333), .A(n9561), .B(n9560), .ZN(
        P1_U3261) );
  OAI21_X1 U10426 ( .B1(n9563), .B2(n9564), .A(n9562), .ZN(n9784) );
  NOR2_X1 U10427 ( .A1(n9564), .A2(n10538), .ZN(n9565) );
  AOI211_X1 U10428 ( .C1(n10498), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9566), .B(
        n9565), .ZN(n9567) );
  OAI21_X1 U10429 ( .B1(n10333), .B2(n9784), .A(n9567), .ZN(P1_U3262) );
  NAND2_X1 U10430 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  NAND2_X1 U10431 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  NAND2_X1 U10432 ( .A1(n9575), .A2(n9574), .ZN(n9580) );
  NAND2_X1 U10433 ( .A1(n9576), .A2(n10516), .ZN(n9577) );
  OAI21_X1 U10434 ( .B1(n9578), .B2(n9745), .A(n9577), .ZN(n9579) );
  AOI21_X1 U10435 ( .B1(n9580), .B2(n10473), .A(n9579), .ZN(n9581) );
  NAND2_X1 U10436 ( .A1(n9795), .A2(n10539), .ZN(n9590) );
  NAND2_X1 U10437 ( .A1(n9790), .A2(n5162), .ZN(n9582) );
  INV_X1 U10438 ( .A(n9584), .ZN(n9585) );
  AOI22_X1 U10439 ( .A1(n9585), .A2(n10544), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10498), .ZN(n9586) );
  OAI21_X1 U10440 ( .B1(n9587), .B2(n10538), .A(n9586), .ZN(n9588) );
  AOI21_X1 U10441 ( .B1(n9791), .B2(n10534), .A(n9588), .ZN(n9589) );
  OAI211_X1 U10442 ( .C1(n9793), .C2(n9757), .A(n9590), .B(n9589), .ZN(
        P1_U3263) );
  XNOR2_X1 U10443 ( .A(n9591), .B(n9595), .ZN(n9800) );
  AOI21_X1 U10444 ( .B1(n9796), .B2(n5163), .A(n5159), .ZN(n9797) );
  AOI22_X1 U10445 ( .A1(n9592), .A2(n10544), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10498), .ZN(n9593) );
  OAI21_X1 U10446 ( .B1(n9594), .B2(n10538), .A(n9593), .ZN(n9603) );
  AOI21_X1 U10447 ( .B1(n9596), .B2(n9595), .A(n10518), .ZN(n9601) );
  OAI22_X1 U10448 ( .A1(n9598), .A2(n9745), .B1(n9597), .B2(n9743), .ZN(n9599)
         );
  AOI21_X1 U10449 ( .B1(n9601), .B2(n9600), .A(n9599), .ZN(n9799) );
  NOR2_X1 U10450 ( .A1(n9799), .A2(n10498), .ZN(n9602) );
  AOI211_X1 U10451 ( .C1(n10534), .C2(n9797), .A(n9603), .B(n9602), .ZN(n9604)
         );
  OAI21_X1 U10452 ( .B1(n9800), .B2(n9718), .A(n9604), .ZN(P1_U3264) );
  NAND2_X1 U10453 ( .A1(n9639), .A2(n9605), .ZN(n9607) );
  AND2_X1 U10454 ( .A1(n9607), .A2(n9606), .ZN(n9608) );
  XNOR2_X1 U10455 ( .A(n9608), .B(n9617), .ZN(n9810) );
  INV_X1 U10456 ( .A(n9633), .ZN(n9611) );
  INV_X1 U10457 ( .A(n9609), .ZN(n9610) );
  AOI21_X1 U10458 ( .B1(n9806), .B2(n9611), .A(n9610), .ZN(n9807) );
  AOI22_X1 U10459 ( .A1(n9612), .A2(n10544), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10498), .ZN(n9613) );
  OAI21_X1 U10460 ( .B1(n9614), .B2(n10538), .A(n9613), .ZN(n9621) );
  OAI21_X1 U10461 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(n9619) );
  AOI222_X1 U10462 ( .A1(n10473), .A2(n9619), .B1(n9618), .B2(n10514), .C1(
        n9654), .C2(n10516), .ZN(n9809) );
  NOR2_X1 U10463 ( .A1(n9809), .A2(n10498), .ZN(n9620) );
  AOI211_X1 U10464 ( .C1(n9807), .C2(n10534), .A(n9621), .B(n9620), .ZN(n9622)
         );
  OAI21_X1 U10465 ( .B1(n9810), .B2(n9718), .A(n9622), .ZN(P1_U3266) );
  NAND2_X1 U10466 ( .A1(n9639), .A2(n9623), .ZN(n9624) );
  XNOR2_X1 U10467 ( .A(n9624), .B(n9629), .ZN(n9815) );
  AOI22_X1 U10468 ( .A1(n9812), .A2(n9702), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n10498), .ZN(n9638) );
  OR2_X1 U10469 ( .A1(n9649), .A2(n9625), .ZN(n9650) );
  AND2_X1 U10470 ( .A1(n9650), .A2(n9626), .ZN(n9630) );
  NAND2_X1 U10471 ( .A1(n9650), .A2(n9627), .ZN(n9628) );
  OAI21_X1 U10472 ( .B1(n9630), .B2(n9629), .A(n9628), .ZN(n9632) );
  AOI222_X1 U10473 ( .A1(n10473), .A2(n9632), .B1(n9631), .B2(n10514), .C1(
        n9670), .C2(n10516), .ZN(n9814) );
  AOI211_X1 U10474 ( .C1(n9812), .C2(n9642), .A(n10565), .B(n9633), .ZN(n9811)
         );
  AOI22_X1 U10475 ( .A1(n9811), .A2(n9697), .B1(n10544), .B2(n9634), .ZN(n9635) );
  AOI21_X1 U10476 ( .B1(n9814), .B2(n9635), .A(n10498), .ZN(n9636) );
  INV_X1 U10477 ( .A(n9636), .ZN(n9637) );
  OAI211_X1 U10478 ( .C1(n9815), .C2(n9718), .A(n9638), .B(n9637), .ZN(
        P1_U3267) );
  INV_X1 U10479 ( .A(n9639), .ZN(n9640) );
  AOI21_X1 U10480 ( .B1(n9651), .B2(n9641), .A(n9640), .ZN(n9820) );
  INV_X1 U10481 ( .A(n9662), .ZN(n9644) );
  INV_X1 U10482 ( .A(n9642), .ZN(n9643) );
  AOI21_X1 U10483 ( .B1(n9816), .B2(n9644), .A(n9643), .ZN(n9817) );
  INV_X1 U10484 ( .A(n9645), .ZN(n9646) );
  AOI22_X1 U10485 ( .A1(n9646), .A2(n10544), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10498), .ZN(n9647) );
  OAI21_X1 U10486 ( .B1(n9648), .B2(n10538), .A(n9647), .ZN(n9658) );
  INV_X1 U10487 ( .A(n9649), .ZN(n9652) );
  OAI211_X1 U10488 ( .C1(n9652), .C2(n9651), .A(n9650), .B(n10473), .ZN(n9656)
         );
  AOI22_X1 U10489 ( .A1(n9654), .A2(n10514), .B1(n10516), .B2(n9653), .ZN(
        n9655) );
  AND2_X1 U10490 ( .A1(n9656), .A2(n9655), .ZN(n9819) );
  NOR2_X1 U10491 ( .A1(n9819), .A2(n10498), .ZN(n9657) );
  AOI211_X1 U10492 ( .C1(n9817), .C2(n10534), .A(n9658), .B(n9657), .ZN(n9659)
         );
  OAI21_X1 U10493 ( .B1(n9820), .B2(n9718), .A(n9659), .ZN(P1_U3268) );
  XNOR2_X1 U10494 ( .A(n9661), .B(n9660), .ZN(n9825) );
  AOI21_X1 U10495 ( .B1(n9821), .B2(n9682), .A(n9662), .ZN(n9822) );
  INV_X1 U10496 ( .A(n9821), .ZN(n9666) );
  INV_X1 U10497 ( .A(n9663), .ZN(n9664) );
  AOI22_X1 U10498 ( .A1(n9664), .A2(n10544), .B1(n10498), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9665) );
  OAI21_X1 U10499 ( .B1(n9666), .B2(n10538), .A(n9665), .ZN(n9672) );
  XNOR2_X1 U10500 ( .A(n9668), .B(n9667), .ZN(n9669) );
  AOI222_X1 U10501 ( .A1(n9693), .A2(n10516), .B1(n9670), .B2(n10514), .C1(
        n10473), .C2(n9669), .ZN(n9824) );
  NOR2_X1 U10502 ( .A1(n9824), .A2(n10498), .ZN(n9671) );
  AOI211_X1 U10503 ( .C1(n9822), .C2(n10534), .A(n9672), .B(n9671), .ZN(n9673)
         );
  OAI21_X1 U10504 ( .B1(n9718), .B2(n9825), .A(n9673), .ZN(P1_U3269) );
  XNOR2_X1 U10505 ( .A(n9674), .B(n9678), .ZN(n9830) );
  AOI22_X1 U10506 ( .A1(n9828), .A2(n9702), .B1(n10498), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U10507 ( .A1(n9675), .A2(n9676), .ZN(n9677) );
  XOR2_X1 U10508 ( .A(n9678), .B(n9677), .Z(n9679) );
  OAI222_X1 U10509 ( .A1(n9745), .A2(n9681), .B1(n9743), .B2(n9680), .C1(
        n10518), .C2(n9679), .ZN(n9826) );
  INV_X1 U10510 ( .A(n9682), .ZN(n9683) );
  AOI211_X1 U10511 ( .C1(n9828), .C2(n9690), .A(n10565), .B(n9683), .ZN(n9827)
         );
  INV_X1 U10512 ( .A(n9827), .ZN(n9686) );
  INV_X1 U10513 ( .A(n9684), .ZN(n9685) );
  OAI22_X1 U10514 ( .A1(n9686), .A2(n10493), .B1(n10488), .B2(n9685), .ZN(
        n9687) );
  OAI21_X1 U10515 ( .B1(n9826), .B2(n9687), .A(n10539), .ZN(n9688) );
  OAI211_X1 U10516 ( .C1(n9830), .C2(n9718), .A(n9689), .B(n9688), .ZN(
        P1_U3270) );
  INV_X1 U10517 ( .A(n9690), .ZN(n9691) );
  AOI211_X1 U10518 ( .C1(n9833), .C2(n5169), .A(n10565), .B(n9691), .ZN(n9832)
         );
  XNOR2_X1 U10519 ( .A(n9692), .B(n9694), .ZN(n9836) );
  AOI22_X1 U10520 ( .A1(n9693), .A2(n10514), .B1(n10516), .B2(n9723), .ZN(
        n9696) );
  OAI211_X1 U10521 ( .C1(n9694), .C2(n4912), .A(n9675), .B(n10473), .ZN(n9695)
         );
  OAI211_X1 U10522 ( .C1(n9836), .C2(n10526), .A(n9696), .B(n9695), .ZN(n9831)
         );
  AOI21_X1 U10523 ( .B1(n9832), .B2(n9697), .A(n9831), .ZN(n9704) );
  INV_X1 U10524 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9699) );
  OAI22_X1 U10525 ( .A1(n10539), .A2(n9699), .B1(n9698), .B2(n10488), .ZN(
        n9701) );
  NOR2_X1 U10526 ( .A1(n9836), .A2(n9757), .ZN(n9700) );
  AOI211_X1 U10527 ( .C1(n9702), .C2(n9833), .A(n9701), .B(n9700), .ZN(n9703)
         );
  OAI21_X1 U10528 ( .B1(n9704), .B2(n10498), .A(n9703), .ZN(P1_U3271) );
  XNOR2_X1 U10529 ( .A(n9706), .B(n9705), .ZN(n9841) );
  AOI21_X1 U10530 ( .B1(n9837), .B2(n9730), .A(n9707), .ZN(n9838) );
  INV_X1 U10531 ( .A(n9708), .ZN(n9709) );
  AOI22_X1 U10532 ( .A1(n10498), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9709), 
        .B2(n10544), .ZN(n9710) );
  OAI21_X1 U10533 ( .B1(n5167), .B2(n10538), .A(n9710), .ZN(n9716) );
  OAI21_X1 U10534 ( .B1(n4889), .B2(n5415), .A(n9711), .ZN(n9714) );
  AOI222_X1 U10535 ( .A1(n10473), .A2(n9714), .B1(n9713), .B2(n10514), .C1(
        n9712), .C2(n10516), .ZN(n9840) );
  NOR2_X1 U10536 ( .A1(n9840), .A2(n10498), .ZN(n9715) );
  AOI211_X1 U10537 ( .C1(n9838), .C2(n10534), .A(n9716), .B(n9715), .ZN(n9717)
         );
  OAI21_X1 U10538 ( .B1(n9718), .B2(n9841), .A(n9717), .ZN(P1_U3272) );
  OAI21_X1 U10539 ( .B1(n9721), .B2(n9720), .A(n9719), .ZN(n9847) );
  AOI22_X1 U10540 ( .A1(n9723), .A2(n10514), .B1(n9722), .B2(n10516), .ZN(
        n9729) );
  OR2_X1 U10541 ( .A1(n9741), .A2(n9742), .ZN(n9739) );
  NAND2_X1 U10542 ( .A1(n9739), .A2(n9724), .ZN(n9726) );
  OAI211_X1 U10543 ( .C1(n9727), .C2(n9726), .A(n9725), .B(n10473), .ZN(n9728)
         );
  OAI211_X1 U10544 ( .C1(n9847), .C2(n10526), .A(n9729), .B(n9728), .ZN(n9842)
         );
  NAND2_X1 U10545 ( .A1(n9842), .A2(n10539), .ZN(n9737) );
  INV_X1 U10546 ( .A(n9730), .ZN(n9731) );
  AOI21_X1 U10547 ( .B1(n9843), .B2(n9750), .A(n9731), .ZN(n9844) );
  INV_X1 U10548 ( .A(n9843), .ZN(n9732) );
  NOR2_X1 U10549 ( .A1(n9732), .A2(n10538), .ZN(n9735) );
  OAI22_X1 U10550 ( .A1(n10539), .A2(n6353), .B1(n9733), .B2(n10488), .ZN(
        n9734) );
  AOI211_X1 U10551 ( .C1(n9844), .C2(n10534), .A(n9735), .B(n9734), .ZN(n9736)
         );
  OAI211_X1 U10552 ( .C1(n9847), .C2(n9757), .A(n9737), .B(n9736), .ZN(
        P1_U3273) );
  OAI21_X1 U10553 ( .B1(n4923), .B2(n9742), .A(n9738), .ZN(n9756) );
  INV_X1 U10554 ( .A(n9739), .ZN(n9740) );
  AOI211_X1 U10555 ( .C1(n9742), .C2(n9741), .A(n10518), .B(n9740), .ZN(n9748)
         );
  OAI22_X1 U10556 ( .A1(n9746), .A2(n9745), .B1(n9744), .B2(n9743), .ZN(n9747)
         );
  AOI211_X1 U10557 ( .C1(n9756), .C2(n9764), .A(n9748), .B(n9747), .ZN(n9851)
         );
  INV_X1 U10558 ( .A(n9749), .ZN(n9752) );
  INV_X1 U10559 ( .A(n9750), .ZN(n9751) );
  AOI21_X1 U10560 ( .B1(n9848), .B2(n9752), .A(n9751), .ZN(n9849) );
  AOI22_X1 U10561 ( .A1(n10498), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9753), 
        .B2(n10544), .ZN(n9754) );
  OAI21_X1 U10562 ( .B1(n9755), .B2(n10538), .A(n9754), .ZN(n9759) );
  INV_X1 U10563 ( .A(n9756), .ZN(n9852) );
  NOR2_X1 U10564 ( .A1(n9852), .A2(n9757), .ZN(n9758) );
  AOI211_X1 U10565 ( .C1(n9849), .C2(n10534), .A(n9759), .B(n9758), .ZN(n9760)
         );
  OAI21_X1 U10566 ( .B1(n10498), .B2(n9851), .A(n9760), .ZN(P1_U3274) );
  XNOR2_X1 U10567 ( .A(n9504), .B(n9762), .ZN(n9768) );
  OAI21_X1 U10568 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n10388) );
  NAND2_X1 U10569 ( .A1(n10388), .A2(n9764), .ZN(n9767) );
  AOI22_X1 U10570 ( .A1(n10514), .A2(n6779), .B1(n10516), .B2(n9765), .ZN(
        n9766) );
  OAI211_X1 U10571 ( .C1(n10518), .C2(n9768), .A(n9767), .B(n9766), .ZN(n10386) );
  MUX2_X1 U10572 ( .A(n10386), .B(P1_REG2_REG_2__SCAN_IN), .S(n10498), .Z(
        n9769) );
  INV_X1 U10573 ( .A(n9769), .ZN(n9777) );
  NAND2_X1 U10574 ( .A1(n10349), .A2(n6697), .ZN(n9770) );
  AND2_X1 U10575 ( .A1(n9771), .A2(n9770), .ZN(n10383) );
  NAND2_X1 U10576 ( .A1(n10534), .A2(n10383), .ZN(n9773) );
  NAND2_X1 U10577 ( .A1(n10544), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9772) );
  OAI211_X1 U10578 ( .C1(n10385), .C2(n10538), .A(n9773), .B(n9772), .ZN(n9774) );
  INV_X1 U10579 ( .A(n9774), .ZN(n9776) );
  NAND2_X1 U10580 ( .A1(n10535), .A2(n10388), .ZN(n9775) );
  NAND3_X1 U10581 ( .A1(n9777), .A2(n9776), .A3(n9775), .ZN(P1_U3289) );
  NAND2_X1 U10582 ( .A1(n9778), .A2(n10549), .ZN(n9779) );
  OAI211_X1 U10583 ( .C1(n9780), .C2(n10565), .A(n9783), .B(n9779), .ZN(n9882)
         );
  MUX2_X1 U10584 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9882), .S(n10591), .Z(
        P1_U3554) );
  NAND2_X1 U10585 ( .A1(n9781), .A2(n10549), .ZN(n9782) );
  OAI211_X1 U10586 ( .C1(n9784), .C2(n10565), .A(n9783), .B(n9782), .ZN(n9883)
         );
  MUX2_X1 U10587 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9883), .S(n10591), .Z(
        P1_U3553) );
  AOI22_X1 U10588 ( .A1(n9791), .A2(n10477), .B1(n10549), .B2(n9790), .ZN(
        n9792) );
  OAI21_X1 U10589 ( .B1(n9793), .B2(n10552), .A(n9792), .ZN(n9794) );
  OR2_X2 U10590 ( .A1(n9795), .A2(n9794), .ZN(n9884) );
  AOI22_X1 U10591 ( .A1(n9797), .A2(n10477), .B1(n10549), .B2(n9796), .ZN(
        n9798) );
  OAI211_X1 U10592 ( .C1(n9800), .C2(n9863), .A(n9799), .B(n9798), .ZN(n9885)
         );
  MUX2_X1 U10593 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9885), .S(n10591), .Z(
        P1_U3550) );
  AOI22_X1 U10594 ( .A1(n9802), .A2(n10477), .B1(n10549), .B2(n9801), .ZN(
        n9803) );
  OAI211_X1 U10595 ( .C1(n9805), .C2(n10552), .A(n9804), .B(n9803), .ZN(n9886)
         );
  MUX2_X1 U10596 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9886), .S(n10591), .Z(
        P1_U3549) );
  AOI22_X1 U10597 ( .A1(n9807), .A2(n10477), .B1(n10549), .B2(n9806), .ZN(
        n9808) );
  OAI211_X1 U10598 ( .C1(n9810), .C2(n9863), .A(n9809), .B(n9808), .ZN(n9887)
         );
  MUX2_X1 U10599 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9887), .S(n10591), .Z(
        P1_U3548) );
  AOI21_X1 U10600 ( .B1(n10549), .B2(n9812), .A(n9811), .ZN(n9813) );
  OAI211_X1 U10601 ( .C1(n9815), .C2(n9863), .A(n9814), .B(n9813), .ZN(n9888)
         );
  MUX2_X1 U10602 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9888), .S(n10591), .Z(
        P1_U3547) );
  AOI22_X1 U10603 ( .A1(n9817), .A2(n10477), .B1(n10549), .B2(n9816), .ZN(
        n9818) );
  OAI211_X1 U10604 ( .C1(n9820), .C2(n9863), .A(n9819), .B(n9818), .ZN(n9889)
         );
  MUX2_X1 U10605 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9889), .S(n10591), .Z(
        P1_U3546) );
  AOI22_X1 U10606 ( .A1(n9822), .A2(n10477), .B1(n10549), .B2(n9821), .ZN(
        n9823) );
  OAI211_X1 U10607 ( .C1(n9825), .C2(n9863), .A(n9824), .B(n9823), .ZN(n9890)
         );
  MUX2_X1 U10608 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9890), .S(n10591), .Z(
        P1_U3545) );
  AOI211_X1 U10609 ( .C1(n10549), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9829)
         );
  OAI21_X1 U10610 ( .B1(n9863), .B2(n9830), .A(n9829), .ZN(n9891) );
  MUX2_X1 U10611 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9891), .S(n10591), .Z(
        P1_U3544) );
  INV_X1 U10612 ( .A(n9831), .ZN(n9835) );
  AOI21_X1 U10613 ( .B1(n10549), .B2(n9833), .A(n9832), .ZN(n9834) );
  OAI211_X1 U10614 ( .C1(n9836), .C2(n10552), .A(n9835), .B(n9834), .ZN(n9892)
         );
  MUX2_X1 U10615 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9892), .S(n10591), .Z(
        P1_U3543) );
  AOI22_X1 U10616 ( .A1(n9838), .A2(n10477), .B1(n10549), .B2(n9837), .ZN(
        n9839) );
  OAI211_X1 U10617 ( .C1(n9841), .C2(n9863), .A(n9840), .B(n9839), .ZN(n9893)
         );
  MUX2_X1 U10618 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9893), .S(n10591), .Z(
        P1_U3542) );
  INV_X1 U10619 ( .A(n9842), .ZN(n9846) );
  AOI22_X1 U10620 ( .A1(n9844), .A2(n10477), .B1(n10549), .B2(n9843), .ZN(
        n9845) );
  OAI211_X1 U10621 ( .C1(n10552), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9894)
         );
  MUX2_X1 U10622 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9894), .S(n10591), .Z(
        P1_U3541) );
  AOI22_X1 U10623 ( .A1(n9849), .A2(n10477), .B1(n10549), .B2(n9848), .ZN(
        n9850) );
  OAI211_X1 U10624 ( .C1(n9852), .C2(n10552), .A(n9851), .B(n9850), .ZN(n9895)
         );
  MUX2_X1 U10625 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9895), .S(n10591), .Z(
        P1_U3540) );
  AOI211_X1 U10626 ( .C1(n10549), .C2(n9855), .A(n9854), .B(n9853), .ZN(n9856)
         );
  OAI21_X1 U10627 ( .B1(n9857), .B2(n9863), .A(n9856), .ZN(n9896) );
  MUX2_X1 U10628 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9896), .S(n10591), .Z(
        P1_U3539) );
  AOI22_X1 U10629 ( .A1(n9859), .A2(n10477), .B1(n10549), .B2(n9858), .ZN(
        n9860) );
  OAI211_X1 U10630 ( .C1(n10552), .C2(n9862), .A(n9861), .B(n9860), .ZN(n9897)
         );
  MUX2_X1 U10631 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9897), .S(n10591), .Z(
        P1_U3538) );
  INV_X1 U10632 ( .A(n9863), .ZN(n10480) );
  NAND2_X1 U10633 ( .A1(n9864), .A2(n10480), .ZN(n9870) );
  OAI21_X1 U10634 ( .B1(n9866), .B2(n10582), .A(n9865), .ZN(n9867) );
  NOR2_X1 U10635 ( .A1(n9868), .A2(n9867), .ZN(n9869) );
  NAND2_X1 U10636 ( .A1(n9870), .A2(n9869), .ZN(n9898) );
  MUX2_X1 U10637 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9898), .S(n10591), .Z(
        P1_U3537) );
  AOI22_X1 U10638 ( .A1(n9872), .A2(n10477), .B1(n10549), .B2(n9871), .ZN(
        n9873) );
  OAI211_X1 U10639 ( .C1(n9875), .C2(n10552), .A(n9874), .B(n9873), .ZN(n9899)
         );
  MUX2_X1 U10640 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9899), .S(n10591), .Z(
        P1_U3536) );
  AOI21_X1 U10641 ( .B1(n10549), .B2(n9877), .A(n9876), .ZN(n9878) );
  OAI211_X1 U10642 ( .C1(n10552), .C2(n9880), .A(n9879), .B(n9878), .ZN(n9900)
         );
  MUX2_X1 U10643 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9900), .S(n10591), .Z(
        P1_U3535) );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9881), .S(n10591), .Z(
        P1_U3523) );
  MUX2_X1 U10645 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9882), .S(n10595), .Z(
        P1_U3522) );
  MUX2_X1 U10646 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9883), .S(n10595), .Z(
        P1_U3521) );
  MUX2_X1 U10647 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9885), .S(n10595), .Z(
        P1_U3518) );
  MUX2_X1 U10648 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9886), .S(n10595), .Z(
        P1_U3517) );
  MUX2_X1 U10649 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9887), .S(n10595), .Z(
        P1_U3516) );
  MUX2_X1 U10650 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9888), .S(n10595), .Z(
        P1_U3515) );
  MUX2_X1 U10651 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9889), .S(n10595), .Z(
        P1_U3514) );
  MUX2_X1 U10652 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9890), .S(n10595), .Z(
        P1_U3513) );
  MUX2_X1 U10653 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9891), .S(n10595), .Z(
        P1_U3512) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9892), .S(n10595), .Z(
        P1_U3511) );
  MUX2_X1 U10655 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9893), .S(n10595), .Z(
        P1_U3510) );
  MUX2_X1 U10656 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9894), .S(n10595), .Z(
        P1_U3508) );
  MUX2_X1 U10657 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9895), .S(n10595), .Z(
        P1_U3505) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9896), .S(n10595), .Z(
        P1_U3502) );
  MUX2_X1 U10659 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9897), .S(n10595), .Z(
        P1_U3499) );
  MUX2_X1 U10660 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9898), .S(n10595), .Z(
        P1_U3496) );
  MUX2_X1 U10661 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9899), .S(n10595), .Z(
        P1_U3493) );
  MUX2_X1 U10662 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9900), .S(n10595), .Z(
        P1_U3490) );
  NOR2_X1 U10663 ( .A1(n9902), .A2(n9901), .ZN(n9922) );
  CLKBUF_X1 U10664 ( .A(n9922), .Z(n9936) );
  MUX2_X1 U10665 ( .A(P1_D_REG_0__SCAN_IN), .B(n9903), .S(n9936), .Z(P1_U3440)
         );
  MUX2_X1 U10666 ( .A(n9904), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10667 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9905) );
  NOR2_X1 U10668 ( .A1(n9922), .A2(n9905), .ZN(P1_U3321) );
  INV_X1 U10669 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9906) );
  NOR2_X1 U10670 ( .A1(n9922), .A2(n9906), .ZN(P1_U3320) );
  INV_X1 U10671 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U10672 ( .A1(n9936), .A2(n9907), .ZN(P1_U3319) );
  INV_X1 U10673 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U10674 ( .A1(n9936), .A2(n9908), .ZN(P1_U3318) );
  INV_X1 U10675 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9909) );
  NOR2_X1 U10676 ( .A1(n9936), .A2(n9909), .ZN(P1_U3317) );
  INV_X1 U10677 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9910) );
  NOR2_X1 U10678 ( .A1(n9936), .A2(n9910), .ZN(P1_U3316) );
  INV_X1 U10679 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9911) );
  NOR2_X1 U10680 ( .A1(n9936), .A2(n9911), .ZN(P1_U3315) );
  INV_X1 U10681 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U10682 ( .A1(n9936), .A2(n9912), .ZN(P1_U3314) );
  INV_X1 U10683 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9913) );
  NOR2_X1 U10684 ( .A1(n9936), .A2(n9913), .ZN(P1_U3313) );
  INV_X1 U10685 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9914) );
  NOR2_X1 U10686 ( .A1(n9922), .A2(n9914), .ZN(P1_U3312) );
  INV_X1 U10687 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9915) );
  NOR2_X1 U10688 ( .A1(n9922), .A2(n9915), .ZN(P1_U3311) );
  INV_X1 U10689 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9916) );
  NOR2_X1 U10690 ( .A1(n9922), .A2(n9916), .ZN(P1_U3310) );
  INV_X1 U10691 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U10692 ( .A1(n9922), .A2(n9917), .ZN(P1_U3309) );
  INV_X1 U10693 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U10694 ( .A1(n9922), .A2(n9918), .ZN(P1_U3308) );
  INV_X1 U10695 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9919) );
  NOR2_X1 U10696 ( .A1(n9922), .A2(n9919), .ZN(P1_U3307) );
  INV_X1 U10697 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U10698 ( .A1(n9922), .A2(n9920), .ZN(P1_U3306) );
  INV_X1 U10699 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9921) );
  NOR2_X1 U10700 ( .A1(n9922), .A2(n9921), .ZN(P1_U3305) );
  INV_X1 U10701 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9923) );
  NOR2_X1 U10702 ( .A1(n9936), .A2(n9923), .ZN(P1_U3304) );
  INV_X1 U10703 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9924) );
  NOR2_X1 U10704 ( .A1(n9936), .A2(n9924), .ZN(P1_U3303) );
  INV_X1 U10705 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U10706 ( .A1(n9936), .A2(n9925), .ZN(P1_U3302) );
  INV_X1 U10707 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9926) );
  NOR2_X1 U10708 ( .A1(n9936), .A2(n9926), .ZN(P1_U3301) );
  INV_X1 U10709 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9927) );
  NOR2_X1 U10710 ( .A1(n9936), .A2(n9927), .ZN(P1_U3300) );
  INV_X1 U10711 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U10712 ( .A1(n9936), .A2(n9928), .ZN(P1_U3299) );
  INV_X1 U10713 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9929) );
  NOR2_X1 U10714 ( .A1(n9936), .A2(n9929), .ZN(P1_U3298) );
  INV_X1 U10715 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9930) );
  NOR2_X1 U10716 ( .A1(n9936), .A2(n9930), .ZN(P1_U3297) );
  INV_X1 U10717 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9931) );
  NOR2_X1 U10718 ( .A1(n9936), .A2(n9931), .ZN(P1_U3296) );
  INV_X1 U10719 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U10720 ( .A1(n9936), .A2(n9932), .ZN(P1_U3295) );
  INV_X1 U10721 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9933) );
  NOR2_X1 U10722 ( .A1(n9936), .A2(n9933), .ZN(P1_U3294) );
  INV_X1 U10723 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9934) );
  NOR2_X1 U10724 ( .A1(n9936), .A2(n9934), .ZN(P1_U3293) );
  INV_X1 U10725 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9935) );
  NOR2_X1 U10726 ( .A1(n9936), .A2(n9935), .ZN(P1_U3292) );
  INV_X1 U10727 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U10728 ( .A1(n10274), .A2(n9937), .ZN(n10271) );
  AOI22_X1 U10729 ( .A1(n9939), .A2(n10271), .B1(n10274), .B2(n9938), .ZN(
        P2_U3438) );
  AND2_X1 U10730 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10271), .ZN(P2_U3326) );
  AND2_X1 U10731 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10271), .ZN(P2_U3325) );
  AND2_X1 U10732 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10271), .ZN(P2_U3324) );
  AND2_X1 U10733 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10271), .ZN(P2_U3323) );
  AND2_X1 U10734 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10271), .ZN(P2_U3322) );
  AND2_X1 U10735 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10271), .ZN(P2_U3321) );
  AND2_X1 U10736 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10271), .ZN(P2_U3320) );
  AND2_X1 U10737 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10271), .ZN(P2_U3319) );
  AND2_X1 U10738 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10271), .ZN(P2_U3318) );
  AND2_X1 U10739 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10271), .ZN(P2_U3317) );
  AND2_X1 U10740 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10271), .ZN(P2_U3316) );
  AND2_X1 U10741 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10271), .ZN(P2_U3315) );
  AND2_X1 U10742 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10271), .ZN(P2_U3314) );
  AND2_X1 U10743 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10271), .ZN(P2_U3313) );
  AND2_X1 U10744 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10271), .ZN(P2_U3312) );
  AND2_X1 U10745 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10271), .ZN(P2_U3311) );
  AND2_X1 U10746 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10271), .ZN(P2_U3310) );
  AND2_X1 U10747 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10271), .ZN(P2_U3309) );
  AND2_X1 U10748 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10271), .ZN(P2_U3308) );
  AND2_X1 U10749 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10271), .ZN(P2_U3307) );
  AND2_X1 U10750 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10271), .ZN(P2_U3306) );
  AND2_X1 U10751 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10271), .ZN(P2_U3305) );
  AND2_X1 U10752 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10271), .ZN(P2_U3304) );
  AND2_X1 U10753 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10271), .ZN(P2_U3303) );
  AND2_X1 U10754 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10271), .ZN(P2_U3302) );
  AND2_X1 U10755 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10271), .ZN(P2_U3301) );
  AND2_X1 U10756 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10271), .ZN(P2_U3300) );
  AND2_X1 U10757 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10271), .ZN(P2_U3299) );
  AND2_X1 U10758 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10271), .ZN(P2_U3298) );
  AND2_X1 U10759 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10271), .ZN(P2_U3297) );
  XNOR2_X1 U10760 ( .A(n10140), .B(keyinput_62), .ZN(n10147) );
  INV_X1 U10761 ( .A(keyinput_61), .ZN(n10031) );
  INV_X1 U10762 ( .A(keyinput_60), .ZN(n10029) );
  OAI22_X1 U10763 ( .A1(n5785), .A2(keyinput_58), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(keyinput_57), .ZN(n9940) );
  AOI221_X1 U10764 ( .B1(n5785), .B2(keyinput_58), .C1(keyinput_57), .C2(
        P2_REG3_REG_22__SCAN_IN), .A(n9940), .ZN(n10026) );
  OAI22_X1 U10765 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_55), .B1(
        keyinput_54), .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n9941) );
  AOI221_X1 U10766 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(
        P2_REG3_REG_0__SCAN_IN), .C2(keyinput_54), .A(n9941), .ZN(n10023) );
  INV_X1 U10767 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9944) );
  OAI22_X1 U10768 ( .A1(n9944), .A2(keyinput_52), .B1(n9943), .B2(keyinput_51), 
        .ZN(n9942) );
  AOI221_X1 U10769 ( .B1(n9944), .B2(keyinput_52), .C1(keyinput_51), .C2(n9943), .A(n9942), .ZN(n10020) );
  INV_X1 U10770 ( .A(keyinput_46), .ZN(n10012) );
  OAI22_X1 U10771 ( .A1(n10112), .A2(keyinput_45), .B1(keyinput_44), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n9945) );
  AOI221_X1 U10772 ( .B1(n10112), .B2(keyinput_45), .C1(P2_REG3_REG_1__SCAN_IN), .C2(keyinput_44), .A(n9945), .ZN(n10009) );
  INV_X1 U10773 ( .A(SI_5_), .ZN(n10092) );
  INV_X1 U10774 ( .A(keyinput_27), .ZN(n9986) );
  INV_X1 U10775 ( .A(SI_6_), .ZN(n9984) );
  INV_X1 U10776 ( .A(SI_7_), .ZN(n9947) );
  OAI22_X1 U10777 ( .A1(n9947), .A2(keyinput_25), .B1(SI_8_), .B2(keyinput_24), 
        .ZN(n9946) );
  AOI221_X1 U10778 ( .B1(n9947), .B2(keyinput_25), .C1(keyinput_24), .C2(SI_8_), .A(n9946), .ZN(n9982) );
  INV_X1 U10779 ( .A(keyinput_23), .ZN(n9980) );
  INV_X1 U10780 ( .A(keyinput_22), .ZN(n9978) );
  OAI22_X1 U10781 ( .A1(n9949), .A2(keyinput_19), .B1(keyinput_20), .B2(SI_12_), .ZN(n9948) );
  AOI221_X1 U10782 ( .B1(n9949), .B2(keyinput_19), .C1(SI_12_), .C2(
        keyinput_20), .A(n9948), .ZN(n9975) );
  INV_X1 U10783 ( .A(SI_18_), .ZN(n10045) );
  AOI22_X1 U10784 ( .A1(n10045), .A2(keyinput_14), .B1(n10048), .B2(
        keyinput_13), .ZN(n9950) );
  OAI221_X1 U10785 ( .B1(n10045), .B2(keyinput_14), .C1(n10048), .C2(
        keyinput_13), .A(n9950), .ZN(n9973) );
  OAI22_X1 U10786 ( .A1(SI_22_), .A2(keyinput_10), .B1(keyinput_11), .B2(
        SI_21_), .ZN(n9951) );
  AOI221_X1 U10787 ( .B1(SI_22_), .B2(keyinput_10), .C1(SI_21_), .C2(
        keyinput_11), .A(n9951), .ZN(n9966) );
  OAI22_X1 U10788 ( .A1(n10042), .A2(keyinput_12), .B1(keyinput_9), .B2(SI_23_), .ZN(n9952) );
  AOI221_X1 U10789 ( .B1(n10042), .B2(keyinput_12), .C1(SI_23_), .C2(
        keyinput_9), .A(n9952), .ZN(n9965) );
  OAI22_X1 U10790 ( .A1(SI_31_), .A2(keyinput_1), .B1(P2_WR_REG_SCAN_IN), .B2(
        keyinput_0), .ZN(n9953) );
  AOI221_X1 U10791 ( .B1(SI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P2_WR_REG_SCAN_IN), .A(n9953), .ZN(n9959) );
  AOI22_X1 U10792 ( .A1(n9955), .A2(keyinput_5), .B1(keyinput_2), .B2(n10056), 
        .ZN(n9954) );
  OAI221_X1 U10793 ( .B1(n9955), .B2(keyinput_5), .C1(n10056), .C2(keyinput_2), 
        .A(n9954), .ZN(n9958) );
  AOI22_X1 U10794 ( .A1(SI_29_), .A2(keyinput_3), .B1(n10058), .B2(keyinput_4), 
        .ZN(n9956) );
  OAI221_X1 U10795 ( .B1(SI_29_), .B2(keyinput_3), .C1(n10058), .C2(keyinput_4), .A(n9956), .ZN(n9957) );
  NOR3_X1 U10796 ( .A1(n9959), .A2(n9958), .A3(n9957), .ZN(n9962) );
  INV_X1 U10797 ( .A(SI_24_), .ZN(n10068) );
  AOI22_X1 U10798 ( .A1(SI_25_), .A2(keyinput_7), .B1(n10068), .B2(keyinput_8), 
        .ZN(n9960) );
  OAI221_X1 U10799 ( .B1(SI_25_), .B2(keyinput_7), .C1(n10068), .C2(keyinput_8), .A(n9960), .ZN(n9961) );
  AOI211_X1 U10800 ( .C1(SI_26_), .C2(keyinput_6), .A(n9962), .B(n9961), .ZN(
        n9963) );
  OAI21_X1 U10801 ( .B1(SI_26_), .B2(keyinput_6), .A(n9963), .ZN(n9964) );
  NAND3_X1 U10802 ( .A1(n9966), .A2(n9965), .A3(n9964), .ZN(n9972) );
  OAI22_X1 U10803 ( .A1(n9968), .A2(keyinput_17), .B1(keyinput_18), .B2(SI_14_), .ZN(n9967) );
  AOI221_X1 U10804 ( .B1(n9968), .B2(keyinput_17), .C1(SI_14_), .C2(
        keyinput_18), .A(n9967), .ZN(n9971) );
  OAI22_X1 U10805 ( .A1(SI_17_), .A2(keyinput_15), .B1(keyinput_16), .B2(
        SI_16_), .ZN(n9969) );
  AOI221_X1 U10806 ( .B1(SI_17_), .B2(keyinput_15), .C1(SI_16_), .C2(
        keyinput_16), .A(n9969), .ZN(n9970) );
  OAI211_X1 U10807 ( .C1(n9973), .C2(n9972), .A(n9971), .B(n9970), .ZN(n9974)
         );
  AOI22_X1 U10808 ( .A1(n9975), .A2(n9974), .B1(keyinput_21), .B2(SI_11_), 
        .ZN(n9976) );
  OAI21_X1 U10809 ( .B1(keyinput_21), .B2(SI_11_), .A(n9976), .ZN(n9977) );
  OAI221_X1 U10810 ( .B1(SI_10_), .B2(keyinput_22), .C1(n10082), .C2(n9978), 
        .A(n9977), .ZN(n9979) );
  OAI221_X1 U10811 ( .B1(SI_9_), .B2(keyinput_23), .C1(n10086), .C2(n9980), 
        .A(n9979), .ZN(n9981) );
  AOI22_X1 U10812 ( .A1(keyinput_26), .A2(n9984), .B1(n9982), .B2(n9981), .ZN(
        n9983) );
  OAI21_X1 U10813 ( .B1(n9984), .B2(keyinput_26), .A(n9983), .ZN(n9985) );
  OAI221_X1 U10814 ( .B1(SI_5_), .B2(keyinput_27), .C1(n10092), .C2(n9986), 
        .A(n9985), .ZN(n9995) );
  OAI22_X1 U10815 ( .A1(n9988), .A2(keyinput_29), .B1(keyinput_28), .B2(SI_4_), 
        .ZN(n9987) );
  AOI221_X1 U10816 ( .B1(n9988), .B2(keyinput_29), .C1(SI_4_), .C2(keyinput_28), .A(n9987), .ZN(n9994) );
  AOI22_X1 U10817 ( .A1(SI_1_), .A2(keyinput_31), .B1(SI_0_), .B2(keyinput_32), 
        .ZN(n9989) );
  OAI221_X1 U10818 ( .B1(SI_1_), .B2(keyinput_31), .C1(SI_0_), .C2(keyinput_32), .A(n9989), .ZN(n9993) );
  XOR2_X1 U10819 ( .A(n5722), .B(keyinput_35), .Z(n9991) );
  XNOR2_X1 U10820 ( .A(SI_2_), .B(keyinput_30), .ZN(n9990) );
  NAND2_X1 U10821 ( .A1(n9991), .A2(n9990), .ZN(n9992) );
  AOI211_X1 U10822 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n9992), .ZN(n9999)
         );
  OAI22_X1 U10823 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_33), .B1(keyinput_34), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n9996) );
  AOI221_X1 U10824 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_33), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_34), .A(n9996), .ZN(n9998) );
  NOR2_X1 U10825 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_36), .ZN(n9997)
         );
  AOI221_X1 U10826 ( .B1(n9999), .B2(n9998), .C1(keyinput_36), .C2(
        P2_REG3_REG_27__SCAN_IN), .A(n9997), .ZN(n10007) );
  AOI22_X1 U10827 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_38), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .ZN(n10000) );
  OAI221_X1 U10828 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_37), .A(n10000), .ZN(n10006) );
  OAI22_X1 U10829 ( .A1(n10002), .A2(keyinput_42), .B1(keyinput_41), .B2(
        P2_REG3_REG_19__SCAN_IN), .ZN(n10001) );
  AOI221_X1 U10830 ( .B1(n10002), .B2(keyinput_42), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_41), .A(n10001), .ZN(n10005) );
  OAI22_X1 U10831 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_40), .B1(
        keyinput_39), .B2(P2_REG3_REG_10__SCAN_IN), .ZN(n10003) );
  AOI221_X1 U10832 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_39), .A(n10003), .ZN(n10004) );
  OAI211_X1 U10833 ( .C1(n10007), .C2(n10006), .A(n10005), .B(n10004), .ZN(
        n10008) );
  OAI211_X1 U10834 ( .C1(P2_REG3_REG_8__SCAN_IN), .C2(keyinput_43), .A(n10009), 
        .B(n10008), .ZN(n10010) );
  AOI21_X1 U10835 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .A(n10010), 
        .ZN(n10011) );
  AOI221_X1 U10836 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .C1(
        n10117), .C2(n10012), .A(n10011), .ZN(n10018) );
  AOI22_X1 U10837 ( .A1(n8816), .A2(keyinput_47), .B1(n10014), .B2(keyinput_48), .ZN(n10013) );
  OAI221_X1 U10838 ( .B1(n8816), .B2(keyinput_47), .C1(n10014), .C2(
        keyinput_48), .A(n10013), .ZN(n10017) );
  OAI22_X1 U10839 ( .A1(n5904), .A2(keyinput_50), .B1(keyinput_49), .B2(
        P2_REG3_REG_5__SCAN_IN), .ZN(n10015) );
  AOI221_X1 U10840 ( .B1(n5904), .B2(keyinput_50), .C1(P2_REG3_REG_5__SCAN_IN), 
        .C2(keyinput_49), .A(n10015), .ZN(n10016) );
  OAI21_X1 U10841 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(n10019) );
  AOI22_X1 U10842 ( .A1(keyinput_53), .A2(n5756), .B1(n10020), .B2(n10019), 
        .ZN(n10021) );
  OAI21_X1 U10843 ( .B1(n5756), .B2(keyinput_53), .A(n10021), .ZN(n10022) );
  AOI22_X1 U10844 ( .A1(n10023), .A2(n10022), .B1(keyinput_56), .B2(
        P2_REG3_REG_13__SCAN_IN), .ZN(n10024) );
  OAI21_X1 U10845 ( .B1(keyinput_56), .B2(P2_REG3_REG_13__SCAN_IN), .A(n10024), 
        .ZN(n10025) );
  AOI22_X1 U10846 ( .A1(keyinput_59), .A2(n10403), .B1(n10026), .B2(n10025), 
        .ZN(n10027) );
  OAI21_X1 U10847 ( .B1(n10403), .B2(keyinput_59), .A(n10027), .ZN(n10028) );
  OAI221_X1 U10848 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(n10029), .C1(n10134), 
        .C2(keyinput_60), .A(n10028), .ZN(n10030) );
  OAI221_X1 U10849 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(n10031), .C1(n10137), 
        .C2(keyinput_61), .A(n10030), .ZN(n10146) );
  INV_X1 U10850 ( .A(keyinput_126), .ZN(n10139) );
  INV_X1 U10851 ( .A(keyinput_125), .ZN(n10136) );
  INV_X1 U10852 ( .A(keyinput_124), .ZN(n10133) );
  OAI22_X1 U10853 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_122), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .ZN(n10032) );
  AOI221_X1 U10854 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        keyinput_121), .C2(P2_REG3_REG_22__SCAN_IN), .A(n10032), .ZN(n10130)
         );
  OAI22_X1 U10855 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_119), .B1(
        keyinput_118), .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n10033) );
  AOI221_X1 U10856 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        P2_REG3_REG_0__SCAN_IN), .C2(keyinput_118), .A(n10033), .ZN(n10127) );
  AOI22_X1 U10857 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_115), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_116), .ZN(n10034) );
  OAI221_X1 U10858 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_116), .A(n10034), .ZN(n10125) );
  OAI22_X1 U10859 ( .A1(n8816), .A2(keyinput_111), .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_112), .ZN(n10035) );
  AOI221_X1 U10860 ( .B1(n8816), .B2(keyinput_111), .C1(keyinput_112), .C2(
        P2_REG3_REG_16__SCAN_IN), .A(n10035), .ZN(n10122) );
  INV_X1 U10861 ( .A(keyinput_110), .ZN(n10118) );
  OAI22_X1 U10862 ( .A1(n10037), .A2(keyinput_101), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .ZN(n10036) );
  AOI221_X1 U10863 ( .B1(n10037), .B2(keyinput_101), .C1(keyinput_102), .C2(
        P2_REG3_REG_23__SCAN_IN), .A(n10036), .ZN(n10110) );
  INV_X1 U10864 ( .A(keyinput_100), .ZN(n10103) );
  INV_X1 U10865 ( .A(keyinput_91), .ZN(n10091) );
  AOI22_X1 U10866 ( .A1(SI_7_), .A2(keyinput_89), .B1(n10039), .B2(keyinput_88), .ZN(n10038) );
  OAI221_X1 U10867 ( .B1(SI_7_), .B2(keyinput_89), .C1(n10039), .C2(
        keyinput_88), .A(n10038), .ZN(n10088) );
  INV_X1 U10868 ( .A(keyinput_87), .ZN(n10085) );
  INV_X1 U10869 ( .A(keyinput_86), .ZN(n10083) );
  AOI22_X1 U10870 ( .A1(SI_12_), .A2(keyinput_84), .B1(SI_13_), .B2(
        keyinput_83), .ZN(n10040) );
  OAI221_X1 U10871 ( .B1(SI_12_), .B2(keyinput_84), .C1(SI_13_), .C2(
        keyinput_83), .A(n10040), .ZN(n10078) );
  AOI22_X1 U10872 ( .A1(n10043), .A2(keyinput_75), .B1(keyinput_76), .B2(
        n10042), .ZN(n10041) );
  OAI221_X1 U10873 ( .B1(n10043), .B2(keyinput_75), .C1(n10042), .C2(
        keyinput_76), .A(n10041), .ZN(n10052) );
  AOI22_X1 U10874 ( .A1(n10046), .A2(keyinput_73), .B1(keyinput_78), .B2(
        n10045), .ZN(n10044) );
  OAI221_X1 U10875 ( .B1(n10046), .B2(keyinput_73), .C1(n10045), .C2(
        keyinput_78), .A(n10044), .ZN(n10051) );
  AOI22_X1 U10876 ( .A1(n10049), .A2(keyinput_74), .B1(keyinput_77), .B2(
        n10048), .ZN(n10047) );
  OAI221_X1 U10877 ( .B1(n10049), .B2(keyinput_74), .C1(n10048), .C2(
        keyinput_77), .A(n10047), .ZN(n10050) );
  NOR3_X1 U10878 ( .A1(n10052), .A2(n10051), .A3(n10050), .ZN(n10076) );
  OAI22_X1 U10879 ( .A1(SI_31_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n10053) );
  AOI221_X1 U10880 ( .B1(SI_31_), .B2(keyinput_65), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_64), .A(n10053), .ZN(n10061) );
  AOI22_X1 U10881 ( .A1(n10056), .A2(keyinput_66), .B1(keyinput_67), .B2(
        n10055), .ZN(n10054) );
  OAI221_X1 U10882 ( .B1(n10056), .B2(keyinput_66), .C1(n10055), .C2(
        keyinput_67), .A(n10054), .ZN(n10060) );
  AOI22_X1 U10883 ( .A1(SI_27_), .A2(keyinput_69), .B1(n10058), .B2(
        keyinput_68), .ZN(n10057) );
  OAI221_X1 U10884 ( .B1(SI_27_), .B2(keyinput_69), .C1(n10058), .C2(
        keyinput_68), .A(n10057), .ZN(n10059) );
  NOR3_X1 U10885 ( .A1(n10061), .A2(n10060), .A3(n10059), .ZN(n10066) );
  AOI22_X1 U10886 ( .A1(n10064), .A2(keyinput_71), .B1(n10063), .B2(
        keyinput_70), .ZN(n10062) );
  OAI221_X1 U10887 ( .B1(n10064), .B2(keyinput_71), .C1(n10063), .C2(
        keyinput_70), .A(n10062), .ZN(n10065) );
  AOI211_X1 U10888 ( .C1(n10068), .C2(keyinput_72), .A(n10066), .B(n10065), 
        .ZN(n10067) );
  OAI21_X1 U10889 ( .B1(n10068), .B2(keyinput_72), .A(n10067), .ZN(n10075) );
  AOI22_X1 U10890 ( .A1(n10071), .A2(keyinput_80), .B1(n10070), .B2(
        keyinput_79), .ZN(n10069) );
  OAI221_X1 U10891 ( .B1(n10071), .B2(keyinput_80), .C1(n10070), .C2(
        keyinput_79), .A(n10069), .ZN(n10074) );
  AOI22_X1 U10892 ( .A1(SI_14_), .A2(keyinput_82), .B1(SI_15_), .B2(
        keyinput_81), .ZN(n10072) );
  OAI221_X1 U10893 ( .B1(SI_14_), .B2(keyinput_82), .C1(SI_15_), .C2(
        keyinput_81), .A(n10072), .ZN(n10073) );
  AOI211_X1 U10894 ( .C1(n10076), .C2(n10075), .A(n10074), .B(n10073), .ZN(
        n10077) );
  OAI22_X1 U10895 ( .A1(keyinput_85), .A2(n10080), .B1(n10078), .B2(n10077), 
        .ZN(n10079) );
  AOI21_X1 U10896 ( .B1(keyinput_85), .B2(n10080), .A(n10079), .ZN(n10081) );
  AOI221_X1 U10897 ( .B1(SI_10_), .B2(n10083), .C1(n10082), .C2(keyinput_86), 
        .A(n10081), .ZN(n10084) );
  AOI221_X1 U10898 ( .B1(SI_9_), .B2(keyinput_87), .C1(n10086), .C2(n10085), 
        .A(n10084), .ZN(n10087) );
  OAI22_X1 U10899 ( .A1(n10088), .A2(n10087), .B1(keyinput_90), .B2(SI_6_), 
        .ZN(n10089) );
  AOI21_X1 U10900 ( .B1(keyinput_90), .B2(SI_6_), .A(n10089), .ZN(n10090) );
  AOI221_X1 U10901 ( .B1(SI_5_), .B2(keyinput_91), .C1(n10092), .C2(n10091), 
        .A(n10090), .ZN(n10099) );
  AOI22_X1 U10902 ( .A1(SI_3_), .A2(keyinput_93), .B1(SI_4_), .B2(keyinput_92), 
        .ZN(n10093) );
  OAI221_X1 U10903 ( .B1(SI_3_), .B2(keyinput_93), .C1(SI_4_), .C2(keyinput_92), .A(n10093), .ZN(n10098) );
  OAI22_X1 U10904 ( .A1(P2_U3152), .A2(keyinput_98), .B1(keyinput_95), .B2(
        SI_1_), .ZN(n10094) );
  AOI221_X1 U10905 ( .B1(P2_U3152), .B2(keyinput_98), .C1(SI_1_), .C2(
        keyinput_95), .A(n10094), .ZN(n10097) );
  OAI22_X1 U10906 ( .A1(n5722), .A2(keyinput_99), .B1(keyinput_96), .B2(SI_0_), 
        .ZN(n10095) );
  AOI221_X1 U10907 ( .B1(n5722), .B2(keyinput_99), .C1(SI_0_), .C2(keyinput_96), .A(n10095), .ZN(n10096) );
  OAI211_X1 U10908 ( .C1(n10099), .C2(n10098), .A(n10097), .B(n10096), .ZN(
        n10102) );
  AOI22_X1 U10909 ( .A1(SI_2_), .A2(keyinput_94), .B1(P2_RD_REG_SCAN_IN), .B2(
        keyinput_97), .ZN(n10100) );
  OAI221_X1 U10910 ( .B1(SI_2_), .B2(keyinput_94), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_97), .A(n10100), .ZN(n10101) );
  OAI222_X1 U10911 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(n10103), .B1(n8785), 
        .B2(keyinput_100), .C1(n10102), .C2(n10101), .ZN(n10109) );
  AOI22_X1 U10912 ( .A1(n10105), .A2(keyinput_103), .B1(keyinput_105), .B2(
        n5931), .ZN(n10104) );
  OAI221_X1 U10913 ( .B1(n10105), .B2(keyinput_103), .C1(n5931), .C2(
        keyinput_105), .A(n10104), .ZN(n10108) );
  AOI22_X1 U10914 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_106), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .ZN(n10106) );
  OAI221_X1 U10915 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_106), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_104), .A(n10106), .ZN(n10107) );
  AOI211_X1 U10916 ( .C1(n10110), .C2(n10109), .A(n10108), .B(n10107), .ZN(
        n10114) );
  AOI22_X1 U10917 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(n10112), .B2(keyinput_109), .ZN(n10111) );
  OAI221_X1 U10918 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        n10112), .C2(keyinput_109), .A(n10111), .ZN(n10113) );
  AOI211_X1 U10919 ( .C1(n10372), .C2(keyinput_108), .A(n10114), .B(n10113), 
        .ZN(n10115) );
  OAI21_X1 U10920 ( .B1(n10372), .B2(keyinput_108), .A(n10115), .ZN(n10116) );
  OAI221_X1 U10921 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(n10118), .C1(n10117), 
        .C2(keyinput_110), .A(n10116), .ZN(n10121) );
  AOI22_X1 U10922 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_113), .B1(n5904), 
        .B2(keyinput_114), .ZN(n10119) );
  OAI221_X1 U10923 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .C1(n5904), .C2(keyinput_114), .A(n10119), .ZN(n10120) );
  AOI21_X1 U10924 ( .B1(n10122), .B2(n10121), .A(n10120), .ZN(n10124) );
  NAND2_X1 U10925 ( .A1(n5756), .A2(keyinput_117), .ZN(n10123) );
  OAI221_X1 U10926 ( .B1(n10125), .B2(n10124), .C1(n5756), .C2(keyinput_117), 
        .A(n10123), .ZN(n10126) );
  AOI22_X1 U10927 ( .A1(n10127), .A2(n10126), .B1(keyinput_120), .B2(
        P2_REG3_REG_13__SCAN_IN), .ZN(n10128) );
  OAI21_X1 U10928 ( .B1(keyinput_120), .B2(P2_REG3_REG_13__SCAN_IN), .A(n10128), .ZN(n10129) );
  AOI22_X1 U10929 ( .A1(keyinput_123), .A2(n10403), .B1(n10130), .B2(n10129), 
        .ZN(n10131) );
  OAI21_X1 U10930 ( .B1(n10403), .B2(keyinput_123), .A(n10131), .ZN(n10132) );
  OAI221_X1 U10931 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(
        n10134), .C2(n10133), .A(n10132), .ZN(n10135) );
  OAI221_X1 U10932 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .C1(
        n10137), .C2(n10136), .A(n10135), .ZN(n10138) );
  OAI221_X1 U10933 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_126), .C1(
        n10140), .C2(n10139), .A(n10138), .ZN(n10142) );
  AOI21_X1 U10934 ( .B1(keyinput_127), .B2(n10142), .A(keyinput_63), .ZN(
        n10144) );
  INV_X1 U10935 ( .A(keyinput_127), .ZN(n10141) );
  AOI21_X1 U10936 ( .B1(n10142), .B2(n10141), .A(n5868), .ZN(n10143) );
  AOI22_X1 U10937 ( .A1(n5868), .A2(n10144), .B1(keyinput_63), .B2(n10143), 
        .ZN(n10145) );
  AOI21_X1 U10938 ( .B1(n10147), .B2(n10146), .A(n10145), .ZN(n10156) );
  INV_X1 U10939 ( .A(n10148), .ZN(n10154) );
  AOI22_X1 U10940 ( .A1(n10151), .A2(n10449), .B1(n10150), .B2(n10149), .ZN(
        n10152) );
  OAI211_X1 U10941 ( .C1(n10154), .C2(n10620), .A(n10153), .B(n10152), .ZN(
        n10619) );
  AOI22_X1 U10942 ( .A1(n10646), .A2(n10619), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n10645), .ZN(n10155) );
  XNOR2_X1 U10943 ( .A(n10156), .B(n10155), .ZN(P2_U3532) );
  XOR2_X1 U10944 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U10945 ( .A(n10157), .ZN(n10158) );
  NAND2_X1 U10946 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  XNOR2_X1 U10947 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10160), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U10948 ( .A(n10162), .B(n10161), .Z(ADD_1071_U54) );
  XOR2_X1 U10949 ( .A(n10164), .B(n10163), .Z(ADD_1071_U53) );
  XNOR2_X1 U10950 ( .A(n10166), .B(n10165), .ZN(ADD_1071_U52) );
  NOR2_X1 U10951 ( .A1(n10168), .A2(n10167), .ZN(n10170) );
  XNOR2_X1 U10952 ( .A(n10170), .B(n10169), .ZN(ADD_1071_U51) );
  XNOR2_X1 U10953 ( .A(n10172), .B(n10171), .ZN(ADD_1071_U50) );
  XNOR2_X1 U10954 ( .A(n10174), .B(n10173), .ZN(ADD_1071_U49) );
  XNOR2_X1 U10955 ( .A(n10176), .B(n10175), .ZN(ADD_1071_U48) );
  XNOR2_X1 U10956 ( .A(n10178), .B(n10177), .ZN(ADD_1071_U47) );
  XOR2_X1 U10957 ( .A(n10180), .B(n10179), .Z(ADD_1071_U63) );
  XOR2_X1 U10958 ( .A(n10182), .B(n10181), .Z(ADD_1071_U62) );
  XNOR2_X1 U10959 ( .A(n10184), .B(n10183), .ZN(ADD_1071_U61) );
  XNOR2_X1 U10960 ( .A(n10186), .B(n10185), .ZN(ADD_1071_U60) );
  XNOR2_X1 U10961 ( .A(n10188), .B(n10187), .ZN(ADD_1071_U59) );
  XNOR2_X1 U10962 ( .A(n10190), .B(n10189), .ZN(ADD_1071_U58) );
  XNOR2_X1 U10963 ( .A(n10192), .B(n10191), .ZN(ADD_1071_U57) );
  XNOR2_X1 U10964 ( .A(n10194), .B(n10193), .ZN(ADD_1071_U56) );
  NOR2_X1 U10965 ( .A1(n10196), .A2(n10195), .ZN(n10197) );
  XOR2_X1 U10966 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10197), .Z(ADD_1071_U55)
         );
  INV_X1 U10967 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10338) );
  NOR2_X1 U10968 ( .A1(n10198), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10199) );
  OAI21_X1 U10969 ( .B1(n10201), .B2(n10199), .A(n10200), .ZN(n10205) );
  INV_X1 U10970 ( .A(n10221), .ZN(n10203) );
  OAI211_X1 U10971 ( .C1(n10201), .C2(n10200), .A(P1_STATE_REG_SCAN_IN), .B(
        n6694), .ZN(n10202) );
  OAI22_X1 U10972 ( .A1(n10236), .A2(P1_REG1_REG_0__SCAN_IN), .B1(n10203), 
        .B2(n10202), .ZN(n10204) );
  AOI22_X1 U10973 ( .A1(n10205), .A2(n10204), .B1(n10259), .B2(
        P1_ADDR_REG_0__SCAN_IN), .ZN(n10206) );
  OAI21_X1 U10974 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n10338), .A(n10206), .ZN(
        P1_U3241) );
  AOI22_X1 U10975 ( .A1(n10259), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n10207), 
        .B2(n10257), .ZN(n10218) );
  INV_X1 U10976 ( .A(n10208), .ZN(n10217) );
  OAI211_X1 U10977 ( .C1(n10211), .C2(n10210), .A(n10226), .B(n10209), .ZN(
        n10216) );
  OAI211_X1 U10978 ( .C1(n10214), .C2(n10213), .A(n10329), .B(n10212), .ZN(
        n10215) );
  NAND4_X1 U10979 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        P1_U3247) );
  INV_X1 U10980 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10225) );
  NOR4_X1 U10981 ( .A1(n10220), .A2(n10225), .A3(P1_U3084), .A4(n10230), .ZN(
        n10222) );
  AND3_X1 U10982 ( .A1(n10229), .A2(n10222), .A3(n10221), .ZN(n10223) );
  AOI211_X1 U10983 ( .C1(n10259), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10224), 
        .B(n10223), .ZN(n10243) );
  NAND2_X1 U10984 ( .A1(n10230), .A2(n10225), .ZN(n10228) );
  OAI211_X1 U10985 ( .C1(n10229), .C2(n10228), .A(n10227), .B(n10226), .ZN(
        n10242) );
  NAND3_X1 U10986 ( .A1(n10232), .A2(n10231), .A3(n10230), .ZN(n10233) );
  NAND3_X1 U10987 ( .A1(n10234), .A2(n10329), .A3(n10233), .ZN(n10241) );
  INV_X1 U10988 ( .A(n10235), .ZN(n10237) );
  OAI21_X1 U10989 ( .B1(n10237), .B2(n10236), .A(n10318), .ZN(n10239) );
  NAND2_X1 U10990 ( .A1(n10239), .A2(n10238), .ZN(n10240) );
  NAND4_X1 U10991 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        P1_U3252) );
  INV_X1 U10992 ( .A(n10244), .ZN(n10249) );
  AOI211_X1 U10993 ( .C1(n10247), .C2(n10246), .A(n10245), .B(n10321), .ZN(
        n10248) );
  AOI211_X1 U10994 ( .C1(n10250), .C2(n10257), .A(n10249), .B(n10248), .ZN(
        n10256) );
  OAI21_X1 U10995 ( .B1(n10253), .B2(n10252), .A(n10251), .ZN(n10254) );
  AOI22_X1 U10996 ( .A1(n10254), .A2(n10329), .B1(n10259), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U10997 ( .A1(n10256), .A2(n10255), .ZN(P1_U3259) );
  AOI22_X1 U10998 ( .A1(n10259), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n10258), 
        .B2(n10257), .ZN(n10269) );
  AOI21_X1 U10999 ( .B1(n10261), .B2(n10260), .A(n4935), .ZN(n10262) );
  OR2_X1 U11000 ( .A1(n10321), .A2(n10262), .ZN(n10267) );
  OAI211_X1 U11001 ( .C1(n10265), .C2(n10264), .A(n10329), .B(n10263), .ZN(
        n10266) );
  NAND4_X1 U11002 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        P1_U3246) );
  INV_X1 U11003 ( .A(n10270), .ZN(n10273) );
  INV_X1 U11004 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U11005 ( .A1(n10274), .A2(n10273), .B1(n10272), .B2(n10271), .ZN(
        P2_U3437) );
  OAI22_X1 U11006 ( .A1(n10301), .A2(n5621), .B1(n10277), .B2(n10297), .ZN(
        n10276) );
  AOI22_X1 U11007 ( .A1(n10276), .A2(n10275), .B1(P2_ADDR_REG_0__SCAN_IN), 
        .B2(n10296), .ZN(n10282) );
  AOI21_X1 U11008 ( .B1(n10278), .B2(n10277), .A(n10308), .ZN(n10279) );
  OAI21_X1 U11009 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n10301), .A(n10279), .ZN(
        n10280) );
  NAND2_X1 U11010 ( .A1(n10280), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10281) );
  OAI211_X1 U11011 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10283), .A(n10282), .B(
        n10281), .ZN(P2_U3245) );
  AOI22_X1 U11012 ( .A1(n10296), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10294) );
  NAND2_X1 U11013 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10286) );
  AOI211_X1 U11014 ( .C1(n10286), .C2(n10285), .A(n10284), .B(n10297), .ZN(
        n10291) );
  NAND2_X1 U11015 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10289) );
  AOI211_X1 U11016 ( .C1(n10289), .C2(n10288), .A(n10287), .B(n10301), .ZN(
        n10290) );
  AOI211_X1 U11017 ( .C1(n10308), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        n10293) );
  NAND2_X1 U11018 ( .A1(n10294), .A2(n10293), .ZN(P2_U3246) );
  AOI22_X1 U11019 ( .A1(n10296), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10310) );
  AOI211_X1 U11020 ( .C1(n10300), .C2(n10299), .A(n10298), .B(n10297), .ZN(
        n10306) );
  AOI211_X1 U11021 ( .C1(n10304), .C2(n10303), .A(n10302), .B(n10301), .ZN(
        n10305) );
  AOI211_X1 U11022 ( .C1(n10308), .C2(n10307), .A(n10306), .B(n10305), .ZN(
        n10309) );
  NAND2_X1 U11023 ( .A1(n10310), .A2(n10309), .ZN(P2_U3247) );
  XNOR2_X1 U11024 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11025 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10332) );
  INV_X1 U11026 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10311) );
  NOR2_X1 U11027 ( .A1(n10312), .A2(n10311), .ZN(n10323) );
  MUX2_X1 U11028 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6323), .S(n10319), .Z(
        n10315) );
  NAND3_X1 U11029 ( .A1(n10315), .A2(n10314), .A3(n10313), .ZN(n10316) );
  NAND2_X1 U11030 ( .A1(n10317), .A2(n10316), .ZN(n10320) );
  OAI22_X1 U11031 ( .A1(n10321), .A2(n10320), .B1(n10319), .B2(n10318), .ZN(
        n10322) );
  NOR2_X1 U11032 ( .A1(n10323), .A2(n10322), .ZN(n10324) );
  AND2_X1 U11033 ( .A1(n10325), .A2(n10324), .ZN(n10331) );
  XOR2_X1 U11034 ( .A(n10327), .B(n10326), .Z(n10328) );
  NAND2_X1 U11035 ( .A1(n10329), .A2(n10328), .ZN(n10330) );
  OAI211_X1 U11036 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n10332), .A(n10331), .B(
        n10330), .ZN(P1_U3243) );
  AOI21_X1 U11037 ( .B1(n10333), .B2(n10538), .A(n10350), .ZN(n10336) );
  NOR2_X1 U11038 ( .A1(n10334), .A2(n10498), .ZN(n10335) );
  AOI211_X1 U11039 ( .C1(n10498), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10336), .B(
        n10335), .ZN(n10337) );
  OAI21_X1 U11040 ( .B1(n10488), .B2(n10338), .A(n10337), .ZN(P1_U3291) );
  AOI22_X1 U11041 ( .A1(n10341), .A2(n10644), .B1(n10340), .B2(n10339), .ZN(
        n10342) );
  AND2_X1 U11042 ( .A1(n10343), .A2(n10342), .ZN(n10345) );
  AOI22_X1 U11043 ( .A1(n10646), .A2(n10345), .B1(n10277), .B2(n10645), .ZN(
        P2_U3520) );
  INV_X1 U11044 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U11045 ( .A1(n10650), .A2(n10345), .B1(n10344), .B2(n10647), .ZN(
        P2_U3451) );
  OAI21_X1 U11046 ( .B1(n10348), .B2(n10347), .A(n10346), .ZN(n10359) );
  INV_X1 U11047 ( .A(n10359), .ZN(n10369) );
  OAI211_X1 U11048 ( .C1(n10351), .C2(n10350), .A(n10477), .B(n10349), .ZN(
        n10366) );
  OAI21_X1 U11049 ( .B1(n10582), .B2(n10351), .A(n10366), .ZN(n10360) );
  XNOR2_X1 U11050 ( .A(n10353), .B(n10352), .ZN(n10354) );
  NAND2_X1 U11051 ( .A1(n10354), .A2(n10473), .ZN(n10358) );
  AOI22_X1 U11052 ( .A1(n10514), .A2(n10356), .B1(n10516), .B2(n10355), .ZN(
        n10357) );
  OAI211_X1 U11053 ( .C1(n10359), .C2(n10526), .A(n10358), .B(n10357), .ZN(
        n10367) );
  AOI211_X1 U11054 ( .C1(n10585), .C2(n10369), .A(n10360), .B(n10367), .ZN(
        n10363) );
  AOI22_X1 U11055 ( .A1(n10591), .A2(n10363), .B1(n10361), .B2(n10589), .ZN(
        P1_U3524) );
  INV_X1 U11056 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U11057 ( .A1(n10595), .A2(n10363), .B1(n10362), .B2(n10592), .ZN(
        P1_U3457) );
  AOI22_X1 U11058 ( .A1(n10544), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n10364), 
        .B2(n6708), .ZN(n10365) );
  OAI21_X1 U11059 ( .B1(n10493), .B2(n10366), .A(n10365), .ZN(n10368) );
  AOI211_X1 U11060 ( .C1(n10370), .C2(n10369), .A(n10368), .B(n10367), .ZN(
        n10371) );
  AOI22_X1 U11061 ( .A1(n10498), .A2(n6325), .B1(n10371), .B2(n10539), .ZN(
        P1_U3290) );
  NOR2_X1 U11062 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  AOI21_X1 U11063 ( .B1(n10461), .B2(n10375), .A(n10374), .ZN(n10382) );
  OAI21_X1 U11064 ( .B1(n10378), .B2(n10377), .A(n10376), .ZN(n10379) );
  AOI22_X1 U11065 ( .A1(n10457), .A2(n10380), .B1(n4833), .B2(n10379), .ZN(
        n10381) );
  OAI211_X1 U11066 ( .C1(n6360), .C2(n4833), .A(n10382), .B(n10381), .ZN(
        P2_U3295) );
  NAND2_X1 U11067 ( .A1(n10383), .A2(n10477), .ZN(n10384) );
  OAI21_X1 U11068 ( .B1(n10582), .B2(n10385), .A(n10384), .ZN(n10387) );
  AOI211_X1 U11069 ( .C1(n10585), .C2(n10388), .A(n10387), .B(n10386), .ZN(
        n10391) );
  INV_X1 U11070 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U11071 ( .A1(n10591), .A2(n10391), .B1(n10389), .B2(n10589), .ZN(
        P1_U3525) );
  INV_X1 U11072 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U11073 ( .A1(n10595), .A2(n10391), .B1(n10390), .B2(n10592), .ZN(
        P1_U3460) );
  OAI22_X1 U11074 ( .A1(n10440), .A2(n10394), .B1(n10393), .B2(n10392), .ZN(
        n10401) );
  XNOR2_X1 U11075 ( .A(n10396), .B(n10395), .ZN(n10398) );
  OAI22_X1 U11076 ( .A1(n10399), .A2(n10405), .B1(n10398), .B2(n10397), .ZN(
        n10400) );
  NOR2_X1 U11077 ( .A1(n10401), .A2(n10400), .ZN(n10402) );
  OAI21_X1 U11078 ( .B1(n10404), .B2(n10403), .A(n10402), .ZN(P2_U3239) );
  OAI22_X1 U11079 ( .A1(n10406), .A2(n10639), .B1(n10405), .B2(n10638), .ZN(
        n10408) );
  AOI211_X1 U11080 ( .C1(n10609), .C2(n10409), .A(n10408), .B(n10407), .ZN(
        n10411) );
  AOI22_X1 U11081 ( .A1(n10646), .A2(n10411), .B1(n6373), .B2(n10645), .ZN(
        P2_U3522) );
  INV_X1 U11082 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U11083 ( .A1(n10650), .A2(n10411), .B1(n10410), .B2(n10647), .ZN(
        P2_U3457) );
  INV_X1 U11084 ( .A(n10412), .ZN(n10417) );
  OAI22_X1 U11085 ( .A1(n10414), .A2(n10565), .B1(n10413), .B2(n10582), .ZN(
        n10416) );
  AOI211_X1 U11086 ( .C1(n10585), .C2(n10417), .A(n10416), .B(n10415), .ZN(
        n10419) );
  AOI22_X1 U11087 ( .A1(n10591), .A2(n10419), .B1(n6576), .B2(n10589), .ZN(
        P1_U3526) );
  INV_X1 U11088 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U11089 ( .A1(n10595), .A2(n10419), .B1(n10418), .B2(n10592), .ZN(
        P1_U3463) );
  OAI22_X1 U11090 ( .A1(n10421), .A2(n10639), .B1(n10420), .B2(n10638), .ZN(
        n10423) );
  AOI211_X1 U11091 ( .C1(n10609), .C2(n10424), .A(n10423), .B(n10422), .ZN(
        n10426) );
  AOI22_X1 U11092 ( .A1(n10646), .A2(n10426), .B1(n6374), .B2(n10645), .ZN(
        P2_U3523) );
  INV_X1 U11093 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U11094 ( .A1(n10650), .A2(n10426), .B1(n10425), .B2(n10647), .ZN(
        P2_U3460) );
  INV_X1 U11095 ( .A(n10427), .ZN(n10431) );
  OAI22_X1 U11096 ( .A1(n10428), .A2(n10565), .B1(n4835), .B2(n10582), .ZN(
        n10430) );
  AOI211_X1 U11097 ( .C1(n10585), .C2(n10431), .A(n10430), .B(n10429), .ZN(
        n10434) );
  AOI22_X1 U11098 ( .A1(n10591), .A2(n10434), .B1(n10432), .B2(n10589), .ZN(
        P1_U3527) );
  INV_X1 U11099 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U11100 ( .A1(n10595), .A2(n10434), .B1(n10433), .B2(n10592), .ZN(
        P1_U3466) );
  XNOR2_X1 U11101 ( .A(n10435), .B(n10438), .ZN(n10456) );
  AOI21_X1 U11102 ( .B1(n10436), .B2(n10438), .A(n10437), .ZN(n10445) );
  OAI22_X1 U11103 ( .A1(n10442), .A2(n10441), .B1(n10440), .B2(n10439), .ZN(
        n10443) );
  AOI21_X1 U11104 ( .B1(n10445), .B2(n10444), .A(n10443), .ZN(n10468) );
  AND2_X1 U11105 ( .A1(n10446), .A2(n10465), .ZN(n10447) );
  NOR2_X1 U11106 ( .A1(n10448), .A2(n10447), .ZN(n10460) );
  NAND2_X1 U11107 ( .A1(n10460), .A2(n10449), .ZN(n10450) );
  OAI211_X1 U11108 ( .C1(n10451), .C2(n10638), .A(n10468), .B(n10450), .ZN(
        n10452) );
  AOI21_X1 U11109 ( .B1(n10456), .B2(n10644), .A(n10452), .ZN(n10455) );
  INV_X1 U11110 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U11111 ( .A1(n10646), .A2(n10455), .B1(n10453), .B2(n10645), .ZN(
        P2_U3524) );
  INV_X1 U11112 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U11113 ( .A1(n10650), .A2(n10455), .B1(n10454), .B2(n10647), .ZN(
        P2_U3463) );
  NAND2_X1 U11114 ( .A1(n10457), .A2(n10456), .ZN(n10463) );
  AOI22_X1 U11115 ( .A1(n10461), .A2(n10460), .B1(n10459), .B2(n10458), .ZN(
        n10462) );
  OAI211_X1 U11116 ( .C1(n5003), .C2(n4833), .A(n10463), .B(n10462), .ZN(
        n10464) );
  AOI21_X1 U11117 ( .B1(n10466), .B2(n10465), .A(n10464), .ZN(n10467) );
  OAI21_X1 U11118 ( .B1(n10469), .B2(n10468), .A(n10467), .ZN(P2_U3292) );
  XNOR2_X1 U11119 ( .A(n10470), .B(n7248), .ZN(n10495) );
  XNOR2_X1 U11120 ( .A(n9391), .B(n10471), .ZN(n10472) );
  AOI222_X1 U11121 ( .A1(n10475), .A2(n10516), .B1(n10474), .B2(n10514), .C1(
        n10473), .C2(n10472), .ZN(n10491) );
  INV_X1 U11122 ( .A(n10476), .ZN(n10478) );
  OAI211_X1 U11123 ( .C1(n10478), .C2(n10486), .A(n10477), .B(n10510), .ZN(
        n10492) );
  OAI211_X1 U11124 ( .C1(n10486), .C2(n10582), .A(n10491), .B(n10492), .ZN(
        n10479) );
  AOI21_X1 U11125 ( .B1(n10480), .B2(n10495), .A(n10479), .ZN(n10483) );
  INV_X1 U11126 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U11127 ( .A1(n10591), .A2(n10483), .B1(n10481), .B2(n10589), .ZN(
        P1_U3528) );
  INV_X1 U11128 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U11129 ( .A1(n10595), .A2(n10483), .B1(n10482), .B2(n10592), .ZN(
        P1_U3469) );
  INV_X1 U11130 ( .A(n10484), .ZN(n10487) );
  OAI22_X1 U11131 ( .A1(n10488), .A2(n10487), .B1(n10486), .B2(n10485), .ZN(
        n10489) );
  INV_X1 U11132 ( .A(n10489), .ZN(n10490) );
  OAI211_X1 U11133 ( .C1(n10493), .C2(n10492), .A(n10491), .B(n10490), .ZN(
        n10494) );
  AOI21_X1 U11134 ( .B1(n10496), .B2(n10495), .A(n10494), .ZN(n10497) );
  AOI22_X1 U11135 ( .A1(n10498), .A2(n6332), .B1(n10497), .B2(n10539), .ZN(
        P1_U3286) );
  INV_X1 U11136 ( .A(n10499), .ZN(n10500) );
  OAI21_X1 U11137 ( .B1(n10501), .B2(n10638), .A(n10500), .ZN(n10504) );
  INV_X1 U11138 ( .A(n10502), .ZN(n10503) );
  AOI211_X1 U11139 ( .C1(n10644), .C2(n10505), .A(n10504), .B(n10503), .ZN(
        n10507) );
  AOI22_X1 U11140 ( .A1(n10646), .A2(n10507), .B1(n6375), .B2(n10645), .ZN(
        P2_U3525) );
  INV_X1 U11141 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U11142 ( .A1(n10650), .A2(n10507), .B1(n10506), .B2(n10647), .ZN(
        P2_U3466) );
  OAI21_X1 U11143 ( .B1(n10509), .B2(n10519), .A(n10508), .ZN(n10536) );
  INV_X1 U11144 ( .A(n10510), .ZN(n10512) );
  OAI21_X1 U11145 ( .B1(n10537), .B2(n10512), .A(n10511), .ZN(n10532) );
  OAI22_X1 U11146 ( .A1(n10532), .A2(n10565), .B1(n10537), .B2(n10582), .ZN(
        n10528) );
  INV_X1 U11147 ( .A(n10536), .ZN(n10527) );
  AOI22_X1 U11148 ( .A1(n10516), .A2(n10515), .B1(n10514), .B2(n10513), .ZN(
        n10525) );
  INV_X1 U11149 ( .A(n10517), .ZN(n10522) );
  AOI21_X1 U11150 ( .B1(n10520), .B2(n10519), .A(n10518), .ZN(n10521) );
  OAI21_X1 U11151 ( .B1(n10523), .B2(n10522), .A(n10521), .ZN(n10524) );
  OAI211_X1 U11152 ( .C1(n10527), .C2(n10526), .A(n10525), .B(n10524), .ZN(
        n10540) );
  AOI211_X1 U11153 ( .C1(n10585), .C2(n10536), .A(n10528), .B(n10540), .ZN(
        n10531) );
  AOI22_X1 U11154 ( .A1(n10591), .A2(n10531), .B1(n10529), .B2(n10589), .ZN(
        P1_U3529) );
  INV_X1 U11155 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U11156 ( .A1(n10595), .A2(n10531), .B1(n10530), .B2(n10592), .ZN(
        P1_U3472) );
  INV_X1 U11157 ( .A(n10532), .ZN(n10533) );
  AOI22_X1 U11158 ( .A1(n10536), .A2(n10535), .B1(n10534), .B2(n10533), .ZN(
        n10546) );
  NOR2_X1 U11159 ( .A1(n10538), .A2(n10537), .ZN(n10542) );
  MUX2_X1 U11160 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10540), .S(n10539), .Z(
        n10541) );
  AOI211_X1 U11161 ( .C1(n10544), .C2(n10543), .A(n10542), .B(n10541), .ZN(
        n10545) );
  NAND2_X1 U11162 ( .A1(n10546), .A2(n10545), .ZN(P1_U3285) );
  AOI21_X1 U11163 ( .B1(n10549), .B2(n10548), .A(n10547), .ZN(n10550) );
  OAI211_X1 U11164 ( .C1(n10553), .C2(n10552), .A(n10551), .B(n10550), .ZN(
        n10554) );
  INV_X1 U11165 ( .A(n10554), .ZN(n10557) );
  AOI22_X1 U11166 ( .A1(n10591), .A2(n10557), .B1(n10555), .B2(n10589), .ZN(
        P1_U3530) );
  INV_X1 U11167 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U11168 ( .A1(n10595), .A2(n10557), .B1(n10556), .B2(n10592), .ZN(
        P1_U3475) );
  OAI22_X1 U11169 ( .A1(n10559), .A2(n10639), .B1(n10558), .B2(n10638), .ZN(
        n10561) );
  AOI211_X1 U11170 ( .C1(n10644), .C2(n10562), .A(n10561), .B(n10560), .ZN(
        n10563) );
  AOI22_X1 U11171 ( .A1(n10646), .A2(n10563), .B1(n6419), .B2(n10645), .ZN(
        P2_U3527) );
  AOI22_X1 U11172 ( .A1(n10650), .A2(n10563), .B1(n5725), .B2(n10647), .ZN(
        P2_U3472) );
  OAI22_X1 U11173 ( .A1(n10566), .A2(n10565), .B1(n10564), .B2(n10582), .ZN(
        n10568) );
  AOI211_X1 U11174 ( .C1(n10585), .C2(n10569), .A(n10568), .B(n10567), .ZN(
        n10572) );
  AOI22_X1 U11175 ( .A1(n10591), .A2(n10572), .B1(n10570), .B2(n10589), .ZN(
        P1_U3531) );
  INV_X1 U11176 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U11177 ( .A1(n10595), .A2(n10572), .B1(n10571), .B2(n10592), .ZN(
        P1_U3478) );
  NAND3_X1 U11178 ( .A1(n10574), .A2(n10573), .A3(n10644), .ZN(n10576) );
  OAI211_X1 U11179 ( .C1(n5131), .C2(n10638), .A(n10576), .B(n10575), .ZN(
        n10577) );
  NOR2_X1 U11180 ( .A1(n10578), .A2(n10577), .ZN(n10580) );
  AOI22_X1 U11181 ( .A1(n10646), .A2(n10580), .B1(n6445), .B2(n10645), .ZN(
        P2_U3528) );
  INV_X1 U11182 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U11183 ( .A1(n10650), .A2(n10580), .B1(n10579), .B2(n10647), .ZN(
        P2_U3475) );
  OAI21_X1 U11184 ( .B1(n10583), .B2(n10582), .A(n10581), .ZN(n10584) );
  AOI21_X1 U11185 ( .B1(n10586), .B2(n10585), .A(n10584), .ZN(n10587) );
  AND2_X1 U11186 ( .A1(n10588), .A2(n10587), .ZN(n10594) );
  AOI22_X1 U11187 ( .A1(n10591), .A2(n10594), .B1(n10590), .B2(n10589), .ZN(
        P1_U3532) );
  INV_X1 U11188 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U11189 ( .A1(n10595), .A2(n10594), .B1(n10593), .B2(n10592), .ZN(
        P1_U3481) );
  INV_X1 U11190 ( .A(n10596), .ZN(n10597) );
  OAI22_X1 U11191 ( .A1(n10598), .A2(n10639), .B1(n10597), .B2(n10638), .ZN(
        n10600) );
  AOI211_X1 U11192 ( .C1(n10609), .C2(n10601), .A(n10600), .B(n10599), .ZN(
        n10602) );
  AOI22_X1 U11193 ( .A1(n10646), .A2(n10602), .B1(n6460), .B2(n10645), .ZN(
        P2_U3529) );
  AOI22_X1 U11194 ( .A1(n10650), .A2(n10602), .B1(n5755), .B2(n10647), .ZN(
        P2_U3478) );
  INV_X1 U11195 ( .A(n10603), .ZN(n10608) );
  OAI22_X1 U11196 ( .A1(n10605), .A2(n10639), .B1(n10604), .B2(n10638), .ZN(
        n10607) );
  AOI211_X1 U11197 ( .C1(n10609), .C2(n10608), .A(n10607), .B(n10606), .ZN(
        n10611) );
  AOI22_X1 U11198 ( .A1(n10646), .A2(n10611), .B1(n6473), .B2(n10645), .ZN(
        P2_U3530) );
  INV_X1 U11199 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U11200 ( .A1(n10650), .A2(n10611), .B1(n10610), .B2(n10647), .ZN(
        P2_U3481) );
  INV_X1 U11201 ( .A(n10612), .ZN(n10615) );
  OAI211_X1 U11202 ( .C1(n10615), .C2(n10638), .A(n10614), .B(n10613), .ZN(
        n10616) );
  AOI21_X1 U11203 ( .B1(n10617), .B2(n10644), .A(n10616), .ZN(n10618) );
  AOI22_X1 U11204 ( .A1(n10646), .A2(n10618), .B1(n7196), .B2(n10645), .ZN(
        P2_U3531) );
  AOI22_X1 U11205 ( .A1(n10650), .A2(n10618), .B1(n5788), .B2(n10647), .ZN(
        P2_U3484) );
  MUX2_X1 U11206 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n10619), .S(n10650), .Z(
        P2_U3487) );
  NOR2_X1 U11207 ( .A1(n10621), .A2(n10620), .ZN(n10626) );
  OAI22_X1 U11208 ( .A1(n10623), .A2(n10639), .B1(n10622), .B2(n10638), .ZN(
        n10625) );
  AOI211_X1 U11209 ( .C1(n10626), .C2(n7877), .A(n10625), .B(n10624), .ZN(
        n10628) );
  AOI22_X1 U11210 ( .A1(n10646), .A2(n10628), .B1(n7544), .B2(n10645), .ZN(
        P2_U3533) );
  INV_X1 U11211 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U11212 ( .A1(n10650), .A2(n10628), .B1(n10627), .B2(n10647), .ZN(
        P2_U3490) );
  INV_X1 U11213 ( .A(n10629), .ZN(n10634) );
  OAI22_X1 U11214 ( .A1(n10631), .A2(n10639), .B1(n10630), .B2(n10638), .ZN(
        n10633) );
  AOI211_X1 U11215 ( .C1(n10644), .C2(n10634), .A(n10633), .B(n10632), .ZN(
        n10636) );
  AOI22_X1 U11216 ( .A1(n10646), .A2(n10636), .B1(n7651), .B2(n10645), .ZN(
        P2_U3534) );
  INV_X1 U11217 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U11218 ( .A1(n10650), .A2(n10636), .B1(n10635), .B2(n10647), .ZN(
        P2_U3493) );
  OAI22_X1 U11219 ( .A1(n10640), .A2(n10639), .B1(n5135), .B2(n10638), .ZN(
        n10642) );
  AOI211_X1 U11220 ( .C1(n10644), .C2(n10643), .A(n10642), .B(n10641), .ZN(
        n10649) );
  AOI22_X1 U11221 ( .A1(n10646), .A2(n10649), .B1(n5871), .B2(n10645), .ZN(
        P2_U3535) );
  INV_X1 U11222 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U11223 ( .A1(n10650), .A2(n10649), .B1(n10648), .B2(n10647), .ZN(
        P2_U3496) );
  XNOR2_X1 U11224 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X4 U6505 ( .A(n5648), .ZN(n5657) );
  CLKBUF_X1 U4895 ( .A(n5620), .Z(n6089) );
  CLKBUF_X1 U4909 ( .A(n6584), .Z(n4831) );
  CLKBUF_X1 U4940 ( .A(n6950), .Z(n8744) );
endmodule

