

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721;

  NAND2_X1 U3402 ( .A1(n3329), .A2(n3328), .ZN(n4977) );
  CLKBUF_X2 U3403 ( .A(n3131), .Z(n4046) );
  CLKBUF_X2 U3404 ( .A(n3239), .Z(n4054) );
  AND2_X1 U3405 ( .A1(n3823), .A2(n4491), .ZN(n3246) );
  CLKBUF_X1 U3406 ( .A(n3180), .Z(n4491) );
  AND4_X1 U3407 ( .A1(n3159), .A2(n3158), .A3(n3157), .A4(n3156), .ZN(n3175)
         );
  INV_X1 U3408 ( .A(n4497), .ZN(n3183) );
  AND4_X1 U3409 ( .A1(n3082), .A2(n3081), .A3(n3080), .A4(n3079), .ZN(n3093)
         );
  AND2_X2 U3410 ( .A1(n5107), .A2(n3053), .ZN(n3140) );
  AND2_X2 U3411 ( .A1(n5107), .A2(n4434), .ZN(n3251) );
  AND2_X1 U3412 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4434) );
  OR2_X1 U3413 ( .A1(n3187), .A2(n6423), .ZN(n3357) );
  AND2_X1 U3414 ( .A1(n3187), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3823) );
  INV_X1 U3415 ( .A(n3180), .ZN(n4372) );
  OR2_X1 U3416 ( .A1(n3544), .A2(n3543), .ZN(n3557) );
  INV_X1 U3417 ( .A(n3188), .ZN(n3826) );
  INV_X2 U3418 ( .A(n4348), .ZN(n4134) );
  AND2_X2 U3419 ( .A1(n3826), .A2(n3187), .ZN(n4283) );
  BUF_X1 U3420 ( .A(n6221), .Z(n2956) );
  INV_X1 U3421 ( .A(n4892), .ZN(n5870) );
  OAI21_X2 U3422 ( .B1(n4518), .B2(n4158), .A(n4170), .ZN(n6007) );
  NAND2_X1 U3424 ( .A1(n3397), .A2(n3375), .ZN(n4517) );
  XNOR2_X1 U3425 ( .A(n3249), .B(n3248), .ZN(n3294) );
  NOR2_X1 U3426 ( .A1(n3210), .A2(n4497), .ZN(n3211) );
  NAND4_X1 U3429 ( .A1(n3154), .A2(n3153), .A3(n3152), .A4(n3151), .ZN(n3188)
         );
  NAND2_X1 U3430 ( .A1(n2963), .A2(n3128), .ZN(n4469) );
  AND4_X1 U3431 ( .A1(n3062), .A2(n3061), .A3(n3060), .A4(n3059), .ZN(n3063)
         );
  AND4_X1 U3432 ( .A1(n3070), .A2(n3069), .A3(n3068), .A4(n3067), .ZN(n3106)
         );
  BUF_X2 U3433 ( .A(n3251), .Z(n4045) );
  BUF_X2 U3434 ( .A(n3307), .Z(n4052) );
  CLKBUF_X2 U3435 ( .A(n3155), .Z(n4033) );
  CLKBUF_X2 U3436 ( .A(n3271), .Z(n4053) );
  AND2_X4 U3437 ( .A1(n4437), .A2(n3052), .ZN(n3310) );
  CLKBUF_X2 U3438 ( .A(n3275), .Z(n4055) );
  AND2_X2 U3439 ( .A1(n3041), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3047)
         );
  INV_X2 U3440 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3039) );
  AND2_X1 U3441 ( .A1(n4026), .A2(n3819), .ZN(n5353) );
  NOR2_X1 U3442 ( .A1(n4251), .A2(n4248), .ZN(n5345) );
  XNOR2_X1 U3443 ( .A(n4078), .B(n4077), .ZN(n4149) );
  NAND2_X1 U3444 ( .A1(n5361), .A2(n4247), .ZN(n4251) );
  NAND2_X1 U34450 ( .A1(n4246), .A2(n4245), .ZN(n5361) );
  INV_X1 U34460 ( .A(n4229), .ZN(n3001) );
  AOI21_X1 U34470 ( .B1(n2999), .B2(n2997), .A(n2971), .ZN(n2996) );
  INV_X1 U34480 ( .A(n2999), .ZN(n2998) );
  OAI21_X1 U3449 ( .B1(n2995), .B2(n4233), .A(n4232), .ZN(n3003) );
  AND2_X1 U3450 ( .A1(n4557), .A2(n4561), .ZN(n4558) );
  NAND2_X1 U34510 ( .A1(n4192), .A2(n4191), .ZN(n4194) );
  AOI21_X1 U34520 ( .B1(n4179), .B2(n3583), .A(n3409), .ZN(n4565) );
  AND2_X1 U34530 ( .A1(n3398), .A2(n3426), .ZN(n4179) );
  CLKBUF_X1 U3454 ( .A(n4457), .Z(n6112) );
  NAND2_X1 U34550 ( .A1(n3294), .A2(n3295), .ZN(n3374) );
  NAND2_X1 U34560 ( .A1(n3372), .A2(n3371), .ZN(n4458) );
  XNOR2_X1 U3457 ( .A(n3350), .B(n6326), .ZN(n4418) );
  OR2_X1 U3458 ( .A1(n6221), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3329) );
  OR2_X2 U34590 ( .A1(n3233), .A2(n3232), .ZN(n3350) );
  NAND2_X2 U34600 ( .A1(n5878), .A2(n3894), .ZN(n5300) );
  AND2_X2 U34610 ( .A1(n5992), .A2(n4144), .ZN(n6006) );
  AOI21_X1 U34620 ( .B1(n3228), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3231), .ZN(n3232) );
  CLKBUF_X1 U34630 ( .A(n3227), .Z(n3228) );
  NAND2_X1 U34640 ( .A1(n3207), .A2(n3206), .ZN(n3291) );
  OAI21_X1 U34650 ( .B1(n3205), .B2(n3185), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3190) );
  CLKBUF_X1 U3466 ( .A(n4080), .Z(n4296) );
  AND4_X1 U3467 ( .A1(n3204), .A2(n3887), .A3(n3203), .A4(n3202), .ZN(n3207)
         );
  AND2_X2 U34680 ( .A1(n3212), .A2(n3211), .ZN(n4133) );
  NAND2_X1 U34690 ( .A1(n4134), .A2(n5128), .ZN(n5272) );
  AND2_X1 U34700 ( .A1(n3182), .A2(n3181), .ZN(n3878) );
  AOI22_X1 U34710 ( .A1(n3246), .A2(n4337), .B1(n3284), .B2(n4487), .ZN(n3189)
         );
  INV_X1 U34720 ( .A(n3357), .ZN(n3284) );
  OR2_X1 U34730 ( .A1(n4141), .A2(n3905), .ZN(n4381) );
  CLKBUF_X1 U34740 ( .A(n3200), .Z(n3891) );
  NAND2_X2 U3475 ( .A1(n3106), .A2(n3107), .ZN(n3214) );
  AND4_X1 U3476 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n3154)
         );
  AND4_X1 U3477 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n3152)
         );
  NAND4_X1 U3478 ( .A1(n3066), .A2(n3065), .A3(n3064), .A4(n3063), .ZN(n3180)
         );
  NAND2_X1 U3479 ( .A1(n2962), .A2(n3104), .ZN(n4497) );
  AND4_X1 U3480 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3174)
         );
  AND4_X1 U3481 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n3104)
         );
  AND4_X1 U3482 ( .A1(n3171), .A2(n3170), .A3(n3169), .A4(n3168), .ZN(n3172)
         );
  AND4_X1 U3483 ( .A1(n3167), .A2(n3166), .A3(n3165), .A4(n3164), .ZN(n3173)
         );
  AND4_X1 U3484 ( .A1(n3045), .A2(n3044), .A3(n3043), .A4(n3042), .ZN(n3066)
         );
  AND4_X1 U3485 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n3153)
         );
  AND4_X1 U3486 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .ZN(n3151)
         );
  AND4_X1 U3487 ( .A1(n3127), .A2(n3126), .A3(n3125), .A4(n3124), .ZN(n3128)
         );
  AND4_X1 U3488 ( .A1(n3057), .A2(n3056), .A3(n3055), .A4(n3054), .ZN(n3064)
         );
  AND4_X1 U3489 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(n3116)
         );
  AND4_X1 U3490 ( .A1(n3078), .A2(n3077), .A3(n3076), .A4(n3075), .ZN(n3094)
         );
  AND4_X1 U3491 ( .A1(n3051), .A2(n3050), .A3(n3049), .A4(n3048), .ZN(n3065)
         );
  INV_X2 U3492 ( .A(n6547), .ZN(n6497) );
  AND2_X2 U3493 ( .A1(n3052), .A2(n3047), .ZN(n3307) );
  AND2_X2 U3494 ( .A1(n3047), .A2(n4434), .ZN(n3155) );
  BUF_X2 U3495 ( .A(n3146), .Z(n4047) );
  AND2_X2 U3496 ( .A1(n4437), .A2(n4434), .ZN(n3146) );
  AND2_X2 U3497 ( .A1(n3039), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5107)
         );
  INV_X2 U3498 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U3499 ( .A1(n3095), .A2(n3214), .ZN(n2954) );
  NAND2_X1 U3500 ( .A1(n3095), .A2(n3214), .ZN(n3176) );
  AOI21_X1 U3501 ( .B1(n3209), .B2(n3213), .A(n4152), .ZN(n3184) );
  NAND2_X1 U3503 ( .A1(n4770), .A2(n4195), .ZN(n4903) );
  NAND2_X1 U3505 ( .A1(n4510), .A2(n4178), .ZN(n6000) );
  XNOR2_X1 U3506 ( .A(n3300), .B(n3299), .ZN(n4150) );
  NAND2_X1 U3508 ( .A1(n3195), .A2(n3194), .ZN(n3289) );
  AND2_X1 U3509 ( .A1(n3052), .A2(n4295), .ZN(n2955) );
  AND2_X1 U3510 ( .A1(n3107), .A2(n3106), .ZN(n3119) );
  OAI21_X1 U3511 ( .B1(n3291), .B2(n3289), .A(n3290), .ZN(n6221) );
  NOR2_X2 U3512 ( .A1(n5261), .A2(n3023), .ZN(n5187) );
  NAND2_X2 U3513 ( .A1(n5209), .A2(n5400), .ZN(n5261) );
  NAND2_X1 U3514 ( .A1(n3373), .A2(n2960), .ZN(n3426) );
  NAND2_X1 U3515 ( .A1(n4372), .A2(n4479), .ZN(n4141) );
  NAND2_X1 U3516 ( .A1(n4418), .A2(n6423), .ZN(n3372) );
  OAI21_X1 U3517 ( .B1(n4517), .B2(n3572), .A(n3383), .ZN(n3384) );
  NOR2_X2 U3519 ( .A1(n5235), .A2(n5288), .ZN(n5221) );
  NOR2_X2 U3520 ( .A1(n5222), .A2(n3027), .ZN(n5209) );
  NAND2_X2 U3522 ( .A1(n3817), .A2(n3033), .ZN(n5141) );
  NOR2_X4 U3523 ( .A1(n5175), .A2(n5176), .ZN(n3817) );
  XNOR2_X2 U3524 ( .A(n5141), .B(n4258), .ZN(n5118) );
  INV_X1 U3525 ( .A(n3246), .ZN(n3452) );
  NAND2_X1 U3526 ( .A1(n2954), .A2(n3177), .ZN(n3208) );
  NAND2_X1 U3527 ( .A1(n6380), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4069) );
  NOR2_X1 U3528 ( .A1(n3894), .A2(n6414), .ZN(n3337) );
  INV_X1 U3529 ( .A(n2961), .ZN(n2997) );
  OR2_X1 U3530 ( .A1(n4364), .A2(n4135), .ZN(n5936) );
  AND2_X1 U3531 ( .A1(n3034), .A2(n5142), .ZN(n3033) );
  NAND2_X1 U3532 ( .A1(n6415), .A2(n6420), .ZN(n4364) );
  NAND2_X1 U3533 ( .A1(n3130), .A2(n3129), .ZN(n3019) );
  AND2_X1 U3534 ( .A1(n3201), .A2(n3894), .ZN(n3129) );
  INV_X1 U3535 ( .A(n3396), .ZN(n3006) );
  NOR2_X1 U3536 ( .A1(n3017), .A2(n3016), .ZN(n3015) );
  AND2_X1 U3537 ( .A1(n2953), .A2(n4243), .ZN(n3016) );
  INV_X1 U3538 ( .A(n4242), .ZN(n3017) );
  NAND2_X1 U3539 ( .A1(n2975), .A2(EBX_REG_1__SCAN_IN), .ZN(n2980) );
  OR2_X1 U3540 ( .A1(n3281), .A2(n3280), .ZN(n4220) );
  OR2_X1 U3541 ( .A1(n3245), .A2(n3244), .ZN(n3247) );
  NAND2_X1 U3542 ( .A1(n3183), .A2(n4469), .ZN(n4152) );
  OR2_X1 U3543 ( .A1(n4491), .A2(n6423), .ZN(n3356) );
  NOR2_X1 U3544 ( .A1(n5153), .A2(n3818), .ZN(n3034) );
  OR2_X1 U3545 ( .A1(n5279), .A2(n5269), .ZN(n3029) );
  AND2_X1 U3546 ( .A1(n2972), .A2(n5034), .ZN(n3030) );
  NOR2_X1 U3547 ( .A1(n4777), .A2(n4780), .ZN(n4778) );
  NAND2_X1 U3548 ( .A1(n5571), .A2(n2989), .ZN(n2994) );
  NOR2_X1 U3549 ( .A1(n2990), .A2(n5201), .ZN(n2989) );
  INV_X1 U3550 ( .A(n2991), .ZN(n2990) );
  INV_X1 U3551 ( .A(n5081), .ZN(n2986) );
  AND2_X1 U3552 ( .A1(n5040), .A2(n2988), .ZN(n2987) );
  INV_X1 U3553 ( .A(n5069), .ZN(n2988) );
  INV_X1 U3554 ( .A(n4233), .ZN(n3005) );
  INV_X1 U3555 ( .A(n4563), .ZN(n2982) );
  NAND2_X1 U3556 ( .A1(n2975), .A2(n4348), .ZN(n3972) );
  NAND2_X1 U3557 ( .A1(n4134), .A2(n5274), .ZN(n3979) );
  INV_X1 U3558 ( .A(n3247), .ZN(n4172) );
  NOR2_X1 U3559 ( .A1(n4469), .A2(n4497), .ZN(n3895) );
  AND2_X1 U3560 ( .A1(n4479), .A2(n4487), .ZN(n4207) );
  AND2_X1 U3562 ( .A1(n5785), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4953) );
  OR2_X1 U3563 ( .A1(n3796), .A2(n3795), .ZN(n5176) );
  INV_X1 U3564 ( .A(n4015), .ZN(n4076) );
  AND2_X1 U3565 ( .A1(n6414), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4075) );
  INV_X1 U3566 ( .A(n4258), .ZN(n3032) );
  AOI21_X1 U3567 ( .B1(n4072), .B2(n5145), .A(n4044), .ZN(n5142) );
  NAND2_X1 U3568 ( .A1(n4020), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4071)
         );
  OR2_X1 U3569 ( .A1(n3026), .A2(n2973), .ZN(n3023) );
  INV_X1 U3570 ( .A(n5198), .ZN(n3026) );
  INV_X1 U3571 ( .A(n5261), .ZN(n3025) );
  NOR2_X1 U3572 ( .A1(n3471), .A2(n3454), .ZN(n3476) );
  NOR2_X1 U3573 ( .A1(n4450), .A2(n4565), .ZN(n4557) );
  INV_X1 U3574 ( .A(n3905), .ZN(n5128) );
  NAND2_X1 U3575 ( .A1(n4226), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4248) );
  INV_X1 U3576 ( .A(n5363), .ZN(n4245) );
  NAND2_X1 U3577 ( .A1(n5571), .A2(n2991), .ZN(n5257) );
  NAND2_X1 U3578 ( .A1(n5449), .A2(n3009), .ZN(n3008) );
  NAND2_X1 U3579 ( .A1(n3037), .A2(n4237), .ZN(n3009) );
  NAND2_X1 U3580 ( .A1(n5291), .A2(n5290), .ZN(n5293) );
  NAND2_X1 U3581 ( .A1(n5055), .A2(n3004), .ZN(n2995) );
  NAND2_X1 U3582 ( .A1(n3001), .A2(n2961), .ZN(n3000) );
  NAND2_X1 U3583 ( .A1(n5819), .A2(n3932), .ZN(n5820) );
  NAND2_X1 U3584 ( .A1(n4366), .A2(n4365), .ZN(n4385) );
  AND2_X1 U3585 ( .A1(n6520), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3898) );
  OR2_X1 U3586 ( .A1(n3866), .A2(n3865), .ZN(n3868) );
  NAND2_X1 U3587 ( .A1(n3246), .A2(n4207), .ZN(n3874) );
  AND2_X1 U3588 ( .A1(n3861), .A2(n3860), .ZN(n4084) );
  OR3_X1 U3589 ( .A1(n3866), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6398), 
        .ZN(n3861) );
  NAND2_X1 U3590 ( .A1(n4281), .A2(n4262), .ZN(n6536) );
  AND2_X1 U3591 ( .A1(n5120), .A2(n5119), .ZN(n5886) );
  AND2_X1 U3592 ( .A1(n5120), .A2(n4343), .ZN(n5322) );
  NAND2_X1 U3593 ( .A1(n5178), .A2(n3818), .ZN(n3819) );
  NAND2_X1 U3594 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6415), .ZN(n6514) );
  OR2_X1 U3595 ( .A1(n3419), .A2(n3418), .ZN(n4198) );
  OR2_X1 U3596 ( .A1(n3438), .A2(n3437), .ZN(n4209) );
  OR2_X1 U3597 ( .A1(n3395), .A2(n3394), .ZN(n4197) );
  NAND2_X1 U3598 ( .A1(n3186), .A2(n4469), .ZN(n3201) );
  AND2_X2 U3599 ( .A1(n3046), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3058)
         );
  AND2_X1 U3600 ( .A1(n4133), .A2(n3187), .ZN(n4079) );
  AND2_X1 U3601 ( .A1(n3542), .A2(n3541), .ZN(n3543) );
  OAI21_X1 U3602 ( .B1(n3452), .B2(n3451), .A(n3450), .ZN(n3453) );
  NOR2_X1 U3603 ( .A1(n3377), .A2(n3376), .ZN(n3401) );
  NAND2_X1 U3604 ( .A1(n3014), .A2(n2974), .ZN(n4246) );
  NAND2_X1 U3605 ( .A1(n5371), .A2(n3015), .ZN(n3014) );
  NOR2_X1 U3606 ( .A1(n3975), .A2(n2992), .ZN(n2991) );
  INV_X1 U3607 ( .A(n5570), .ZN(n2992) );
  NOR2_X1 U3608 ( .A1(n4238), .A2(n3013), .ZN(n3010) );
  INV_X1 U3609 ( .A(n4228), .ZN(n3004) );
  INV_X1 U3610 ( .A(n4566), .ZN(n2984) );
  NAND2_X1 U3611 ( .A1(n2979), .A2(n2968), .ZN(n3904) );
  AND3_X1 U3612 ( .A1(n3972), .A2(n3901), .A3(n2980), .ZN(n2979) );
  NAND2_X1 U3613 ( .A1(n5128), .A2(n2978), .ZN(n2977) );
  OR2_X1 U3614 ( .A1(n3891), .A2(n3591), .ZN(n4126) );
  INV_X1 U3615 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6387) );
  OAI21_X1 U3616 ( .B1(n6542), .B2(n4444), .A(n6514), .ZN(n4467) );
  NAND2_X1 U3617 ( .A1(n3357), .A2(n3356), .ZN(n3843) );
  CLKBUF_X1 U3618 ( .A(n4079), .Z(n4266) );
  OR4_X1 U3619 ( .A1(n6473), .A2(n6471), .A3(n4113), .A4(n5039), .ZN(n5763) );
  NAND2_X1 U3620 ( .A1(n5191), .A2(n3991), .ZN(n5156) );
  AND2_X1 U3621 ( .A1(n3909), .A2(n3908), .ZN(n4415) );
  CLKBUF_X1 U3622 ( .A(n3306), .Z(n4332) );
  OR2_X1 U3623 ( .A1(n4071), .A2(n5146), .ZN(n4090) );
  AND2_X1 U3624 ( .A1(n4019), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4020)
         );
  OR2_X1 U3625 ( .A1(n4025), .A2(n4024), .ZN(n5153) );
  INV_X1 U3626 ( .A(n3817), .ZN(n5178) );
  NAND2_X1 U3627 ( .A1(n3792), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4018)
         );
  AND2_X1 U3628 ( .A1(n5368), .A2(n4072), .ZN(n3770) );
  NOR2_X1 U3629 ( .A1(n3748), .A2(n5643), .ZN(n3749) );
  INV_X1 U3630 ( .A(n5254), .ZN(n3024) );
  INV_X1 U3631 ( .A(n3703), .ZN(n3704) );
  AND2_X1 U3632 ( .A1(n3688), .A2(n3687), .ZN(n5400) );
  NAND2_X1 U3633 ( .A1(n3028), .A2(n5210), .ZN(n3027) );
  INV_X1 U3634 ( .A(n3029), .ZN(n3028) );
  NAND2_X1 U3635 ( .A1(n3655), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3703)
         );
  NOR2_X1 U3636 ( .A1(n3619), .A2(n5435), .ZN(n3620) );
  AND2_X1 U3637 ( .A1(n3620), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3654)
         );
  CLKBUF_X1 U3638 ( .A(n5222), .Z(n5223) );
  NAND2_X1 U3639 ( .A1(n3574), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3590)
         );
  NOR2_X1 U3640 ( .A1(n5237), .A2(n3022), .ZN(n3021) );
  INV_X1 U3641 ( .A(n5079), .ZN(n3022) );
  AND2_X1 U3642 ( .A1(n3539), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3540)
         );
  NAND2_X1 U3643 ( .A1(n3540), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3573)
         );
  OAI211_X1 U3644 ( .C1(n3572), .C2(n3538), .A(n3537), .B(n3536), .ZN(n5034)
         );
  OR2_X1 U3645 ( .A1(n3493), .A2(n5828), .ZN(n3494) );
  NOR2_X1 U3646 ( .A1(n6660), .A2(n3494), .ZN(n3535) );
  NAND2_X1 U3647 ( .A1(n3476), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3493)
         );
  NAND2_X1 U3648 ( .A1(n4917), .A2(n4215), .ZN(n4962) );
  AND4_X1 U3649 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n4780)
         );
  CLKBUF_X1 U3650 ( .A(n4778), .Z(n4779) );
  AND2_X1 U3651 ( .A1(n3441), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3442)
         );
  NAND2_X1 U3652 ( .A1(n3442), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3471)
         );
  CLKBUF_X1 U3653 ( .A(n4558), .Z(n4559) );
  AND2_X1 U3654 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3401), .ZN(n3441)
         );
  INV_X1 U3655 ( .A(n3382), .ZN(n3383) );
  NAND2_X1 U3656 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3377) );
  AOI21_X1 U3657 ( .B1(n4457), .B2(n3583), .A(n4075), .ZN(n4412) );
  NAND2_X1 U3658 ( .A1(n3304), .A2(n3303), .ZN(n4345) );
  NAND2_X1 U3659 ( .A1(n3976), .A2(n5274), .ZN(n4104) );
  OR2_X1 U3660 ( .A1(n5156), .A2(n5155), .ZN(n5158) );
  NOR2_X1 U3661 ( .A1(n5158), .A2(n4102), .ZN(n5126) );
  NOR2_X1 U3662 ( .A1(n2994), .A2(n2993), .ZN(n5191) );
  INV_X1 U3663 ( .A(n5189), .ZN(n2993) );
  AND2_X1 U3664 ( .A1(n5213), .A2(n3964), .ZN(n5571) );
  NAND2_X1 U3665 ( .A1(n5571), .A2(n5570), .ZN(n5573) );
  NOR2_X1 U3666 ( .A1(n5281), .A2(n5276), .ZN(n5213) );
  OR2_X1 U3668 ( .A1(n5293), .A2(n5226), .ZN(n5281) );
  AOI21_X1 U3669 ( .B1(n4236), .B2(n3012), .A(n3011), .ZN(n5421) );
  AND2_X1 U3670 ( .A1(n5802), .A2(n2976), .ZN(n5291) );
  INV_X1 U3671 ( .A(n5241), .ZN(n2985) );
  NAND2_X1 U3672 ( .A1(n5802), .A2(n2970), .ZN(n5242) );
  NAND2_X1 U3673 ( .A1(n5802), .A2(n5040), .ZN(n5070) );
  NAND2_X1 U3674 ( .A1(n5802), .A2(n2987), .ZN(n5082) );
  NOR2_X1 U3675 ( .A1(n3003), .A2(n5086), .ZN(n2999) );
  AND3_X1 U3676 ( .A1(n3934), .A2(n3972), .A3(n3933), .ZN(n4930) );
  OR2_X1 U3677 ( .A1(n5820), .A2(n4930), .ZN(n5800) );
  AND2_X1 U3678 ( .A1(n3931), .A2(n3930), .ZN(n5817) );
  AND2_X1 U3679 ( .A1(n4764), .A2(n4693), .ZN(n5819) );
  AND2_X1 U3680 ( .A1(n3920), .A2(n3919), .ZN(n4762) );
  AND2_X1 U3681 ( .A1(n2981), .A2(n2958), .ZN(n4764) );
  NOR2_X1 U3682 ( .A1(n4454), .A2(n4762), .ZN(n2981) );
  NAND2_X1 U3683 ( .A1(n2983), .A2(n2958), .ZN(n4763) );
  NAND2_X1 U3684 ( .A1(n2983), .A2(n2957), .ZN(n4569) );
  XNOR2_X1 U3685 ( .A(n4177), .B(n6672), .ZN(n4512) );
  NOR2_X1 U3686 ( .A1(n4454), .A2(n4453), .ZN(n4567) );
  OR2_X1 U3687 ( .A1(n6030), .A2(n4907), .ZN(n5583) );
  AND2_X1 U3688 ( .A1(n4397), .A2(n5706), .ZN(n6030) );
  INV_X1 U3689 ( .A(n4518), .ZN(n4457) );
  INV_X1 U3690 ( .A(n4126), .ZN(n6380) );
  INV_X1 U3691 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4430) );
  AND2_X1 U3692 ( .A1(n6217), .A2(n4573), .ZN(n4580) );
  AND2_X1 U3693 ( .A1(n4663), .A2(n6218), .ZN(n4665) );
  AND2_X1 U3694 ( .A1(n4828), .A2(n6146), .ZN(n4787) );
  AND2_X1 U3695 ( .A1(n4825), .A2(n4824), .ZN(n6109) );
  INV_X1 U3696 ( .A(n6110), .ZN(n6113) );
  NAND2_X1 U3697 ( .A1(n6423), .A2(n4467), .ZN(n4744) );
  NOR2_X1 U3698 ( .A1(n4531), .A2(n5622), .ZN(n4537) );
  AND2_X1 U3699 ( .A1(n4468), .A2(n4467), .ZN(n4498) );
  INV_X1 U3700 ( .A(n4977), .ZN(n4824) );
  NOR2_X1 U3701 ( .A1(n4531), .A2(n4573), .ZN(n4463) );
  NOR2_X1 U3702 ( .A1(n6473), .A2(n5777), .ZN(n5766) );
  INV_X1 U3703 ( .A(n5845), .ZN(n5856) );
  INV_X1 U3704 ( .A(n5848), .ZN(n5858) );
  AND2_X1 U3705 ( .A1(n4883), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4884) );
  AND2_X1 U3706 ( .A1(n4953), .A2(n4880), .ZN(n5848) );
  AND2_X1 U3707 ( .A1(n4891), .A2(n5810), .ZN(n5843) );
  INV_X1 U3708 ( .A(n5353), .ZN(n5308) );
  NAND2_X1 U3709 ( .A1(n4136), .A2(n5936), .ZN(n5120) );
  CLKBUF_X1 U3710 ( .A(n5898), .Z(n6539) );
  INV_X1 U3711 ( .A(n5924), .ZN(n5978) );
  XNOR2_X1 U3712 ( .A(n4091), .B(n6638), .ZN(n4883) );
  OR2_X1 U3713 ( .A1(n4090), .A2(n4256), .ZN(n4091) );
  AND2_X1 U3714 ( .A1(n3817), .A2(n3031), .ZN(n4078) );
  AND2_X1 U3715 ( .A1(n3032), .A2(n3033), .ZN(n3031) );
  NAND2_X1 U3717 ( .A1(n5054), .A2(n5055), .ZN(n5983) );
  CLKBUF_X1 U3718 ( .A(n4691), .Z(n4692) );
  AOI21_X1 U3719 ( .B1(n4254), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4253), 
        .ZN(n4255) );
  AND2_X1 U3720 ( .A1(n5579), .A2(n5467), .ZN(n5543) );
  NOR2_X1 U3721 ( .A1(n5690), .A2(n5470), .ZN(n5579) );
  INV_X1 U3722 ( .A(n3003), .ZN(n3002) );
  NOR2_X1 U3723 ( .A1(n5708), .A2(n5094), .ZN(n6016) );
  AND2_X1 U3724 ( .A1(n4912), .A2(n4911), .ZN(n6066) );
  NAND2_X1 U3725 ( .A1(n4385), .A2(n4379), .ZN(n6099) );
  INV_X1 U3726 ( .A(n6097), .ZN(n6079) );
  INV_X1 U3727 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4660) );
  INV_X1 U3729 ( .A(n4573), .ZN(n5622) );
  AND2_X1 U3730 ( .A1(n6112), .A2(n4572), .ZN(n6217) );
  CLKBUF_X1 U3731 ( .A(n4418), .Z(n6146) );
  CLKBUF_X1 U3732 ( .A(n4517), .Z(n6110) );
  INV_X1 U3733 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4330) );
  INV_X1 U3734 ( .A(n6253), .ZN(n6555) );
  INV_X1 U3735 ( .A(n6281), .ZN(n6342) );
  INV_X1 U3736 ( .A(n6291), .ZN(n6354) );
  AND2_X1 U3737 ( .A1(n4537), .A2(n4977), .ZN(n6375) );
  AND2_X1 U3738 ( .A1(n3898), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U3739 ( .A1(n3876), .A2(n3875), .ZN(n6415) );
  OR2_X1 U3740 ( .A1(n3874), .A2(n4085), .ZN(n3875) );
  OR2_X1 U3741 ( .A1(n3873), .A2(n3872), .ZN(n3876) );
  INV_X1 U3742 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6520) );
  AND2_X1 U3743 ( .A1(n6413), .A2(n6412), .ZN(n6508) );
  NAND2_X1 U3744 ( .A1(n5353), .A2(n3900), .ZN(n3999) );
  NAND2_X1 U3745 ( .A1(n3025), .A2(n3708), .ZN(n5253) );
  NOR2_X1 U3746 ( .A1(n4453), .A2(n2984), .ZN(n2957) );
  OR2_X1 U3747 ( .A1(n5222), .A2(n5279), .ZN(n5268) );
  AND2_X1 U3748 ( .A1(n2957), .A2(n2982), .ZN(n2958) );
  NOR2_X1 U3749 ( .A1(n5261), .A2(n2973), .ZN(n2959) );
  AND2_X2 U3750 ( .A1(n4434), .A2(n4295), .ZN(n3275) );
  AND2_X1 U3751 ( .A1(n4458), .A2(n3006), .ZN(n2960) );
  INV_X1 U3752 ( .A(n4246), .ZN(n5335) );
  NAND2_X1 U3753 ( .A1(n4487), .A2(n3187), .ZN(n4348) );
  AND2_X1 U3754 ( .A1(n4821), .A2(n2972), .ZN(n4991) );
  AND2_X1 U3755 ( .A1(n4821), .A2(n4925), .ZN(n4926) );
  AND2_X1 U3756 ( .A1(n3005), .A2(n5055), .ZN(n2961) );
  NAND3_X1 U3757 ( .A1(n3877), .A2(n3179), .A3(n4381), .ZN(n3205) );
  AND4_X1 U3758 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n2962)
         );
  AND4_X1 U3759 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n2963)
         );
  NOR2_X1 U3760 ( .A1(n5222), .A2(n3029), .ZN(n2964) );
  AND4_X1 U3761 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n2965)
         );
  NAND2_X1 U3762 ( .A1(n4236), .A2(n4235), .ZN(n5457) );
  XNOR2_X1 U3763 ( .A(n4216), .B(n3453), .ZN(n4206) );
  OR2_X1 U3764 ( .A1(n4977), .A2(n4158), .ZN(n2966) );
  INV_X1 U3765 ( .A(n4237), .ZN(n3011) );
  NAND2_X1 U3766 ( .A1(n4226), .A2(n5458), .ZN(n2967) );
  OR2_X1 U3767 ( .A1(n4348), .A2(n2977), .ZN(n2968) );
  INV_X1 U3768 ( .A(n3013), .ZN(n3012) );
  NAND2_X1 U3769 ( .A1(n4235), .A2(n2967), .ZN(n3013) );
  INV_X1 U3770 ( .A(n5449), .ZN(n4238) );
  OR2_X1 U3771 ( .A1(n4172), .A2(n3356), .ZN(n2969) );
  NOR2_X2 U3772 ( .A1(n3214), .A2(n6414), .ZN(n3583) );
  NAND2_X1 U3773 ( .A1(n5076), .A2(n5079), .ZN(n5078) );
  AND2_X1 U3774 ( .A1(n4778), .A2(n3492), .ZN(n4821) );
  AND2_X1 U3775 ( .A1(n2987), .A2(n2986), .ZN(n2970) );
  AND2_X1 U3776 ( .A1(n4226), .A2(n5704), .ZN(n2971) );
  NAND2_X1 U3777 ( .A1(n4229), .A2(n4228), .ZN(n5054) );
  NAND2_X1 U3778 ( .A1(n3000), .A2(n3002), .ZN(n5085) );
  AND2_X1 U3779 ( .A1(n4925), .A2(n4992), .ZN(n2972) );
  NAND2_X1 U3780 ( .A1(n3024), .A2(n3708), .ZN(n2973) );
  OR2_X1 U3781 ( .A1(n2953), .A2(n4244), .ZN(n2974) );
  AND2_X1 U3782 ( .A1(n3884), .A2(n3187), .ZN(n2975) );
  AND2_X1 U3783 ( .A1(n3557), .A2(n3545), .ZN(n5063) );
  AND2_X1 U3784 ( .A1(n2970), .A2(n2985), .ZN(n2976) );
  NAND2_X1 U3785 ( .A1(n3374), .A2(n3298), .ZN(n4518) );
  NAND2_X1 U3786 ( .A1(n3446), .A2(n3445), .ZN(n4761) );
  NAND3_X1 U3787 ( .A1(n4890), .A2(n3209), .A3(n3895), .ZN(n3889) );
  INV_X1 U3788 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6423) );
  NAND2_X1 U3789 ( .A1(n3019), .A2(n4890), .ZN(n3877) );
  OR2_X1 U3790 ( .A1(n4414), .A2(n4415), .ZN(n4454) );
  INV_X1 U3791 ( .A(n4454), .ZN(n2983) );
  INV_X1 U3792 ( .A(EBX_REG_1__SCAN_IN), .ZN(n2978) );
  INV_X1 U3793 ( .A(n2994), .ZN(n5200) );
  NOR2_X4 U3794 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4437) );
  OAI21_X2 U3795 ( .B1(n3001), .B2(n2998), .A(n2996), .ZN(n5681) );
  NAND2_X1 U3796 ( .A1(n3373), .A2(n4458), .ZN(n3397) );
  NAND2_X1 U3797 ( .A1(n3007), .A2(n3008), .ZN(n5441) );
  NAND2_X1 U3798 ( .A1(n4236), .A2(n3010), .ZN(n3007) );
  INV_X1 U3799 ( .A(n5421), .ZN(n5448) );
  OAI21_X1 U3800 ( .B1(n5493), .B2(n5992), .A(n4250), .ZN(U2955) );
  XNOR2_X1 U3801 ( .A(n3018), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5493)
         );
  OAI22_X1 U3802 ( .A1(n5325), .A2(n5484), .B1(n5361), .B2(n4249), .ZN(n3018)
         );
  AND2_X4 U3803 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4295) );
  NOR2_X1 U3804 ( .A1(n3036), .A2(n3019), .ZN(n4080) );
  NAND2_X1 U3805 ( .A1(n3020), .A2(n2969), .ZN(n3249) );
  NAND3_X1 U3806 ( .A1(n3350), .A2(n3234), .A3(n6423), .ZN(n3020) );
  NAND2_X1 U3807 ( .A1(n3350), .A2(n3234), .ZN(n4315) );
  NAND2_X1 U3808 ( .A1(n5076), .A2(n3021), .ZN(n5235) );
  NAND2_X2 U3809 ( .A1(n5068), .A2(n3557), .ZN(n5076) );
  NAND2_X1 U3810 ( .A1(n4821), .A2(n3030), .ZN(n3544) );
  NAND2_X1 U3811 ( .A1(n3544), .A2(n3543), .ZN(n3545) );
  AND2_X1 U3812 ( .A1(n3817), .A2(n3034), .ZN(n5140) );
  NAND2_X1 U3813 ( .A1(n3817), .A2(n3816), .ZN(n4026) );
  NAND2_X1 U3815 ( .A1(n4149), .A2(n4138), .ZN(n4140) );
  AND2_X2 U3817 ( .A1(n3052), .A2(n5107), .ZN(n3131) );
  AND2_X2 U3818 ( .A1(n5107), .A2(n3058), .ZN(n3239) );
  NAND4_X2 U3819 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3178)
         );
  NAND2_X1 U3820 ( .A1(n3119), .A2(n3894), .ZN(n3200) );
  AOI22_X1 U3821 ( .A1(n3316), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U3822 ( .A1(n3119), .A2(n3178), .ZN(n3186) );
  INV_X1 U3823 ( .A(n3178), .ZN(n3095) );
  AND2_X1 U3824 ( .A1(n5785), .A2(n4884), .ZN(n4892) );
  NAND2_X1 U3825 ( .A1(n5785), .A2(n4092), .ZN(n5810) );
  NAND2_X1 U3826 ( .A1(n5878), .A2(n4137), .ZN(n5872) );
  INV_X1 U3827 ( .A(n5872), .ZN(n3996) );
  INV_X1 U3828 ( .A(n5300), .ZN(n3900) );
  NOR2_X1 U3829 ( .A1(n6007), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3035)
         );
  OR2_X1 U3830 ( .A1(n4141), .A2(n3187), .ZN(n3036) );
  XNOR2_X1 U3831 ( .A(n3447), .B(n3448), .ZN(n4196) );
  OR2_X1 U3832 ( .A1(n4226), .A2(n5420), .ZN(n3037) );
  INV_X1 U3833 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5828) );
  INV_X1 U3834 ( .A(n5521), .ZN(n3997) );
  OR2_X2 U3835 ( .A1(n5118), .A2(n5987), .ZN(n3038) );
  OAI21_X1 U3836 ( .B1(n3452), .B2(n3440), .A(n3439), .ZN(n3448) );
  NAND2_X1 U3837 ( .A1(n4079), .A2(n3213), .ZN(n3216) );
  INV_X1 U3838 ( .A(n3457), .ZN(n3458) );
  AOI22_X1 U3839 ( .A1(n3271), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        INSTQUEUE_REG_1__6__SCAN_IN), .B2(n3140), .ZN(n3074) );
  NAND2_X1 U3840 ( .A1(n3209), .A2(n4469), .ZN(n3210) );
  INV_X1 U3841 ( .A(n5263), .ZN(n3708) );
  INV_X1 U3842 ( .A(n4820), .ZN(n3492) );
  OR2_X1 U3843 ( .A1(n3262), .A2(n3261), .ZN(n4151) );
  OR2_X1 U3844 ( .A1(n3221), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3222)
         );
  OR2_X1 U3845 ( .A1(n3370), .A2(n3369), .ZN(n4180) );
  INV_X1 U3846 ( .A(n3818), .ZN(n3816) );
  OAI21_X1 U3847 ( .B1(n3452), .B2(n3421), .A(n3420), .ZN(n3427) );
  AND2_X1 U3848 ( .A1(n3791), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3792)
         );
  INV_X1 U3849 ( .A(n3337), .ZN(n4015) );
  INV_X1 U3850 ( .A(n3573), .ZN(n3574) );
  INV_X1 U3851 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3376) );
  AND2_X1 U3852 ( .A1(n5467), .A2(n5594), .ZN(n4244) );
  NAND2_X1 U3853 ( .A1(n3188), .A2(n4469), .ZN(n3905) );
  AND2_X1 U3854 ( .A1(n5982), .A2(n4231), .ZN(n4232) );
  INV_X1 U3855 ( .A(n2975), .ZN(n3976) );
  AND2_X1 U3856 ( .A1(n3230), .A2(n6111), .ZN(n4593) );
  AND2_X1 U3857 ( .A1(n3654), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3655)
         );
  AND2_X1 U3858 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3704), .ZN(n3705)
         );
  INV_X1 U3859 ( .A(n4069), .ZN(n4042) );
  AND2_X1 U3860 ( .A1(n3925), .A2(n3924), .ZN(n4693) );
  AND2_X1 U3861 ( .A1(n4623), .A2(n6218), .ZN(n4625) );
  OAI211_X1 U3862 ( .C1(n6549), .C2(n6512), .A(n4986), .B(n4985), .ZN(n6548)
         );
  INV_X1 U3863 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U3864 ( .A1(n3355), .A2(n3354), .ZN(n6326) );
  AND2_X1 U3865 ( .A1(n5186), .A2(n4118), .ZN(n5154) );
  NAND2_X1 U3866 ( .A1(n3705), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3748)
         );
  NOR2_X1 U3867 ( .A1(n3590), .A2(n5238), .ZN(n3605) );
  INV_X1 U3868 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U3869 ( .A1(n4953), .A2(n4110), .ZN(n5787) );
  INV_X1 U3870 ( .A(n3187), .ZN(n3306) );
  NAND2_X1 U3871 ( .A1(n3749), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3790)
         );
  NAND2_X1 U3872 ( .A1(n3605), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3619)
         );
  AND2_X1 U3873 ( .A1(n3535), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3539)
         );
  INV_X1 U3874 ( .A(n5325), .ZN(n4254) );
  INV_X1 U3875 ( .A(n5158), .ZN(n5144) );
  OR2_X1 U3876 ( .A1(n4364), .A2(n4363), .ZN(n4365) );
  OR2_X1 U3877 ( .A1(n4629), .A2(n4977), .ZN(n4864) );
  INV_X1 U3878 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4985) );
  INV_X1 U3879 ( .A(n6146), .ZN(n6317) );
  INV_X1 U3880 ( .A(n4150), .ZN(n4573) );
  INV_X1 U3881 ( .A(n5810), .ZN(n4093) );
  AND2_X1 U3882 ( .A1(n5785), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5845) );
  AND2_X1 U3883 ( .A1(n4953), .A2(n4107), .ZN(n5825) );
  OR2_X1 U3884 ( .A1(n6536), .A2(n4089), .ZN(n5785) );
  AND2_X1 U3885 ( .A1(n5120), .A2(n4137), .ZN(n4138) );
  INV_X1 U3886 ( .A(n5936), .ZN(n5977) );
  OR2_X1 U3887 ( .A1(n6525), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4143) );
  AND2_X1 U3888 ( .A1(n4385), .A2(n6383), .ZN(n5719) );
  INV_X1 U3889 ( .A(n6032), .ZN(n6076) );
  INV_X1 U3890 ( .A(n6086), .ZN(n6102) );
  AND2_X1 U3891 ( .A1(n4385), .A2(n4375), .ZN(n6097) );
  INV_X1 U3892 ( .A(n4868), .ZN(n6139) );
  AND2_X1 U3893 ( .A1(n4580), .A2(n4977), .ZN(n6208) );
  AND2_X1 U3894 ( .A1(n4575), .A2(n6206), .ZN(n4578) );
  OR2_X1 U3895 ( .A1(n4746), .A2(n4745), .ZN(n6271) );
  NOR2_X1 U3896 ( .A1(n4668), .A2(n4977), .ZN(n4816) );
  OR2_X1 U3897 ( .A1(n6331), .A2(n6330), .ZN(n6376) );
  AND2_X1 U3898 ( .A1(DATAI_1_), .A2(n4702), .ZN(n6336) );
  INV_X1 U3899 ( .A(n6307), .ZN(n6550) );
  INV_X1 U3900 ( .A(n4698), .ZN(n4733) );
  AND2_X1 U3901 ( .A1(n4463), .A2(n4824), .ZN(n4619) );
  OR2_X1 U3902 ( .A1(n4364), .A2(n4270), .ZN(n4281) );
  INV_X1 U3903 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6322) );
  AND2_X1 U3904 ( .A1(n5636), .A2(n4116), .ZN(n5186) );
  INV_X1 U3905 ( .A(n5825), .ZN(n5861) );
  AOI21_X1 U3906 ( .B1(n3997), .B2(n3996), .A(n3995), .ZN(n3998) );
  INV_X1 U3907 ( .A(n5322), .ZN(n4782) );
  OR2_X1 U3908 ( .A1(n4364), .A2(n4261), .ZN(n5919) );
  INV_X1 U3909 ( .A(n5965), .ZN(n5924) );
  OR2_X1 U3910 ( .A1(n4364), .A2(n6411), .ZN(n5980) );
  OR2_X1 U3911 ( .A1(n6431), .A2(n6325), .ZN(n5987) );
  OR2_X1 U3912 ( .A1(n6006), .A2(n4404), .ZN(n6015) );
  NAND2_X1 U3913 ( .A1(n4385), .A2(n4371), .ZN(n6086) );
  OR2_X1 U3914 ( .A1(n4629), .A2(n4824), .ZN(n4658) );
  NAND2_X1 U3915 ( .A1(n6110), .A2(n6109), .ZN(n6176) );
  NAND2_X1 U3916 ( .A1(n4580), .A2(n4824), .ZN(n6558) );
  NAND2_X1 U3917 ( .A1(n6217), .A2(n4978), .ZN(n6253) );
  NAND2_X1 U3918 ( .A1(n6217), .A2(n4739), .ZN(n6274) );
  INV_X1 U3919 ( .A(n4816), .ZN(n4688) );
  NAND2_X1 U3920 ( .A1(n6109), .A2(n6113), .ZN(n6379) );
  NAND2_X1 U3921 ( .A1(n4463), .A2(n4977), .ZN(n4736) );
  INV_X1 U3922 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U3923 ( .A1(n3999), .A2(n3998), .ZN(U2832) );
  NAND2_X1 U3924 ( .A1(n3251), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3045)
         );
  INV_X1 U3925 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3040) );
  AND2_X2 U3926 ( .A1(n3040), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3052)
         );
  NAND2_X1 U3927 ( .A1(n3131), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3044) );
  INV_X1 U3928 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3041) );
  NAND2_X1 U3929 ( .A1(n3307), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U3930 ( .A1(n3155), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3042)
         );
  INV_X1 U3931 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3046) );
  AND2_X4 U3932 ( .A1(n3047), .A2(n3058), .ZN(n3256) );
  NAND2_X1 U3933 ( .A1(n3256), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3051)
         );
  AND2_X4 U3934 ( .A1(n3058), .A2(n4437), .ZN(n3316) );
  NAND2_X1 U3935 ( .A1(n3316), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3050) );
  NOR2_X4 U3936 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3053) );
  NAND2_X1 U3938 ( .A1(n3271), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3049) );
  NAND2_X1 U3939 ( .A1(n3140), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3048) );
  NAND2_X1 U3940 ( .A1(n3310), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3057) );
  AND2_X4 U3941 ( .A1(n3052), .A2(n4295), .ZN(n3145) );
  NAND2_X1 U3942 ( .A1(n3145), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3056) );
  AND2_X4 U3943 ( .A1(n4437), .A2(n3053), .ZN(n3265) );
  NAND2_X1 U3944 ( .A1(n3265), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3055) );
  AND2_X4 U3945 ( .A1(n3053), .A2(n4295), .ZN(n3272) );
  NAND2_X1 U3946 ( .A1(n3272), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3054) );
  NAND2_X1 U3947 ( .A1(n3239), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3062) );
  AND2_X4 U3948 ( .A1(n3058), .A2(n4295), .ZN(n3362) );
  NAND2_X1 U3949 ( .A1(n3362), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3061)
         );
  NAND2_X1 U3950 ( .A1(n3146), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3060)
         );
  NAND2_X1 U3951 ( .A1(n3275), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3059)
         );
  AOI22_X1 U3952 ( .A1(n3131), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3251), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3070) );
  AOI22_X1 U3953 ( .A1(n3307), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U3954 ( .A1(n3310), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3068) );
  AOI22_X1 U3955 ( .A1(n3145), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3067) );
  AOI22_X1 U3956 ( .A1(n3239), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3073) );
  AOI22_X1 U3957 ( .A1(n3256), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3072) );
  AOI22_X1 U3958 ( .A1(n3362), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3146), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3071) );
  NAND2_X1 U3960 ( .A1(n3155), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3078)
         );
  NAND2_X1 U3961 ( .A1(n3307), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3077) );
  NAND2_X1 U3962 ( .A1(n3251), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3076)
         );
  NAND2_X1 U3963 ( .A1(n3265), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U3964 ( .A1(n3316), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3082) );
  NAND2_X1 U3965 ( .A1(n3362), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3081)
         );
  NAND2_X1 U3966 ( .A1(n3271), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3080) );
  NAND2_X1 U3967 ( .A1(n3140), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3079) );
  NAND2_X1 U3968 ( .A1(n3239), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3086) );
  NAND2_X1 U3969 ( .A1(n3256), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3085)
         );
  NAND2_X1 U3970 ( .A1(n3272), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U3971 ( .A1(n3275), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3083)
         );
  NAND2_X1 U3973 ( .A1(n3310), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3974 ( .A1(n3131), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U3975 ( .A1(n2955), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3976 ( .A1(n3146), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3087)
         );
  OAI21_X1 U3977 ( .B1(n4372), .B2(n3214), .A(n3176), .ZN(n3105) );
  AOI22_X1 U3978 ( .A1(n3251), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3099) );
  AOI22_X1 U3979 ( .A1(n3145), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3098) );
  AOI22_X1 U3980 ( .A1(n3239), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3097) );
  AOI22_X1 U3981 ( .A1(n3256), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3096) );
  AOI22_X1 U3982 ( .A1(n3131), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3103) );
  AOI22_X1 U3983 ( .A1(n3271), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3102) );
  AOI22_X1 U3984 ( .A1(n3310), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3101) );
  AOI22_X1 U3985 ( .A1(n3272), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3146), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3100) );
  NAND2_X1 U3986 ( .A1(n3105), .A2(n3183), .ZN(n3118) );
  AOI22_X1 U3987 ( .A1(n3131), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3111) );
  AOI22_X1 U3988 ( .A1(n3310), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U3989 ( .A1(n3239), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3146), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U3990 ( .A1(n3256), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U3991 ( .A1(n3307), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3251), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U3992 ( .A1(n3145), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U3993 ( .A1(n3362), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3112) );
  NAND2_X2 U3994 ( .A1(n2965), .A2(n3116), .ZN(n3894) );
  NAND4_X1 U3995 ( .A1(n3176), .A2(n4497), .A3(n3200), .A4(n4372), .ZN(n3117)
         );
  NAND2_X1 U3996 ( .A1(n3118), .A2(n3117), .ZN(n3130) );
  AOI22_X1 U3997 ( .A1(n3131), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3251), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U3998 ( .A1(n3307), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3122) );
  AOI22_X1 U3999 ( .A1(n3310), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3121) );
  AOI22_X1 U4000 ( .A1(n3145), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U4001 ( .A1(n3239), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U4002 ( .A1(n3362), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3146), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U4003 ( .A1(n3256), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U4004 ( .A1(n3271), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3140), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3124) );
  NAND2_X1 U4005 ( .A1(n3251), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3135)
         );
  NAND2_X1 U4006 ( .A1(n3131), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U4007 ( .A1(n3307), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U4008 ( .A1(n3155), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3132)
         );
  NAND2_X1 U4009 ( .A1(n3239), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3139) );
  NAND2_X1 U4010 ( .A1(n3362), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3138)
         );
  NAND2_X1 U4011 ( .A1(n3256), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3137)
         );
  NAND2_X1 U4012 ( .A1(n3316), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U4013 ( .A1(n3310), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U4014 ( .A1(n3271), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U4015 ( .A1(n3140), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U4016 ( .A1(n3275), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3141)
         );
  NAND2_X1 U4017 ( .A1(n3145), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U4018 ( .A1(n3272), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4019 ( .A1(n3265), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4020 ( .A1(n3146), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3147)
         );
  NAND2_X1 U4021 ( .A1(n3251), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3159)
         );
  NAND2_X1 U4022 ( .A1(n3131), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U4023 ( .A1(n3307), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U4024 ( .A1(n3155), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3156)
         );
  NAND2_X1 U4025 ( .A1(n3256), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3163)
         );
  NAND2_X1 U4026 ( .A1(n3316), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3162) );
  NAND2_X1 U4027 ( .A1(n3271), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U4028 ( .A1(n3140), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U4029 ( .A1(n3310), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U4030 ( .A1(n3145), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4031 ( .A1(n3265), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U4032 ( .A1(n3272), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U4033 ( .A1(n3239), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4034 ( .A1(n3362), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3170)
         );
  NAND2_X1 U4035 ( .A1(n3146), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3169)
         );
  NAND2_X1 U4036 ( .A1(n3275), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3168)
         );
  NAND4_X4 U4037 ( .A1(n3175), .A2(n3174), .A3(n3173), .A4(n3172), .ZN(n3187)
         );
  AND2_X1 U4038 ( .A1(n4372), .A2(n3894), .ZN(n3177) );
  NAND2_X1 U4039 ( .A1(n3208), .A2(n4283), .ZN(n3179) );
  BUF_X4 U4040 ( .A(n3178), .Z(n4479) );
  AND2_X1 U4041 ( .A1(n2954), .A2(n3894), .ZN(n3182) );
  OR2_X1 U4042 ( .A1(n3186), .A2(n4491), .ZN(n3181) );
  NAND2_X1 U4043 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6435) );
  OAI21_X1 U4044 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6435), .ZN(n4108) );
  NAND2_X1 U4045 ( .A1(n3826), .A2(n4108), .ZN(n3213) );
  NAND2_X1 U4046 ( .A1(n3878), .A2(n3184), .ZN(n3185) );
  NAND2_X1 U4047 ( .A1(n3190), .A2(n3189), .ZN(n3227) );
  NAND2_X1 U4048 ( .A1(n3227), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3195) );
  INV_X1 U4049 ( .A(n3898), .ZN(n3192) );
  NAND2_X1 U4050 ( .A1(n6512), .A2(n6520), .ZN(n6525) );
  INV_X1 U4051 ( .A(n4143), .ZN(n3191) );
  MUX2_X1 U4052 ( .A(n3192), .B(n3191), .S(n4660), .Z(n3193) );
  INV_X1 U4053 ( .A(n3193), .ZN(n3194) );
  INV_X1 U4054 ( .A(n3878), .ZN(n3198) );
  NAND2_X1 U4055 ( .A1(n4337), .A2(n4491), .ZN(n3196) );
  NAND2_X1 U4056 ( .A1(n3196), .A2(n4469), .ZN(n3197) );
  OAI21_X1 U4057 ( .B1(n3198), .B2(n3197), .A(n4487), .ZN(n3204) );
  NAND2_X1 U4058 ( .A1(n4141), .A2(n4487), .ZN(n3199) );
  MUX2_X1 U4059 ( .A(n3199), .B(n3183), .S(n3187), .Z(n3887) );
  INV_X1 U4060 ( .A(n3891), .ZN(n3330) );
  OR2_X1 U4061 ( .A1(n6525), .A2(n6423), .ZN(n6425) );
  AOI21_X1 U4062 ( .B1(n3330), .B2(n3895), .A(n6425), .ZN(n3203) );
  NAND2_X1 U4063 ( .A1(n3201), .A2(n4283), .ZN(n3202) );
  INV_X1 U4064 ( .A(n3205), .ZN(n3206) );
  NAND2_X2 U4065 ( .A1(n3289), .A2(n3291), .ZN(n3290) );
  INV_X1 U4066 ( .A(n3290), .ZN(n3226) );
  NAND2_X1 U4067 ( .A1(n3227), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4068 ( .A1(n4080), .A2(n3826), .ZN(n4128) );
  INV_X1 U4069 ( .A(n3208), .ZN(n3212) );
  INV_X1 U4070 ( .A(n4479), .ZN(n3209) );
  NAND2_X1 U4071 ( .A1(n3214), .A2(n3894), .ZN(n4360) );
  INV_X1 U4073 ( .A(n4373), .ZN(n3215) );
  NAND3_X1 U4074 ( .A1(n4128), .A2(n3216), .A3(n3215), .ZN(n3217) );
  NAND2_X1 U4075 ( .A1(n3217), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3220) );
  XNOR2_X1 U4076 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4979) );
  OAI22_X1 U4077 ( .A1(n4143), .A2(n4979), .B1(n3898), .B2(n6387), .ZN(n3221)
         );
  INV_X1 U4078 ( .A(n3221), .ZN(n3218) );
  INV_X1 U4080 ( .A(n3220), .ZN(n3223) );
  NAND2_X1 U4081 ( .A1(n3223), .A2(n3222), .ZN(n3224) );
  NAND2_X1 U4083 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4084 ( .A1(n3229), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3230) );
  NOR2_X1 U4085 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6387), .ZN(n4823)
         );
  NAND2_X1 U4086 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4823), .ZN(n6111) );
  OAI22_X1 U4087 ( .A1(n4143), .A2(n4593), .B1(n3898), .B2(n6391), .ZN(n3231)
         );
  NAND2_X1 U4088 ( .A1(n3233), .A2(n3232), .ZN(n3234) );
  AOI22_X1 U4089 ( .A1(n4046), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3238) );
  INV_X1 U4090 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6699) );
  AOI22_X1 U4091 ( .A1(n4052), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4093 ( .A1(n3273), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3236) );
  BUF_X1 U4094 ( .A(n3145), .Z(n3274) );
  AOI22_X1 U4095 ( .A1(n3145), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3235) );
  NAND4_X1 U4096 ( .A1(n3238), .A2(n3237), .A3(n3236), .A4(n3235), .ZN(n3245)
         );
  BUF_X1 U4097 ( .A(n3316), .Z(n3264) );
  AOI22_X1 U4098 ( .A1(n3309), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3243) );
  CLKBUF_X2 U4099 ( .A(n3140), .Z(n3308) );
  AOI22_X1 U4100 ( .A1(n3271), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4101 ( .A1(n3266), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4102 ( .A1(n4054), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3240) );
  NAND4_X1 U4103 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3244)
         );
  AOI22_X1 U4104 ( .A1(n3246), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3284), 
        .B2(n3247), .ZN(n3248) );
  XNOR2_X1 U4105 ( .A(n3290), .B(n3250), .ZN(n4459) );
  INV_X1 U4106 ( .A(n3356), .ZN(n3283) );
  AOI22_X1 U4107 ( .A1(n3131), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4108 ( .A1(n4033), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4109 ( .A1(n4054), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4110 ( .A1(n3266), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3252) );
  NAND4_X1 U4111 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3262)
         );
  AOI22_X1 U4113 ( .A1(n3309), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4114 ( .A1(n4052), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4115 ( .A1(n3145), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4116 ( .A1(n3264), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3257) );
  NAND4_X1 U4117 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .ZN(n3261)
         );
  NAND2_X1 U4118 ( .A1(n3283), .A2(n4151), .ZN(n3263) );
  OAI21_X2 U4119 ( .B1(n4459), .B2(STATE2_REG_0__SCAN_IN), .A(n3263), .ZN(
        n3292) );
  INV_X1 U4120 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4121 ( .A1(n3131), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4122 ( .A1(n4052), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3155), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4123 ( .A1(n3264), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3268) );
  BUF_X1 U4124 ( .A(n3362), .Z(n3266) );
  AOI22_X1 U4125 ( .A1(n3266), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3267) );
  NAND4_X1 U4126 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3281)
         );
  AOI22_X1 U4127 ( .A1(n3256), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3279) );
  BUF_X1 U4128 ( .A(n3310), .Z(n3273) );
  BUF_X1 U4129 ( .A(n3272), .Z(n3364) );
  AOI22_X1 U4130 ( .A1(n3273), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4131 ( .A1(n3145), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4132 ( .A1(n4054), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3276) );
  NAND4_X1 U4133 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), .ZN(n3280)
         );
  INV_X1 U4134 ( .A(n4220), .ZN(n3282) );
  NAND2_X1 U4135 ( .A1(n3283), .A2(n3282), .ZN(n3305) );
  NAND2_X1 U4136 ( .A1(n3284), .A2(n4151), .ZN(n3285) );
  OAI211_X1 U4137 ( .C1(n3452), .C2(n3286), .A(n3305), .B(n3285), .ZN(n3287)
         );
  INV_X1 U4138 ( .A(n3287), .ZN(n3288) );
  NAND2_X1 U4139 ( .A1(n4372), .A2(n4220), .ZN(n4217) );
  MUX2_X2 U4140 ( .A(n4217), .B(n2956), .S(n6423), .Z(n3299) );
  INV_X1 U4141 ( .A(n3292), .ZN(n3293) );
  INV_X1 U4142 ( .A(n3294), .ZN(n3297) );
  INV_X1 U4143 ( .A(n3295), .ZN(n3296) );
  NAND2_X1 U4144 ( .A1(n3297), .A2(n3296), .ZN(n3298) );
  NAND2_X1 U4145 ( .A1(n4150), .A2(n3583), .ZN(n3304) );
  AOI22_X1 U4146 ( .A1(n3337), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6414), .ZN(n3302) );
  INV_X1 U4147 ( .A(n4360), .ZN(n3879) );
  NAND2_X1 U4148 ( .A1(n3879), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3381) );
  INV_X1 U4149 ( .A(n3381), .ZN(n3399) );
  NAND2_X1 U4150 ( .A1(n3399), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3301) );
  AND2_X1 U4151 ( .A1(n3302), .A2(n3301), .ZN(n3303) );
  INV_X1 U4152 ( .A(n3305), .ZN(n3323) );
  AOI22_X1 U4153 ( .A1(n4052), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4154 ( .A1(n3145), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4155 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3309), .B1(n3308), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4156 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3273), .B1(n3363), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4157 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3322)
         );
  AOI22_X1 U4158 ( .A1(n4046), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4159 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n3271), .B1(n3264), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4160 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4047), .B1(n3364), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4161 ( .A1(n4054), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3317) );
  NAND4_X1 U4162 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3321)
         );
  OR2_X1 U4163 ( .A1(n3322), .A2(n3321), .ZN(n4160) );
  OAI21_X1 U4164 ( .B1(n3323), .B2(n4332), .A(n4160), .ZN(n3327) );
  INV_X1 U4165 ( .A(n4217), .ZN(n3324) );
  AOI21_X1 U4166 ( .B1(n3324), .B2(n4160), .A(n6423), .ZN(n3326) );
  NAND2_X1 U4167 ( .A1(n3246), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3325) );
  NAND3_X1 U4168 ( .A1(n3327), .A2(n3326), .A3(n3325), .ZN(n3328) );
  AOI21_X1 U4169 ( .B1(n4977), .B2(n3330), .A(n6414), .ZN(n4339) );
  INV_X1 U4170 ( .A(n3583), .ZN(n3572) );
  OR2_X1 U4171 ( .A1(n2956), .A2(n3572), .ZN(n3334) );
  AOI22_X1 U4172 ( .A1(n3337), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6414), .ZN(n3332) );
  NAND2_X1 U4173 ( .A1(n3399), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3331) );
  AND2_X1 U4174 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  NAND2_X1 U4175 ( .A1(n3334), .A2(n3333), .ZN(n4338) );
  NAND2_X1 U4176 ( .A1(n4339), .A2(n4338), .ZN(n4341) );
  INV_X1 U4177 ( .A(n4338), .ZN(n3335) );
  NAND2_X1 U4178 ( .A1(n6414), .A2(n6322), .ZN(n3338) );
  NAND2_X1 U4179 ( .A1(n3335), .A2(n4072), .ZN(n3336) );
  NAND2_X1 U4180 ( .A1(n4341), .A2(n3336), .ZN(n4344) );
  NAND2_X1 U4181 ( .A1(n4345), .A2(n4344), .ZN(n3347) );
  INV_X1 U4182 ( .A(n3347), .ZN(n3345) );
  NAND2_X1 U4183 ( .A1(n3399), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3343) );
  INV_X1 U4184 ( .A(n3338), .ZN(n4072) );
  OAI21_X1 U4185 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3377), .ZN(n6014) );
  INV_X1 U4186 ( .A(n6014), .ZN(n3340) );
  INV_X1 U4187 ( .A(n4075), .ZN(n3422) );
  INV_X1 U4188 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3339) );
  OAI22_X1 U4189 ( .A1(n3338), .A2(n3340), .B1(n3422), .B2(n3339), .ZN(n3341)
         );
  AOI21_X1 U4190 ( .B1(n4076), .B2(EAX_REG_2__SCAN_IN), .A(n3341), .ZN(n3342)
         );
  AND2_X1 U4191 ( .A1(n3343), .A2(n3342), .ZN(n4411) );
  INV_X1 U4192 ( .A(n4411), .ZN(n3344) );
  NAND2_X1 U4193 ( .A1(n3345), .A2(n3344), .ZN(n3346) );
  NAND2_X1 U4194 ( .A1(n4412), .A2(n3346), .ZN(n3349) );
  NAND2_X1 U4195 ( .A1(n3347), .A2(n4411), .ZN(n3348) );
  NAND2_X1 U4196 ( .A1(n3349), .A2(n3348), .ZN(n4410) );
  INV_X1 U4197 ( .A(n4410), .ZN(n3385) );
  INV_X1 U4198 ( .A(n3374), .ZN(n3373) );
  NAND2_X1 U4199 ( .A1(n3228), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3355) );
  NAND3_X1 U4200 ( .A1(n4985), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6228) );
  INV_X1 U4201 ( .A(n6228), .ZN(n3351) );
  NAND2_X1 U4202 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3351), .ZN(n6252) );
  NAND2_X1 U4203 ( .A1(n4985), .A2(n6252), .ZN(n3352) );
  NAND3_X1 U4204 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4697) );
  INV_X1 U4205 ( .A(n4697), .ZN(n4465) );
  NAND2_X1 U4206 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4465), .ZN(n4499) );
  NAND2_X1 U4207 ( .A1(n3352), .A2(n4499), .ZN(n4589) );
  OAI22_X1 U4208 ( .A1(n4143), .A2(n4589), .B1(n3898), .B2(n4985), .ZN(n3353)
         );
  INV_X1 U4209 ( .A(n3353), .ZN(n3354) );
  AOI22_X1 U4210 ( .A1(n4045), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4211 ( .A1(n4052), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4212 ( .A1(n3309), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4213 ( .A1(n4053), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3358) );
  NAND4_X1 U4214 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n3370)
         );
  AOI22_X1 U4215 ( .A1(n4054), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4216 ( .A1(n4046), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4217 ( .A1(n3364), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4218 ( .A1(n3264), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4219 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3369)
         );
  AOI22_X1 U4220 ( .A1(n3246), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3843), 
        .B2(n4180), .ZN(n3371) );
  INV_X1 U4221 ( .A(n4458), .ZN(n4572) );
  NAND2_X1 U4222 ( .A1(n3374), .A2(n4572), .ZN(n3375) );
  INV_X1 U4223 ( .A(n3377), .ZN(n3378) );
  INV_X1 U4224 ( .A(n3401), .ZN(n3402) );
  OAI21_X1 U4225 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3378), .A(n3402), 
        .ZN(n5022) );
  AOI22_X1 U4226 ( .A1(n4072), .A2(n5022), .B1(n4075), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3380) );
  NAND2_X1 U4227 ( .A1(n4076), .A2(EAX_REG_3__SCAN_IN), .ZN(n3379) );
  OAI211_X1 U4228 ( .C1(n3381), .C2(n4430), .A(n3380), .B(n3379), .ZN(n3382)
         );
  INV_X1 U4229 ( .A(n3384), .ZN(n4452) );
  NAND2_X1 U4230 ( .A1(n3385), .A2(n3384), .ZN(n4450) );
  AOI22_X1 U4231 ( .A1(n4046), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4232 ( .A1(n4052), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4233 ( .A1(n3273), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4234 ( .A1(n3145), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3386) );
  NAND4_X1 U4235 ( .A1(n3389), .A2(n3388), .A3(n3387), .A4(n3386), .ZN(n3395)
         );
  AOI22_X1 U4236 ( .A1(n3309), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4237 ( .A1(n4053), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4238 ( .A1(n3266), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4239 ( .A1(n4054), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3390) );
  NAND4_X1 U4240 ( .A1(n3393), .A2(n3392), .A3(n3391), .A4(n3390), .ZN(n3394)
         );
  AOI22_X1 U4241 ( .A1(n3246), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3843), 
        .B2(n4197), .ZN(n3396) );
  NAND2_X1 U4242 ( .A1(n3397), .A2(n3396), .ZN(n3398) );
  NAND2_X1 U4243 ( .A1(n3399), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3408) );
  INV_X1 U4244 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3403) );
  AOI21_X1 U4245 ( .B1(n3403), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3400) );
  AOI21_X1 U4246 ( .B1(n4076), .B2(EAX_REG_4__SCAN_IN), .A(n3400), .ZN(n3407)
         );
  INV_X1 U4247 ( .A(n3441), .ZN(n3405) );
  NAND2_X1 U4248 ( .A1(n3403), .A2(n3402), .ZN(n3404) );
  NAND2_X1 U4249 ( .A1(n3405), .A2(n3404), .ZN(n6005) );
  NOR2_X1 U4250 ( .A1(n6005), .A2(n3338), .ZN(n3406) );
  AOI21_X1 U4251 ( .B1(n3408), .B2(n3407), .A(n3406), .ZN(n3409) );
  INV_X1 U4252 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4253 ( .A1(n3273), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4254 ( .A1(n4054), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4255 ( .A1(n3309), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4256 ( .A1(n4033), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3410) );
  NAND4_X1 U4257 ( .A1(n3413), .A2(n3412), .A3(n3411), .A4(n3410), .ZN(n3419)
         );
  AOI22_X1 U4258 ( .A1(n4046), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4259 ( .A1(n3264), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4260 ( .A1(n4052), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4261 ( .A1(n4047), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3414) );
  NAND4_X1 U4262 ( .A1(n3417), .A2(n3416), .A3(n3415), .A4(n3414), .ZN(n3418)
         );
  NAND2_X1 U4263 ( .A1(n3843), .A2(n4198), .ZN(n3420) );
  XNOR2_X1 U4264 ( .A(n3426), .B(n3427), .ZN(n4187) );
  NAND2_X1 U4265 ( .A1(n4187), .A2(n3583), .ZN(n3425) );
  INV_X1 U4266 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4773) );
  XNOR2_X1 U4267 ( .A(n3441), .B(n4773), .ZN(n4898) );
  OAI22_X1 U4268 ( .A1(n4898), .A2(n3338), .B1(n3422), .B2(n4773), .ZN(n3423)
         );
  AOI21_X1 U4269 ( .B1(n4076), .B2(EAX_REG_5__SCAN_IN), .A(n3423), .ZN(n3424)
         );
  NAND2_X1 U4270 ( .A1(n3425), .A2(n3424), .ZN(n4561) );
  INV_X1 U4271 ( .A(n3426), .ZN(n3428) );
  NAND2_X1 U4272 ( .A1(n3428), .A2(n3427), .ZN(n3447) );
  INV_X1 U4273 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4274 ( .A1(n4046), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4275 ( .A1(n4052), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4276 ( .A1(n3273), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4277 ( .A1(n3145), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3429) );
  NAND4_X1 U4278 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3438)
         );
  AOI22_X1 U4279 ( .A1(n3309), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4280 ( .A1(n4053), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4281 ( .A1(n3266), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4282 ( .A1(n4054), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3433) );
  NAND4_X1 U4283 ( .A1(n3436), .A2(n3435), .A3(n3434), .A4(n3433), .ZN(n3437)
         );
  NAND2_X1 U4284 ( .A1(n3843), .A2(n4209), .ZN(n3439) );
  NAND2_X1 U4285 ( .A1(n4196), .A2(n3583), .ZN(n3446) );
  OAI21_X1 U4286 ( .B1(n3442), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3471), 
        .ZN(n5997) );
  INV_X1 U4287 ( .A(n5997), .ZN(n3444) );
  AOI22_X1 U4288 ( .A1(n4076), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6414), .ZN(n3443) );
  MUX2_X1 U4289 ( .A(n3444), .B(n3443), .S(n3338), .Z(n3445) );
  NAND2_X1 U4290 ( .A1(n4558), .A2(n4761), .ZN(n4691) );
  INV_X1 U4291 ( .A(n4691), .ZN(n3460) );
  INV_X1 U4292 ( .A(n3447), .ZN(n3449) );
  NAND2_X1 U4293 ( .A1(n3449), .A2(n3448), .ZN(n4216) );
  INV_X1 U4294 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3451) );
  NAND2_X1 U4295 ( .A1(n3843), .A2(n4220), .ZN(n3450) );
  NAND2_X1 U4296 ( .A1(n4206), .A2(n3583), .ZN(n3459) );
  INV_X1 U4297 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3456) );
  INV_X1 U4298 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3454) );
  XNOR2_X1 U4299 ( .A(n3471), .B(n3454), .ZN(n4921) );
  AOI22_X1 U4300 ( .A1(n4921), .A2(n4072), .B1(n4075), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3455) );
  OAI21_X1 U4301 ( .B1(n4015), .B2(n3456), .A(n3455), .ZN(n3457) );
  NAND2_X1 U4302 ( .A1(n3459), .A2(n3458), .ZN(n4689) );
  NAND2_X1 U4303 ( .A1(n3460), .A2(n4689), .ZN(n4777) );
  AOI22_X1 U4304 ( .A1(n4046), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4305 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4054), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4306 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n4053), .B1(n3308), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4307 ( .A1(n3309), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3461) );
  NAND4_X1 U4308 ( .A1(n3464), .A2(n3463), .A3(n3462), .A4(n3461), .ZN(n3470)
         );
  AOI22_X1 U4309 ( .A1(n4052), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4310 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3362), .B1(n3264), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4311 ( .A1(n3363), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4312 ( .A1(n3274), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3465) );
  NAND4_X1 U4313 ( .A1(n3468), .A2(n3467), .A3(n3466), .A4(n3465), .ZN(n3469)
         );
  OAI21_X1 U4314 ( .B1(n3470), .B2(n3469), .A(n3583), .ZN(n3475) );
  NAND2_X1 U4315 ( .A1(n4076), .A2(EAX_REG_8__SCAN_IN), .ZN(n3474) );
  XNOR2_X1 U4316 ( .A(n3476), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U4317 ( .A1(n4964), .A2(n4072), .ZN(n3473) );
  NAND2_X1 U4318 ( .A1(n4075), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3472)
         );
  XNOR2_X1 U4319 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3493), .ZN(n5816) );
  INV_X1 U4320 ( .A(n5816), .ZN(n3491) );
  AOI22_X1 U4321 ( .A1(n4046), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4322 ( .A1(n3145), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4323 ( .A1(n4054), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4324 ( .A1(n3264), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3477) );
  NAND4_X1 U4325 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n3486)
         );
  AOI22_X1 U4326 ( .A1(n4045), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4327 ( .A1(n3309), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4328 ( .A1(n4053), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4329 ( .A1(n3273), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3481) );
  NAND4_X1 U4330 ( .A1(n3484), .A2(n3483), .A3(n3482), .A4(n3481), .ZN(n3485)
         );
  OAI21_X1 U4331 ( .B1(n3486), .B2(n3485), .A(n3583), .ZN(n3489) );
  NAND2_X1 U4332 ( .A1(n4076), .A2(EAX_REG_9__SCAN_IN), .ZN(n3488) );
  NAND2_X1 U4333 ( .A1(n4075), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3487)
         );
  NAND3_X1 U4334 ( .A1(n3489), .A2(n3488), .A3(n3487), .ZN(n3490) );
  AOI21_X1 U4335 ( .B1(n3491), .B2(n4072), .A(n3490), .ZN(n4820) );
  NAND2_X1 U4336 ( .A1(n3494), .A2(n6660), .ZN(n3496) );
  INV_X1 U4337 ( .A(n3535), .ZN(n3495) );
  NAND2_X1 U4338 ( .A1(n3496), .A2(n3495), .ZN(n5058) );
  NAND2_X1 U4339 ( .A1(n5058), .A2(n4072), .ZN(n3511) );
  AOI22_X1 U4340 ( .A1(n4045), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4341 ( .A1(n3309), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4342 ( .A1(n3266), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4343 ( .A1(n4054), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4344 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3506)
         );
  AOI22_X1 U4345 ( .A1(n4046), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4346 ( .A1(n3264), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4347 ( .A1(n4052), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4348 ( .A1(n3274), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3501) );
  NAND4_X1 U4349 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3505)
         );
  OAI21_X1 U4350 ( .B1(n3506), .B2(n3505), .A(n3583), .ZN(n3509) );
  NAND2_X1 U4351 ( .A1(n4076), .A2(EAX_REG_10__SCAN_IN), .ZN(n3508) );
  NAND2_X1 U4352 ( .A1(n4075), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3507)
         );
  AND3_X1 U4353 ( .A1(n3509), .A2(n3508), .A3(n3507), .ZN(n3510) );
  NAND2_X1 U4354 ( .A1(n3511), .A2(n3510), .ZN(n4925) );
  INV_X1 U4355 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5806) );
  XNOR2_X1 U4356 ( .A(n5806), .B(n3535), .ZN(n5809) );
  AOI22_X1 U4357 ( .A1(n4045), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4358 ( .A1(n4054), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4359 ( .A1(n3309), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4360 ( .A1(n4053), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3512) );
  NAND4_X1 U4361 ( .A1(n3515), .A2(n3514), .A3(n3513), .A4(n3512), .ZN(n3521)
         );
  AOI22_X1 U4362 ( .A1(n4046), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4363 ( .A1(n4052), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4364 ( .A1(n3364), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4365 ( .A1(n3266), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3516) );
  NAND4_X1 U4366 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3520)
         );
  OR2_X1 U4367 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  AOI22_X1 U4368 ( .A1(n3583), .A2(n3522), .B1(n4075), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3524) );
  NAND2_X1 U4369 ( .A1(n4076), .A2(EAX_REG_11__SCAN_IN), .ZN(n3523) );
  OAI211_X1 U4370 ( .C1(n5809), .C2(n3338), .A(n3524), .B(n3523), .ZN(n4992)
         );
  AOI22_X1 U4371 ( .A1(n4046), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4372 ( .A1(n4054), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4373 ( .A1(n4033), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4374 ( .A1(n3274), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3525) );
  NAND4_X1 U4375 ( .A1(n3528), .A2(n3527), .A3(n3526), .A4(n3525), .ZN(n3534)
         );
  AOI22_X1 U4376 ( .A1(n3273), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4377 ( .A1(n4053), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4378 ( .A1(n4052), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4379 ( .A1(n3309), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3529) );
  NAND4_X1 U4380 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(n3533)
         );
  NOR2_X1 U4381 ( .A1(n3534), .A2(n3533), .ZN(n3538) );
  XNOR2_X1 U4382 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3539), .ZN(n5102)
         );
  AOI22_X1 U4383 ( .A1(n4072), .A2(n5102), .B1(n4075), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U4384 ( .A1(n4076), .A2(EAX_REG_12__SCAN_IN), .ZN(n3536) );
  NAND2_X1 U4385 ( .A1(n4076), .A2(EAX_REG_13__SCAN_IN), .ZN(n3542) );
  OAI21_X1 U4386 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3540), .A(n3573), 
        .ZN(n5792) );
  AOI22_X1 U4387 ( .A1(n4072), .A2(n5792), .B1(n4075), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4388 ( .A1(n4046), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4389 ( .A1(n4052), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4390 ( .A1(n3309), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4391 ( .A1(n3264), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3546) );
  NAND4_X1 U4392 ( .A1(n3549), .A2(n3548), .A3(n3547), .A4(n3546), .ZN(n3555)
         );
  AOI22_X1 U4393 ( .A1(n3266), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4394 ( .A1(n4033), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4395 ( .A1(n3273), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4396 ( .A1(n3274), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3550) );
  NAND4_X1 U4397 ( .A1(n3553), .A2(n3552), .A3(n3551), .A4(n3550), .ZN(n3554)
         );
  OR2_X1 U4398 ( .A1(n3555), .A2(n3554), .ZN(n3556) );
  AND2_X1 U4399 ( .A1(n3583), .A2(n3556), .ZN(n5064) );
  NAND2_X1 U4400 ( .A1(n5063), .A2(n5064), .ZN(n5068) );
  AOI22_X1 U4401 ( .A1(n4052), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4402 ( .A1(n3264), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4403 ( .A1(n3273), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4404 ( .A1(n4054), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4405 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3567)
         );
  AOI22_X1 U4406 ( .A1(n4046), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4407 ( .A1(n3309), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4408 ( .A1(n3274), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4409 ( .A1(n3362), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3562) );
  NAND4_X1 U4410 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3566)
         );
  NOR2_X1 U4411 ( .A1(n3567), .A2(n3566), .ZN(n3571) );
  XNOR2_X1 U4412 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3573), .ZN(n5780)
         );
  INV_X1 U4413 ( .A(n5780), .ZN(n3568) );
  AOI22_X1 U4414 ( .A1(n4072), .A2(n3568), .B1(n4075), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3570) );
  NAND2_X1 U4415 ( .A1(n4076), .A2(EAX_REG_14__SCAN_IN), .ZN(n3569) );
  OAI211_X1 U4416 ( .C1(n3572), .C2(n3571), .A(n3570), .B(n3569), .ZN(n5079)
         );
  XNOR2_X1 U4417 ( .A(n3590), .B(n5238), .ZN(n5452) );
  AOI22_X1 U4418 ( .A1(n3264), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4419 ( .A1(n4045), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4420 ( .A1(n3266), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4421 ( .A1(n4054), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3575) );
  NAND4_X1 U4422 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(n3585)
         );
  AOI22_X1 U4423 ( .A1(n4046), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4424 ( .A1(n4052), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4425 ( .A1(n3309), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4426 ( .A1(n3274), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4427 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3584)
         );
  OAI21_X1 U4428 ( .B1(n3585), .B2(n3584), .A(n3583), .ZN(n3588) );
  NAND2_X1 U4429 ( .A1(n4076), .A2(EAX_REG_15__SCAN_IN), .ZN(n3587) );
  NAND2_X1 U4430 ( .A1(n4075), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3586)
         );
  NAND3_X1 U4431 ( .A1(n3588), .A2(n3587), .A3(n3586), .ZN(n3589) );
  AOI21_X1 U4432 ( .B1(n5452), .B2(n4072), .A(n3589), .ZN(n5237) );
  INV_X1 U4433 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5238) );
  XOR2_X1 U4434 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3605), .Z(n5771) );
  INV_X1 U4435 ( .A(n5771), .ZN(n5444) );
  NAND2_X1 U4436 ( .A1(n4479), .A2(n4491), .ZN(n3591) );
  AOI22_X1 U4437 ( .A1(n3273), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4438 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3309), .B1(n3308), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4439 ( .A1(n4052), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4440 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3362), .B1(n4047), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3592) );
  NAND4_X1 U4441 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3601)
         );
  AOI22_X1 U4442 ( .A1(n4046), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4443 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n4053), .B1(n3316), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4444 ( .A1(n4033), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4445 ( .A1(n4054), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4446 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3600)
         );
  NOR2_X1 U4447 ( .A1(n3601), .A2(n3600), .ZN(n3603) );
  AOI22_X1 U4448 ( .A1(n4076), .A2(EAX_REG_16__SCAN_IN), .B1(n4075), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3602) );
  OAI21_X1 U4449 ( .B1(n4069), .B2(n3603), .A(n3602), .ZN(n3604) );
  AOI21_X1 U4450 ( .B1(n5444), .B2(n4072), .A(n3604), .ZN(n5288) );
  XNOR2_X1 U4451 ( .A(n3619), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5437)
         );
  INV_X1 U4452 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5435) );
  AOI21_X1 U4453 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5435), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3606) );
  AOI21_X1 U4454 ( .B1(n4076), .B2(EAX_REG_17__SCAN_IN), .A(n3606), .ZN(n3618)
         );
  AOI22_X1 U4455 ( .A1(n4045), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4456 ( .A1(n4054), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4457 ( .A1(n4053), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4458 ( .A1(n3274), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3607) );
  NAND4_X1 U4459 ( .A1(n3610), .A2(n3609), .A3(n3608), .A4(n3607), .ZN(n3616)
         );
  AOI22_X1 U4460 ( .A1(n4046), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4461 ( .A1(n3309), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4462 ( .A1(n3273), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4463 ( .A1(n4047), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3611) );
  NAND4_X1 U4464 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(n3615)
         );
  OAI21_X1 U4465 ( .B1(n3616), .B2(n3615), .A(n4042), .ZN(n3617) );
  AOI22_X1 U4466 ( .A1(n5437), .A2(n4072), .B1(n3618), .B2(n3617), .ZN(n5224)
         );
  NAND2_X1 U4467 ( .A1(n5221), .A2(n5224), .ZN(n5222) );
  NOR2_X1 U4468 ( .A1(n3620), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3621)
         );
  OR2_X1 U4469 ( .A1(n3654), .A2(n3621), .ZN(n5757) );
  AOI22_X1 U4470 ( .A1(n4045), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4471 ( .A1(n4054), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4472 ( .A1(n3309), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4473 ( .A1(n3274), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3622) );
  NAND4_X1 U4474 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3631)
         );
  AOI22_X1 U4475 ( .A1(n4046), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4476 ( .A1(n3273), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4477 ( .A1(n3266), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4478 ( .A1(n3308), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3626) );
  NAND4_X1 U4479 ( .A1(n3629), .A2(n3628), .A3(n3627), .A4(n3626), .ZN(n3630)
         );
  NOR2_X1 U4480 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  NOR2_X1 U4481 ( .A1(n4069), .A2(n3632), .ZN(n3636) );
  INV_X1 U4482 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3634) );
  NAND2_X1 U4483 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3633)
         );
  OAI211_X1 U4484 ( .C1(n4015), .C2(n3634), .A(n3338), .B(n3633), .ZN(n3635)
         );
  OAI22_X1 U4485 ( .A1(n5757), .A2(n3338), .B1(n3636), .B2(n3635), .ZN(n5279)
         );
  INV_X1 U4486 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3637) );
  XNOR2_X1 U4487 ( .A(n3654), .B(n3637), .ZN(n5660) );
  NAND2_X1 U4488 ( .A1(n5660), .A2(n4072), .ZN(n3653) );
  AOI22_X1 U4489 ( .A1(n4045), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4490 ( .A1(n3266), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4491 ( .A1(n3309), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4492 ( .A1(n3273), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4493 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3647)
         );
  AOI22_X1 U4494 ( .A1(n4046), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4495 ( .A1(n3274), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4496 ( .A1(n4054), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4497 ( .A1(n3308), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3642) );
  NAND4_X1 U4498 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3646)
         );
  NOR2_X1 U4499 ( .A1(n3647), .A2(n3646), .ZN(n3651) );
  NAND2_X1 U4500 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3648)
         );
  NAND2_X1 U4501 ( .A1(n3338), .A2(n3648), .ZN(n3649) );
  AOI21_X1 U4502 ( .B1(n4076), .B2(EAX_REG_19__SCAN_IN), .A(n3649), .ZN(n3650)
         );
  OAI21_X1 U4503 ( .B1(n4069), .B2(n3651), .A(n3650), .ZN(n3652) );
  NAND2_X1 U4504 ( .A1(n3653), .A2(n3652), .ZN(n5269) );
  OR2_X1 U4505 ( .A1(n3655), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3656)
         );
  NAND2_X1 U4506 ( .A1(n3656), .A2(n3703), .ZN(n5409) );
  INV_X1 U4507 ( .A(n5409), .ZN(n3672) );
  AOI22_X1 U4508 ( .A1(n4046), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4509 ( .A1(n4052), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4510 ( .A1(n4054), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4511 ( .A1(n3274), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3657) );
  NAND4_X1 U4512 ( .A1(n3660), .A2(n3659), .A3(n3658), .A4(n3657), .ZN(n3666)
         );
  AOI22_X1 U4513 ( .A1(n3309), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4514 ( .A1(n4045), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4515 ( .A1(n3266), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4516 ( .A1(n3316), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3661) );
  NAND4_X1 U4517 ( .A1(n3664), .A2(n3663), .A3(n3662), .A4(n3661), .ZN(n3665)
         );
  OR2_X1 U4518 ( .A1(n3666), .A2(n3665), .ZN(n3670) );
  INV_X1 U4519 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3668) );
  NAND2_X1 U4520 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3667)
         );
  OAI211_X1 U4521 ( .C1(n4015), .C2(n3668), .A(n3338), .B(n3667), .ZN(n3669)
         );
  AOI21_X1 U4522 ( .B1(n4042), .B2(n3670), .A(n3669), .ZN(n3671) );
  AOI21_X1 U4523 ( .B1(n3672), .B2(n4072), .A(n3671), .ZN(n5210) );
  AOI22_X1 U4524 ( .A1(n4046), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4525 ( .A1(n4052), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4526 ( .A1(n3310), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4527 ( .A1(n3274), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3673) );
  NAND4_X1 U4528 ( .A1(n3676), .A2(n3675), .A3(n3674), .A4(n3673), .ZN(n3682)
         );
  AOI22_X1 U4529 ( .A1(n3256), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4530 ( .A1(n4053), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4531 ( .A1(n3266), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4532 ( .A1(n4054), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3677) );
  NAND4_X1 U4533 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(n3681)
         );
  NOR2_X1 U4534 ( .A1(n3682), .A2(n3681), .ZN(n3686) );
  INV_X1 U4535 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3683) );
  AOI21_X1 U4536 ( .B1(n3683), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3684) );
  AOI21_X1 U4537 ( .B1(n3337), .B2(EAX_REG_21__SCAN_IN), .A(n3684), .ZN(n3685)
         );
  OAI21_X1 U4538 ( .B1(n4069), .B2(n3686), .A(n3685), .ZN(n3688) );
  XNOR2_X1 U4539 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3703), .ZN(n5655)
         );
  NAND2_X1 U4540 ( .A1(n4072), .A2(n5655), .ZN(n3687) );
  AOI22_X1 U4541 ( .A1(n4046), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4542 ( .A1(n3310), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4543 ( .A1(n4054), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4544 ( .A1(n3256), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3689) );
  NAND4_X1 U4545 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3698)
         );
  AOI22_X1 U4546 ( .A1(n4045), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4547 ( .A1(n3264), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4548 ( .A1(n3363), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4549 ( .A1(n4047), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3693) );
  NAND4_X1 U4550 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3697)
         );
  NOR2_X1 U4551 ( .A1(n3698), .A2(n3697), .ZN(n3702) );
  NAND2_X1 U4552 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3699)
         );
  NAND2_X1 U4553 ( .A1(n3338), .A2(n3699), .ZN(n3700) );
  AOI21_X1 U4554 ( .B1(n3337), .B2(EAX_REG_22__SCAN_IN), .A(n3700), .ZN(n3701)
         );
  OAI21_X1 U4555 ( .B1(n4069), .B2(n3702), .A(n3701), .ZN(n3707) );
  OAI21_X1 U4556 ( .B1(n3705), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3748), 
        .ZN(n5644) );
  OR2_X1 U4557 ( .A1(n5644), .A2(n3338), .ZN(n3706) );
  NAND2_X1 U4558 ( .A1(n3707), .A2(n3706), .ZN(n5263) );
  AOI22_X1 U4559 ( .A1(n4046), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4560 ( .A1(n4054), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4561 ( .A1(n4033), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4562 ( .A1(n4053), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3709) );
  NAND4_X1 U4563 ( .A1(n3712), .A2(n3711), .A3(n3710), .A4(n3709), .ZN(n3718)
         );
  AOI22_X1 U4564 ( .A1(n3362), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4565 ( .A1(n3309), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4566 ( .A1(n4052), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4567 ( .A1(n3273), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3713) );
  NAND4_X1 U4568 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3717)
         );
  NOR2_X1 U4569 ( .A1(n3718), .A2(n3717), .ZN(n3736) );
  AOI22_X1 U4570 ( .A1(n4046), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4571 ( .A1(n4052), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4572 ( .A1(n3273), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4573 ( .A1(n3274), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4574 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3728)
         );
  AOI22_X1 U4575 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3309), .B1(n3264), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4576 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3308), .B1(n4053), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4577 ( .A1(n3266), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4578 ( .A1(n4054), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3723) );
  NAND4_X1 U4579 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3727)
         );
  NOR2_X1 U4580 ( .A1(n3728), .A2(n3727), .ZN(n3737) );
  XOR2_X1 U4581 ( .A(n3736), .B(n3737), .Z(n3729) );
  NAND2_X1 U4582 ( .A1(n3729), .A2(n4042), .ZN(n3733) );
  NAND2_X1 U4583 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3730)
         );
  NAND2_X1 U4584 ( .A1(n3338), .A2(n3730), .ZN(n3731) );
  AOI21_X1 U4585 ( .B1(n3337), .B2(EAX_REG_23__SCAN_IN), .A(n3731), .ZN(n3732)
         );
  NAND2_X1 U4586 ( .A1(n3733), .A2(n3732), .ZN(n3735) );
  XNOR2_X1 U4587 ( .A(n3748), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5635)
         );
  NAND2_X1 U4588 ( .A1(n5635), .A2(n4072), .ZN(n3734) );
  NAND2_X1 U4589 ( .A1(n3735), .A2(n3734), .ZN(n5254) );
  OR2_X1 U4590 ( .A1(n3737), .A2(n3736), .ZN(n3756) );
  AOI22_X1 U4591 ( .A1(n3316), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4592 ( .A1(n4046), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3740) );
  INV_X1 U4593 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6686) );
  AOI22_X1 U4594 ( .A1(n3273), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4595 ( .A1(n3309), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3738) );
  NAND4_X1 U4596 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3747)
         );
  AOI22_X1 U4597 ( .A1(n4052), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4598 ( .A1(n4054), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4599 ( .A1(n3364), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4600 ( .A1(n4033), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3742) );
  NAND4_X1 U4601 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3746)
         );
  NOR2_X1 U4602 ( .A1(n3747), .A2(n3746), .ZN(n3755) );
  XNOR2_X1 U4603 ( .A(n3756), .B(n3755), .ZN(n3754) );
  INV_X1 U4604 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5643) );
  INV_X1 U4605 ( .A(n3749), .ZN(n3750) );
  INV_X1 U4606 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U4607 ( .A1(n3750), .A2(n5202), .ZN(n3751) );
  NAND2_X1 U4608 ( .A1(n3790), .A2(n3751), .ZN(n5379) );
  AOI22_X1 U4609 ( .A1(n5379), .A2(n4072), .B1(n4075), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3753) );
  NAND2_X1 U4610 ( .A1(n3337), .A2(EAX_REG_24__SCAN_IN), .ZN(n3752) );
  OAI211_X1 U4611 ( .C1(n3754), .C2(n4069), .A(n3753), .B(n3752), .ZN(n5198)
         );
  OR2_X1 U4612 ( .A1(n3756), .A2(n3755), .ZN(n3773) );
  AOI22_X1 U4613 ( .A1(n4053), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4614 ( .A1(n4046), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4615 ( .A1(n3274), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4616 ( .A1(n4047), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3757) );
  NAND4_X1 U4617 ( .A1(n3760), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3766)
         );
  AOI22_X1 U4618 ( .A1(n4045), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4619 ( .A1(n4052), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4620 ( .A1(n4054), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4621 ( .A1(n3256), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3761) );
  NAND4_X1 U4622 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3765)
         );
  NOR2_X1 U4623 ( .A1(n3766), .A2(n3765), .ZN(n3774) );
  XOR2_X1 U4624 ( .A(n3773), .B(n3774), .Z(n3767) );
  NAND2_X1 U4625 ( .A1(n3767), .A2(n4042), .ZN(n3772) );
  NAND2_X1 U4626 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3768)
         );
  NAND2_X1 U4627 ( .A1(n3338), .A2(n3768), .ZN(n3769) );
  AOI21_X1 U4628 ( .B1(n3337), .B2(EAX_REG_25__SCAN_IN), .A(n3769), .ZN(n3771)
         );
  XNOR2_X1 U4629 ( .A(n3790), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5368)
         );
  AOI21_X1 U4630 ( .B1(n3772), .B2(n3771), .A(n3770), .ZN(n5188) );
  NAND2_X1 U4631 ( .A1(n5187), .A2(n5188), .ZN(n5175) );
  NOR2_X1 U4632 ( .A1(n3774), .A2(n3773), .ZN(n3798) );
  AOI22_X1 U4633 ( .A1(n4046), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4634 ( .A1(n4052), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4635 ( .A1(n3310), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4636 ( .A1(n3274), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4637 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3784)
         );
  AOI22_X1 U4638 ( .A1(n3256), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4639 ( .A1(n4053), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4640 ( .A1(n3266), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4641 ( .A1(n4054), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3779) );
  NAND4_X1 U4642 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3783)
         );
  OR2_X1 U4643 ( .A1(n3784), .A2(n3783), .ZN(n3797) );
  INV_X1 U4644 ( .A(n3797), .ZN(n3785) );
  XNOR2_X1 U4645 ( .A(n3798), .B(n3785), .ZN(n3789) );
  INV_X1 U4646 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3787) );
  NAND2_X1 U4647 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3786)
         );
  OAI211_X1 U4648 ( .C1(n4015), .C2(n3787), .A(n3338), .B(n3786), .ZN(n3788)
         );
  AOI21_X1 U4649 ( .B1(n3789), .B2(n4042), .A(n3788), .ZN(n3796) );
  INV_X1 U4650 ( .A(n3790), .ZN(n3791) );
  INV_X1 U4651 ( .A(n3792), .ZN(n3793) );
  INV_X1 U4652 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U4653 ( .A1(n3793), .A2(n5179), .ZN(n3794) );
  NAND2_X1 U4654 ( .A1(n4018), .A2(n3794), .ZN(n5357) );
  NOR2_X1 U4655 ( .A1(n5357), .A2(n3338), .ZN(n3795) );
  NAND2_X1 U4656 ( .A1(n3798), .A2(n3797), .ZN(n4000) );
  AOI22_X1 U4657 ( .A1(n4046), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4658 ( .A1(n3310), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4659 ( .A1(n3264), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4660 ( .A1(n4054), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3799) );
  NAND4_X1 U4661 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n3808)
         );
  AOI22_X1 U4662 ( .A1(n4045), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4663 ( .A1(n3256), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4664 ( .A1(n3363), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4665 ( .A1(n3362), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4666 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3807)
         );
  NOR2_X1 U4667 ( .A1(n3808), .A2(n3807), .ZN(n4001) );
  XOR2_X1 U4668 ( .A(n4000), .B(n4001), .Z(n3809) );
  NAND2_X1 U4669 ( .A1(n3809), .A2(n4042), .ZN(n3813) );
  NAND2_X1 U4670 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3810)
         );
  NAND2_X1 U4671 ( .A1(n3338), .A2(n3810), .ZN(n3811) );
  AOI21_X1 U4672 ( .B1(n3337), .B2(EAX_REG_27__SCAN_IN), .A(n3811), .ZN(n3812)
         );
  NAND2_X1 U4673 ( .A1(n3813), .A2(n3812), .ZN(n3815) );
  XNOR2_X1 U4674 ( .A(n4018), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5349)
         );
  NAND2_X1 U4675 ( .A1(n5349), .A2(n4072), .ZN(n3814) );
  NAND2_X1 U4676 ( .A1(n3815), .A2(n3814), .ZN(n3818) );
  NAND2_X1 U4677 ( .A1(n3843), .A2(n4487), .ZN(n3820) );
  NAND2_X1 U4678 ( .A1(n3820), .A2(n4479), .ZN(n3835) );
  XNOR2_X1 U4679 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3839) );
  NAND2_X1 U4680 ( .A1(n4660), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3838) );
  XNOR2_X1 U4681 ( .A(n3839), .B(n3838), .ZN(n4081) );
  AND2_X1 U4682 ( .A1(n4081), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3831) );
  INV_X1 U4683 ( .A(n3843), .ZN(n3869) );
  NAND2_X1 U4684 ( .A1(n3041), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3821) );
  NAND2_X1 U4685 ( .A1(n3838), .A2(n3821), .ZN(n3822) );
  OAI21_X1 U4686 ( .B1(n3869), .B2(n3822), .A(n3874), .ZN(n3830) );
  INV_X1 U4687 ( .A(n3822), .ZN(n3825) );
  INV_X1 U4688 ( .A(n3823), .ZN(n3824) );
  AOI21_X1 U4689 ( .B1(n4141), .B2(n3825), .A(n3824), .ZN(n3828) );
  INV_X1 U4690 ( .A(n4890), .ZN(n4267) );
  NAND2_X1 U4691 ( .A1(n3826), .A2(n4479), .ZN(n3827) );
  NAND2_X1 U4692 ( .A1(n4267), .A2(n3827), .ZN(n3844) );
  OR2_X1 U4693 ( .A1(n3828), .A2(n3844), .ZN(n3829) );
  OAI211_X1 U4694 ( .C1(n3835), .C2(n3831), .A(n3830), .B(n3829), .ZN(n3837)
         );
  INV_X1 U4695 ( .A(n4081), .ZN(n3834) );
  INV_X1 U4696 ( .A(n3831), .ZN(n3832) );
  NAND2_X1 U4697 ( .A1(n3874), .A2(n3832), .ZN(n3833) );
  OAI21_X1 U4698 ( .B1(n3835), .B2(n3834), .A(n3833), .ZN(n3836) );
  NAND2_X1 U4699 ( .A1(n3837), .A2(n3836), .ZN(n3849) );
  INV_X1 U4700 ( .A(n3838), .ZN(n3840) );
  NAND2_X1 U4701 ( .A1(n3840), .A2(n3839), .ZN(n3842) );
  NAND2_X1 U4702 ( .A1(n6387), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U4703 ( .A1(n3842), .A2(n3841), .ZN(n3852) );
  XNOR2_X1 U4704 ( .A(n4330), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3850)
         );
  XNOR2_X1 U4705 ( .A(n3852), .B(n3850), .ZN(n4082) );
  OAI211_X1 U4706 ( .C1(n3849), .C2(n3844), .A(n4082), .B(n3843), .ZN(n3864)
         );
  INV_X1 U4707 ( .A(n3844), .ZN(n3847) );
  INV_X1 U4708 ( .A(n4082), .ZN(n3845) );
  NAND2_X1 U4709 ( .A1(n3246), .A2(n3845), .ZN(n3846) );
  NAND2_X1 U4710 ( .A1(n3847), .A2(n3846), .ZN(n3848) );
  NAND2_X1 U4711 ( .A1(n3849), .A2(n3848), .ZN(n3863) );
  INV_X1 U4712 ( .A(n3850), .ZN(n3851) );
  NAND2_X1 U4713 ( .A1(n3852), .A2(n3851), .ZN(n3854) );
  NAND2_X1 U4714 ( .A1(n6391), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3853) );
  NAND2_X1 U4715 ( .A1(n3854), .A2(n3853), .ZN(n3859) );
  XNOR2_X1 U4716 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3857) );
  NAND2_X1 U4717 ( .A1(n3859), .A2(n3857), .ZN(n3856) );
  NAND2_X1 U4718 ( .A1(n4985), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3855) );
  NAND2_X1 U4719 ( .A1(n3856), .A2(n3855), .ZN(n3866) );
  INV_X1 U4720 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6398) );
  INV_X1 U4721 ( .A(n3857), .ZN(n3858) );
  XNOR2_X1 U4722 ( .A(n3859), .B(n3858), .ZN(n3860) );
  NOR2_X1 U4723 ( .A1(n3246), .A2(n4084), .ZN(n3862) );
  AOI21_X1 U4724 ( .B1(n3864), .B2(n3863), .A(n3862), .ZN(n3873) );
  AND2_X1 U4725 ( .A1(n6398), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3865)
         );
  INV_X1 U4726 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U4727 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5730), .ZN(n3867) );
  NAND2_X1 U4728 ( .A1(n3868), .A2(n3867), .ZN(n4085) );
  NOR2_X1 U4729 ( .A1(n3869), .A2(n4085), .ZN(n3870) );
  AOI21_X1 U4730 ( .B1(n6423), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n3870), 
        .ZN(n3871) );
  OAI21_X1 U4731 ( .B1(n3874), .B2(n4084), .A(n3871), .ZN(n3872) );
  OAI22_X1 U4732 ( .A1(n3878), .A2(n5274), .B1(n3183), .B2(n3879), .ZN(n3880)
         );
  INV_X1 U4733 ( .A(n3880), .ZN(n3888) );
  NAND3_X1 U4734 ( .A1(n3208), .A2(n3187), .A3(n4337), .ZN(n3883) );
  INV_X1 U4735 ( .A(n4337), .ZN(n3881) );
  NAND2_X1 U4736 ( .A1(n3881), .A2(n4283), .ZN(n3882) );
  AND2_X1 U4737 ( .A1(n3883), .A2(n3882), .ZN(n4297) );
  NAND2_X1 U4738 ( .A1(n4332), .A2(n4487), .ZN(n4951) );
  NOR2_X1 U4739 ( .A1(n4951), .A2(n4497), .ZN(n4306) );
  INV_X1 U4740 ( .A(n4469), .ZN(n3884) );
  OAI21_X1 U4741 ( .B1(n4306), .B2(n4104), .A(n4152), .ZN(n3885) );
  AND2_X1 U4742 ( .A1(n4297), .A2(n3885), .ZN(n3886) );
  NAND4_X1 U4743 ( .A1(n3877), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n4318)
         );
  AND2_X1 U4744 ( .A1(n3895), .A2(n4332), .ZN(n3890) );
  NAND2_X1 U4745 ( .A1(n6380), .A2(n3890), .ZN(n4424) );
  OAI21_X1 U4746 ( .B1(n3889), .B2(n3891), .A(n4424), .ZN(n3892) );
  NOR2_X1 U4747 ( .A1(n4318), .A2(n3892), .ZN(n4380) );
  NOR2_X1 U4748 ( .A1(n4126), .A2(n4348), .ZN(n3893) );
  NAND2_X1 U4749 ( .A1(n4380), .A2(n3893), .ZN(n4321) );
  OR2_X1 U4750 ( .A1(n6415), .A2(n4321), .ZN(n4309) );
  INV_X1 U4751 ( .A(n2954), .ZN(n3896) );
  INV_X1 U4752 ( .A(n3894), .ZN(n4137) );
  NAND4_X1 U4753 ( .A1(n3896), .A2(n4372), .A3(n4137), .A4(n3895), .ZN(n4131)
         );
  OR2_X1 U4754 ( .A1(n4131), .A2(n4348), .ZN(n3897) );
  NAND2_X1 U4755 ( .A1(n4309), .A2(n3897), .ZN(n3899) );
  AND2_X2 U4756 ( .A1(n3899), .A2(n6420), .ZN(n5878) );
  NAND2_X1 U4757 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4348), .ZN(n3901)
         );
  NAND2_X1 U4758 ( .A1(n3976), .A2(EBX_REG_0__SCAN_IN), .ZN(n3903) );
  INV_X1 U4759 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4401) );
  NAND2_X1 U4760 ( .A1(n5274), .A2(n4401), .ZN(n3902) );
  NAND2_X1 U4761 ( .A1(n3903), .A2(n3902), .ZN(n4376) );
  XNOR2_X1 U4762 ( .A(n3904), .B(n4376), .ZN(n4347) );
  NAND2_X1 U4763 ( .A1(n4347), .A2(n4134), .ZN(n4350) );
  NAND2_X1 U4764 ( .A1(n4350), .A2(n3904), .ZN(n4414) );
  OR2_X1 U4765 ( .A1(n5272), .A2(EBX_REG_2__SCAN_IN), .ZN(n3909) );
  INV_X1 U4766 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U4767 ( .A1(n3976), .A2(n6106), .ZN(n3907) );
  INV_X1 U4768 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U4769 ( .A1(n4134), .A2(n5857), .ZN(n3906) );
  NAND3_X1 U4770 ( .A1(n3907), .A2(n5274), .A3(n3906), .ZN(n3908) );
  MUX2_X1 U4771 ( .A(n3979), .B(n5274), .S(EBX_REG_3__SCAN_IN), .Z(n3910) );
  OAI21_X1 U4772 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4104), .A(n3910), 
        .ZN(n4453) );
  MUX2_X1 U4773 ( .A(n5272), .B(n3976), .S(EBX_REG_4__SCAN_IN), .Z(n3913) );
  NAND2_X1 U4774 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n4348), .ZN(n3911)
         );
  AND2_X1 U4775 ( .A1(n3972), .A2(n3911), .ZN(n3912) );
  NAND2_X1 U4776 ( .A1(n3913), .A2(n3912), .ZN(n4566) );
  INV_X1 U4777 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U4778 ( .A1(n4134), .A2(n4894), .ZN(n3915) );
  NAND2_X1 U4779 ( .A1(n5274), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3914)
         );
  NAND3_X1 U4780 ( .A1(n3915), .A2(n3976), .A3(n3914), .ZN(n3916) );
  OAI21_X1 U4781 ( .B1(n3979), .B2(EBX_REG_5__SCAN_IN), .A(n3916), .ZN(n4563)
         );
  OR2_X1 U4782 ( .A1(n5272), .A2(EBX_REG_6__SCAN_IN), .ZN(n3920) );
  INV_X1 U4783 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U4784 ( .A1(n3976), .A2(n5090), .ZN(n3918) );
  INV_X1 U4785 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U4786 ( .A1(n4134), .A2(n5834), .ZN(n3917) );
  NAND3_X1 U4787 ( .A1(n3918), .A2(n5274), .A3(n3917), .ZN(n3919) );
  INV_X1 U4788 ( .A(n3979), .ZN(n3986) );
  INV_X1 U4789 ( .A(EBX_REG_7__SCAN_IN), .ZN(n3921) );
  NAND2_X1 U4790 ( .A1(n3986), .A2(n3921), .ZN(n3925) );
  NAND2_X1 U4791 ( .A1(n4134), .A2(n3921), .ZN(n3923) );
  NAND2_X1 U4792 ( .A1(n5274), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3922)
         );
  NAND3_X1 U4793 ( .A1(n3923), .A2(n3976), .A3(n3922), .ZN(n3924) );
  MUX2_X1 U4794 ( .A(n3979), .B(n5274), .S(EBX_REG_9__SCAN_IN), .Z(n3926) );
  OAI21_X1 U4795 ( .B1(n4104), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n3926), 
        .ZN(n5823) );
  OR2_X1 U4796 ( .A1(n5272), .A2(EBX_REG_8__SCAN_IN), .ZN(n3931) );
  INV_X1 U4797 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4223) );
  NAND2_X1 U4798 ( .A1(n3976), .A2(n4223), .ZN(n3929) );
  INV_X1 U4799 ( .A(EBX_REG_8__SCAN_IN), .ZN(n3927) );
  NAND2_X1 U4800 ( .A1(n4134), .A2(n3927), .ZN(n3928) );
  NAND3_X1 U4801 ( .A1(n3929), .A2(n5274), .A3(n3928), .ZN(n3930) );
  NOR2_X1 U4802 ( .A1(n5823), .A2(n5817), .ZN(n3932) );
  MUX2_X1 U4803 ( .A(n5272), .B(n3976), .S(EBX_REG_10__SCAN_IN), .Z(n3934) );
  NAND2_X1 U4804 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4348), .ZN(n3933) );
  INV_X1 U4805 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U4806 ( .A1(n4134), .A2(n5875), .ZN(n3936) );
  NAND2_X1 U4807 ( .A1(n5274), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3935) );
  NAND3_X1 U4808 ( .A1(n3936), .A2(n3976), .A3(n3935), .ZN(n3937) );
  OAI21_X1 U4809 ( .B1(n3979), .B2(EBX_REG_11__SCAN_IN), .A(n3937), .ZN(n5799)
         );
  NOR2_X2 U4810 ( .A1(n5800), .A2(n5799), .ZN(n5802) );
  MUX2_X1 U4811 ( .A(n5272), .B(n3976), .S(EBX_REG_12__SCAN_IN), .Z(n3940) );
  NAND2_X1 U4812 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4348), .ZN(n3938) );
  AND2_X1 U4813 ( .A1(n3972), .A2(n3938), .ZN(n3939) );
  NAND2_X1 U4814 ( .A1(n3940), .A2(n3939), .ZN(n5040) );
  INV_X1 U4815 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U4816 ( .A1(n4134), .A2(n5798), .ZN(n3942) );
  NAND2_X1 U4817 ( .A1(n5274), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3941) );
  NAND3_X1 U4818 ( .A1(n3942), .A2(n3976), .A3(n3941), .ZN(n3943) );
  OAI21_X1 U4819 ( .B1(n3979), .B2(EBX_REG_13__SCAN_IN), .A(n3943), .ZN(n5069)
         );
  MUX2_X1 U4820 ( .A(n5272), .B(n3976), .S(EBX_REG_14__SCAN_IN), .Z(n3945) );
  NAND2_X1 U4821 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4348), .ZN(n3944) );
  AND3_X1 U4822 ( .A1(n3945), .A2(n3972), .A3(n3944), .ZN(n5081) );
  INV_X1 U4823 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U4824 ( .A1(n4134), .A2(n5297), .ZN(n3947) );
  NAND2_X1 U4825 ( .A1(n5274), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3946) );
  NAND3_X1 U4826 ( .A1(n3947), .A2(n3976), .A3(n3946), .ZN(n3948) );
  OAI21_X1 U4827 ( .B1(n3979), .B2(EBX_REG_15__SCAN_IN), .A(n3948), .ZN(n5241)
         );
  OR2_X1 U4828 ( .A1(n5272), .A2(EBX_REG_16__SCAN_IN), .ZN(n3952) );
  INV_X1 U4829 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U4830 ( .A1(n3976), .A2(n6595), .ZN(n3950) );
  INV_X1 U4831 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U4832 ( .A1(n4134), .A2(n5294), .ZN(n3949) );
  NAND3_X1 U4833 ( .A1(n3950), .A2(n5274), .A3(n3949), .ZN(n3951) );
  NAND2_X1 U4834 ( .A1(n3952), .A2(n3951), .ZN(n5290) );
  MUX2_X1 U4835 ( .A(n3979), .B(n5274), .S(EBX_REG_17__SCAN_IN), .Z(n3953) );
  OAI21_X1 U4836 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n4104), .A(n3953), 
        .ZN(n5226) );
  MUX2_X1 U4837 ( .A(n5272), .B(n3976), .S(EBX_REG_19__SCAN_IN), .Z(n3955) );
  NAND2_X1 U4838 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n4348), .ZN(n3954) );
  AND3_X1 U4839 ( .A1(n3955), .A2(n3972), .A3(n3954), .ZN(n5276) );
  OR2_X1 U4840 ( .A1(n4104), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3958)
         );
  INV_X1 U4841 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3956) );
  NAND2_X1 U4842 ( .A1(n4134), .A2(n3956), .ZN(n3957) );
  AND2_X1 U4843 ( .A1(n3958), .A2(n3957), .ZN(n5214) );
  OR2_X1 U4844 ( .A1(n4104), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3960)
         );
  INV_X1 U4845 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U4846 ( .A1(n4134), .A2(n5284), .ZN(n3959) );
  NAND2_X1 U4847 ( .A1(n3960), .A2(n3959), .ZN(n5271) );
  NAND2_X1 U4848 ( .A1(n5128), .A2(EBX_REG_20__SCAN_IN), .ZN(n3962) );
  NAND2_X1 U4849 ( .A1(n5271), .A2(n5274), .ZN(n3961) );
  OAI211_X1 U4850 ( .C1(n5214), .C2(n5271), .A(n3962), .B(n3961), .ZN(n3963)
         );
  INV_X1 U4851 ( .A(n3963), .ZN(n3964) );
  INV_X1 U4852 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U4853 ( .A1(n3986), .A2(n6644), .ZN(n3968) );
  NAND2_X1 U4854 ( .A1(n4134), .A2(n6644), .ZN(n3966) );
  NAND2_X1 U4855 ( .A1(n5274), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3965) );
  NAND3_X1 U4856 ( .A1(n3966), .A2(n3976), .A3(n3965), .ZN(n3967) );
  AND2_X1 U4857 ( .A1(n3968), .A2(n3967), .ZN(n5570) );
  MUX2_X1 U4858 ( .A(n3979), .B(n5274), .S(EBX_REG_23__SCAN_IN), .Z(n3969) );
  OAI21_X1 U4859 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n4104), .A(n3969), 
        .ZN(n3970) );
  INV_X1 U4860 ( .A(n3970), .ZN(n5255) );
  MUX2_X1 U4861 ( .A(n5272), .B(n3976), .S(EBX_REG_22__SCAN_IN), .Z(n3974) );
  NAND2_X1 U4862 ( .A1(n4348), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3971) );
  AND2_X1 U4863 ( .A1(n3972), .A2(n3971), .ZN(n3973) );
  NAND2_X1 U4864 ( .A1(n3974), .A2(n3973), .ZN(n5264) );
  NAND2_X1 U4865 ( .A1(n5255), .A2(n5264), .ZN(n3975) );
  MUX2_X1 U4866 ( .A(n5272), .B(n3976), .S(EBX_REG_24__SCAN_IN), .Z(n3978) );
  NAND2_X1 U4867 ( .A1(n4348), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3977) );
  AND2_X1 U4868 ( .A1(n3978), .A2(n3977), .ZN(n5201) );
  MUX2_X1 U4869 ( .A(n3979), .B(n5274), .S(EBX_REG_25__SCAN_IN), .Z(n3981) );
  OR2_X1 U4870 ( .A1(n4104), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3980)
         );
  AND2_X1 U4871 ( .A1(n3981), .A2(n3980), .ZN(n5189) );
  OR2_X1 U4872 ( .A1(n5272), .A2(EBX_REG_26__SCAN_IN), .ZN(n3985) );
  INV_X1 U4873 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U4874 ( .A1(n3976), .A2(n5529), .ZN(n3983) );
  INV_X1 U4875 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U4876 ( .A1(n4134), .A2(n5250), .ZN(n3982) );
  NAND3_X1 U4877 ( .A1(n3983), .A2(n5274), .A3(n3982), .ZN(n3984) );
  NAND2_X1 U4878 ( .A1(n3985), .A2(n3984), .ZN(n5180) );
  AND2_X1 U4879 ( .A1(n5191), .A2(n5180), .ZN(n3993) );
  INV_X1 U4880 ( .A(EBX_REG_27__SCAN_IN), .ZN(n3994) );
  NAND2_X1 U4881 ( .A1(n3986), .A2(n3994), .ZN(n3990) );
  NAND2_X1 U4882 ( .A1(n4134), .A2(n3994), .ZN(n3988) );
  NAND2_X1 U4883 ( .A1(n5274), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3987) );
  NAND3_X1 U4884 ( .A1(n3988), .A2(n3976), .A3(n3987), .ZN(n3989) );
  AND2_X1 U4885 ( .A1(n3990), .A2(n3989), .ZN(n3992) );
  AND2_X1 U4886 ( .A1(n3992), .A2(n5180), .ZN(n3991) );
  OAI21_X1 U4887 ( .B1(n3993), .B2(n3992), .A(n5156), .ZN(n5521) );
  NOR2_X1 U4888 ( .A1(n5878), .A2(n3994), .ZN(n3995) );
  NOR2_X1 U4889 ( .A1(n4001), .A2(n4000), .ZN(n4028) );
  AOI22_X1 U4890 ( .A1(n4046), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4891 ( .A1(n4052), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4892 ( .A1(n3310), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4893 ( .A1(n3274), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4002) );
  NAND4_X1 U4894 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4011)
         );
  AOI22_X1 U4895 ( .A1(n3256), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4896 ( .A1(n4053), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4897 ( .A1(n3266), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4898 ( .A1(n4054), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U4899 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4010)
         );
  OR2_X1 U4900 ( .A1(n4011), .A2(n4010), .ZN(n4027) );
  INV_X1 U4901 ( .A(n4027), .ZN(n4012) );
  XNOR2_X1 U4902 ( .A(n4028), .B(n4012), .ZN(n4017) );
  INV_X1 U4903 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4014) );
  NAND2_X1 U4904 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4013)
         );
  OAI211_X1 U4905 ( .C1(n4015), .C2(n4014), .A(n3338), .B(n4013), .ZN(n4016)
         );
  AOI21_X1 U4906 ( .B1(n4017), .B2(n4042), .A(n4016), .ZN(n4025) );
  INV_X1 U4907 ( .A(n4018), .ZN(n4019) );
  INV_X1 U4908 ( .A(n4020), .ZN(n4022) );
  INV_X1 U4909 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4021) );
  NAND2_X1 U4910 ( .A1(n4022), .A2(n4021), .ZN(n4023) );
  NAND2_X1 U4911 ( .A1(n4071), .A2(n4023), .ZN(n5341) );
  NOR2_X1 U4912 ( .A1(n5341), .A2(n3338), .ZN(n4024) );
  XNOR2_X1 U4913 ( .A(n4071), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5145)
         );
  NAND2_X1 U4914 ( .A1(n4028), .A2(n4027), .ZN(n4062) );
  AOI22_X1 U4915 ( .A1(n4053), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4916 ( .A1(n4045), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4917 ( .A1(n3310), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4918 ( .A1(n3256), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U4919 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4039)
         );
  AOI22_X1 U4920 ( .A1(n4046), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4921 ( .A1(n4052), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4922 ( .A1(n4054), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4923 ( .A1(n3362), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4034) );
  NAND4_X1 U4924 ( .A1(n4037), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(n4038)
         );
  NOR2_X1 U4925 ( .A1(n4039), .A2(n4038), .ZN(n4063) );
  XOR2_X1 U4926 ( .A(n4062), .B(n4063), .Z(n4043) );
  INV_X1 U4927 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U4928 ( .A1(n3337), .A2(EAX_REG_29__SCAN_IN), .ZN(n4040) );
  OAI211_X1 U4929 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n5146), .A(n4040), .B(
        n3338), .ZN(n4041) );
  AOI21_X1 U4930 ( .B1(n4043), .B2(n4042), .A(n4041), .ZN(n4044) );
  AOI22_X1 U4931 ( .A1(n4046), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4045), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4932 ( .A1(n3362), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4933 ( .A1(n3310), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4934 ( .A1(n3274), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4047), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4048) );
  NAND4_X1 U4935 ( .A1(n4051), .A2(n4050), .A3(n4049), .A4(n4048), .ZN(n4061)
         );
  AOI22_X1 U4936 ( .A1(n4052), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4033), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U4937 ( .A1(n3256), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4053), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U4938 ( .A1(n4054), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U4939 ( .A1(n3316), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4056) );
  NAND4_X1 U4940 ( .A1(n4059), .A2(n4058), .A3(n4057), .A4(n4056), .ZN(n4060)
         );
  NOR2_X1 U4941 ( .A1(n4061), .A2(n4060), .ZN(n4065) );
  NOR2_X1 U4942 ( .A1(n4063), .A2(n4062), .ZN(n4064) );
  XOR2_X1 U4943 ( .A(n4065), .B(n4064), .Z(n4070) );
  NAND2_X1 U4944 ( .A1(n6414), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4066)
         );
  NAND2_X1 U4945 ( .A1(n3338), .A2(n4066), .ZN(n4067) );
  AOI21_X1 U4946 ( .B1(n3337), .B2(EAX_REG_30__SCAN_IN), .A(n4067), .ZN(n4068)
         );
  OAI21_X1 U4947 ( .B1(n4070), .B2(n4069), .A(n4068), .ZN(n4074) );
  XNOR2_X1 U4948 ( .A(n4090), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5131)
         );
  NAND2_X1 U4949 ( .A1(n5131), .A2(n4072), .ZN(n4073) );
  NAND2_X1 U4950 ( .A1(n4074), .A2(n4073), .ZN(n4258) );
  AOI22_X1 U4951 ( .A1(n4076), .A2(EAX_REG_31__SCAN_IN), .B1(n4075), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4077) );
  INV_X1 U4952 ( .A(n4266), .ZN(n4270) );
  AND2_X1 U4953 ( .A1(n4082), .A2(n4081), .ZN(n4083) );
  NAND2_X1 U4954 ( .A1(n4084), .A2(n4083), .ZN(n4086) );
  NAND2_X1 U4955 ( .A1(n4086), .A2(n4085), .ZN(n4269) );
  INV_X1 U4956 ( .A(n4269), .ZN(n4087) );
  AND2_X1 U4957 ( .A1(n4296), .A2(n4087), .ZN(n4265) );
  NAND2_X1 U4958 ( .A1(n4265), .A2(n6420), .ZN(n4262) );
  OR2_X1 U4959 ( .A1(n4143), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6032) );
  NOR3_X1 U4960 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6520), .A3(n3338), .ZN(
        n6429) );
  OR2_X1 U4961 ( .A1(n6076), .A2(n6429), .ZN(n4088) );
  NAND2_X1 U4962 ( .A1(n6520), .A2(n6414), .ZN(n6430) );
  NOR3_X1 U4963 ( .A1(n6512), .A2(n6423), .A3(n6430), .ZN(n6418) );
  OR2_X1 U4964 ( .A1(n4088), .A2(n6418), .ZN(n4089) );
  INV_X1 U4965 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4256) );
  INV_X1 U4966 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6638) );
  NOR2_X1 U4967 ( .A1(n4883), .A2(n6520), .ZN(n4092) );
  NAND2_X1 U4968 ( .A1(n4149), .A2(n4093), .ZN(n4125) );
  OR2_X1 U4969 ( .A1(n5272), .A2(EBX_REG_28__SCAN_IN), .ZN(n4098) );
  INV_X1 U4970 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4094) );
  NAND2_X1 U4971 ( .A1(n3976), .A2(n4094), .ZN(n4096) );
  INV_X1 U4972 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U4973 ( .A1(n4134), .A2(n6630), .ZN(n4095) );
  NAND3_X1 U4974 ( .A1(n4096), .A2(n5274), .A3(n4095), .ZN(n4097) );
  AND2_X1 U4975 ( .A1(n4098), .A2(n4097), .ZN(n5155) );
  OR2_X1 U4976 ( .A1(n4104), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4101)
         );
  INV_X1 U4977 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U4978 ( .A1(n4134), .A2(n4099), .ZN(n4100) );
  NAND2_X1 U4979 ( .A1(n4101), .A2(n4100), .ZN(n4102) );
  MUX2_X1 U4980 ( .A(n4102), .B(EBX_REG_29__SCAN_IN), .S(n5128), .Z(n5143) );
  INV_X1 U4981 ( .A(n4104), .ZN(n4378) );
  INV_X1 U4982 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5139) );
  INV_X1 U4983 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5494) );
  OAI22_X1 U4984 ( .A1(n4378), .A2(n5139), .B1(n4134), .B2(n5494), .ZN(n5127)
         );
  NOR2_X1 U4985 ( .A1(n5143), .A2(n5127), .ZN(n4103) );
  NOR2_X1 U4986 ( .A1(n5126), .A2(n5128), .ZN(n5123) );
  AOI21_X1 U4987 ( .B1(n5144), .B2(n4103), .A(n5123), .ZN(n4106) );
  OAI22_X1 U4988 ( .A1(n4104), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4348), .B2(EBX_REG_31__SCAN_IN), .ZN(n4105) );
  XNOR2_X1 U4989 ( .A(n4106), .B(n4105), .ZN(n5490) );
  INV_X1 U4990 ( .A(READY_N), .ZN(n6538) );
  NAND2_X1 U4991 ( .A1(n6538), .A2(n6322), .ZN(n4877) );
  AND3_X1 U4992 ( .A1(n4134), .A2(EBX_REG_31__SCAN_IN), .A3(n4877), .ZN(n4107)
         );
  INV_X1 U4993 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6475) );
  INV_X1 U4994 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6473) );
  OR2_X1 U4995 ( .A1(n4108), .A2(STATE_REG_0__SCAN_IN), .ZN(n6442) );
  INV_X1 U4996 ( .A(n6442), .ZN(n4301) );
  OR2_X1 U4997 ( .A1(n4487), .A2(n4301), .ZN(n4359) );
  INV_X1 U4998 ( .A(n4877), .ZN(n4119) );
  AND2_X1 U4999 ( .A1(n3187), .A2(n4119), .ZN(n4109) );
  AND2_X1 U5000 ( .A1(n4359), .A2(n4109), .ZN(n4110) );
  INV_X1 U5001 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6467) );
  INV_X1 U5002 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6458) );
  INV_X1 U5003 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6456) );
  NAND3_X1 U5004 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5021) );
  NOR3_X1 U5005 ( .A1(n6458), .A2(n6456), .A3(n5021), .ZN(n4873) );
  INV_X1 U5006 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U5007 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n4943) );
  NOR2_X1 U5008 ( .A1(n6463), .A2(n4943), .ZN(n4937) );
  NAND4_X1 U5009 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n4873), .A4(n4937), .ZN(n5803) );
  NOR2_X1 U5010 ( .A1(n6467), .A2(n5803), .ZN(n5038) );
  NAND2_X1 U5011 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5038), .ZN(n4113) );
  NOR2_X1 U5012 ( .A1(n5787), .A2(n4113), .ZN(n5791) );
  NAND2_X1 U5013 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5791), .ZN(n5777) );
  NAND2_X1 U5014 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5766), .ZN(n5769) );
  NOR2_X1 U5015 ( .A1(n6475), .A2(n5769), .ZN(n5230) );
  NAND2_X1 U5016 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5230), .ZN(n5762) );
  NAND3_X1 U5017 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4111) );
  NOR2_X1 U5018 ( .A1(n5762), .A2(n4111), .ZN(n5648) );
  NAND4_X1 U5019 ( .A1(n5648), .A2(REIP_REG_23__SCAN_IN), .A3(
        REIP_REG_22__SCAN_IN), .A4(REIP_REG_21__SCAN_IN), .ZN(n5173) );
  AND2_X1 U5020 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5174) );
  NAND2_X1 U5021 ( .A1(n5174), .A2(REIP_REG_26__SCAN_IN), .ZN(n4115) );
  NOR2_X1 U5022 ( .A1(n5173), .A2(n4115), .ZN(n5171) );
  NAND3_X1 U5023 ( .A1(n5171), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5149) );
  INV_X1 U5024 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4112) );
  INV_X1 U5025 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6495) );
  NOR4_X1 U5026 ( .A1(n5149), .A2(REIP_REG_31__SCAN_IN), .A3(n4112), .A4(n6495), .ZN(n4123) );
  INV_X1 U5027 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5765) );
  INV_X1 U5028 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6471) );
  INV_X1 U5029 ( .A(n5785), .ZN(n5039) );
  NOR4_X1 U5030 ( .A1(n5434), .A2(n6475), .A3(n5765), .A4(n5763), .ZN(n5228)
         );
  NAND4_X1 U5031 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5228), .ZN(n5212) );
  NAND3_X1 U5032 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4114) );
  NAND2_X1 U5033 ( .A1(n5787), .A2(n5785), .ZN(n5764) );
  OAI21_X1 U5034 ( .B1(n5212), .B2(n4114), .A(n5764), .ZN(n5636) );
  INV_X1 U5035 ( .A(n5787), .ZN(n5865) );
  NAND2_X1 U5036 ( .A1(n5865), .A2(n4115), .ZN(n4116) );
  NAND2_X1 U5037 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4117) );
  NAND2_X1 U5038 ( .A1(n5865), .A2(n4117), .ZN(n4118) );
  OAI211_X1 U5039 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5787), .A(n5154), .B(
        REIP_REG_30__SCAN_IN), .ZN(n5134) );
  NAND3_X1 U5040 ( .A1(n5134), .A2(REIP_REG_31__SCAN_IN), .A3(n5764), .ZN(
        n4121) );
  NAND2_X1 U5041 ( .A1(n4301), .A2(n4119), .ZN(n6410) );
  AND2_X1 U5042 ( .A1(n4283), .A2(n6410), .ZN(n4876) );
  NAND3_X1 U5043 ( .A1(n4953), .A2(EBX_REG_31__SCAN_IN), .A3(n4876), .ZN(n4120) );
  OAI211_X1 U5044 ( .C1(n6638), .C2(n5856), .A(n4121), .B(n4120), .ZN(n4122)
         );
  AOI211_X1 U5045 ( .C1(n5490), .C2(n5825), .A(n4123), .B(n4122), .ZN(n4124)
         );
  NAND2_X1 U5046 ( .A1(n4125), .A2(n4124), .ZN(U2796) );
  AOI21_X1 U5047 ( .B1(n4126), .B2(n4332), .A(n4152), .ZN(n4127) );
  AND2_X1 U5048 ( .A1(n3878), .A2(n4127), .ZN(n4298) );
  AND2_X1 U5049 ( .A1(n4298), .A2(n4890), .ZN(n4320) );
  NAND2_X1 U5050 ( .A1(n6415), .A2(n4320), .ZN(n4130) );
  INV_X1 U5051 ( .A(n4128), .ZN(n5727) );
  NOR2_X1 U5052 ( .A1(READY_N), .A2(n4269), .ZN(n4353) );
  NAND2_X1 U5053 ( .A1(n5727), .A2(n4353), .ZN(n4129) );
  NAND2_X1 U5054 ( .A1(n4130), .A2(n4129), .ZN(n4310) );
  NOR2_X1 U5055 ( .A1(n4131), .A2(n4267), .ZN(n4132) );
  OAI21_X1 U5056 ( .B1(n4310), .B2(n4132), .A(n6420), .ZN(n4136) );
  AND2_X1 U5057 ( .A1(n4133), .A2(n4134), .ZN(n4367) );
  NAND2_X1 U5058 ( .A1(n4367), .A2(n6538), .ZN(n4135) );
  INV_X2 U5059 ( .A(n5120), .ZN(n5885) );
  NOR2_X2 U5060 ( .A1(n5885), .A2(n4360), .ZN(n5882) );
  AOI22_X1 U5061 ( .A1(n5882), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5885), .ZN(n4139) );
  NAND2_X1 U5062 ( .A1(n4140), .A2(n4139), .ZN(U2860) );
  NAND3_X1 U5063 ( .A1(n6423), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U5064 ( .A1(n6512), .A2(n6414), .ZN(n6325) );
  INV_X2 U5065 ( .A(n5987), .ZN(n5446) );
  INV_X1 U5066 ( .A(n4141), .ZN(n4142) );
  NAND2_X1 U5067 ( .A1(n4298), .A2(n4142), .ZN(n6400) );
  OR2_X2 U5068 ( .A1(n4364), .A2(n6400), .ZN(n5992) );
  NAND2_X1 U5069 ( .A1(n4143), .A2(n6325), .ZN(n6537) );
  NAND2_X1 U5070 ( .A1(n6537), .A2(n6423), .ZN(n4144) );
  NAND2_X1 U5071 ( .A1(n6423), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4146) );
  NAND2_X1 U5072 ( .A1(n6322), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4145) );
  AND2_X1 U5073 ( .A1(n4146), .A2(n4145), .ZN(n4404) );
  INV_X1 U5074 ( .A(n6032), .ZN(n6095) );
  AND2_X1 U5075 ( .A1(n6095), .A2(REIP_REG_31__SCAN_IN), .ZN(n5488) );
  AOI21_X1 U5076 ( .B1(n6006), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5488), 
        .ZN(n4147) );
  OAI21_X1 U5077 ( .B1(n6015), .B2(n4883), .A(n4147), .ZN(n4148) );
  AOI21_X1 U5078 ( .B1(n4149), .B2(n5446), .A(n4148), .ZN(n4250) );
  NAND2_X1 U5079 ( .A1(n4150), .A2(n4207), .ZN(n4157) );
  NAND2_X1 U5080 ( .A1(n4151), .A2(n4160), .ZN(n4173) );
  OAI21_X1 U5081 ( .B1(n4160), .B2(n4151), .A(n4173), .ZN(n4154) );
  INV_X1 U5082 ( .A(n4283), .ZN(n6541) );
  INV_X1 U5083 ( .A(n4152), .ZN(n4153) );
  OAI211_X1 U5084 ( .C1(n4154), .C2(n6541), .A(n4153), .B(n4479), .ZN(n4155)
         );
  INV_X1 U5085 ( .A(n4155), .ZN(n4156) );
  NAND2_X1 U5086 ( .A1(n4157), .A2(n4156), .ZN(n4396) );
  INV_X1 U5087 ( .A(n4207), .ZN(n4158) );
  AND2_X1 U5088 ( .A1(n4332), .A2(n4469), .ZN(n4168) );
  INV_X1 U5089 ( .A(n4168), .ZN(n4159) );
  OAI21_X1 U5090 ( .B1(n6541), .B2(n4160), .A(n4159), .ZN(n4161) );
  INV_X1 U5091 ( .A(n4161), .ZN(n4162) );
  NAND2_X1 U5092 ( .A1(n2966), .A2(n4162), .ZN(n4352) );
  AND2_X1 U5093 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U5094 ( .A1(n4352), .A2(n4163), .ZN(n4166) );
  NAND2_X1 U5095 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4164)
         );
  INV_X1 U5096 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U5097 ( .A1(n4164), .A2(n4905), .ZN(n4165) );
  AND2_X1 U5098 ( .A1(n4166), .A2(n4165), .ZN(n4395) );
  INV_X1 U5099 ( .A(n4166), .ZN(n4167) );
  AOI21_X1 U5100 ( .B1(n4396), .B2(n4395), .A(n4167), .ZN(n6009) );
  XNOR2_X1 U5101 ( .A(n4173), .B(n4172), .ZN(n4169) );
  AOI21_X1 U5102 ( .B1(n4169), .B2(n4283), .A(n4168), .ZN(n4170) );
  NAND2_X1 U5103 ( .A1(n6007), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4171)
         );
  AOI21_X1 U5104 ( .B1(n6009), .B2(n4171), .A(n3035), .ZN(n4511) );
  NAND2_X1 U5105 ( .A1(n4173), .A2(n4172), .ZN(n4181) );
  INV_X1 U5106 ( .A(n4180), .ZN(n4174) );
  XNOR2_X1 U5107 ( .A(n4181), .B(n4174), .ZN(n4175) );
  NAND2_X1 U5108 ( .A1(n4175), .A2(n4283), .ZN(n4176) );
  INV_X1 U5110 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U5111 ( .A1(n4511), .A2(n4512), .ZN(n4510) );
  NAND2_X1 U5112 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4178)
         );
  NAND2_X1 U5113 ( .A1(n4179), .A2(n4207), .ZN(n4184) );
  NAND2_X1 U5114 ( .A1(n4181), .A2(n4180), .ZN(n4200) );
  XNOR2_X1 U5115 ( .A(n4200), .B(n4197), .ZN(n4182) );
  NAND2_X1 U5116 ( .A1(n4182), .A2(n4283), .ZN(n4183) );
  NAND2_X1 U5117 ( .A1(n4184), .A2(n4183), .ZN(n4185) );
  INV_X1 U5118 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6561) );
  XNOR2_X1 U5119 ( .A(n4185), .B(n6561), .ZN(n5999) );
  NAND2_X1 U5120 ( .A1(n6000), .A2(n5999), .ZN(n5998) );
  NAND2_X1 U5121 ( .A1(n4185), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4186)
         );
  NAND2_X1 U5122 ( .A1(n5998), .A2(n4186), .ZN(n4772) );
  NAND2_X1 U5123 ( .A1(n4187), .A2(n4207), .ZN(n4192) );
  INV_X1 U5124 ( .A(n4197), .ZN(n4188) );
  OR2_X1 U5125 ( .A1(n4200), .A2(n4188), .ZN(n4189) );
  XNOR2_X1 U5126 ( .A(n4189), .B(n4198), .ZN(n4190) );
  NAND2_X1 U5127 ( .A1(n4190), .A2(n4283), .ZN(n4191) );
  INV_X1 U5128 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4193) );
  XNOR2_X1 U5129 ( .A(n4194), .B(n4193), .ZN(n4771) );
  NAND2_X1 U5130 ( .A1(n4772), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U5131 ( .A1(n4194), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4195)
         );
  NAND2_X1 U5132 ( .A1(n4196), .A2(n4207), .ZN(n4203) );
  NAND2_X1 U5133 ( .A1(n4198), .A2(n4197), .ZN(n4199) );
  OR2_X1 U5134 ( .A1(n4200), .A2(n4199), .ZN(n4208) );
  XNOR2_X1 U5135 ( .A(n4208), .B(n4209), .ZN(n4201) );
  NAND2_X1 U5136 ( .A1(n4201), .A2(n4283), .ZN(n4202) );
  NAND2_X1 U5137 ( .A1(n4203), .A2(n4202), .ZN(n4204) );
  XNOR2_X1 U5138 ( .A(n4204), .B(n5090), .ZN(n4902) );
  NAND2_X1 U5139 ( .A1(n4903), .A2(n4902), .ZN(n4901) );
  NAND2_X1 U5140 ( .A1(n4204), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4205)
         );
  NAND2_X1 U5141 ( .A1(n4901), .A2(n4205), .ZN(n4919) );
  NAND2_X1 U5142 ( .A1(n4206), .A2(n4207), .ZN(n4213) );
  INV_X1 U5143 ( .A(n4208), .ZN(n4210) );
  NAND2_X1 U5144 ( .A1(n4210), .A2(n4209), .ZN(n4219) );
  XNOR2_X1 U5145 ( .A(n4219), .B(n4220), .ZN(n4211) );
  NAND2_X1 U5146 ( .A1(n4211), .A2(n4283), .ZN(n4212) );
  NAND2_X1 U5147 ( .A1(n4213), .A2(n4212), .ZN(n4214) );
  INV_X1 U5148 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6646) );
  XNOR2_X1 U5149 ( .A(n4214), .B(n6646), .ZN(n4918) );
  NAND2_X1 U5150 ( .A1(n4919), .A2(n4918), .ZN(n4917) );
  NAND2_X1 U5151 ( .A1(n4214), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4215)
         );
  NOR3_X1 U5152 ( .A1(n4217), .A2(n4158), .A3(n6423), .ZN(n4218) );
  NAND2_X4 U5153 ( .A1(n4216), .A2(n4218), .ZN(n4226) );
  INV_X1 U5154 ( .A(n4219), .ZN(n4221) );
  NAND3_X1 U5155 ( .A1(n4221), .A2(n4283), .A3(n4220), .ZN(n4222) );
  NAND2_X1 U5156 ( .A1(n4226), .A2(n4222), .ZN(n4224) );
  XNOR2_X1 U5157 ( .A(n4224), .B(n4223), .ZN(n4961) );
  NAND2_X1 U5158 ( .A1(n4962), .A2(n4961), .ZN(n4960) );
  NAND2_X1 U5159 ( .A1(n4224), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4225)
         );
  NAND2_X1 U5160 ( .A1(n4960), .A2(n4225), .ZN(n5046) );
  INV_X1 U5161 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U5162 ( .A1(n4226), .A2(n5047), .ZN(n4227) );
  NAND2_X1 U5163 ( .A1(n5046), .A2(n4227), .ZN(n4229) );
  NAND2_X1 U5164 ( .A1(n2953), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4228)
         );
  INV_X1 U5165 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4230) );
  NAND2_X1 U5166 ( .A1(n4226), .A2(n4230), .ZN(n5055) );
  INV_X1 U5167 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6022) );
  AND2_X1 U5168 ( .A1(n4226), .A2(n6022), .ZN(n4233) );
  NAND2_X1 U5169 ( .A1(n2953), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U5170 ( .A1(n2953), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4231) );
  INV_X1 U5171 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5704) );
  NOR2_X1 U5172 ( .A1(n4226), .A2(n5704), .ZN(n5086) );
  XNOR2_X1 U5173 ( .A(n4226), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5682)
         );
  NAND2_X1 U5174 ( .A1(n5681), .A2(n5682), .ZN(n4236) );
  INV_X1 U5175 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4234) );
  NAND2_X1 U5176 ( .A1(n4226), .A2(n4234), .ZN(n4235) );
  INV_X1 U5177 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U5178 ( .A1(n2953), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4237) );
  INV_X1 U5179 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U5180 ( .A1(n4226), .A2(n5420), .ZN(n5449) );
  NAND2_X1 U5181 ( .A1(n4226), .A2(n6595), .ZN(n4239) );
  NAND2_X1 U5183 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U5184 ( .A1(n4226), .A2(n5593), .ZN(n4240) );
  INV_X1 U5186 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5617) );
  INV_X1 U5187 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5615) );
  NAND3_X1 U5188 ( .A1(n5617), .A2(n5615), .A3(n6595), .ZN(n4241) );
  NAND2_X1 U5189 ( .A1(n2953), .A2(n4241), .ZN(n4242) );
  NOR2_X1 U5190 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5562) );
  NOR2_X1 U5191 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5595) );
  INV_X1 U5192 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5558) );
  INV_X1 U5193 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5547) );
  NAND4_X1 U5194 ( .A1(n5562), .A2(n5595), .A3(n5558), .A4(n5547), .ZN(n4243)
         );
  NAND2_X1 U5195 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U5196 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5476) );
  NOR2_X1 U5197 ( .A1(n5474), .A2(n5476), .ZN(n5467) );
  AND2_X1 U5198 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5594) );
  INV_X1 U5199 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5542) );
  XNOR2_X1 U5200 ( .A(n4226), .B(n5542), .ZN(n5363) );
  NAND2_X1 U5201 ( .A1(n4226), .A2(n5542), .ZN(n4247) );
  AND2_X1 U5202 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U5203 ( .A1(n5345), .A2(n5512), .ZN(n5325) );
  NAND2_X1 U5204 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5484) );
  NOR2_X1 U5205 ( .A1(n4226), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5336)
         );
  NOR2_X1 U5206 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U5207 ( .A1(n5336), .A2(n5513), .ZN(n5326) );
  NOR2_X1 U5208 ( .A1(n5326), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4252)
         );
  NAND2_X1 U5209 ( .A1(n4252), .A2(n5494), .ZN(n4249) );
  AND2_X1 U5210 ( .A1(n4251), .A2(n4252), .ZN(n4253) );
  XNOR2_X1 U5211 ( .A(n4255), .B(n5494), .ZN(n5502) );
  INV_X1 U5212 ( .A(n6015), .ZN(n5464) );
  INV_X1 U5213 ( .A(n6006), .ZN(n5461) );
  NAND2_X1 U5214 ( .A1(n6095), .A2(REIP_REG_30__SCAN_IN), .ZN(n5496) );
  OAI21_X1 U5215 ( .B1(n5461), .B2(n4256), .A(n5496), .ZN(n4257) );
  AOI21_X1 U5216 ( .B1(n5131), .B2(n5464), .A(n4257), .ZN(n4259) );
  OAI211_X1 U5217 ( .C1(n5502), .C2(n5992), .A(n4259), .B(n3038), .ZN(U2956)
         );
  AND2_X1 U5218 ( .A1(n4296), .A2(n4487), .ZN(n6383) );
  NAND2_X1 U5219 ( .A1(n4133), .A2(n4283), .ZN(n6411) );
  INV_X1 U5220 ( .A(n6411), .ZN(n4260) );
  OAI21_X1 U5221 ( .B1(n6383), .B2(n4260), .A(n4301), .ZN(n4261) );
  NOR2_X1 U5222 ( .A1(n6520), .A2(n6414), .ZN(n4444) );
  NAND2_X1 U5223 ( .A1(n6423), .A2(n4444), .ZN(n5915) );
  AND2_X2 U5224 ( .A1(n5919), .A2(n5915), .ZN(n5917) );
  AND2_X1 U5225 ( .A1(n5917), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U5226 ( .A(n4262), .ZN(n4264) );
  INV_X1 U5227 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6590) );
  NOR2_X1 U5228 ( .A1(n6325), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4875) );
  INV_X1 U5229 ( .A(n4875), .ZN(n4263) );
  OAI211_X1 U5230 ( .C1(n4264), .C2(n6590), .A(n4281), .B(n4263), .ZN(U2788)
         );
  OAI22_X1 U5231 ( .A1(n6415), .A2(n4890), .B1(n4266), .B2(n4265), .ZN(n5735)
         );
  NAND2_X1 U5232 ( .A1(n4348), .A2(n4267), .ZN(n4278) );
  OR2_X1 U5233 ( .A1(n4278), .A2(n4301), .ZN(n4268) );
  AND2_X1 U5234 ( .A1(n4268), .A2(n6538), .ZN(n6540) );
  OR2_X1 U5235 ( .A1(n5735), .A2(n6540), .ZN(n6403) );
  AND2_X1 U5236 ( .A1(n6403), .A2(n6420), .ZN(n5741) );
  INV_X1 U5237 ( .A(MORE_REG_SCAN_IN), .ZN(n6605) );
  INV_X1 U5238 ( .A(n4321), .ZN(n4379) );
  NAND2_X1 U5239 ( .A1(n4379), .A2(n6415), .ZN(n4275) );
  NAND2_X1 U5240 ( .A1(n4296), .A2(n4269), .ZN(n4274) );
  NAND2_X1 U5241 ( .A1(n4270), .A2(n6400), .ZN(n4271) );
  NOR2_X1 U5242 ( .A1(n4271), .A2(n4320), .ZN(n4272) );
  OR2_X1 U5243 ( .A1(n6415), .A2(n4272), .ZN(n4273) );
  AND3_X1 U5244 ( .A1(n4275), .A2(n4274), .A3(n4273), .ZN(n6401) );
  INV_X1 U5245 ( .A(n6401), .ZN(n4276) );
  NAND2_X1 U5246 ( .A1(n5741), .A2(n4276), .ZN(n4277) );
  OAI21_X1 U5247 ( .B1(n5741), .B2(n6605), .A(n4277), .ZN(U3471) );
  NOR2_X1 U5248 ( .A1(n4875), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4280) );
  NAND2_X1 U5249 ( .A1(n6536), .A2(n4278), .ZN(n4279) );
  OAI21_X1 U5250 ( .B1(n6536), .B2(n4280), .A(n4279), .ZN(U3474) );
  INV_X1 U5251 ( .A(n4281), .ZN(n4282) );
  OAI21_X1 U5252 ( .B1(n4283), .B2(n6538), .A(n4282), .ZN(n5965) );
  INV_X1 U5253 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n6571) );
  INV_X1 U5254 ( .A(n5980), .ZN(n5971) );
  AND2_X1 U5255 ( .A1(n5977), .A2(DATAI_6_), .ZN(n5951) );
  AOI21_X1 U5256 ( .B1(n5971), .B2(EAX_REG_22__SCAN_IN), .A(n5951), .ZN(n4284)
         );
  OAI21_X1 U5257 ( .B1(n5924), .B2(n6571), .A(n4284), .ZN(U2930) );
  INV_X1 U5258 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n6610) );
  INV_X1 U5259 ( .A(DATAI_14_), .ZN(n4285) );
  NOR2_X1 U5260 ( .A1(n5936), .A2(n4285), .ZN(n5974) );
  AOI21_X1 U5261 ( .B1(n5971), .B2(EAX_REG_30__SCAN_IN), .A(n5974), .ZN(n4286)
         );
  OAI21_X1 U5262 ( .B1(n5924), .B2(n6610), .A(n4286), .ZN(U2938) );
  INV_X1 U5263 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n6582) );
  AND2_X1 U5264 ( .A1(n5977), .A2(DATAI_2_), .ZN(n5942) );
  AOI21_X1 U5265 ( .B1(n5971), .B2(EAX_REG_18__SCAN_IN), .A(n5942), .ZN(n4287)
         );
  OAI21_X1 U5266 ( .B1(n5924), .B2(n6582), .A(n4287), .ZN(U2926) );
  INV_X1 U5267 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6669) );
  INV_X1 U5268 ( .A(DATAI_11_), .ZN(n4288) );
  NOR2_X1 U5269 ( .A1(n5936), .A2(n4288), .ZN(n5964) );
  AOI21_X1 U5270 ( .B1(n5971), .B2(EAX_REG_27__SCAN_IN), .A(n5964), .ZN(n4289)
         );
  OAI21_X1 U5271 ( .B1(n5924), .B2(n6669), .A(n4289), .ZN(U2935) );
  INV_X1 U5272 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n5916) );
  INV_X1 U5273 ( .A(DATAI_1_), .ZN(n4290) );
  NOR2_X1 U5274 ( .A1(n5936), .A2(n4290), .ZN(n5922) );
  AOI21_X1 U5275 ( .B1(n5971), .B2(EAX_REG_1__SCAN_IN), .A(n5922), .ZN(n4291)
         );
  OAI21_X1 U5276 ( .B1(n5924), .B2(n5916), .A(n4291), .ZN(U2940) );
  INV_X1 U5277 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U5278 ( .A1(n5971), .A2(EAX_REG_5__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U5279 ( .A1(n5977), .A2(DATAI_5_), .ZN(n4293) );
  OAI211_X1 U5280 ( .C1(n5924), .C2(n5909), .A(n4292), .B(n4293), .ZN(U2944)
         );
  INV_X1 U5281 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U5282 ( .A1(n5971), .A2(EAX_REG_21__SCAN_IN), .ZN(n4294) );
  OAI211_X1 U5283 ( .C1(n5924), .C2(n6666), .A(n4294), .B(n4293), .ZN(U2929)
         );
  INV_X1 U5284 ( .A(n4295), .ZN(n4314) );
  INV_X1 U5285 ( .A(n6514), .ZN(n5114) );
  INV_X1 U5286 ( .A(n4296), .ZN(n4300) );
  NAND2_X1 U5287 ( .A1(n4298), .A2(n4297), .ZN(n4299) );
  NAND2_X1 U5288 ( .A1(n4300), .A2(n4299), .ZN(n4356) );
  OAI21_X1 U5289 ( .B1(n6383), .B2(n4133), .A(n4301), .ZN(n4303) );
  INV_X1 U5290 ( .A(n4367), .ZN(n4302) );
  NAND2_X1 U5291 ( .A1(n4303), .A2(n4302), .ZN(n4305) );
  AND2_X1 U5292 ( .A1(n6415), .A2(n6538), .ZN(n4304) );
  NAND2_X1 U5293 ( .A1(n4305), .A2(n4304), .ZN(n4308) );
  INV_X1 U5294 ( .A(n4306), .ZN(n4307) );
  AND4_X1 U5295 ( .A1(n4309), .A2(n4356), .A3(n4308), .A4(n4307), .ZN(n4312)
         );
  INV_X1 U5296 ( .A(n4310), .ZN(n4311) );
  NAND2_X1 U5297 ( .A1(n4312), .A2(n4311), .ZN(n6384) );
  INV_X1 U5298 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5740) );
  NAND2_X1 U5299 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4444), .ZN(n6509) );
  NOR2_X1 U5300 ( .A1(n5740), .A2(n6509), .ZN(n4313) );
  AOI21_X1 U5301 ( .B1(n6420), .B2(n6384), .A(n4313), .ZN(n5732) );
  NOR2_X1 U5302 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6512), .ZN(n4468) );
  INV_X1 U5303 ( .A(n4468), .ZN(n6510) );
  NAND2_X1 U5304 ( .A1(n5732), .A2(n6510), .ZN(n6521) );
  INV_X1 U5305 ( .A(n6521), .ZN(n5115) );
  AOI21_X1 U5306 ( .B1(n4314), .B2(n5114), .A(n5115), .ZN(n4331) );
  INV_X1 U5307 ( .A(n4133), .ZN(n4316) );
  NAND3_X1 U5308 ( .A1(n4316), .A2(n4381), .A3(n3889), .ZN(n4317) );
  NOR2_X1 U5309 ( .A1(n4318), .A2(n4317), .ZN(n4319) );
  AND2_X1 U5310 ( .A1(n4128), .A2(n4319), .ZN(n5111) );
  INV_X1 U5311 ( .A(n4320), .ZN(n4369) );
  NAND2_X1 U5312 ( .A1(n4321), .A2(n4369), .ZN(n4427) );
  XNOR2_X1 U5313 ( .A(n4295), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4325)
         );
  XNOR2_X1 U5314 ( .A(n3039), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4322)
         );
  NAND2_X1 U5315 ( .A1(n6383), .A2(n4322), .ZN(n4323) );
  OAI21_X1 U5316 ( .B1(n4325), .B2(n4424), .A(n4323), .ZN(n4324) );
  AOI21_X1 U5317 ( .B1(n4427), .B2(n4325), .A(n4324), .ZN(n4326) );
  OAI21_X1 U5318 ( .B1(n4315), .B2(n5111), .A(n4326), .ZN(n4432) );
  INV_X1 U5319 ( .A(n6525), .ZN(n5728) );
  INV_X1 U5320 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5485) );
  AOI22_X1 U5321 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5485), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4905), .ZN(n5113) );
  NAND2_X1 U5322 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5108) );
  NAND3_X1 U5323 ( .A1(n4295), .A2(n4330), .A3(n5114), .ZN(n4327) );
  OAI21_X1 U5324 ( .B1(n5113), .B2(n5108), .A(n4327), .ZN(n4328) );
  AOI21_X1 U5325 ( .B1(n4432), .B2(n5728), .A(n4328), .ZN(n4329) );
  OAI22_X1 U5326 ( .A1(n4331), .A2(n4330), .B1(n4329), .B2(n5115), .ZN(U3459)
         );
  INV_X1 U5327 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5930) );
  OR2_X1 U5328 ( .A1(n5919), .A2(n4332), .ZN(n5889) );
  INV_X1 U5329 ( .A(n5915), .ZN(n5898) );
  AOI22_X1 U5330 ( .A1(n5898), .A2(UWORD_REG_8__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4333) );
  OAI21_X1 U5331 ( .B1(n5930), .B2(n5889), .A(n4333), .ZN(U2899) );
  INV_X1 U5332 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5921) );
  AOI22_X1 U5333 ( .A1(n5898), .A2(UWORD_REG_0__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4334) );
  OAI21_X1 U5334 ( .B1(n5921), .B2(n5889), .A(n4334), .ZN(U2907) );
  AOI22_X1 U5335 ( .A1(n5898), .A2(UWORD_REG_4__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4335) );
  OAI21_X1 U5336 ( .B1(n3668), .B2(n5889), .A(n4335), .ZN(U2903) );
  INV_X1 U5337 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5926) );
  AOI22_X1 U5338 ( .A1(n5898), .A2(UWORD_REG_3__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4336) );
  OAI21_X1 U5339 ( .B1(n5926), .B2(n5889), .A(n4336), .ZN(U2904) );
  NAND2_X1 U5340 ( .A1(n4337), .A2(n3894), .ZN(n4342) );
  NAND2_X2 U5341 ( .A1(n5120), .A2(n4342), .ZN(n5671) );
  OR2_X1 U5342 ( .A1(n4339), .A2(n4338), .ZN(n4340) );
  NAND2_X1 U5343 ( .A1(n4341), .A2(n4340), .ZN(n4959) );
  INV_X1 U5344 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5941) );
  INV_X1 U5345 ( .A(n4342), .ZN(n4343) );
  INV_X1 U5346 ( .A(DATAI_0_), .ZN(n4483) );
  OAI222_X1 U5347 ( .A1(n5671), .A2(n4959), .B1(n5120), .B2(n5941), .C1(n4782), 
        .C2(n4483), .ZN(U2891) );
  OAI21_X1 U5348 ( .B1(n4345), .B2(n4344), .A(n3347), .ZN(n4976) );
  AOI22_X1 U5349 ( .A1(n5322), .A2(DATAI_1_), .B1(n5885), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4346) );
  OAI21_X1 U5350 ( .B1(n4976), .B2(n5671), .A(n4346), .ZN(U2890) );
  INV_X1 U5351 ( .A(n4347), .ZN(n4349) );
  NAND2_X1 U5352 ( .A1(n4349), .A2(n4348), .ZN(n4351) );
  AND2_X1 U5353 ( .A1(n4351), .A2(n4350), .ZN(n4968) );
  OAI222_X1 U5354 ( .A1(n4976), .A2(n5300), .B1(n2978), .B2(n5878), .C1(n5872), 
        .C2(n4968), .ZN(U2858) );
  XNOR2_X1 U5355 ( .A(n4352), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4409)
         );
  NAND2_X1 U5356 ( .A1(n6380), .A2(n4487), .ZN(n4357) );
  NAND2_X1 U5357 ( .A1(n4487), .A2(n6442), .ZN(n4354) );
  NAND3_X1 U5358 ( .A1(n4354), .A2(n4353), .A3(n4497), .ZN(n4355) );
  OAI211_X1 U5359 ( .C1(n6415), .C2(n4357), .A(n4356), .B(n4355), .ZN(n4358)
         );
  NAND2_X1 U5360 ( .A1(n4358), .A2(n6420), .ZN(n4366) );
  NAND3_X1 U5361 ( .A1(n4133), .A2(n4359), .A3(n6538), .ZN(n4361) );
  NAND3_X1 U5362 ( .A1(n4361), .A2(n3187), .A3(n4360), .ZN(n4362) );
  NAND2_X1 U5363 ( .A1(n4362), .A2(n3183), .ZN(n4363) );
  AND2_X1 U5364 ( .A1(n4373), .A2(n4491), .ZN(n4368) );
  NOR2_X1 U5365 ( .A1(n4368), .A2(n4367), .ZN(n4370) );
  NAND4_X1 U5366 ( .A1(n4128), .A2(n4370), .A3(n4369), .A4(n6400), .ZN(n4371)
         );
  NAND2_X1 U5367 ( .A1(n4373), .A2(n4372), .ZN(n4374) );
  NAND2_X1 U5368 ( .A1(n4374), .A2(n6411), .ZN(n4375) );
  INV_X1 U5369 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4386) );
  INV_X1 U5370 ( .A(n4376), .ZN(n4377) );
  AOI21_X1 U5371 ( .B1(n4378), .B2(n4386), .A(n4377), .ZN(n4954) );
  AND2_X1 U5372 ( .A1(n6095), .A2(REIP_REG_0__SCAN_IN), .ZN(n4406) );
  OAI21_X1 U5373 ( .B1(n3187), .B2(n4381), .A(n4380), .ZN(n4382) );
  NAND2_X1 U5374 ( .A1(n4385), .A2(n4382), .ZN(n5706) );
  AND2_X1 U5375 ( .A1(n6099), .A2(n5706), .ZN(n5710) );
  OR2_X1 U5376 ( .A1(n5710), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4384)
         );
  OR2_X1 U5377 ( .A1(n4385), .A2(n6095), .ZN(n4383) );
  NAND2_X1 U5378 ( .A1(n4384), .A2(n4383), .ZN(n4906) );
  INV_X1 U5379 ( .A(n4906), .ZN(n4387) );
  INV_X1 U5380 ( .A(n5719), .ZN(n4397) );
  AOI22_X1 U5381 ( .A1(n4387), .A2(n4397), .B1(n5710), .B2(n4386), .ZN(n4388)
         );
  AOI211_X1 U5382 ( .C1(n6097), .C2(n4954), .A(n4406), .B(n4388), .ZN(n4389)
         );
  OAI21_X1 U5383 ( .B1(n4409), .B2(n6086), .A(n4389), .ZN(U3018) );
  INV_X1 U5384 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6626) );
  AOI22_X1 U5385 ( .A1(n5898), .A2(UWORD_REG_1__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4390) );
  OAI21_X1 U5386 ( .B1(n6626), .B2(n5889), .A(n4390), .ZN(U2906) );
  INV_X1 U5387 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U5388 ( .A1(n5898), .A2(UWORD_REG_7__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4391) );
  OAI21_X1 U5389 ( .B1(n6670), .B2(n5889), .A(n4391), .ZN(U2900) );
  AOI22_X1 U5390 ( .A1(n6539), .A2(UWORD_REG_12__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4392) );
  OAI21_X1 U5391 ( .B1(n4014), .B2(n5889), .A(n4392), .ZN(U2895) );
  INV_X1 U5392 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5933) );
  AOI22_X1 U5393 ( .A1(n6539), .A2(UWORD_REG_9__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4393) );
  OAI21_X1 U5394 ( .B1(n5933), .B2(n5889), .A(n4393), .ZN(U2898) );
  AOI22_X1 U5395 ( .A1(n6539), .A2(UWORD_REG_10__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4394) );
  OAI21_X1 U5396 ( .B1(n3787), .B2(n5889), .A(n4394), .ZN(U2897) );
  XNOR2_X1 U5397 ( .A(n4396), .B(n4395), .ZN(n4509) );
  INV_X1 U5398 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6527) );
  OAI22_X1 U5399 ( .A1(n6079), .A2(n4968), .B1(n6527), .B2(n6032), .ZN(n4399)
         );
  NAND2_X1 U5400 ( .A1(n6030), .A2(n6099), .ZN(n6031) );
  INV_X1 U5401 ( .A(n6031), .ZN(n5691) );
  NOR2_X1 U5402 ( .A1(n5719), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4907)
         );
  NOR3_X1 U5403 ( .A1(n5691), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4907), 
        .ZN(n4398) );
  AOI211_X1 U5404 ( .C1(INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n4906), .A(n4399), 
        .B(n4398), .ZN(n4400) );
  OAI21_X1 U5405 ( .B1(n4509), .B2(n6086), .A(n4400), .ZN(U3017) );
  INV_X1 U5406 ( .A(n4954), .ZN(n4402) );
  OAI222_X1 U5407 ( .A1(n4402), .A2(n5872), .B1(n4401), .B2(n5878), .C1(n4959), 
        .C2(n5300), .ZN(U2859) );
  INV_X1 U5408 ( .A(n4959), .ZN(n4407) );
  INV_X1 U5409 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4403) );
  AOI21_X1 U5410 ( .B1(n5461), .B2(n4404), .A(n4403), .ZN(n4405) );
  AOI211_X1 U5411 ( .C1(n4407), .C2(n5446), .A(n4406), .B(n4405), .ZN(n4408)
         );
  OAI21_X1 U5412 ( .B1(n4409), .B2(n5992), .A(n4408), .ZN(U2986) );
  NAND3_X1 U5413 ( .A1(n4412), .A2(n4411), .A3(n3347), .ZN(n4413) );
  AND2_X1 U5414 ( .A1(n4410), .A2(n4413), .ZN(n6010) );
  INV_X1 U5415 ( .A(n6010), .ZN(n4417) );
  AOI21_X1 U5416 ( .B1(n4415), .B2(n4414), .A(n2983), .ZN(n6096) );
  INV_X1 U5417 ( .A(n5878), .ZN(n5286) );
  AOI22_X1 U5418 ( .A1(n3996), .A2(n6096), .B1(EBX_REG_2__SCAN_IN), .B2(n5286), 
        .ZN(n4416) );
  OAI21_X1 U5419 ( .B1(n4417), .B2(n5300), .A(n4416), .ZN(U2857) );
  INV_X1 U5420 ( .A(DATAI_2_), .ZN(n4496) );
  INV_X1 U5421 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5944) );
  OAI222_X1 U5422 ( .A1(n4417), .A2(n5671), .B1(n4782), .B2(n4496), .C1(n5120), 
        .C2(n5944), .ZN(U2889) );
  INV_X1 U5423 ( .A(n5111), .ZN(n6381) );
  NAND2_X1 U5424 ( .A1(n6146), .A2(n6381), .ZN(n4429) );
  NOR2_X1 U5425 ( .A1(n4295), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4419)
         );
  XNOR2_X1 U5426 ( .A(n4419), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4426)
         );
  AOI21_X1 U5427 ( .B1(n4295), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4430), 
        .ZN(n4420) );
  NOR2_X1 U5428 ( .A1(n3274), .A2(n4420), .ZN(n6515) );
  NAND2_X1 U5429 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4421) );
  XNOR2_X1 U5430 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n4421), .ZN(n4422)
         );
  NAND2_X1 U5431 ( .A1(n6383), .A2(n4422), .ZN(n4423) );
  OAI21_X1 U5432 ( .B1(n6515), .B2(n4424), .A(n4423), .ZN(n4425) );
  AOI21_X1 U5433 ( .B1(n4427), .B2(n4426), .A(n4425), .ZN(n4428) );
  NAND2_X1 U5434 ( .A1(n4429), .A2(n4428), .ZN(n6513) );
  NOR2_X1 U5435 ( .A1(n6384), .A2(n4430), .ZN(n4431) );
  AOI21_X1 U5436 ( .B1(n6513), .B2(n6384), .A(n4431), .ZN(n6396) );
  INV_X1 U5437 ( .A(n6396), .ZN(n4433) );
  MUX2_X1 U5438 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4432), .S(n6384), 
        .Z(n6394) );
  NAND3_X1 U5439 ( .A1(n4433), .A2(n6394), .A3(n6520), .ZN(n4436) );
  NOR2_X1 U5440 ( .A1(n6520), .A2(FLUSH_REG_SCAN_IN), .ZN(n4440) );
  NAND2_X1 U5441 ( .A1(n4434), .A2(n4440), .ZN(n4435) );
  AND2_X1 U5442 ( .A1(n4436), .A2(n4435), .ZN(n6406) );
  NOR2_X1 U5443 ( .A1(n6406), .A2(n4437), .ZN(n4446) );
  INV_X1 U5444 ( .A(n6326), .ZN(n4574) );
  NOR2_X1 U5445 ( .A1(n3350), .A2(n4574), .ZN(n4438) );
  XNOR2_X1 U5446 ( .A(n4438), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5852)
         );
  OAI22_X1 U5447 ( .A1(n5852), .A2(n4128), .B1(n5730), .B2(n6384), .ZN(n4439)
         );
  NAND2_X1 U5448 ( .A1(n4439), .A2(n6520), .ZN(n4442) );
  NAND2_X1 U5449 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4440), .ZN(n4441) );
  NAND2_X1 U5450 ( .A1(n4442), .A2(n4441), .ZN(n6405) );
  NOR3_X1 U5451 ( .A1(n4446), .A2(n6405), .A3(FLUSH_REG_SCAN_IN), .ZN(n4443)
         );
  INV_X1 U5452 ( .A(n6430), .ZN(n6542) );
  OAI21_X1 U5453 ( .B1(n4443), .B2(n6509), .A(n4744), .ZN(n6108) );
  INV_X1 U5454 ( .A(n4444), .ZN(n4445) );
  OR3_X1 U5455 ( .A1(n4446), .A2(n6405), .A3(n4445), .ZN(n6422) );
  INV_X1 U5456 ( .A(n6422), .ZN(n4448) );
  NAND2_X1 U5457 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6512), .ZN(n5629) );
  INV_X1 U5458 ( .A(n5629), .ZN(n5626) );
  OAI22_X1 U5459 ( .A1(n4977), .A2(n6325), .B1(n2956), .B2(n5626), .ZN(n4447)
         );
  OAI21_X1 U5460 ( .B1(n4448), .B2(n4447), .A(n6108), .ZN(n4449) );
  OAI21_X1 U5461 ( .B1(n6108), .B2(n4660), .A(n4449), .ZN(U3465) );
  INV_X1 U5462 ( .A(n4450), .ZN(n4451) );
  AOI21_X1 U5463 ( .B1(n4452), .B2(n4410), .A(n4451), .ZN(n4515) );
  INV_X1 U5464 ( .A(n4515), .ZN(n5033) );
  AND2_X1 U5465 ( .A1(n4454), .A2(n4453), .ZN(n4455) );
  NOR2_X1 U5466 ( .A1(n4567), .A2(n4455), .ZN(n6084) );
  AOI22_X1 U5467 ( .A1(n3996), .A2(n6084), .B1(EBX_REG_3__SCAN_IN), .B2(n5286), 
        .ZN(n4456) );
  OAI21_X1 U5468 ( .B1(n5033), .B2(n5300), .A(n4456), .ZN(U2856) );
  NAND2_X1 U5469 ( .A1(n6112), .A2(n4458), .ZN(n4531) );
  NAND2_X1 U5470 ( .A1(n5446), .A2(DATAI_27_), .ZN(n6353) );
  AOI21_X1 U5471 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4660), .A(n4744), .ZN(
        n6116) );
  NOR2_X1 U5472 ( .A1(n6317), .A2(n2956), .ZN(n4662) );
  NOR2_X1 U5473 ( .A1(n4315), .A2(n5624), .ZN(n6224) );
  INV_X1 U5474 ( .A(n4499), .ZN(n4460) );
  AOI21_X1 U5475 ( .B1(n4662), .B2(n6224), .A(n4460), .ZN(n4464) );
  OR2_X1 U5476 ( .A1(n6325), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6148) );
  OAI21_X1 U5477 ( .B1(n4463), .B2(n5987), .A(n6148), .ZN(n4461) );
  AOI22_X1 U5478 ( .A1(n4464), .A2(n4461), .B1(n4697), .B2(n6325), .ZN(n4462)
         );
  NAND2_X1 U5479 ( .A1(n6116), .A2(n4462), .ZN(n4495) );
  NAND2_X1 U5480 ( .A1(n4495), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4472)
         );
  NAND2_X1 U5481 ( .A1(n5446), .A2(DATAI_19_), .ZN(n6290) );
  INV_X1 U5482 ( .A(n6290), .ZN(n6350) );
  INV_X1 U5483 ( .A(n4464), .ZN(n4466) );
  INV_X1 U5484 ( .A(n6325), .ZN(n6218) );
  AOI22_X1 U5485 ( .A1(n4466), .A2(n6218), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4465), .ZN(n4500) );
  INV_X1 U5486 ( .A(DATAI_3_), .ZN(n4504) );
  NOR2_X1 U5487 ( .A1(n4504), .A2(n4744), .ZN(n6349) );
  INV_X1 U5488 ( .A(n6349), .ZN(n5008) );
  NAND2_X1 U5489 ( .A1(n4498), .A2(n4469), .ZN(n6286) );
  OAI22_X1 U5490 ( .A1(n4500), .A2(n5008), .B1(n4499), .B2(n6286), .ZN(n4470)
         );
  AOI21_X1 U5491 ( .B1(n6350), .B2(n4619), .A(n4470), .ZN(n4471) );
  OAI211_X1 U5492 ( .C1(n4736), .C2(n6353), .A(n4472), .B(n4471), .ZN(U3143)
         );
  NAND2_X1 U5493 ( .A1(n5446), .A2(DATAI_30_), .ZN(n6371) );
  NAND2_X1 U5494 ( .A1(n4495), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4475)
         );
  NAND2_X1 U5495 ( .A1(n5446), .A2(DATAI_22_), .ZN(n6305) );
  INV_X1 U5496 ( .A(n6305), .ZN(n6368) );
  INV_X1 U5497 ( .A(DATAI_6_), .ZN(n4768) );
  NOR2_X1 U5498 ( .A1(n4768), .A2(n4744), .ZN(n6367) );
  INV_X1 U5499 ( .A(n6367), .ZN(n5012) );
  NAND2_X1 U5500 ( .A1(n4498), .A2(n3214), .ZN(n6301) );
  OAI22_X1 U5501 ( .A1(n4500), .A2(n5012), .B1(n4499), .B2(n6301), .ZN(n4473)
         );
  AOI21_X1 U5502 ( .B1(n6368), .B2(n4619), .A(n4473), .ZN(n4474) );
  OAI211_X1 U5503 ( .C1(n4736), .C2(n6371), .A(n4475), .B(n4474), .ZN(U3146)
         );
  NAND2_X1 U5504 ( .A1(n5446), .A2(DATAI_31_), .ZN(n6559) );
  NAND2_X1 U5505 ( .A1(n4495), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4478)
         );
  NAND2_X1 U5506 ( .A1(n5446), .A2(DATAI_23_), .ZN(n6314) );
  INV_X1 U5507 ( .A(n6314), .ZN(n6556) );
  INV_X1 U5508 ( .A(DATAI_7_), .ZN(n4737) );
  NOR2_X1 U5509 ( .A1(n4737), .A2(n4744), .ZN(n6374) );
  INV_X1 U5510 ( .A(n6374), .ZN(n6553) );
  NAND2_X1 U5511 ( .A1(n4498), .A2(n3894), .ZN(n6307) );
  OAI22_X1 U5512 ( .A1(n4500), .A2(n6553), .B1(n4499), .B2(n6307), .ZN(n4476)
         );
  AOI21_X1 U5513 ( .B1(n6556), .B2(n4619), .A(n4476), .ZN(n4477) );
  OAI211_X1 U5514 ( .C1(n4736), .C2(n6559), .A(n4478), .B(n4477), .ZN(U3147)
         );
  NAND2_X1 U5515 ( .A1(n5446), .A2(DATAI_29_), .ZN(n6365) );
  NAND2_X1 U5516 ( .A1(n4495), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4482)
         );
  NAND2_X1 U5517 ( .A1(n5446), .A2(DATAI_21_), .ZN(n6297) );
  INV_X1 U5518 ( .A(n6297), .ZN(n6362) );
  INV_X1 U5519 ( .A(DATAI_5_), .ZN(n4586) );
  NOR2_X1 U5520 ( .A1(n4586), .A2(n4744), .ZN(n6361) );
  INV_X1 U5521 ( .A(n6361), .ZN(n5000) );
  NAND2_X1 U5522 ( .A1(n4498), .A2(n4479), .ZN(n6296) );
  OAI22_X1 U5523 ( .A1(n4500), .A2(n5000), .B1(n4499), .B2(n6296), .ZN(n4480)
         );
  AOI21_X1 U5524 ( .B1(n6362), .B2(n4619), .A(n4480), .ZN(n4481) );
  OAI211_X1 U5525 ( .C1(n4736), .C2(n6365), .A(n4482), .B(n4481), .ZN(U3145)
         );
  NAND2_X1 U5526 ( .A1(n5446), .A2(DATAI_24_), .ZN(n6335) );
  NAND2_X1 U5527 ( .A1(n4495), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4486)
         );
  NAND2_X1 U5528 ( .A1(n5446), .A2(DATAI_16_), .ZN(n6233) );
  INV_X1 U5529 ( .A(n6233), .ZN(n6332) );
  NOR2_X1 U5530 ( .A1(n4483), .A2(n4744), .ZN(n6321) );
  INV_X1 U5531 ( .A(n6321), .ZN(n5004) );
  NAND2_X1 U5532 ( .A1(n4498), .A2(n3187), .ZN(n6215) );
  OAI22_X1 U5533 ( .A1(n4500), .A2(n5004), .B1(n4499), .B2(n6215), .ZN(n4484)
         );
  AOI21_X1 U5534 ( .B1(n6332), .B2(n4619), .A(n4484), .ZN(n4485) );
  OAI211_X1 U5535 ( .C1(n6335), .C2(n4736), .A(n4486), .B(n4485), .ZN(U3140)
         );
  NAND2_X1 U5536 ( .A1(n5446), .A2(DATAI_25_), .ZN(n6341) );
  NAND2_X1 U5537 ( .A1(n4495), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4490)
         );
  NAND2_X1 U5538 ( .A1(n5446), .A2(DATAI_17_), .ZN(n6280) );
  INV_X1 U5539 ( .A(n6280), .ZN(n6338) );
  INV_X1 U5540 ( .A(n4744), .ZN(n4702) );
  INV_X1 U5541 ( .A(n6336), .ZN(n4988) );
  NAND2_X1 U5542 ( .A1(n4498), .A2(n4487), .ZN(n6275) );
  OAI22_X1 U5543 ( .A1(n4500), .A2(n4988), .B1(n4499), .B2(n6275), .ZN(n4488)
         );
  AOI21_X1 U5544 ( .B1(n6338), .B2(n4619), .A(n4488), .ZN(n4489) );
  OAI211_X1 U5545 ( .C1(n4736), .C2(n6341), .A(n4490), .B(n4489), .ZN(U3141)
         );
  NAND2_X1 U5546 ( .A1(n5446), .A2(DATAI_28_), .ZN(n6359) );
  NAND2_X1 U5547 ( .A1(n4495), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4494)
         );
  NAND2_X1 U5548 ( .A1(n5446), .A2(DATAI_20_), .ZN(n6295) );
  INV_X1 U5549 ( .A(n6295), .ZN(n6356) );
  INV_X1 U5550 ( .A(DATAI_4_), .ZN(n6653) );
  NOR2_X1 U5551 ( .A1(n6653), .A2(n4744), .ZN(n6355) );
  INV_X1 U5552 ( .A(n6355), .ZN(n4996) );
  NAND2_X1 U5553 ( .A1(n4498), .A2(n4491), .ZN(n6291) );
  OAI22_X1 U5554 ( .A1(n4500), .A2(n4996), .B1(n4499), .B2(n6291), .ZN(n4492)
         );
  AOI21_X1 U5555 ( .B1(n6356), .B2(n4619), .A(n4492), .ZN(n4493) );
  OAI211_X1 U5556 ( .C1(n4736), .C2(n6359), .A(n4494), .B(n4493), .ZN(U3144)
         );
  NAND2_X1 U5557 ( .A1(n5446), .A2(DATAI_26_), .ZN(n6347) );
  NAND2_X1 U5558 ( .A1(n4495), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4503)
         );
  NAND2_X1 U5559 ( .A1(n5446), .A2(DATAI_18_), .ZN(n6282) );
  INV_X1 U5560 ( .A(n6282), .ZN(n6344) );
  NOR2_X1 U5561 ( .A1(n4496), .A2(n4744), .ZN(n6343) );
  INV_X1 U5562 ( .A(n6343), .ZN(n5016) );
  NAND2_X1 U5563 ( .A1(n4498), .A2(n4497), .ZN(n6281) );
  OAI22_X1 U5564 ( .A1(n4500), .A2(n5016), .B1(n4499), .B2(n6281), .ZN(n4501)
         );
  AOI21_X1 U5565 ( .B1(n6344), .B2(n4619), .A(n4501), .ZN(n4502) );
  OAI211_X1 U5566 ( .C1(n4736), .C2(n6347), .A(n4503), .B(n4502), .ZN(U3142)
         );
  INV_X1 U5567 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5947) );
  OAI222_X1 U5568 ( .A1(n5033), .A2(n5671), .B1(n4782), .B2(n4504), .C1(n5120), 
        .C2(n5947), .ZN(U2888) );
  INV_X1 U5569 ( .A(n4976), .ZN(n4507) );
  INV_X1 U5570 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4970) );
  AOI22_X1 U5571 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6095), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4505) );
  OAI21_X1 U5572 ( .B1(n6015), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4505), 
        .ZN(n4506) );
  AOI21_X1 U5573 ( .B1(n4507), .B2(n5446), .A(n4506), .ZN(n4508) );
  OAI21_X1 U5574 ( .B1(n4509), .B2(n5992), .A(n4508), .ZN(U2985) );
  OAI21_X1 U5575 ( .B1(n4512), .B2(n4511), .A(n4510), .ZN(n6087) );
  AND2_X1 U5576 ( .A1(n6095), .A2(REIP_REG_3__SCAN_IN), .ZN(n6083) );
  AOI21_X1 U5577 ( .B1(n6006), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6083), 
        .ZN(n4513) );
  OAI21_X1 U5578 ( .B1(n6015), .B2(n5022), .A(n4513), .ZN(n4514) );
  AOI21_X1 U5579 ( .B1(n4515), .B2(n5446), .A(n4514), .ZN(n4516) );
  OAI21_X1 U5580 ( .B1(n5992), .B2(n6087), .A(n4516), .ZN(U2983) );
  NOR2_X1 U5581 ( .A1(n4573), .A2(n6322), .ZN(n5630) );
  NAND3_X1 U5582 ( .A1(n6113), .A2(n5630), .A3(n4518), .ZN(n4519) );
  NAND2_X1 U5583 ( .A1(n4519), .A2(n6218), .ZN(n4523) );
  INV_X1 U5584 ( .A(n5624), .ZN(n4532) );
  AND2_X1 U5585 ( .A1(n4315), .A2(n4532), .ZN(n4828) );
  INV_X1 U5586 ( .A(n2956), .ZN(n6382) );
  NOR2_X1 U5587 ( .A1(n4985), .A2(n6111), .ZN(n4520) );
  AOI21_X1 U5588 ( .B1(n4787), .B2(n6382), .A(n4520), .ZN(n4521) );
  NAND2_X1 U5589 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4823), .ZN(n4785) );
  OAI22_X1 U5590 ( .A1(n4523), .A2(n4521), .B1(n4785), .B2(n6414), .ZN(n6310)
         );
  INV_X1 U5591 ( .A(n6310), .ZN(n4530) );
  NOR2_X1 U5592 ( .A1(n6112), .A2(n4573), .ZN(n4825) );
  INV_X1 U5593 ( .A(n6379), .ZN(n4528) );
  NAND3_X1 U5594 ( .A1(n4825), .A2(n6113), .A3(n4977), .ZN(n6308) );
  INV_X1 U5595 ( .A(n4520), .ZN(n6306) );
  OAI22_X1 U5596 ( .A1(n6308), .A2(n6335), .B1(n6215), .B2(n6306), .ZN(n4527)
         );
  INV_X1 U5597 ( .A(n6116), .ZN(n6225) );
  INV_X1 U5598 ( .A(n4521), .ZN(n4522) );
  NOR2_X1 U5599 ( .A1(n4523), .A2(n4522), .ZN(n4524) );
  AOI211_X1 U5600 ( .C1(n4785), .C2(n6325), .A(n6225), .B(n4524), .ZN(n6277)
         );
  INV_X1 U5601 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4525) );
  NOR2_X1 U5602 ( .A1(n6277), .A2(n4525), .ZN(n4526) );
  AOI211_X1 U5603 ( .C1(n4528), .C2(n6332), .A(n4527), .B(n4526), .ZN(n4529)
         );
  OAI21_X1 U5604 ( .B1(n4530), .B2(n5004), .A(n4529), .ZN(U3108) );
  NAND2_X1 U5605 ( .A1(n4537), .A2(n4824), .ZN(n4698) );
  AOI21_X1 U5606 ( .B1(n4537), .B2(STATEBS16_REG_SCAN_IN), .A(n6325), .ZN(
        n4534) );
  NOR2_X1 U5607 ( .A1(n4315), .A2(n4532), .ZN(n6327) );
  NAND3_X1 U5608 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6387), .ZN(n6319) );
  NOR2_X1 U5609 ( .A1(n4660), .A2(n6319), .ZN(n4554) );
  AOI21_X1 U5610 ( .B1(n4662), .B2(n6327), .A(n4554), .ZN(n4536) );
  AOI22_X1 U5611 ( .A1(n4534), .A2(n4536), .B1(n6325), .B2(n6319), .ZN(n4533)
         );
  NAND2_X1 U5612 ( .A1(n6116), .A2(n4533), .ZN(n4553) );
  INV_X1 U5613 ( .A(n4534), .ZN(n4535) );
  OAI22_X1 U5614 ( .A1(n4536), .A2(n4535), .B1(n6414), .B2(n6319), .ZN(n4552)
         );
  AOI22_X1 U5615 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4553), .B1(n6367), 
        .B2(n4552), .ZN(n4539) );
  INV_X1 U5616 ( .A(n6371), .ZN(n6202) );
  INV_X1 U5617 ( .A(n6301), .ZN(n6366) );
  AOI22_X1 U5618 ( .A1(n6375), .A2(n6202), .B1(n6366), .B2(n4554), .ZN(n4538)
         );
  OAI211_X1 U5619 ( .C1(n6305), .C2(n4698), .A(n4539), .B(n4538), .ZN(U3130)
         );
  AOI22_X1 U5620 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4553), .B1(n6321), 
        .B2(n4552), .ZN(n4541) );
  INV_X1 U5621 ( .A(n6335), .ZN(n6178) );
  INV_X1 U5622 ( .A(n6215), .ZN(n6320) );
  AOI22_X1 U5623 ( .A1(n6375), .A2(n6178), .B1(n6320), .B2(n4554), .ZN(n4540)
         );
  OAI211_X1 U5624 ( .C1(n6233), .C2(n4698), .A(n4541), .B(n4540), .ZN(U3124)
         );
  AOI22_X1 U5625 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4553), .B1(n6336), 
        .B2(n4552), .ZN(n4543) );
  INV_X1 U5626 ( .A(n6341), .ZN(n6182) );
  INV_X1 U5627 ( .A(n6275), .ZN(n6337) );
  AOI22_X1 U5628 ( .A1(n6375), .A2(n6182), .B1(n6337), .B2(n4554), .ZN(n4542)
         );
  OAI211_X1 U5629 ( .C1(n6280), .C2(n4698), .A(n4543), .B(n4542), .ZN(U3125)
         );
  AOI22_X1 U5630 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4553), .B1(n6349), 
        .B2(n4552), .ZN(n4545) );
  INV_X1 U5631 ( .A(n6353), .ZN(n6192) );
  INV_X1 U5632 ( .A(n6286), .ZN(n6348) );
  AOI22_X1 U5633 ( .A1(n6375), .A2(n6192), .B1(n6348), .B2(n4554), .ZN(n4544)
         );
  OAI211_X1 U5634 ( .C1(n6290), .C2(n4698), .A(n4545), .B(n4544), .ZN(U3127)
         );
  AOI22_X1 U5635 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4553), .B1(n6355), 
        .B2(n4552), .ZN(n4547) );
  INV_X1 U5636 ( .A(n6359), .ZN(n6131) );
  AOI22_X1 U5637 ( .A1(n6375), .A2(n6131), .B1(n6354), .B2(n4554), .ZN(n4546)
         );
  OAI211_X1 U5638 ( .C1(n6295), .C2(n4698), .A(n4547), .B(n4546), .ZN(U3128)
         );
  AOI22_X1 U5639 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4553), .B1(n6343), 
        .B2(n4552), .ZN(n4549) );
  INV_X1 U5640 ( .A(n6347), .ZN(n6187) );
  AOI22_X1 U5641 ( .A1(n6375), .A2(n6187), .B1(n6342), .B2(n4554), .ZN(n4548)
         );
  OAI211_X1 U5642 ( .C1(n6282), .C2(n4698), .A(n4549), .B(n4548), .ZN(U3126)
         );
  AOI22_X1 U5643 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4553), .B1(n6374), 
        .B2(n4552), .ZN(n4551) );
  INV_X1 U5644 ( .A(n6559), .ZN(n6209) );
  AOI22_X1 U5645 ( .A1(n6375), .A2(n6209), .B1(n6550), .B2(n4554), .ZN(n4550)
         );
  OAI211_X1 U5646 ( .C1(n6314), .C2(n4698), .A(n4551), .B(n4550), .ZN(U3131)
         );
  AOI22_X1 U5647 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4553), .B1(n6361), 
        .B2(n4552), .ZN(n4556) );
  INV_X1 U5648 ( .A(n6365), .ZN(n6197) );
  INV_X1 U5649 ( .A(n6296), .ZN(n6360) );
  AOI22_X1 U5650 ( .A1(n6375), .A2(n6197), .B1(n6360), .B2(n4554), .ZN(n4555)
         );
  OAI211_X1 U5651 ( .C1(n6297), .C2(n4698), .A(n4556), .B(n4555), .ZN(U3129)
         );
  INV_X1 U5652 ( .A(n4559), .ZN(n4560) );
  OAI21_X1 U5653 ( .B1(n4557), .B2(n4561), .A(n4560), .ZN(n4900) );
  INV_X1 U5654 ( .A(n4763), .ZN(n4562) );
  AOI21_X1 U5655 ( .B1(n4563), .B2(n4569), .A(n4562), .ZN(n6068) );
  AOI22_X1 U5656 ( .A1(n6068), .A2(n3996), .B1(EBX_REG_5__SCAN_IN), .B2(n5286), 
        .ZN(n4564) );
  OAI21_X1 U5657 ( .B1(n4900), .B2(n5300), .A(n4564), .ZN(U2854) );
  INV_X1 U5658 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5950) );
  XOR2_X1 U5659 ( .A(n4450), .B(n4565), .Z(n6002) );
  INV_X1 U5660 ( .A(n6002), .ZN(n4570) );
  OAI222_X1 U5661 ( .A1(n5120), .A2(n5950), .B1(n4782), .B2(n6653), .C1(n5671), 
        .C2(n4570), .ZN(U2887) );
  OR2_X1 U5662 ( .A1(n4567), .A2(n4566), .ZN(n4568) );
  NAND2_X1 U5663 ( .A1(n4569), .A2(n4568), .ZN(n6078) );
  INV_X1 U5664 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4571) );
  OAI222_X1 U5665 ( .A1(n6078), .A2(n5872), .B1(n4571), .B2(n5878), .C1(n5300), 
        .C2(n4570), .ZN(U2855) );
  AOI21_X1 U5666 ( .B1(n4580), .B2(STATEBS16_REG_SCAN_IN), .A(n6325), .ZN(
        n6150) );
  NAND2_X1 U5667 ( .A1(n6327), .A2(n4574), .ZN(n6149) );
  OR2_X1 U5668 ( .A1(n6149), .A2(n2956), .ZN(n4575) );
  NAND3_X1 U5669 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n4985), .A3(n6387), .ZN(n6147) );
  NOR2_X1 U5670 ( .A1(n4660), .A2(n6147), .ZN(n4581) );
  INV_X1 U5671 ( .A(n4581), .ZN(n6206) );
  INV_X1 U5672 ( .A(n6147), .ZN(n4576) );
  OAI21_X1 U5673 ( .B1(n6218), .B2(n4576), .A(n6116), .ZN(n4577) );
  AOI21_X1 U5674 ( .B1(n6150), .B2(n4578), .A(n4577), .ZN(n6214) );
  INV_X1 U5675 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4585) );
  INV_X1 U5676 ( .A(n6150), .ZN(n4579) );
  OAI22_X1 U5677 ( .A1(n4579), .A2(n4578), .B1(n6147), .B2(n6414), .ZN(n6210)
         );
  AOI22_X1 U5678 ( .A1(n6208), .A2(n6131), .B1(n6354), .B2(n4581), .ZN(n4582)
         );
  OAI21_X1 U5679 ( .B1(n6295), .B2(n6558), .A(n4582), .ZN(n4583) );
  AOI21_X1 U5680 ( .B1(n6210), .B2(n6355), .A(n4583), .ZN(n4584) );
  OAI21_X1 U5681 ( .B1(n6214), .B2(n4585), .A(n4584), .ZN(U3064) );
  INV_X1 U5682 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5908) );
  OAI222_X1 U5683 ( .A1(n4900), .A2(n5671), .B1(n4782), .B2(n4586), .C1(n5120), 
        .C2(n5908), .ZN(U2886) );
  NOR2_X1 U5684 ( .A1(n6112), .A2(n5622), .ZN(n4659) );
  NAND2_X1 U5685 ( .A1(n6110), .A2(n4659), .ZN(n4629) );
  INV_X1 U5686 ( .A(n4658), .ZN(n4587) );
  OAI21_X1 U5687 ( .B1(n4587), .B2(n4619), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4588) );
  NAND2_X1 U5688 ( .A1(n4315), .A2(n5624), .ZN(n4740) );
  INV_X1 U5689 ( .A(n4740), .ZN(n4661) );
  NAND2_X1 U5690 ( .A1(n6317), .A2(n4661), .ZN(n4592) );
  NAND3_X1 U5691 ( .A1(n4588), .A2(n6218), .A3(n4592), .ZN(n4591) );
  NAND3_X1 U5692 ( .A1(n4985), .A2(n6391), .A3(n6387), .ZN(n4626) );
  OR2_X1 U5693 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4626), .ZN(n4616)
         );
  NOR2_X1 U5694 ( .A1(n4593), .A2(n6414), .ZN(n4786) );
  INV_X1 U5695 ( .A(n4589), .ZN(n4743) );
  INV_X1 U5696 ( .A(n4979), .ZN(n4833) );
  NOR2_X1 U5697 ( .A1(n4743), .A2(n4833), .ZN(n6144) );
  OAI21_X1 U5698 ( .B1(n6144), .B2(n6414), .A(n4702), .ZN(n6153) );
  AOI211_X1 U5699 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4616), .A(n4786), .B(
        n6153), .ZN(n4590) );
  NAND2_X1 U5700 ( .A1(n4591), .A2(n4590), .ZN(n4615) );
  NAND2_X1 U5701 ( .A1(n4615), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4596) );
  INV_X1 U5702 ( .A(n4592), .ZN(n4622) );
  AND2_X1 U5703 ( .A1(n4593), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6152) );
  AOI22_X1 U5704 ( .A1(n4622), .A2(n6218), .B1(n6152), .B2(n6144), .ZN(n4617)
         );
  OAI22_X1 U5705 ( .A1(n5000), .A2(n4617), .B1(n6296), .B2(n4616), .ZN(n4594)
         );
  AOI21_X1 U5706 ( .B1(n6197), .B2(n4619), .A(n4594), .ZN(n4595) );
  OAI211_X1 U5707 ( .C1(n4658), .C2(n6297), .A(n4596), .B(n4595), .ZN(U3025)
         );
  NAND2_X1 U5708 ( .A1(n4615), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4599) );
  OAI22_X1 U5709 ( .A1(n5012), .A2(n4617), .B1(n6301), .B2(n4616), .ZN(n4597)
         );
  AOI21_X1 U5710 ( .B1(n6202), .B2(n4619), .A(n4597), .ZN(n4598) );
  OAI211_X1 U5711 ( .C1(n4658), .C2(n6305), .A(n4599), .B(n4598), .ZN(U3026)
         );
  NAND2_X1 U5712 ( .A1(n4615), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4602) );
  OAI22_X1 U5713 ( .A1(n6275), .A2(n4616), .B1(n4617), .B2(n4988), .ZN(n4600)
         );
  AOI21_X1 U5714 ( .B1(n4619), .B2(n6182), .A(n4600), .ZN(n4601) );
  OAI211_X1 U5715 ( .C1(n4658), .C2(n6280), .A(n4602), .B(n4601), .ZN(U3021)
         );
  NAND2_X1 U5716 ( .A1(n4615), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4605) );
  OAI22_X1 U5717 ( .A1(n5016), .A2(n4617), .B1(n6281), .B2(n4616), .ZN(n4603)
         );
  AOI21_X1 U5718 ( .B1(n6187), .B2(n4619), .A(n4603), .ZN(n4604) );
  OAI211_X1 U5719 ( .C1(n4658), .C2(n6282), .A(n4605), .B(n4604), .ZN(U3022)
         );
  NAND2_X1 U5720 ( .A1(n4615), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4608) );
  OAI22_X1 U5721 ( .A1(n5004), .A2(n4617), .B1(n6215), .B2(n4616), .ZN(n4606)
         );
  AOI21_X1 U5722 ( .B1(n6178), .B2(n4619), .A(n4606), .ZN(n4607) );
  OAI211_X1 U5723 ( .C1(n4658), .C2(n6233), .A(n4608), .B(n4607), .ZN(U3020)
         );
  NAND2_X1 U5724 ( .A1(n4615), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4611) );
  OAI22_X1 U5725 ( .A1(n4996), .A2(n4617), .B1(n6291), .B2(n4616), .ZN(n4609)
         );
  AOI21_X1 U5726 ( .B1(n6131), .B2(n4619), .A(n4609), .ZN(n4610) );
  OAI211_X1 U5727 ( .C1(n4658), .C2(n6295), .A(n4611), .B(n4610), .ZN(U3024)
         );
  NAND2_X1 U5728 ( .A1(n4615), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4614) );
  OAI22_X1 U5729 ( .A1(n5008), .A2(n4617), .B1(n6286), .B2(n4616), .ZN(n4612)
         );
  AOI21_X1 U5730 ( .B1(n6192), .B2(n4619), .A(n4612), .ZN(n4613) );
  OAI211_X1 U5731 ( .C1(n4658), .C2(n6290), .A(n4614), .B(n4613), .ZN(U3023)
         );
  NAND2_X1 U5732 ( .A1(n4615), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4621) );
  OAI22_X1 U5733 ( .A1(n6553), .A2(n4617), .B1(n6307), .B2(n4616), .ZN(n4618)
         );
  AOI21_X1 U5734 ( .B1(n6209), .B2(n4619), .A(n4618), .ZN(n4620) );
  OAI211_X1 U5735 ( .C1(n4658), .C2(n6314), .A(n4621), .B(n4620), .ZN(U3027)
         );
  NOR2_X1 U5736 ( .A1(n4660), .A2(n4626), .ZN(n4630) );
  AOI21_X1 U5737 ( .B1(n4622), .B2(n6382), .A(n4630), .ZN(n4628) );
  OR2_X1 U5738 ( .A1(n4629), .A2(n6322), .ZN(n4623) );
  AOI22_X1 U5739 ( .A1(n4628), .A2(n4625), .B1(n6325), .B2(n4626), .ZN(n4624)
         );
  NAND2_X1 U5740 ( .A1(n6116), .A2(n4624), .ZN(n4653) );
  INV_X1 U5741 ( .A(n4625), .ZN(n4627) );
  OAI22_X1 U5742 ( .A1(n4628), .A2(n4627), .B1(n6414), .B2(n4626), .ZN(n4652)
         );
  AOI22_X1 U5743 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4653), .B1(n6336), 
        .B2(n4652), .ZN(n4633) );
  INV_X1 U5744 ( .A(n4630), .ZN(n4654) );
  OAI22_X1 U5745 ( .A1(n4864), .A2(n6280), .B1(n6275), .B2(n4654), .ZN(n4631)
         );
  INV_X1 U5746 ( .A(n4631), .ZN(n4632) );
  OAI211_X1 U5747 ( .C1(n6341), .C2(n4658), .A(n4633), .B(n4632), .ZN(U3029)
         );
  AOI22_X1 U5748 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4653), .B1(n6355), 
        .B2(n4652), .ZN(n4636) );
  OAI22_X1 U5749 ( .A1(n4864), .A2(n6295), .B1(n6291), .B2(n4654), .ZN(n4634)
         );
  INV_X1 U5750 ( .A(n4634), .ZN(n4635) );
  OAI211_X1 U5751 ( .C1(n6359), .C2(n4658), .A(n4636), .B(n4635), .ZN(U3032)
         );
  AOI22_X1 U5752 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4653), .B1(n6361), 
        .B2(n4652), .ZN(n4639) );
  OAI22_X1 U5753 ( .A1(n4864), .A2(n6297), .B1(n6296), .B2(n4654), .ZN(n4637)
         );
  INV_X1 U5754 ( .A(n4637), .ZN(n4638) );
  OAI211_X1 U5755 ( .C1(n6365), .C2(n4658), .A(n4639), .B(n4638), .ZN(U3033)
         );
  AOI22_X1 U5756 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4653), .B1(n6367), 
        .B2(n4652), .ZN(n4642) );
  OAI22_X1 U5757 ( .A1(n4864), .A2(n6305), .B1(n6301), .B2(n4654), .ZN(n4640)
         );
  INV_X1 U5758 ( .A(n4640), .ZN(n4641) );
  OAI211_X1 U5759 ( .C1(n6371), .C2(n4658), .A(n4642), .B(n4641), .ZN(U3034)
         );
  AOI22_X1 U5760 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4653), .B1(n6321), 
        .B2(n4652), .ZN(n4645) );
  OAI22_X1 U5761 ( .A1(n4864), .A2(n6233), .B1(n6215), .B2(n4654), .ZN(n4643)
         );
  INV_X1 U5762 ( .A(n4643), .ZN(n4644) );
  OAI211_X1 U5763 ( .C1(n6335), .C2(n4658), .A(n4645), .B(n4644), .ZN(U3028)
         );
  AOI22_X1 U5764 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4653), .B1(n6374), 
        .B2(n4652), .ZN(n4648) );
  OAI22_X1 U5765 ( .A1(n4864), .A2(n6314), .B1(n6307), .B2(n4654), .ZN(n4646)
         );
  INV_X1 U5766 ( .A(n4646), .ZN(n4647) );
  OAI211_X1 U5767 ( .C1(n6559), .C2(n4658), .A(n4648), .B(n4647), .ZN(U3035)
         );
  AOI22_X1 U5768 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4653), .B1(n6349), 
        .B2(n4652), .ZN(n4651) );
  OAI22_X1 U5769 ( .A1(n4864), .A2(n6290), .B1(n6286), .B2(n4654), .ZN(n4649)
         );
  INV_X1 U5770 ( .A(n4649), .ZN(n4650) );
  OAI211_X1 U5771 ( .C1(n6353), .C2(n4658), .A(n4651), .B(n4650), .ZN(U3031)
         );
  AOI22_X1 U5772 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4653), .B1(n6343), 
        .B2(n4652), .ZN(n4657) );
  OAI22_X1 U5773 ( .A1(n4864), .A2(n6282), .B1(n6281), .B2(n4654), .ZN(n4655)
         );
  INV_X1 U5774 ( .A(n4655), .ZN(n4656) );
  OAI211_X1 U5775 ( .C1(n6347), .C2(n4658), .A(n4657), .B(n4656), .ZN(U3030)
         );
  NAND2_X1 U5776 ( .A1(n4659), .A2(n6113), .ZN(n4668) );
  NAND3_X1 U5777 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6391), .A3(n6387), .ZN(n4742) );
  NOR2_X1 U5778 ( .A1(n4660), .A2(n4742), .ZN(n4685) );
  AOI21_X1 U5779 ( .B1(n4662), .B2(n4661), .A(n4685), .ZN(n4667) );
  OR2_X1 U5780 ( .A1(n4668), .A2(n6322), .ZN(n4663) );
  AOI22_X1 U5781 ( .A1(n4667), .A2(n4665), .B1(n6325), .B2(n4742), .ZN(n4664)
         );
  NAND2_X1 U5782 ( .A1(n6116), .A2(n4664), .ZN(n4684) );
  INV_X1 U5783 ( .A(n4665), .ZN(n4666) );
  OAI22_X1 U5784 ( .A1(n4667), .A2(n4666), .B1(n6414), .B2(n4742), .ZN(n4683)
         );
  AOI22_X1 U5785 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4684), .B1(n6336), 
        .B2(n4683), .ZN(n4670) );
  NOR2_X2 U5786 ( .A1(n4668), .A2(n4824), .ZN(n6270) );
  AOI22_X1 U5787 ( .A1(n6270), .A2(n6182), .B1(n6337), .B2(n4685), .ZN(n4669)
         );
  OAI211_X1 U5788 ( .C1(n4688), .C2(n6280), .A(n4670), .B(n4669), .ZN(U3093)
         );
  AOI22_X1 U5789 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4684), .B1(n6361), 
        .B2(n4683), .ZN(n4672) );
  AOI22_X1 U5790 ( .A1(n6270), .A2(n6197), .B1(n6360), .B2(n4685), .ZN(n4671)
         );
  OAI211_X1 U5791 ( .C1(n4688), .C2(n6297), .A(n4672), .B(n4671), .ZN(U3097)
         );
  AOI22_X1 U5792 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4684), .B1(n6349), 
        .B2(n4683), .ZN(n4674) );
  AOI22_X1 U5793 ( .A1(n6270), .A2(n6192), .B1(n6348), .B2(n4685), .ZN(n4673)
         );
  OAI211_X1 U5794 ( .C1(n4688), .C2(n6290), .A(n4674), .B(n4673), .ZN(U3095)
         );
  AOI22_X1 U5795 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4684), .B1(n6367), 
        .B2(n4683), .ZN(n4676) );
  AOI22_X1 U5796 ( .A1(n6270), .A2(n6202), .B1(n6366), .B2(n4685), .ZN(n4675)
         );
  OAI211_X1 U5797 ( .C1(n4688), .C2(n6305), .A(n4676), .B(n4675), .ZN(U3098)
         );
  AOI22_X1 U5798 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4684), .B1(n6355), 
        .B2(n4683), .ZN(n4678) );
  AOI22_X1 U5799 ( .A1(n6270), .A2(n6131), .B1(n6354), .B2(n4685), .ZN(n4677)
         );
  OAI211_X1 U5800 ( .C1(n4688), .C2(n6295), .A(n4678), .B(n4677), .ZN(U3096)
         );
  AOI22_X1 U5801 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4684), .B1(n6343), 
        .B2(n4683), .ZN(n4680) );
  AOI22_X1 U5802 ( .A1(n6270), .A2(n6187), .B1(n6342), .B2(n4685), .ZN(n4679)
         );
  OAI211_X1 U5803 ( .C1(n4688), .C2(n6282), .A(n4680), .B(n4679), .ZN(U3094)
         );
  AOI22_X1 U5804 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4684), .B1(n6321), 
        .B2(n4683), .ZN(n4682) );
  AOI22_X1 U5805 ( .A1(n6270), .A2(n6178), .B1(n6320), .B2(n4685), .ZN(n4681)
         );
  OAI211_X1 U5806 ( .C1(n4688), .C2(n6233), .A(n4682), .B(n4681), .ZN(U3092)
         );
  AOI22_X1 U5807 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4684), .B1(n6374), 
        .B2(n4683), .ZN(n4687) );
  AOI22_X1 U5808 ( .A1(n6270), .A2(n6209), .B1(n6550), .B2(n4685), .ZN(n4686)
         );
  OAI211_X1 U5809 ( .C1(n4688), .C2(n6314), .A(n4687), .B(n4686), .ZN(U3099)
         );
  INV_X1 U5810 ( .A(n4689), .ZN(n4690) );
  XOR2_X1 U5811 ( .A(n4690), .B(n4692), .Z(n4923) );
  INV_X1 U5812 ( .A(n4923), .ZN(n4738) );
  INV_X1 U5813 ( .A(n4693), .ZN(n4695) );
  INV_X1 U5814 ( .A(n4764), .ZN(n4694) );
  AOI21_X1 U5815 ( .B1(n4695), .B2(n4694), .A(n5819), .ZN(n6059) );
  AOI22_X1 U5816 ( .A1(n6059), .A2(n3996), .B1(EBX_REG_7__SCAN_IN), .B2(n5286), 
        .ZN(n4696) );
  OAI21_X1 U5817 ( .B1(n4738), .B2(n5300), .A(n4696), .ZN(U2852) );
  NOR2_X1 U5818 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4697), .ZN(n4707)
         );
  INV_X1 U5819 ( .A(n6224), .ZN(n4705) );
  INV_X1 U5820 ( .A(n4736), .ZN(n4699) );
  OAI21_X1 U5821 ( .B1(n4733), .B2(n4699), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4700) );
  NAND3_X1 U5822 ( .A1(n4705), .A2(n6218), .A3(n4700), .ZN(n4704) );
  NAND2_X1 U5823 ( .A1(n4979), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U5824 ( .A1(n4702), .A2(n4701), .ZN(n4983) );
  NOR3_X1 U5825 ( .A1(n4983), .A2(n4985), .A3(n6152), .ZN(n4703) );
  OAI211_X1 U5826 ( .C1(n4707), .C2(n6512), .A(n4704), .B(n4703), .ZN(n4729)
         );
  NAND2_X1 U5827 ( .A1(n4729), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4710)
         );
  NOR2_X1 U5828 ( .A1(n4705), .A2(n6325), .ZN(n4981) );
  INV_X1 U5829 ( .A(n4786), .ZN(n6316) );
  NOR3_X1 U5830 ( .A1(n6316), .A2(n4979), .A3(n4985), .ZN(n4706) );
  AOI21_X1 U5831 ( .B1(n4981), .B2(n6146), .A(n4706), .ZN(n4731) );
  INV_X1 U5832 ( .A(n4707), .ZN(n4730) );
  OAI22_X1 U5833 ( .A1(n5012), .A2(n4731), .B1(n6301), .B2(n4730), .ZN(n4708)
         );
  AOI21_X1 U5834 ( .B1(n4733), .B2(n6202), .A(n4708), .ZN(n4709) );
  OAI211_X1 U5835 ( .C1(n4736), .C2(n6305), .A(n4710), .B(n4709), .ZN(U3138)
         );
  NAND2_X1 U5836 ( .A1(n4729), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4713)
         );
  OAI22_X1 U5837 ( .A1(n5000), .A2(n4731), .B1(n6296), .B2(n4730), .ZN(n4711)
         );
  AOI21_X1 U5838 ( .B1(n4733), .B2(n6197), .A(n4711), .ZN(n4712) );
  OAI211_X1 U5839 ( .C1(n4736), .C2(n6297), .A(n4713), .B(n4712), .ZN(U3137)
         );
  NAND2_X1 U5840 ( .A1(n4729), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4716)
         );
  OAI22_X1 U5841 ( .A1(n4996), .A2(n4731), .B1(n6291), .B2(n4730), .ZN(n4714)
         );
  AOI21_X1 U5842 ( .B1(n4733), .B2(n6131), .A(n4714), .ZN(n4715) );
  OAI211_X1 U5843 ( .C1(n4736), .C2(n6295), .A(n4716), .B(n4715), .ZN(U3136)
         );
  NAND2_X1 U5844 ( .A1(n4729), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4719)
         );
  OAI22_X1 U5845 ( .A1(n5008), .A2(n4731), .B1(n6286), .B2(n4730), .ZN(n4717)
         );
  AOI21_X1 U5846 ( .B1(n4733), .B2(n6192), .A(n4717), .ZN(n4718) );
  OAI211_X1 U5847 ( .C1(n4736), .C2(n6290), .A(n4719), .B(n4718), .ZN(U3135)
         );
  NAND2_X1 U5848 ( .A1(n4729), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4722)
         );
  OAI22_X1 U5849 ( .A1(n5016), .A2(n4731), .B1(n6281), .B2(n4730), .ZN(n4720)
         );
  AOI21_X1 U5850 ( .B1(n4733), .B2(n6187), .A(n4720), .ZN(n4721) );
  OAI211_X1 U5851 ( .C1(n4736), .C2(n6282), .A(n4722), .B(n4721), .ZN(U3134)
         );
  NAND2_X1 U5852 ( .A1(n4729), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4725)
         );
  OAI22_X1 U5853 ( .A1(n4731), .A2(n4988), .B1(n6275), .B2(n4730), .ZN(n4723)
         );
  AOI21_X1 U5854 ( .B1(n4733), .B2(n6182), .A(n4723), .ZN(n4724) );
  OAI211_X1 U5855 ( .C1(n4736), .C2(n6280), .A(n4725), .B(n4724), .ZN(U3133)
         );
  NAND2_X1 U5856 ( .A1(n4729), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4728)
         );
  OAI22_X1 U5857 ( .A1(n5004), .A2(n4731), .B1(n6215), .B2(n4730), .ZN(n4726)
         );
  AOI21_X1 U5858 ( .B1(n4733), .B2(n6178), .A(n4726), .ZN(n4727) );
  OAI211_X1 U5859 ( .C1(n4736), .C2(n6233), .A(n4728), .B(n4727), .ZN(U3132)
         );
  NAND2_X1 U5860 ( .A1(n4729), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4735)
         );
  OAI22_X1 U5861 ( .A1(n6553), .A2(n4731), .B1(n6307), .B2(n4730), .ZN(n4732)
         );
  AOI21_X1 U5862 ( .B1(n4733), .B2(n6209), .A(n4732), .ZN(n4734) );
  OAI211_X1 U5863 ( .C1(n4736), .C2(n6314), .A(n4735), .B(n4734), .ZN(U3139)
         );
  OAI222_X1 U5864 ( .A1(n5671), .A2(n4738), .B1(n4782), .B2(n4737), .C1(n5120), 
        .C2(n3456), .ZN(U2884) );
  INV_X1 U5865 ( .A(n6270), .ZN(n4760) );
  AND2_X1 U5866 ( .A1(n5622), .A2(n4824), .ZN(n4739) );
  AOI21_X1 U5867 ( .B1(n4760), .B2(n6274), .A(n6322), .ZN(n4741) );
  NOR2_X1 U5868 ( .A1(n6317), .A2(n4740), .ZN(n4748) );
  NOR3_X1 U5869 ( .A1(n4741), .A2(n4748), .A3(n6325), .ZN(n4746) );
  NOR2_X1 U5870 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4742), .ZN(n6268)
         );
  NAND2_X1 U5871 ( .A1(n4743), .A2(n4979), .ZN(n6315) );
  AOI21_X1 U5872 ( .B1(n6315), .B2(STATE2_REG_2__SCAN_IN), .A(n4744), .ZN(
        n6328) );
  OAI211_X1 U5873 ( .C1(n6512), .C2(n6268), .A(n6316), .B(n6328), .ZN(n4745)
         );
  NAND2_X1 U5874 ( .A1(n6271), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4751) );
  INV_X1 U5875 ( .A(n6274), .ZN(n4757) );
  INV_X1 U5876 ( .A(n6315), .ZN(n4747) );
  AOI22_X1 U5877 ( .A1(n4748), .A2(n6218), .B1(n6152), .B2(n4747), .ZN(n6259)
         );
  INV_X1 U5878 ( .A(n6268), .ZN(n4755) );
  OAI22_X1 U5879 ( .A1(n5004), .A2(n6259), .B1(n6215), .B2(n4755), .ZN(n4749)
         );
  AOI21_X1 U5880 ( .B1(n6178), .B2(n4757), .A(n4749), .ZN(n4750) );
  OAI211_X1 U5881 ( .C1(n4760), .C2(n6233), .A(n4751), .B(n4750), .ZN(U3084)
         );
  NAND2_X1 U5882 ( .A1(n6271), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4754) );
  OAI22_X1 U5883 ( .A1(n5008), .A2(n6259), .B1(n6286), .B2(n4755), .ZN(n4752)
         );
  AOI21_X1 U5884 ( .B1(n6192), .B2(n4757), .A(n4752), .ZN(n4753) );
  OAI211_X1 U5885 ( .C1(n4760), .C2(n6290), .A(n4754), .B(n4753), .ZN(U3087)
         );
  NAND2_X1 U5886 ( .A1(n6271), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4759) );
  OAI22_X1 U5887 ( .A1(n5012), .A2(n6259), .B1(n6301), .B2(n4755), .ZN(n4756)
         );
  AOI21_X1 U5888 ( .B1(n6202), .B2(n4757), .A(n4756), .ZN(n4758) );
  OAI211_X1 U5889 ( .C1(n4760), .C2(n6305), .A(n4759), .B(n4758), .ZN(U3090)
         );
  XOR2_X1 U5890 ( .A(n4761), .B(n4559), .Z(n5993) );
  AND2_X1 U5891 ( .A1(n4763), .A2(n4762), .ZN(n4765) );
  OR2_X1 U5892 ( .A1(n4765), .A2(n4764), .ZN(n5833) );
  OAI22_X1 U5893 ( .A1(n5833), .A2(n5872), .B1(n5834), .B2(n5878), .ZN(n4766)
         );
  AOI21_X1 U5894 ( .B1(n5993), .B2(n3900), .A(n4766), .ZN(n4767) );
  INV_X1 U5895 ( .A(n4767), .ZN(U2853) );
  INV_X1 U5896 ( .A(n5993), .ZN(n4769) );
  INV_X1 U5897 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5953) );
  OAI222_X1 U5898 ( .A1(n5671), .A2(n4769), .B1(n4782), .B2(n4768), .C1(n5120), 
        .C2(n5953), .ZN(U2885) );
  OAI21_X1 U5899 ( .B1(n4772), .B2(n4771), .A(n4770), .ZN(n6067) );
  OAI22_X1 U5900 ( .A1(n5461), .A2(n4773), .B1(n6032), .B2(n6458), .ZN(n4775)
         );
  NOR2_X1 U5901 ( .A1(n4900), .A2(n5987), .ZN(n4774) );
  AOI211_X1 U5902 ( .C1(n5464), .C2(n4898), .A(n4775), .B(n4774), .ZN(n4776)
         );
  OAI21_X1 U5903 ( .B1(n5992), .B2(n6067), .A(n4776), .ZN(U2981) );
  AOI21_X1 U5904 ( .B1(n4780), .B2(n4777), .A(n4779), .ZN(n4966) );
  INV_X1 U5905 ( .A(n4966), .ZN(n4950) );
  XNOR2_X1 U5906 ( .A(n5819), .B(n5817), .ZN(n6051) );
  AOI22_X1 U5907 ( .A1(n6051), .A2(n3996), .B1(EBX_REG_8__SCAN_IN), .B2(n5286), 
        .ZN(n4781) );
  OAI21_X1 U5908 ( .B1(n4950), .B2(n5300), .A(n4781), .ZN(U2851) );
  INV_X1 U5909 ( .A(DATAI_8_), .ZN(n6592) );
  INV_X1 U5910 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6641) );
  OAI222_X1 U5911 ( .A1(n4950), .A2(n5671), .B1(n4782), .B2(n6592), .C1(n5120), 
        .C2(n6641), .ZN(U2883) );
  NAND2_X1 U5912 ( .A1(n6308), .A2(n6218), .ZN(n4783) );
  OAI21_X1 U5913 ( .B1(n4816), .B2(n4783), .A(n6148), .ZN(n4789) );
  INV_X1 U5914 ( .A(n6152), .ZN(n6329) );
  NOR3_X1 U5915 ( .A1(n6329), .A2(n4979), .A3(n4985), .ZN(n4784) );
  AOI21_X1 U5916 ( .B1(n4789), .B2(n4787), .A(n4784), .ZN(n4819) );
  NOR2_X1 U5917 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4785), .ZN(n4791)
         );
  NOR2_X1 U5918 ( .A1(n4786), .A2(n4983), .ZN(n4831) );
  INV_X1 U5919 ( .A(n4787), .ZN(n4788) );
  AOI22_X1 U5920 ( .A1(n4789), .A2(n4788), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4985), .ZN(n4790) );
  OAI211_X1 U5921 ( .C1(n4791), .C2(n6512), .A(n4831), .B(n4790), .ZN(n4813)
         );
  NAND2_X1 U5922 ( .A1(n4813), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4794)
         );
  INV_X1 U5923 ( .A(n4791), .ZN(n4814) );
  OAI22_X1 U5924 ( .A1(n6308), .A2(n6295), .B1(n4814), .B2(n6291), .ZN(n4792)
         );
  AOI21_X1 U5925 ( .B1(n4816), .B2(n6131), .A(n4792), .ZN(n4793) );
  OAI211_X1 U5926 ( .C1(n4819), .C2(n4996), .A(n4794), .B(n4793), .ZN(U3104)
         );
  NAND2_X1 U5927 ( .A1(n4813), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4797)
         );
  OAI22_X1 U5928 ( .A1(n6308), .A2(n6282), .B1(n4814), .B2(n6281), .ZN(n4795)
         );
  AOI21_X1 U5929 ( .B1(n4816), .B2(n6187), .A(n4795), .ZN(n4796) );
  OAI211_X1 U5930 ( .C1(n4819), .C2(n5016), .A(n4797), .B(n4796), .ZN(U3102)
         );
  NAND2_X1 U5931 ( .A1(n4813), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4800)
         );
  OAI22_X1 U5932 ( .A1(n6308), .A2(n6297), .B1(n4814), .B2(n6296), .ZN(n4798)
         );
  AOI21_X1 U5933 ( .B1(n4816), .B2(n6197), .A(n4798), .ZN(n4799) );
  OAI211_X1 U5934 ( .C1(n4819), .C2(n5000), .A(n4800), .B(n4799), .ZN(U3105)
         );
  NAND2_X1 U5935 ( .A1(n4813), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4803)
         );
  OAI22_X1 U5936 ( .A1(n6308), .A2(n6280), .B1(n4814), .B2(n6275), .ZN(n4801)
         );
  AOI21_X1 U5937 ( .B1(n4816), .B2(n6182), .A(n4801), .ZN(n4802) );
  OAI211_X1 U5938 ( .C1(n4819), .C2(n4988), .A(n4803), .B(n4802), .ZN(U3101)
         );
  NAND2_X1 U5939 ( .A1(n4813), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4806)
         );
  OAI22_X1 U5940 ( .A1(n6308), .A2(n6290), .B1(n4814), .B2(n6286), .ZN(n4804)
         );
  AOI21_X1 U5941 ( .B1(n4816), .B2(n6192), .A(n4804), .ZN(n4805) );
  OAI211_X1 U5942 ( .C1(n4819), .C2(n5008), .A(n4806), .B(n4805), .ZN(U3103)
         );
  NAND2_X1 U5943 ( .A1(n4813), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4809)
         );
  OAI22_X1 U5944 ( .A1(n6308), .A2(n6314), .B1(n4814), .B2(n6307), .ZN(n4807)
         );
  AOI21_X1 U5945 ( .B1(n4816), .B2(n6209), .A(n4807), .ZN(n4808) );
  OAI211_X1 U5946 ( .C1(n4819), .C2(n6553), .A(n4809), .B(n4808), .ZN(U3107)
         );
  NAND2_X1 U5947 ( .A1(n4813), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4812)
         );
  OAI22_X1 U5948 ( .A1(n6308), .A2(n6305), .B1(n4814), .B2(n6301), .ZN(n4810)
         );
  AOI21_X1 U5949 ( .B1(n4816), .B2(n6202), .A(n4810), .ZN(n4811) );
  OAI211_X1 U5950 ( .C1(n4819), .C2(n5012), .A(n4812), .B(n4811), .ZN(U3106)
         );
  NAND2_X1 U5951 ( .A1(n4813), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4818)
         );
  OAI22_X1 U5952 ( .A1(n6308), .A2(n6233), .B1(n6215), .B2(n4814), .ZN(n4815)
         );
  AOI21_X1 U5953 ( .B1(n4816), .B2(n6178), .A(n4815), .ZN(n4817) );
  OAI211_X1 U5954 ( .C1(n4819), .C2(n5004), .A(n4818), .B(n4817), .ZN(U3100)
         );
  INV_X1 U5955 ( .A(n4821), .ZN(n4927) );
  OAI21_X1 U5956 ( .B1(n4779), .B2(n3492), .A(n4927), .ZN(n5815) );
  AOI22_X1 U5957 ( .A1(n5322), .A2(DATAI_9_), .B1(n5885), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4822) );
  OAI21_X1 U5958 ( .B1(n5815), .B2(n5671), .A(n4822), .ZN(U2882) );
  NAND2_X1 U5959 ( .A1(n4823), .A2(n4985), .ZN(n6120) );
  NOR2_X1 U5960 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6120), .ZN(n4865)
         );
  INV_X1 U5961 ( .A(n4864), .ZN(n4827) );
  NOR2_X1 U5962 ( .A1(n6113), .A2(n4824), .ZN(n4826) );
  NAND2_X1 U5963 ( .A1(n4826), .A2(n4825), .ZN(n4868) );
  OAI21_X1 U5964 ( .B1(n4827), .B2(n6139), .A(n6148), .ZN(n4830) );
  AND2_X1 U5965 ( .A1(n6317), .A2(n4828), .ZN(n6115) );
  INV_X1 U5966 ( .A(n6115), .ZN(n4829) );
  AOI21_X1 U5967 ( .B1(n4830), .B2(n4829), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4832) );
  OAI21_X1 U5968 ( .B1(n4865), .B2(n4832), .A(n4831), .ZN(n4871) );
  NOR2_X1 U5969 ( .A1(n4864), .A2(n6371), .ZN(n4838) );
  NAND2_X1 U5970 ( .A1(n6115), .A2(n6218), .ZN(n4835) );
  NAND3_X1 U5971 ( .A1(n6152), .A2(n4833), .A3(n4985), .ZN(n4834) );
  NAND2_X1 U5972 ( .A1(n4835), .A2(n4834), .ZN(n4866) );
  AOI22_X1 U5973 ( .A1(n6367), .A2(n4866), .B1(n6366), .B2(n4865), .ZN(n4836)
         );
  OAI21_X1 U5974 ( .B1(n4868), .B2(n6305), .A(n4836), .ZN(n4837) );
  AOI211_X1 U5975 ( .C1(n4871), .C2(INSTQUEUE_REG_2__6__SCAN_IN), .A(n4838), 
        .B(n4837), .ZN(n4839) );
  INV_X1 U5976 ( .A(n4839), .ZN(U3042) );
  NOR2_X1 U5977 ( .A1(n4864), .A2(n6341), .ZN(n4842) );
  AOI22_X1 U5978 ( .A1(n6337), .A2(n4865), .B1(n6336), .B2(n4866), .ZN(n4840)
         );
  OAI21_X1 U5979 ( .B1(n4868), .B2(n6280), .A(n4840), .ZN(n4841) );
  AOI211_X1 U5980 ( .C1(n4871), .C2(INSTQUEUE_REG_2__1__SCAN_IN), .A(n4842), 
        .B(n4841), .ZN(n4843) );
  INV_X1 U5981 ( .A(n4843), .ZN(U3037) );
  NOR2_X1 U5982 ( .A1(n4864), .A2(n6347), .ZN(n4846) );
  AOI22_X1 U5983 ( .A1(n6343), .A2(n4866), .B1(n6342), .B2(n4865), .ZN(n4844)
         );
  OAI21_X1 U5984 ( .B1(n4868), .B2(n6282), .A(n4844), .ZN(n4845) );
  AOI211_X1 U5985 ( .C1(n4871), .C2(INSTQUEUE_REG_2__2__SCAN_IN), .A(n4846), 
        .B(n4845), .ZN(n4847) );
  INV_X1 U5986 ( .A(n4847), .ZN(U3038) );
  NOR2_X1 U5987 ( .A1(n4864), .A2(n6335), .ZN(n4850) );
  AOI22_X1 U5988 ( .A1(n6321), .A2(n4866), .B1(n6320), .B2(n4865), .ZN(n4848)
         );
  OAI21_X1 U5989 ( .B1(n4868), .B2(n6233), .A(n4848), .ZN(n4849) );
  AOI211_X1 U5990 ( .C1(n4871), .C2(INSTQUEUE_REG_2__0__SCAN_IN), .A(n4850), 
        .B(n4849), .ZN(n4851) );
  INV_X1 U5991 ( .A(n4851), .ZN(U3036) );
  NOR2_X1 U5992 ( .A1(n4864), .A2(n6359), .ZN(n4854) );
  AOI22_X1 U5993 ( .A1(n6355), .A2(n4866), .B1(n6354), .B2(n4865), .ZN(n4852)
         );
  OAI21_X1 U5994 ( .B1(n4868), .B2(n6295), .A(n4852), .ZN(n4853) );
  AOI211_X1 U5995 ( .C1(n4871), .C2(INSTQUEUE_REG_2__4__SCAN_IN), .A(n4854), 
        .B(n4853), .ZN(n4855) );
  INV_X1 U5996 ( .A(n4855), .ZN(U3040) );
  NOR2_X1 U5997 ( .A1(n4864), .A2(n6365), .ZN(n4858) );
  AOI22_X1 U5998 ( .A1(n6361), .A2(n4866), .B1(n6360), .B2(n4865), .ZN(n4856)
         );
  OAI21_X1 U5999 ( .B1(n4868), .B2(n6297), .A(n4856), .ZN(n4857) );
  AOI211_X1 U6000 ( .C1(n4871), .C2(INSTQUEUE_REG_2__5__SCAN_IN), .A(n4858), 
        .B(n4857), .ZN(n4859) );
  INV_X1 U6001 ( .A(n4859), .ZN(U3041) );
  NOR2_X1 U6002 ( .A1(n4864), .A2(n6559), .ZN(n4862) );
  AOI22_X1 U6003 ( .A1(n6374), .A2(n4866), .B1(n6550), .B2(n4865), .ZN(n4860)
         );
  OAI21_X1 U6004 ( .B1(n4868), .B2(n6314), .A(n4860), .ZN(n4861) );
  AOI211_X1 U6005 ( .C1(n4871), .C2(INSTQUEUE_REG_2__7__SCAN_IN), .A(n4862), 
        .B(n4861), .ZN(n4863) );
  INV_X1 U6006 ( .A(n4863), .ZN(U3043) );
  NOR2_X1 U6007 ( .A1(n4864), .A2(n6353), .ZN(n4870) );
  AOI22_X1 U6008 ( .A1(n6349), .A2(n4866), .B1(n6348), .B2(n4865), .ZN(n4867)
         );
  OAI21_X1 U6009 ( .B1(n4868), .B2(n6290), .A(n4867), .ZN(n4869) );
  AOI211_X1 U6010 ( .C1(n4871), .C2(INSTQUEUE_REG_2__3__SCAN_IN), .A(n4870), 
        .B(n4869), .ZN(n4872) );
  INV_X1 U6011 ( .A(n4872), .ZN(U3039) );
  NAND2_X1 U6012 ( .A1(n5785), .A2(n4873), .ZN(n4874) );
  NAND2_X1 U6013 ( .A1(n5764), .A2(n4874), .ZN(n5840) );
  INV_X1 U6014 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U6015 ( .A1(n4875), .A2(n5785), .ZN(n5826) );
  INV_X1 U6016 ( .A(n5826), .ZN(n5854) );
  AOI21_X1 U6017 ( .B1(n5845), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5854), 
        .ZN(n4882) );
  INV_X1 U6018 ( .A(n4876), .ZN(n4879) );
  INV_X1 U6019 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5247) );
  NAND3_X1 U6020 ( .A1(n3187), .A2(n5247), .A3(n4877), .ZN(n4878) );
  NAND2_X1 U6021 ( .A1(n4879), .A2(n4878), .ZN(n4880) );
  AOI22_X1 U6022 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5848), .B1(n5825), .B2(n6059), 
        .ZN(n4881) );
  OAI211_X1 U6023 ( .C1(n5840), .C2(n6461), .A(n4882), .B(n4881), .ZN(n4888)
         );
  NOR2_X1 U6024 ( .A1(n5787), .A2(n5021), .ZN(n5849) );
  NOR2_X1 U6025 ( .A1(n6456), .A2(n6458), .ZN(n4885) );
  AND2_X1 U6026 ( .A1(n5849), .A2(n4885), .ZN(n5837) );
  OAI211_X1 U6027 ( .C1(REIP_REG_7__SCAN_IN), .C2(REIP_REG_6__SCAN_IN), .A(
        n5837), .B(n4943), .ZN(n4886) );
  OAI21_X1 U6028 ( .B1(n5870), .B2(n4921), .A(n4886), .ZN(n4887) );
  AOI211_X1 U6029 ( .C1(n4923), .C2(n4093), .A(n4888), .B(n4887), .ZN(n4889)
         );
  INV_X1 U6030 ( .A(n4889), .ZN(U2820) );
  NAND2_X1 U6031 ( .A1(n4953), .A2(n4890), .ZN(n4891) );
  AOI22_X1 U6032 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n5845), .B1(n5825), 
        .B2(n6068), .ZN(n4893) );
  OAI211_X1 U6033 ( .C1(n5858), .C2(n4894), .A(n4893), .B(n5826), .ZN(n4897)
         );
  NAND2_X1 U6034 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5849), .ZN(n4895) );
  AOI21_X1 U6035 ( .B1(n6458), .B2(n4895), .A(n5840), .ZN(n4896) );
  AOI211_X1 U6036 ( .C1(n4892), .C2(n4898), .A(n4897), .B(n4896), .ZN(n4899)
         );
  OAI21_X1 U6037 ( .B1(n5843), .B2(n4900), .A(n4899), .ZN(U2822) );
  OAI21_X1 U6038 ( .B1(n4903), .B2(n4902), .A(n4901), .ZN(n4904) );
  INV_X1 U6039 ( .A(n4904), .ZN(n5994) );
  INV_X1 U6040 ( .A(REIP_REG_6__SCAN_IN), .ZN(n5836) );
  OAI22_X1 U6041 ( .A1(n5833), .A2(n6079), .B1(n6032), .B2(n5836), .ZN(n4915)
         );
  AOI21_X1 U6043 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6093) );
  NOR2_X1 U6044 ( .A1(n6672), .A2(n6561), .ZN(n6689) );
  NAND2_X1 U6045 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6689), .ZN(n5089)
         );
  OR2_X1 U6046 ( .A1(n6093), .A2(n5089), .ZN(n5088) );
  NOR2_X1 U6047 ( .A1(n6106), .A2(n4905), .ZN(n6094) );
  NAND2_X1 U6048 ( .A1(n4906), .A2(n6099), .ZN(n6025) );
  OAI21_X1 U6049 ( .B1(n6030), .B2(n6094), .A(n6025), .ZN(n6092) );
  AOI21_X1 U6050 ( .B1(n5088), .B2(n6031), .A(n6092), .ZN(n6073) );
  INV_X1 U6051 ( .A(n5583), .ZN(n4908) );
  NAND2_X1 U6052 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4908), .ZN(n6107)
         );
  INV_X1 U6053 ( .A(n6107), .ZN(n4909) );
  NAND2_X1 U6054 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n4909), .ZN(n4910)
         );
  NAND2_X1 U6055 ( .A1(n6099), .A2(n4910), .ZN(n4912) );
  INV_X1 U6056 ( .A(n6093), .ZN(n4911) );
  INV_X1 U6057 ( .A(n6066), .ZN(n6085) );
  OAI33_X1 U6058 ( .A1(1'b0), .A2(n6073), .A3(n5090), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n5089), .B3(n6085), .ZN(n4914) );
  AOI211_X1 U6059 ( .C1(n5994), .C2(n6102), .A(n4915), .B(n4914), .ZN(n4916)
         );
  INV_X1 U6060 ( .A(n4916), .ZN(U3012) );
  OAI21_X1 U6061 ( .B1(n4919), .B2(n4918), .A(n4917), .ZN(n6060) );
  NAND2_X1 U6062 ( .A1(n6095), .A2(REIP_REG_7__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U6063 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4920)
         );
  OAI211_X1 U6064 ( .C1(n6015), .C2(n4921), .A(n6057), .B(n4920), .ZN(n4922)
         );
  AOI21_X1 U6065 ( .B1(n4923), .B2(n5446), .A(n4922), .ZN(n4924) );
  OAI21_X1 U6066 ( .B1(n6060), .B2(n5992), .A(n4924), .ZN(U2979) );
  INV_X1 U6067 ( .A(n4925), .ZN(n4928) );
  AOI21_X1 U6068 ( .B1(n4928), .B2(n4927), .A(n4926), .ZN(n5060) );
  INV_X1 U6069 ( .A(n5060), .ZN(n4941) );
  AOI22_X1 U6070 ( .A1(n5322), .A2(DATAI_10_), .B1(n5885), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4929) );
  OAI21_X1 U6071 ( .B1(n4941), .B2(n5671), .A(n4929), .ZN(U2881) );
  INV_X1 U6072 ( .A(n5058), .ZN(n4935) );
  INV_X1 U6073 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U6074 ( .A1(n5820), .A2(n4930), .ZN(n4931) );
  NAND2_X1 U6075 ( .A1(n5800), .A2(n4931), .ZN(n6033) );
  OAI22_X1 U6076 ( .A1(n4940), .A2(n5858), .B1(n5861), .B2(n6033), .ZN(n4934)
         );
  INV_X1 U6077 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6465) );
  NAND4_X1 U6078 ( .A1(REIP_REG_9__SCAN_IN), .A2(n4937), .A3(n5837), .A4(n6465), .ZN(n4932) );
  OAI211_X1 U6079 ( .C1(n5856), .C2(n6660), .A(n5826), .B(n4932), .ZN(n4933)
         );
  AOI211_X1 U6080 ( .C1(n4892), .C2(n4935), .A(n4934), .B(n4933), .ZN(n4939)
         );
  NAND2_X1 U6081 ( .A1(n4937), .A2(n5837), .ZN(n4936) );
  NOR2_X1 U6082 ( .A1(REIP_REG_9__SCAN_IN), .A2(n4936), .ZN(n5830) );
  OAI21_X1 U6083 ( .B1(n4937), .B2(n5787), .A(n5840), .ZN(n5824) );
  OAI21_X1 U6084 ( .B1(n5830), .B2(n5824), .A(REIP_REG_10__SCAN_IN), .ZN(n4938) );
  OAI211_X1 U6085 ( .C1(n4941), .C2(n5810), .A(n4939), .B(n4938), .ZN(U2817)
         );
  OAI222_X1 U6086 ( .A1(n4941), .A2(n5300), .B1(n5878), .B2(n4940), .C1(n6033), 
        .C2(n5872), .ZN(U2849) );
  INV_X1 U6087 ( .A(n5837), .ZN(n4942) );
  OAI21_X1 U6088 ( .B1(n4943), .B2(n4942), .A(n6463), .ZN(n4948) );
  AOI22_X1 U6089 ( .A1(EBX_REG_8__SCAN_IN), .A2(n5848), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n5845), .ZN(n4946) );
  INV_X1 U6090 ( .A(n4964), .ZN(n4944) );
  AOI22_X1 U6091 ( .A1(n6051), .A2(n5825), .B1(n4944), .B2(n4892), .ZN(n4945)
         );
  NAND3_X1 U6092 ( .A1(n4946), .A2(n4945), .A3(n5826), .ZN(n4947) );
  AOI21_X1 U6093 ( .B1(n4948), .B2(n5824), .A(n4947), .ZN(n4949) );
  OAI21_X1 U6094 ( .B1(n4950), .B2(n5810), .A(n4949), .ZN(U2819) );
  INV_X1 U6095 ( .A(n4951), .ZN(n4952) );
  NAND2_X1 U6096 ( .A1(n4953), .A2(n4952), .ZN(n5859) );
  AOI22_X1 U6097 ( .A1(EBX_REG_0__SCAN_IN), .A2(n5848), .B1(n5825), .B2(n4954), 
        .ZN(n4956) );
  OAI21_X1 U6098 ( .B1(n5845), .B2(n4892), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4955) );
  OAI211_X1 U6099 ( .C1(n5859), .C2(n2956), .A(n4956), .B(n4955), .ZN(n4957)
         );
  AOI21_X1 U6100 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5764), .A(n4957), .ZN(n4958)
         );
  OAI21_X1 U6101 ( .B1(n5843), .B2(n4959), .A(n4958), .ZN(U2827) );
  OAI21_X1 U6102 ( .B1(n4962), .B2(n4961), .A(n4960), .ZN(n6052) );
  NAND2_X1 U6103 ( .A1(n6095), .A2(REIP_REG_8__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U6104 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4963)
         );
  OAI211_X1 U6105 ( .C1(n6015), .C2(n4964), .A(n6049), .B(n4963), .ZN(n4965)
         );
  AOI21_X1 U6106 ( .B1(n4966), .B2(n5446), .A(n4965), .ZN(n4967) );
  OAI21_X1 U6107 ( .B1(n6052), .B2(n5992), .A(n4967), .ZN(U2978) );
  OAI22_X1 U6108 ( .A1(n4968), .A2(n5861), .B1(n5785), .B2(n6527), .ZN(n4969)
         );
  AOI21_X1 U6109 ( .B1(EBX_REG_1__SCAN_IN), .B2(n5848), .A(n4969), .ZN(n4975)
         );
  NAND2_X1 U6110 ( .A1(n5865), .A2(n6527), .ZN(n4972) );
  AOI22_X1 U6111 ( .A1(n5845), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n4892), 
        .B2(n4970), .ZN(n4971) );
  OAI211_X1 U6112 ( .C1(n5859), .C2(n5624), .A(n4972), .B(n4971), .ZN(n4973)
         );
  INV_X1 U6113 ( .A(n4973), .ZN(n4974) );
  OAI211_X1 U6114 ( .C1(n5843), .C2(n4976), .A(n4975), .B(n4974), .ZN(U2826)
         );
  AND2_X1 U6115 ( .A1(n5622), .A2(n4977), .ZN(n4978) );
  NOR3_X1 U6116 ( .A1(n6316), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n4979), 
        .ZN(n4980) );
  AOI21_X1 U6117 ( .B1(n4981), .B2(n6317), .A(n4980), .ZN(n6552) );
  NOR2_X1 U6118 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6228), .ZN(n6549)
         );
  AOI21_X1 U6119 ( .B1(n6558), .B2(n6253), .A(n6322), .ZN(n4982) );
  NOR3_X1 U6120 ( .A1(n6325), .A2(n6224), .A3(n4982), .ZN(n4984) );
  NOR3_X1 U6121 ( .A1(n6152), .A2(n4984), .A3(n4983), .ZN(n4986) );
  AOI22_X1 U6122 ( .A1(n6337), .A2(n6549), .B1(INSTQUEUE_REG_6__1__SCAN_IN), 
        .B2(n6548), .ZN(n4987) );
  OAI21_X1 U6123 ( .B1(n6552), .B2(n4988), .A(n4987), .ZN(n4989) );
  AOI21_X1 U6124 ( .B1(n6555), .B2(n6338), .A(n4989), .ZN(n4990) );
  OAI21_X1 U6125 ( .B1(n6341), .B2(n6558), .A(n4990), .ZN(U3069) );
  NOR2_X1 U6126 ( .A1(n4926), .A2(n4992), .ZN(n4993) );
  OR2_X1 U6127 ( .A1(n4991), .A2(n4993), .ZN(n5988) );
  AOI22_X1 U6128 ( .A1(n5322), .A2(DATAI_11_), .B1(n5885), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4994) );
  OAI21_X1 U6129 ( .B1(n5988), .B2(n5671), .A(n4994), .ZN(U2880) );
  AOI22_X1 U6130 ( .A1(n6354), .A2(n6549), .B1(INSTQUEUE_REG_6__4__SCAN_IN), 
        .B2(n6548), .ZN(n4995) );
  OAI21_X1 U6131 ( .B1(n4996), .B2(n6552), .A(n4995), .ZN(n4997) );
  AOI21_X1 U6132 ( .B1(n6356), .B2(n6555), .A(n4997), .ZN(n4998) );
  OAI21_X1 U6133 ( .B1(n6359), .B2(n6558), .A(n4998), .ZN(U3072) );
  AOI22_X1 U6134 ( .A1(n6360), .A2(n6549), .B1(INSTQUEUE_REG_6__5__SCAN_IN), 
        .B2(n6548), .ZN(n4999) );
  OAI21_X1 U6135 ( .B1(n5000), .B2(n6552), .A(n4999), .ZN(n5001) );
  AOI21_X1 U6136 ( .B1(n6362), .B2(n6555), .A(n5001), .ZN(n5002) );
  OAI21_X1 U6137 ( .B1(n6365), .B2(n6558), .A(n5002), .ZN(U3073) );
  AOI22_X1 U6138 ( .A1(n6320), .A2(n6549), .B1(INSTQUEUE_REG_6__0__SCAN_IN), 
        .B2(n6548), .ZN(n5003) );
  OAI21_X1 U6139 ( .B1(n5004), .B2(n6552), .A(n5003), .ZN(n5005) );
  AOI21_X1 U6140 ( .B1(n6332), .B2(n6555), .A(n5005), .ZN(n5006) );
  OAI21_X1 U6141 ( .B1(n6335), .B2(n6558), .A(n5006), .ZN(U3068) );
  AOI22_X1 U6142 ( .A1(n6348), .A2(n6549), .B1(INSTQUEUE_REG_6__3__SCAN_IN), 
        .B2(n6548), .ZN(n5007) );
  OAI21_X1 U6143 ( .B1(n5008), .B2(n6552), .A(n5007), .ZN(n5009) );
  AOI21_X1 U6144 ( .B1(n6350), .B2(n6555), .A(n5009), .ZN(n5010) );
  OAI21_X1 U6145 ( .B1(n6353), .B2(n6558), .A(n5010), .ZN(U3071) );
  AOI22_X1 U6146 ( .A1(n6366), .A2(n6549), .B1(INSTQUEUE_REG_6__6__SCAN_IN), 
        .B2(n6548), .ZN(n5011) );
  OAI21_X1 U6147 ( .B1(n5012), .B2(n6552), .A(n5011), .ZN(n5013) );
  AOI21_X1 U6148 ( .B1(n6368), .B2(n6555), .A(n5013), .ZN(n5014) );
  OAI21_X1 U6149 ( .B1(n6371), .B2(n6558), .A(n5014), .ZN(U3074) );
  AOI22_X1 U6150 ( .A1(n6342), .A2(n6549), .B1(INSTQUEUE_REG_6__2__SCAN_IN), 
        .B2(n6548), .ZN(n5015) );
  OAI21_X1 U6151 ( .B1(n5016), .B2(n6552), .A(n5015), .ZN(n5017) );
  AOI21_X1 U6152 ( .B1(n6344), .B2(n6555), .A(n5017), .ZN(n5018) );
  OAI21_X1 U6153 ( .B1(n6347), .B2(n6558), .A(n5018), .ZN(U3070) );
  INV_X1 U6154 ( .A(n5859), .ZN(n5031) );
  INV_X1 U6155 ( .A(n5021), .ZN(n5019) );
  NAND2_X1 U6156 ( .A1(n5785), .A2(n5019), .ZN(n5020) );
  NAND2_X1 U6157 ( .A1(n5764), .A2(n5020), .ZN(n5844) );
  INV_X1 U6158 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6454) );
  NOR2_X1 U6159 ( .A1(n5844), .A2(n6454), .ZN(n5030) );
  OAI211_X1 U6160 ( .C1(n5787), .C2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .B(n5785), .ZN(n5866) );
  NAND2_X1 U6161 ( .A1(n5865), .A2(n5021), .ZN(n5028) );
  INV_X1 U6162 ( .A(n5022), .ZN(n5023) );
  AOI22_X1 U6163 ( .A1(n5023), .A2(n4892), .B1(n5845), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U6164 ( .A1(n5825), .A2(n6084), .ZN(n5025) );
  NAND2_X1 U6165 ( .A1(n5848), .A2(EBX_REG_3__SCAN_IN), .ZN(n5024) );
  AND3_X1 U6166 ( .A1(n5026), .A2(n5025), .A3(n5024), .ZN(n5027) );
  OAI21_X1 U6167 ( .B1(n5866), .B2(n5028), .A(n5027), .ZN(n5029) );
  AOI211_X1 U6168 ( .C1(n5031), .C2(n6146), .A(n5030), .B(n5029), .ZN(n5032)
         );
  OAI21_X1 U6169 ( .B1(n5033), .B2(n5843), .A(n5032), .ZN(U2824) );
  XOR2_X1 U6170 ( .A(n5034), .B(n4991), .Z(n5104) );
  INV_X1 U6171 ( .A(n5104), .ZN(n5052) );
  AOI22_X1 U6172 ( .A1(n5322), .A2(DATAI_12_), .B1(n5885), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5035) );
  OAI21_X1 U6173 ( .B1(n5052), .B2(n5671), .A(n5035), .ZN(U2879) );
  INV_X1 U6174 ( .A(n5102), .ZN(n5044) );
  AOI22_X1 U6175 ( .A1(EBX_REG_12__SCAN_IN), .A2(n5848), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5845), .ZN(n5037) );
  INV_X1 U6176 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6469) );
  NAND3_X1 U6177 ( .A1(n5865), .A2(n5038), .A3(n6469), .ZN(n5036) );
  NAND3_X1 U6178 ( .A1(n5037), .A2(n5826), .A3(n5036), .ZN(n5043) );
  NOR2_X1 U6179 ( .A1(n5787), .A2(n5038), .ZN(n5804) );
  NOR2_X1 U6180 ( .A1(n5039), .A2(n5804), .ZN(n5807) );
  OR2_X1 U6181 ( .A1(n5802), .A2(n5040), .ZN(n5041) );
  NAND2_X1 U6182 ( .A1(n5070), .A2(n5041), .ZN(n5093) );
  OAI22_X1 U6183 ( .A1(n5807), .A2(n6469), .B1(n5861), .B2(n5093), .ZN(n5042)
         );
  AOI211_X1 U6184 ( .C1(n4892), .C2(n5044), .A(n5043), .B(n5042), .ZN(n5045)
         );
  OAI21_X1 U6185 ( .B1(n5052), .B2(n5810), .A(n5045), .ZN(U2815) );
  XNOR2_X1 U6186 ( .A(n4226), .B(n5047), .ZN(n5048) );
  XNOR2_X1 U6187 ( .A(n5046), .B(n5048), .ZN(n6044) );
  INV_X1 U6188 ( .A(n5992), .ZN(n6011) );
  NAND2_X1 U6189 ( .A1(n6044), .A2(n6011), .ZN(n5051) );
  NAND2_X1 U6190 ( .A1(n6095), .A2(REIP_REG_9__SCAN_IN), .ZN(n6040) );
  OAI21_X1 U6191 ( .B1(n5461), .B2(n5828), .A(n6040), .ZN(n5049) );
  AOI21_X1 U6192 ( .B1(n5464), .B2(n5816), .A(n5049), .ZN(n5050) );
  OAI211_X1 U6193 ( .C1(n5987), .C2(n5815), .A(n5051), .B(n5050), .ZN(U2977)
         );
  INV_X1 U6194 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5053) );
  OAI222_X1 U6195 ( .A1(n5093), .A2(n5872), .B1(n5878), .B2(n5053), .C1(n5300), 
        .C2(n5052), .ZN(U2847) );
  NAND2_X1 U6196 ( .A1(n5982), .A2(n5055), .ZN(n5056) );
  XNOR2_X1 U6197 ( .A(n5054), .B(n5056), .ZN(n6035) );
  INV_X1 U6198 ( .A(n6035), .ZN(n5062) );
  AOI22_X1 U6199 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6095), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5057) );
  OAI21_X1 U6200 ( .B1(n6015), .B2(n5058), .A(n5057), .ZN(n5059) );
  AOI21_X1 U6201 ( .B1(n5060), .B2(n5446), .A(n5059), .ZN(n5061) );
  OAI21_X1 U6202 ( .B1(n5062), .B2(n5992), .A(n5061), .ZN(U2976) );
  INV_X1 U6203 ( .A(n5063), .ZN(n5066) );
  INV_X1 U6204 ( .A(n5064), .ZN(n5065) );
  NAND2_X1 U6205 ( .A1(n5066), .A2(n5065), .ZN(n5067) );
  AND2_X1 U6206 ( .A1(n5068), .A2(n5067), .ZN(n5795) );
  NAND2_X1 U6207 ( .A1(n5070), .A2(n5069), .ZN(n5071) );
  NAND2_X1 U6208 ( .A1(n5082), .A2(n5071), .ZN(n5793) );
  OAI22_X1 U6209 ( .A1(n5793), .A2(n5872), .B1(n5798), .B2(n5878), .ZN(n5072)
         );
  AOI21_X1 U6210 ( .B1(n5795), .B2(n3900), .A(n5072), .ZN(n5073) );
  INV_X1 U6211 ( .A(n5073), .ZN(U2846) );
  INV_X1 U6212 ( .A(n5795), .ZN(n5075) );
  AOI22_X1 U6213 ( .A1(n5322), .A2(DATAI_13_), .B1(n5885), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5074) );
  OAI21_X1 U6214 ( .B1(n5075), .B2(n5671), .A(n5074), .ZN(U2878) );
  OAI21_X1 U6215 ( .B1(n5076), .B2(n5079), .A(n5078), .ZN(n5779) );
  AOI22_X1 U6216 ( .A1(n5322), .A2(DATAI_14_), .B1(n5885), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5080) );
  OAI21_X1 U6217 ( .B1(n5779), .B2(n5671), .A(n5080), .ZN(U2877) );
  INV_X1 U6218 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6219 ( .A1(n5082), .A2(n5081), .ZN(n5083) );
  NAND2_X1 U6220 ( .A1(n5242), .A2(n5083), .ZN(n5784) );
  OAI222_X1 U6221 ( .A1(n5779), .A2(n5300), .B1(n5084), .B2(n5878), .C1(n5872), 
        .C2(n5784), .ZN(U2845) );
  NOR2_X1 U6222 ( .A1(n5086), .A2(n2971), .ZN(n5087) );
  XNOR2_X1 U6223 ( .A(n5085), .B(n5087), .ZN(n5106) );
  INV_X1 U6224 ( .A(n6099), .ZN(n6074) );
  NAND2_X1 U6225 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U6226 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6037) );
  NOR2_X1 U6227 ( .A1(n6048), .A2(n6037), .ZN(n5091) );
  NOR2_X1 U6228 ( .A1(n5090), .A2(n5088), .ZN(n6026) );
  NAND2_X1 U6229 ( .A1(n5091), .A2(n6026), .ZN(n5468) );
  NOR2_X1 U6230 ( .A1(n5090), .A2(n5089), .ZN(n6036) );
  AND2_X1 U6231 ( .A1(n6094), .A2(n6036), .ZN(n6029) );
  NAND2_X1 U6232 ( .A1(n6029), .A2(n5091), .ZN(n5705) );
  INV_X1 U6233 ( .A(n5705), .ZN(n5717) );
  OAI21_X1 U6234 ( .B1(n6030), .B2(n5717), .A(n6025), .ZN(n5587) );
  AOI21_X1 U6235 ( .B1(n6074), .B2(n5468), .A(n5587), .ZN(n6024) );
  NOR2_X1 U6236 ( .A1(n5705), .A2(n5583), .ZN(n5094) );
  OAI21_X1 U6237 ( .B1(n6074), .B2(n5094), .A(n6022), .ZN(n5092) );
  AOI21_X1 U6238 ( .B1(n6024), .B2(n5092), .A(n5704), .ZN(n5098) );
  NAND2_X1 U6239 ( .A1(n6095), .A2(REIP_REG_12__SCAN_IN), .ZN(n5101) );
  INV_X1 U6240 ( .A(n5101), .ZN(n5097) );
  NOR2_X1 U6241 ( .A1(n5093), .A2(n6079), .ZN(n5096) );
  NOR2_X1 U6242 ( .A1(n6099), .A2(n5468), .ZN(n5708) );
  NOR3_X1 U6243 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6016), .A3(n6022), 
        .ZN(n5095) );
  NOR4_X1 U6244 ( .A1(n5098), .A2(n5097), .A3(n5096), .A4(n5095), .ZN(n5099)
         );
  OAI21_X1 U6245 ( .B1(n5106), .B2(n6086), .A(n5099), .ZN(U3006) );
  NAND2_X1 U6246 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5100)
         );
  OAI211_X1 U6247 ( .C1(n6015), .C2(n5102), .A(n5101), .B(n5100), .ZN(n5103)
         );
  AOI21_X1 U6248 ( .B1(n5104), .B2(n5446), .A(n5103), .ZN(n5105) );
  OAI21_X1 U6249 ( .B1(n5106), .B2(n5992), .A(n5105), .ZN(U2974) );
  OAI21_X1 U6250 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6514), .A(n6521), 
        .ZN(n6522) );
  INV_X1 U6251 ( .A(n6522), .ZN(n5117) );
  INV_X1 U6252 ( .A(n5108), .ZN(n5112) );
  NOR2_X1 U6253 ( .A1(n4437), .A2(n4295), .ZN(n5109) );
  AOI22_X1 U6254 ( .A1(n6383), .A2(n3039), .B1(n5109), .B2(n6380), .ZN(n5110)
         );
  OAI21_X1 U6255 ( .B1(n5624), .B2(n5111), .A(n5110), .ZN(n6385) );
  AOI222_X1 U6256 ( .A1(n5114), .A2(n5107), .B1(n5113), .B2(n5112), .C1(n6385), 
        .C2(n5728), .ZN(n5116) );
  OAI22_X1 U6257 ( .A1(n5117), .A2(n3039), .B1(n5116), .B2(n5115), .ZN(U3460)
         );
  AOI22_X1 U6258 ( .A1(n5882), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5885), .ZN(n5122) );
  AND2_X1 U6259 ( .A1(n3209), .A2(n3894), .ZN(n5119) );
  NAND2_X1 U6260 ( .A1(n5886), .A2(DATAI_14_), .ZN(n5121) );
  OAI211_X1 U6261 ( .C1(n5118), .C2(n5671), .A(n5122), .B(n5121), .ZN(U2861)
         );
  INV_X1 U6262 ( .A(n5126), .ZN(n5125) );
  INV_X1 U6263 ( .A(n5127), .ZN(n5124) );
  AOI211_X1 U6264 ( .C1(n5144), .C2(n5125), .A(n5124), .B(n5123), .ZN(n5130)
         );
  AOI211_X1 U6265 ( .C1(n5128), .C2(n5158), .A(n5127), .B(n5126), .ZN(n5129)
         );
  NOR2_X1 U6266 ( .A1(n5130), .A2(n5129), .ZN(n5500) );
  AOI22_X1 U6267 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5845), .B1(n4892), 
        .B2(n5131), .ZN(n5132) );
  OAI21_X1 U6268 ( .B1(n5858), .B2(n5139), .A(n5132), .ZN(n5133) );
  AOI21_X1 U6269 ( .B1(n5500), .B2(n5825), .A(n5133), .ZN(n5137) );
  NOR2_X1 U6270 ( .A1(n5149), .A2(n6495), .ZN(n5135) );
  OAI21_X1 U6271 ( .B1(n5135), .B2(REIP_REG_30__SCAN_IN), .A(n5134), .ZN(n5136) );
  OAI211_X1 U6272 ( .C1(n5118), .C2(n5810), .A(n5137), .B(n5136), .ZN(U2797)
         );
  INV_X1 U6273 ( .A(n5500), .ZN(n5138) );
  OAI222_X1 U6274 ( .A1(n5300), .A2(n5118), .B1(n5139), .B2(n5878), .C1(n5138), 
        .C2(n5872), .ZN(U2829) );
  OAI21_X2 U6275 ( .B1(n5140), .B2(n5142), .A(n5141), .ZN(n5328) );
  XNOR2_X1 U6276 ( .A(n5144), .B(n5143), .ZN(n5509) );
  INV_X1 U6277 ( .A(n5145), .ZN(n5330) );
  OAI22_X1 U6278 ( .A1(n5146), .A2(n5856), .B1(n5870), .B2(n5330), .ZN(n5147)
         );
  AOI21_X1 U6279 ( .B1(n5848), .B2(EBX_REG_29__SCAN_IN), .A(n5147), .ZN(n5148)
         );
  OAI21_X1 U6280 ( .B1(n5154), .B2(n6495), .A(n5148), .ZN(n5151) );
  NOR2_X1 U6281 ( .A1(n5149), .A2(REIP_REG_29__SCAN_IN), .ZN(n5150) );
  AOI211_X1 U6282 ( .C1(n5825), .C2(n5509), .A(n5151), .B(n5150), .ZN(n5152)
         );
  OAI21_X1 U6283 ( .B1(n5328), .B2(n5810), .A(n5152), .ZN(U2798) );
  AOI21_X1 U6284 ( .B1(n5153), .B2(n4026), .A(n5140), .ZN(n5343) );
  INV_X1 U6285 ( .A(n5343), .ZN(n5305) );
  INV_X1 U6286 ( .A(n5154), .ZN(n5165) );
  NAND2_X1 U6287 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  NAND2_X1 U6288 ( .A1(n5158), .A2(n5157), .ZN(n5516) );
  INV_X1 U6289 ( .A(n5341), .ZN(n5159) );
  AOI22_X1 U6290 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n5845), .B1(n4892), 
        .B2(n5159), .ZN(n5161) );
  NAND2_X1 U6291 ( .A1(n5848), .A2(EBX_REG_28__SCAN_IN), .ZN(n5160) );
  OAI211_X1 U6292 ( .C1(n5516), .C2(n5861), .A(n5161), .B(n5160), .ZN(n5164)
         );
  INV_X1 U6293 ( .A(n5171), .ZN(n5162) );
  INV_X1 U6294 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6611) );
  NOR3_X1 U6295 ( .A1(n5162), .A2(REIP_REG_28__SCAN_IN), .A3(n6611), .ZN(n5163) );
  AOI211_X1 U6296 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5165), .A(n5164), .B(n5163), .ZN(n5166) );
  OAI21_X1 U6297 ( .B1(n5305), .B2(n5810), .A(n5166), .ZN(U2799) );
  NOR2_X1 U6298 ( .A1(n5186), .A2(n6611), .ZN(n5170) );
  AOI22_X1 U6299 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n5845), .B1(n4892), 
        .B2(n5349), .ZN(n5168) );
  NAND2_X1 U6300 ( .A1(n5848), .A2(EBX_REG_27__SCAN_IN), .ZN(n5167) );
  OAI211_X1 U6301 ( .C1(n5521), .C2(n5861), .A(n5168), .B(n5167), .ZN(n5169)
         );
  AOI211_X1 U6302 ( .C1(n5171), .C2(n6611), .A(n5170), .B(n5169), .ZN(n5172)
         );
  OAI21_X1 U6303 ( .B1(n5308), .B2(n5810), .A(n5172), .ZN(U2800) );
  INV_X1 U6304 ( .A(n5173), .ZN(n5207) );
  AOI21_X1 U6305 ( .B1(n5207), .B2(n5174), .A(REIP_REG_26__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6306 ( .A1(n5175), .A2(n5176), .ZN(n5177) );
  NAND2_X1 U6307 ( .A1(n5178), .A2(n5177), .ZN(n5311) );
  INV_X1 U6308 ( .A(n5311), .ZN(n5359) );
  NAND2_X1 U6309 ( .A1(n5359), .A2(n4093), .ZN(n5184) );
  OAI22_X1 U6310 ( .A1(n5179), .A2(n5856), .B1(n5870), .B2(n5357), .ZN(n5182)
         );
  XNOR2_X1 U6311 ( .A(n5191), .B(n5180), .ZN(n5533) );
  NOR2_X1 U6312 ( .A1(n5533), .A2(n5861), .ZN(n5181) );
  AOI211_X1 U6313 ( .C1(n5848), .C2(EBX_REG_26__SCAN_IN), .A(n5182), .B(n5181), 
        .ZN(n5183) );
  OAI211_X1 U6314 ( .C1(n5186), .C2(n5185), .A(n5184), .B(n5183), .ZN(U2801)
         );
  XNOR2_X1 U6315 ( .A(n5187), .B(n5188), .ZN(n5365) );
  XOR2_X1 U6316 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .Z(n5196) );
  INV_X1 U6317 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6490) );
  NOR2_X1 U6318 ( .A1(n5636), .A2(n6490), .ZN(n5195) );
  NOR2_X1 U6319 ( .A1(n5200), .A2(n5189), .ZN(n5190) );
  OR2_X1 U6320 ( .A1(n5191), .A2(n5190), .ZN(n5539) );
  AOI22_X1 U6321 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n5845), .B1(n4892), 
        .B2(n5368), .ZN(n5193) );
  NAND2_X1 U6322 ( .A1(n5848), .A2(EBX_REG_25__SCAN_IN), .ZN(n5192) );
  OAI211_X1 U6323 ( .C1(n5539), .C2(n5861), .A(n5193), .B(n5192), .ZN(n5194)
         );
  AOI211_X1 U6324 ( .C1(n5196), .C2(n5207), .A(n5195), .B(n5194), .ZN(n5197)
         );
  OAI21_X1 U6325 ( .B1(n5365), .B2(n5810), .A(n5197), .ZN(U2802) );
  NOR2_X1 U6326 ( .A1(n2959), .A2(n5198), .ZN(n5199) );
  OR2_X1 U6327 ( .A1(n5187), .A2(n5199), .ZN(n5377) );
  INV_X1 U6328 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6487) );
  AOI21_X1 U6329 ( .B1(n5201), .B2(n5257), .A(n5200), .ZN(n5551) );
  NAND2_X1 U6330 ( .A1(n5551), .A2(n5825), .ZN(n5205) );
  OAI22_X1 U6331 ( .A1(n5202), .A2(n5856), .B1(n5870), .B2(n5379), .ZN(n5203)
         );
  AOI21_X1 U6332 ( .B1(n5848), .B2(EBX_REG_24__SCAN_IN), .A(n5203), .ZN(n5204)
         );
  OAI211_X1 U6333 ( .C1(n5636), .C2(n6487), .A(n5205), .B(n5204), .ZN(n5206)
         );
  AOI21_X1 U6334 ( .B1(n5207), .B2(n6487), .A(n5206), .ZN(n5208) );
  OAI21_X1 U6335 ( .B1(n5377), .B2(n5810), .A(n5208), .ZN(U2803) );
  NOR2_X1 U6336 ( .A1(n2964), .A2(n5210), .ZN(n5211) );
  OR2_X1 U6337 ( .A1(n5209), .A2(n5211), .ZN(n5407) );
  NAND2_X1 U6338 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5662) );
  INV_X1 U6339 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6481) );
  OAI21_X1 U6340 ( .B1(n5762), .B2(n5662), .A(n6481), .ZN(n5219) );
  AND2_X1 U6341 ( .A1(n5764), .A2(n5212), .ZN(n5654) );
  MUX2_X1 U6342 ( .A(n5274), .B(n5271), .S(n5213), .Z(n5215) );
  XNOR2_X1 U6343 ( .A(n5215), .B(n5214), .ZN(n5603) );
  INV_X1 U6344 ( .A(n5603), .ZN(n5267) );
  OAI22_X1 U6345 ( .A1(n3956), .A2(n5858), .B1(n5409), .B2(n5870), .ZN(n5216)
         );
  AOI21_X1 U6346 ( .B1(n5845), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5216), 
        .ZN(n5217) );
  OAI21_X1 U6347 ( .B1(n5267), .B2(n5861), .A(n5217), .ZN(n5218) );
  AOI21_X1 U6348 ( .B1(n5219), .B2(n5654), .A(n5218), .ZN(n5220) );
  OAI21_X1 U6349 ( .B1(n5407), .B2(n5810), .A(n5220), .ZN(U2807) );
  OAI21_X1 U6350 ( .B1(n5221), .B2(n5224), .A(n5223), .ZN(n5440) );
  INV_X1 U6351 ( .A(n5281), .ZN(n5225) );
  AOI21_X1 U6352 ( .B1(n5226), .B2(n5293), .A(n5225), .ZN(n5686) );
  AOI22_X1 U6353 ( .A1(EBX_REG_17__SCAN_IN), .A2(n5848), .B1(n5437), .B2(n4892), .ZN(n5227) );
  OAI211_X1 U6354 ( .C1(n5856), .C2(n5435), .A(n5227), .B(n5826), .ZN(n5233)
         );
  INV_X1 U6355 ( .A(n5764), .ZN(n5229) );
  NOR2_X1 U6356 ( .A1(n5229), .A2(n5228), .ZN(n5755) );
  OAI21_X1 U6357 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5230), .A(n5755), .ZN(n5231) );
  INV_X1 U6358 ( .A(n5231), .ZN(n5232) );
  AOI211_X1 U6359 ( .C1(n5686), .C2(n5825), .A(n5233), .B(n5232), .ZN(n5234)
         );
  OAI21_X1 U6360 ( .B1(n5440), .B2(n5810), .A(n5234), .ZN(U2810) );
  INV_X1 U6361 ( .A(n5235), .ZN(n5236) );
  AOI21_X1 U6362 ( .B1(n5237), .B2(n5078), .A(n5236), .ZN(n5454) );
  INV_X1 U6363 ( .A(n5454), .ZN(n5324) );
  OAI21_X1 U6364 ( .B1(n5856), .B2(n5238), .A(n5826), .ZN(n5240) );
  NAND2_X1 U6365 ( .A1(n5764), .A2(n5763), .ZN(n5776) );
  OAI22_X1 U6366 ( .A1(n5297), .A2(n5858), .B1(n5765), .B2(n5776), .ZN(n5239)
         );
  AOI211_X1 U6367 ( .C1(n5766), .C2(n5765), .A(n5240), .B(n5239), .ZN(n5246)
         );
  AND2_X1 U6368 ( .A1(n5242), .A2(n5241), .ZN(n5243) );
  NOR2_X1 U6369 ( .A1(n5291), .A2(n5243), .ZN(n5697) );
  INV_X1 U6370 ( .A(n5452), .ZN(n5244) );
  AOI22_X1 U6371 ( .A1(n5697), .A2(n5825), .B1(n4892), .B2(n5244), .ZN(n5245)
         );
  OAI211_X1 U6372 ( .C1(n5324), .C2(n5810), .A(n5246), .B(n5245), .ZN(U2812)
         );
  INV_X1 U6373 ( .A(n5490), .ZN(n5248) );
  OAI22_X1 U6374 ( .A1(n5248), .A2(n5872), .B1(n5878), .B2(n5247), .ZN(U2828)
         );
  AOI22_X1 U6375 ( .A1(n5509), .A2(n3996), .B1(EBX_REG_29__SCAN_IN), .B2(n5286), .ZN(n5249) );
  OAI21_X1 U6376 ( .B1(n5328), .B2(n5300), .A(n5249), .ZN(U2830) );
  OAI222_X1 U6377 ( .A1(n5300), .A2(n5305), .B1(n6630), .B2(n5878), .C1(n5516), 
        .C2(n5872), .ZN(U2831) );
  OAI222_X1 U6378 ( .A1(n5311), .A2(n5300), .B1(n5250), .B2(n5878), .C1(n5872), 
        .C2(n5533), .ZN(U2833) );
  INV_X1 U6379 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5251) );
  OAI222_X1 U6380 ( .A1(n5365), .A2(n5300), .B1(n5251), .B2(n5878), .C1(n5539), 
        .C2(n5872), .ZN(U2834) );
  AOI22_X1 U6381 ( .A1(n5551), .A2(n3996), .B1(EBX_REG_24__SCAN_IN), .B2(n5286), .ZN(n5252) );
  OAI21_X1 U6382 ( .B1(n5377), .B2(n5300), .A(n5252), .ZN(U2835) );
  XOR2_X1 U6383 ( .A(n5254), .B(n5253), .Z(n5389) );
  INV_X1 U6384 ( .A(n5389), .ZN(n5638) );
  INV_X1 U6385 ( .A(n5573), .ZN(n5256) );
  AOI21_X1 U6386 ( .B1(n5256), .B2(n5264), .A(n5255), .ZN(n5259) );
  INV_X1 U6387 ( .A(n5257), .ZN(n5258) );
  NOR2_X1 U6388 ( .A1(n5259), .A2(n5258), .ZN(n5640) );
  AOI22_X1 U6389 ( .A1(n5640), .A2(n3996), .B1(EBX_REG_23__SCAN_IN), .B2(n5286), .ZN(n5260) );
  OAI21_X1 U6390 ( .B1(n5638), .B2(n5300), .A(n5260), .ZN(U2836) );
  INV_X1 U6391 ( .A(n5253), .ZN(n5262) );
  AOI21_X1 U6392 ( .B1(n5263), .B2(n5261), .A(n5262), .ZN(n5672) );
  INV_X1 U6393 ( .A(n5672), .ZN(n5266) );
  XNOR2_X1 U6394 ( .A(n5573), .B(n5264), .ZN(n5647) );
  AOI22_X1 U6395 ( .A1(n5647), .A2(n3996), .B1(EBX_REG_22__SCAN_IN), .B2(n5286), .ZN(n5265) );
  OAI21_X1 U6396 ( .B1(n5266), .B2(n5300), .A(n5265), .ZN(U2837) );
  OAI222_X1 U6397 ( .A1(n5407), .A2(n5300), .B1(n5878), .B2(n3956), .C1(n5267), 
        .C2(n5872), .ZN(U2839) );
  AND2_X1 U6398 ( .A1(n5268), .A2(n5269), .ZN(n5270) );
  OR2_X1 U6399 ( .A1(n5270), .A2(n2964), .ZN(n5664) );
  INV_X1 U6400 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5277) );
  INV_X1 U6401 ( .A(n5271), .ZN(n5275) );
  INV_X1 U6402 ( .A(n5272), .ZN(n5273) );
  AOI22_X1 U6403 ( .A1(n5275), .A2(n5274), .B1(n5273), .B2(n5284), .ZN(n5282)
         );
  NOR2_X1 U6404 ( .A1(n5281), .A2(n5282), .ZN(n5280) );
  XOR2_X1 U6405 ( .A(n5276), .B(n5280), .Z(n5668) );
  OAI222_X1 U6406 ( .A1(n5664), .A2(n5300), .B1(n5878), .B2(n5277), .C1(n5872), 
        .C2(n5668), .ZN(U2840) );
  INV_X1 U6407 ( .A(n5268), .ZN(n5278) );
  AOI21_X1 U6408 ( .B1(n5279), .B2(n5223), .A(n5278), .ZN(n5879) );
  INV_X1 U6409 ( .A(n5879), .ZN(n5285) );
  AOI21_X1 U6410 ( .B1(n5282), .B2(n5281), .A(n5280), .ZN(n5759) );
  INV_X1 U6411 ( .A(n5759), .ZN(n5283) );
  OAI222_X1 U6412 ( .A1(n5285), .A2(n5300), .B1(n5284), .B2(n5878), .C1(n5872), 
        .C2(n5283), .ZN(U2841) );
  AOI22_X1 U6413 ( .A1(n5686), .A2(n3996), .B1(EBX_REG_17__SCAN_IN), .B2(n5286), .ZN(n5287) );
  OAI21_X1 U6414 ( .B1(n5440), .B2(n5300), .A(n5287), .ZN(U2842) );
  AND2_X1 U6415 ( .A1(n5235), .A2(n5288), .ZN(n5289) );
  NOR2_X1 U6416 ( .A1(n5221), .A2(n5289), .ZN(n5884) );
  OR2_X1 U6417 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  NAND2_X1 U6418 ( .A1(n5293), .A2(n5292), .ZN(n5774) );
  OAI22_X1 U6419 ( .A1(n5774), .A2(n5872), .B1(n5294), .B2(n5878), .ZN(n5295)
         );
  AOI21_X1 U6420 ( .B1(n5884), .B2(n3900), .A(n5295), .ZN(n5296) );
  INV_X1 U6421 ( .A(n5296), .ZN(U2843) );
  NOR2_X1 U6422 ( .A1(n5878), .A2(n5297), .ZN(n5298) );
  AOI21_X1 U6423 ( .B1(n5697), .B2(n3996), .A(n5298), .ZN(n5299) );
  OAI21_X1 U6424 ( .B1(n5324), .B2(n5300), .A(n5299), .ZN(U2844) );
  AOI22_X1 U6425 ( .A1(n5882), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5885), .ZN(n5302) );
  NAND2_X1 U6426 ( .A1(n5886), .A2(DATAI_13_), .ZN(n5301) );
  OAI211_X1 U6427 ( .C1(n5328), .C2(n5671), .A(n5302), .B(n5301), .ZN(U2862)
         );
  AOI22_X1 U6428 ( .A1(n5882), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5885), .ZN(n5304) );
  NAND2_X1 U6429 ( .A1(n5886), .A2(DATAI_12_), .ZN(n5303) );
  OAI211_X1 U6430 ( .C1(n5305), .C2(n5671), .A(n5304), .B(n5303), .ZN(U2863)
         );
  AOI22_X1 U6431 ( .A1(n5882), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5885), .ZN(n5307) );
  NAND2_X1 U6432 ( .A1(n5886), .A2(DATAI_11_), .ZN(n5306) );
  OAI211_X1 U6433 ( .C1(n5308), .C2(n5671), .A(n5307), .B(n5306), .ZN(U2864)
         );
  AOI22_X1 U6434 ( .A1(n5882), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5885), .ZN(n5310) );
  NAND2_X1 U6435 ( .A1(n5886), .A2(DATAI_10_), .ZN(n5309) );
  OAI211_X1 U6436 ( .C1(n5311), .C2(n5671), .A(n5310), .B(n5309), .ZN(U2865)
         );
  AOI22_X1 U6437 ( .A1(n5882), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5885), .ZN(n5313) );
  NAND2_X1 U6438 ( .A1(n5886), .A2(DATAI_9_), .ZN(n5312) );
  OAI211_X1 U6439 ( .C1(n5365), .C2(n5671), .A(n5313), .B(n5312), .ZN(U2866)
         );
  AOI22_X1 U6440 ( .A1(n5882), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5885), .ZN(n5315) );
  NAND2_X1 U6441 ( .A1(n5886), .A2(DATAI_8_), .ZN(n5314) );
  OAI211_X1 U6442 ( .C1(n5377), .C2(n5671), .A(n5315), .B(n5314), .ZN(U2867)
         );
  AOI22_X1 U6443 ( .A1(n5886), .A2(DATAI_7_), .B1(n5885), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6444 ( .A1(n5882), .A2(DATAI_23_), .ZN(n5316) );
  OAI211_X1 U6445 ( .C1(n5638), .C2(n5671), .A(n5317), .B(n5316), .ZN(U2868)
         );
  AOI22_X1 U6446 ( .A1(n5886), .A2(DATAI_3_), .B1(n5885), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6447 ( .A1(n5882), .A2(DATAI_19_), .ZN(n5318) );
  OAI211_X1 U6448 ( .C1(n5664), .C2(n5671), .A(n5319), .B(n5318), .ZN(U2872)
         );
  AOI22_X1 U6449 ( .A1(n5882), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5885), .ZN(n5321) );
  NAND2_X1 U6450 ( .A1(n5886), .A2(DATAI_1_), .ZN(n5320) );
  OAI211_X1 U6451 ( .C1(n5440), .C2(n5671), .A(n5321), .B(n5320), .ZN(U2874)
         );
  AOI22_X1 U6452 ( .A1(n5322), .A2(DATAI_15_), .B1(n5885), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5323) );
  OAI21_X1 U6453 ( .B1(n5324), .B2(n5671), .A(n5323), .ZN(U2876) );
  INV_X1 U6454 ( .A(n4251), .ZN(n5334) );
  OAI21_X1 U6455 ( .B1(n5334), .B2(n5326), .A(n5325), .ZN(n5327) );
  XNOR2_X1 U6456 ( .A(n5327), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5511)
         );
  INV_X1 U6457 ( .A(n5328), .ZN(n5332) );
  AND2_X1 U6458 ( .A1(n6095), .A2(REIP_REG_29__SCAN_IN), .ZN(n5504) );
  AOI21_X1 U6459 ( .B1(n6006), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5504), 
        .ZN(n5329) );
  OAI21_X1 U6460 ( .B1(n6015), .B2(n5330), .A(n5329), .ZN(n5331) );
  AOI21_X1 U6461 ( .B1(n5332), .B2(n5446), .A(n5331), .ZN(n5333) );
  OAI21_X1 U6462 ( .B1(n5511), .B2(n5992), .A(n5333), .ZN(U2957) );
  NAND3_X1 U6463 ( .A1(n5334), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n4226), .ZN(n5338) );
  INV_X1 U6464 ( .A(n5336), .ZN(n5337) );
  OR3_X1 U6465 ( .A1(n5335), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n5337), 
        .ZN(n5346) );
  AOI22_X1 U6466 ( .A1(n5338), .A2(n5346), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5529), .ZN(n5339) );
  XNOR2_X1 U6467 ( .A(n5339), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5520)
         );
  AND2_X1 U6468 ( .A1(n6095), .A2(REIP_REG_28__SCAN_IN), .ZN(n5515) );
  AOI21_X1 U6469 ( .B1(n6006), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5515), 
        .ZN(n5340) );
  OAI21_X1 U6470 ( .B1(n6015), .B2(n5341), .A(n5340), .ZN(n5342) );
  AOI21_X1 U6471 ( .B1(n5343), .B2(n5446), .A(n5342), .ZN(n5344) );
  OAI21_X1 U6472 ( .B1(n5992), .B2(n5520), .A(n5344), .ZN(U2958) );
  INV_X1 U6473 ( .A(n5345), .ZN(n5347) );
  NAND2_X1 U6474 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  XNOR2_X1 U6475 ( .A(n5348), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5528)
         );
  INV_X1 U6476 ( .A(n5349), .ZN(n5351) );
  AND2_X1 U6477 ( .A1(n6095), .A2(REIP_REG_27__SCAN_IN), .ZN(n5522) );
  AOI21_X1 U6478 ( .B1(n6006), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5522), 
        .ZN(n5350) );
  OAI21_X1 U6479 ( .B1(n6015), .B2(n5351), .A(n5350), .ZN(n5352) );
  AOI21_X1 U6480 ( .B1(n5353), .B2(n5446), .A(n5352), .ZN(n5354) );
  OAI21_X1 U6481 ( .B1(n5528), .B2(n5992), .A(n5354), .ZN(U2959) );
  XNOR2_X1 U6482 ( .A(n4226), .B(n5529), .ZN(n5355) );
  XNOR2_X1 U6483 ( .A(n4251), .B(n5355), .ZN(n5537) );
  AND2_X1 U6484 ( .A1(n6095), .A2(REIP_REG_26__SCAN_IN), .ZN(n5531) );
  AOI21_X1 U6485 ( .B1(n6006), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5531), 
        .ZN(n5356) );
  OAI21_X1 U6486 ( .B1(n6015), .B2(n5357), .A(n5356), .ZN(n5358) );
  AOI21_X1 U6487 ( .B1(n5359), .B2(n5446), .A(n5358), .ZN(n5360) );
  OAI21_X1 U6488 ( .B1(n5992), .B2(n5537), .A(n5360), .ZN(U2960) );
  INV_X1 U6489 ( .A(n5361), .ZN(n5362) );
  AOI21_X1 U6490 ( .B1(n5363), .B2(n5335), .A(n5362), .ZN(n5545) );
  INV_X1 U6491 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6492 ( .A1(n6095), .A2(REIP_REG_25__SCAN_IN), .ZN(n5538) );
  OAI21_X1 U6493 ( .B1(n5461), .B2(n5364), .A(n5538), .ZN(n5367) );
  NOR2_X1 U6494 ( .A1(n5365), .A2(n5987), .ZN(n5366) );
  AOI211_X1 U6495 ( .C1(n5464), .C2(n5368), .A(n5367), .B(n5366), .ZN(n5369)
         );
  OAI21_X1 U6496 ( .B1(n5545), .B2(n5992), .A(n5369), .ZN(U2961) );
  INV_X1 U6497 ( .A(n5412), .ZN(n5370) );
  INV_X1 U6498 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U6499 ( .A1(n5370), .A2(n5609), .ZN(n5373) );
  INV_X1 U6500 ( .A(n5371), .ZN(n5372) );
  AOI22_X2 U6501 ( .A1(n5373), .A2(n2953), .B1(n5372), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5406) );
  XNOR2_X1 U6502 ( .A(n2953), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5405)
         );
  INV_X1 U6503 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5599) );
  OAI22_X2 U6504 ( .A1(n5406), .A2(n5405), .B1(n4226), .B2(n5599), .ZN(n5398)
         );
  XNOR2_X1 U6505 ( .A(n2953), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5399)
         );
  NOR2_X1 U6507 ( .A1(n4226), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5391)
         );
  NAND2_X1 U6508 ( .A1(n5397), .A2(n5391), .ZN(n5383) );
  NAND3_X1 U6509 ( .A1(n4226), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5375) );
  INV_X1 U6510 ( .A(n5397), .ZN(n5374) );
  OAI22_X1 U6511 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5375), .B2(n5393), .ZN(n5376) );
  XNOR2_X1 U6512 ( .A(n5376), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5553)
         );
  INV_X1 U6513 ( .A(n5377), .ZN(n5381) );
  NOR2_X1 U6514 ( .A1(n6032), .A2(n6487), .ZN(n5550) );
  AOI21_X1 U6515 ( .B1(n6006), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5550), 
        .ZN(n5378) );
  OAI21_X1 U6516 ( .B1(n6015), .B2(n5379), .A(n5378), .ZN(n5380) );
  AOI21_X1 U6517 ( .B1(n5381), .B2(n5446), .A(n5380), .ZN(n5382) );
  OAI21_X1 U6518 ( .B1(n5553), .B2(n5992), .A(n5382), .ZN(U2962) );
  INV_X1 U6519 ( .A(n5474), .ZN(n5563) );
  NAND3_X1 U6520 ( .A1(n4226), .A2(n5563), .A3(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5384) );
  OAI21_X1 U6521 ( .B1(n5406), .B2(n5384), .A(n5383), .ZN(n5385) );
  XNOR2_X1 U6522 ( .A(n5385), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5561)
         );
  INV_X1 U6523 ( .A(n5635), .ZN(n5387) );
  NAND2_X1 U6524 ( .A1(n6095), .A2(REIP_REG_23__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U6525 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5386)
         );
  OAI211_X1 U6526 ( .C1(n6015), .C2(n5387), .A(n5555), .B(n5386), .ZN(n5388)
         );
  AOI21_X1 U6527 ( .B1(n5389), .B2(n5446), .A(n5388), .ZN(n5390) );
  OAI21_X1 U6528 ( .B1(n5561), .B2(n5992), .A(n5390), .ZN(U2963) );
  AOI21_X1 U6529 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4226), .A(n5391), 
        .ZN(n5392) );
  XNOR2_X1 U6530 ( .A(n5393), .B(n5392), .ZN(n5569) );
  AND2_X1 U6531 ( .A1(n6095), .A2(REIP_REG_22__SCAN_IN), .ZN(n5566) );
  AOI21_X1 U6532 ( .B1(n6006), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5566), 
        .ZN(n5394) );
  OAI21_X1 U6533 ( .B1(n6015), .B2(n5644), .A(n5394), .ZN(n5395) );
  AOI21_X1 U6534 ( .B1(n5672), .B2(n5446), .A(n5395), .ZN(n5396) );
  OAI21_X1 U6535 ( .B1(n5569), .B2(n5992), .A(n5396), .ZN(U2964) );
  AOI21_X1 U6536 ( .B1(n5399), .B2(n5398), .A(n5397), .ZN(n5582) );
  XOR2_X1 U6537 ( .A(n5400), .B(n5209), .Z(n5675) );
  INV_X1 U6538 ( .A(n5655), .ZN(n5402) );
  NAND2_X1 U6539 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5401)
         );
  NAND2_X1 U6540 ( .A1(n6095), .A2(REIP_REG_21__SCAN_IN), .ZN(n5575) );
  OAI211_X1 U6541 ( .C1(n6015), .C2(n5402), .A(n5401), .B(n5575), .ZN(n5403)
         );
  AOI21_X1 U6542 ( .B1(n5675), .B2(n5446), .A(n5403), .ZN(n5404) );
  OAI21_X1 U6543 ( .B1(n5582), .B2(n5992), .A(n5404), .ZN(U2965) );
  XNOR2_X1 U6544 ( .A(n5406), .B(n5405), .ZN(n5600) );
  INV_X1 U6545 ( .A(n5407), .ZN(n5678) );
  NAND2_X1 U6546 ( .A1(n6095), .A2(REIP_REG_20__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U6547 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5408)
         );
  OAI211_X1 U6548 ( .C1(n5409), .C2(n6015), .A(n5597), .B(n5408), .ZN(n5410)
         );
  AOI21_X1 U6549 ( .B1(n5678), .B2(n5446), .A(n5410), .ZN(n5411) );
  OAI21_X1 U6550 ( .B1(n5600), .B2(n5992), .A(n5411), .ZN(U2966) );
  XNOR2_X1 U6551 ( .A(n4226), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5413)
         );
  XNOR2_X1 U6552 ( .A(n5412), .B(n5413), .ZN(n5612) );
  NAND2_X1 U6553 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5414)
         );
  NAND2_X1 U6554 ( .A1(n6095), .A2(REIP_REG_19__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U6555 ( .A1(n5414), .A2(n5605), .ZN(n5415) );
  AOI21_X1 U6556 ( .B1(n5660), .B2(n5464), .A(n5415), .ZN(n5418) );
  INV_X1 U6557 ( .A(n5664), .ZN(n5416) );
  NAND2_X1 U6558 ( .A1(n5416), .A2(n5446), .ZN(n5417) );
  OAI211_X1 U6559 ( .C1(n5612), .C2(n5992), .A(n5418), .B(n5417), .ZN(U2967)
         );
  NAND3_X1 U6560 ( .A1(n5419), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n4226), .ZN(n5430) );
  NOR2_X1 U6561 ( .A1(n4226), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5426)
         );
  NAND4_X1 U6562 ( .A1(n5421), .A2(n5426), .A3(n5617), .A4(n5420), .ZN(n5431)
         );
  NAND2_X1 U6563 ( .A1(n5430), .A2(n5431), .ZN(n5422) );
  XNOR2_X1 U6564 ( .A(n5422), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5621)
         );
  NAND2_X1 U6565 ( .A1(n6095), .A2(REIP_REG_18__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U6566 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5423)
         );
  OAI211_X1 U6567 ( .C1(n5757), .C2(n6015), .A(n5614), .B(n5423), .ZN(n5424)
         );
  AOI21_X1 U6568 ( .B1(n5879), .B2(n5446), .A(n5424), .ZN(n5425) );
  OAI21_X1 U6569 ( .B1(n5621), .B2(n5992), .A(n5425), .ZN(U2968) );
  INV_X1 U6570 ( .A(n5419), .ZN(n5427) );
  AOI21_X1 U6571 ( .B1(n5427), .B2(n5426), .A(n5617), .ZN(n5428) );
  AOI21_X1 U6572 ( .B1(n5419), .B2(n4226), .A(n5428), .ZN(n5433) );
  INV_X1 U6573 ( .A(n5430), .ZN(n5432) );
  OAI21_X1 U6574 ( .B1(n5433), .B2(n5432), .A(n5431), .ZN(n5687) );
  NAND2_X1 U6575 ( .A1(n5687), .A2(n6011), .ZN(n5439) );
  INV_X1 U6576 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5434) );
  OAI22_X1 U6577 ( .A1(n5461), .A2(n5435), .B1(n6032), .B2(n5434), .ZN(n5436)
         );
  AOI21_X1 U6578 ( .B1(n5464), .B2(n5437), .A(n5436), .ZN(n5438) );
  OAI211_X1 U6579 ( .C1(n5987), .C2(n5440), .A(n5439), .B(n5438), .ZN(U2969)
         );
  XNOR2_X1 U6580 ( .A(n4226), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5442)
         );
  XNOR2_X1 U6581 ( .A(n5441), .B(n5442), .ZN(n5693) );
  AOI22_X1 U6582 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6095), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5443) );
  OAI21_X1 U6583 ( .B1(n6015), .B2(n5444), .A(n5443), .ZN(n5445) );
  AOI21_X1 U6584 ( .B1(n5884), .B2(n5446), .A(n5445), .ZN(n5447) );
  OAI21_X1 U6585 ( .B1(n5693), .B2(n5992), .A(n5447), .ZN(U2970) );
  NAND2_X1 U6586 ( .A1(n3037), .A2(n5449), .ZN(n5450) );
  XNOR2_X1 U6587 ( .A(n5448), .B(n5450), .ZN(n5698) );
  INV_X1 U6588 ( .A(n5698), .ZN(n5456) );
  AOI22_X1 U6589 ( .A1(n6006), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6095), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5451) );
  OAI21_X1 U6590 ( .B1(n6015), .B2(n5452), .A(n5451), .ZN(n5453) );
  AOI21_X1 U6591 ( .B1(n5454), .B2(n5446), .A(n5453), .ZN(n5455) );
  OAI21_X1 U6592 ( .B1(n5456), .B2(n5992), .A(n5455), .ZN(U2971) );
  XNOR2_X1 U6593 ( .A(n4226), .B(n5458), .ZN(n5459) );
  XNOR2_X1 U6594 ( .A(n5457), .B(n5459), .ZN(n5713) );
  INV_X1 U6595 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5460) );
  OAI22_X1 U6596 ( .A1(n5461), .A2(n5460), .B1(n6032), .B2(n6473), .ZN(n5463)
         );
  NOR2_X1 U6597 ( .A1(n5779), .A2(n5987), .ZN(n5462) );
  AOI211_X1 U6598 ( .C1(n5464), .C2(n5780), .A(n5463), .B(n5462), .ZN(n5465)
         );
  OAI21_X1 U6599 ( .B1(n5992), .B2(n5713), .A(n5465), .ZN(U2972) );
  NAND3_X1 U6600 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5712) );
  NOR2_X1 U6601 ( .A1(n5458), .A2(n5712), .ZN(n5692) );
  INV_X1 U6602 ( .A(n5692), .ZN(n5466) );
  NOR2_X1 U6603 ( .A1(n6016), .A2(n5466), .ZN(n5701) );
  NAND3_X1 U6604 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5701), .ZN(n5690) );
  NAND4_X1 U6605 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_19__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5470) );
  AND2_X1 U6606 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6607 ( .A1(n5543), .A2(n5479), .ZN(n5525) );
  INV_X1 U6608 ( .A(n5512), .ZN(n5482) );
  NOR2_X1 U6609 ( .A1(n5525), .A2(n5482), .ZN(n5503) );
  NOR2_X1 U6610 ( .A1(n5484), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5489)
         );
  NAND3_X1 U6611 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5692), .ZN(n5584) );
  NOR2_X1 U6612 ( .A1(n5584), .A2(n5468), .ZN(n5586) );
  INV_X1 U6613 ( .A(n5586), .ZN(n5469) );
  NOR2_X1 U6614 ( .A1(n5470), .A2(n5469), .ZN(n5473) );
  NOR3_X1 U6615 ( .A1(n5705), .A2(n5584), .A3(n5470), .ZN(n5471) );
  OR2_X1 U6616 ( .A1(n6030), .A2(n5471), .ZN(n5472) );
  OAI211_X1 U6617 ( .C1(n5473), .C2(n6099), .A(n6025), .B(n5472), .ZN(n5574)
         );
  AND2_X1 U6618 ( .A1(n6031), .A2(n5474), .ZN(n5475) );
  OR2_X1 U6619 ( .A1(n5574), .A2(n5475), .ZN(n5554) );
  INV_X1 U6620 ( .A(n5476), .ZN(n5477) );
  AOI21_X1 U6621 ( .B1(n5583), .B2(n6099), .A(n5477), .ZN(n5478) );
  NOR2_X1 U6622 ( .A1(n5554), .A2(n5478), .ZN(n5546) );
  INV_X1 U6623 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U6624 ( .A1(n6031), .A2(n5480), .ZN(n5481) );
  NAND2_X1 U6625 ( .A1(n5546), .A2(n5481), .ZN(n5523) );
  AND2_X1 U6626 ( .A1(n6031), .A2(n5482), .ZN(n5483) );
  OR2_X1 U6627 ( .A1(n5523), .A2(n5483), .ZN(n5505) );
  OAI21_X1 U6628 ( .B1(n5505), .B2(n5484), .A(n6031), .ZN(n5486) );
  AOI21_X1 U6629 ( .B1(n5486), .B2(n5546), .A(n5485), .ZN(n5487) );
  AOI211_X1 U6630 ( .C1(n5503), .C2(n5489), .A(n5488), .B(n5487), .ZN(n5492)
         );
  NAND2_X1 U6631 ( .A1(n5490), .A2(n6097), .ZN(n5491) );
  OAI211_X1 U6632 ( .C1(n5493), .C2(n6086), .A(n5492), .B(n5491), .ZN(U2987)
         );
  AOI21_X1 U6633 ( .B1(n5503), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5498) );
  INV_X1 U6634 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5495) );
  AOI211_X1 U6635 ( .C1(n5495), .C2(n6031), .A(n5494), .B(n5505), .ZN(n5497)
         );
  OAI21_X1 U6636 ( .B1(n5498), .B2(n5497), .A(n5496), .ZN(n5499) );
  AOI21_X1 U6637 ( .B1(n5500), .B2(n6097), .A(n5499), .ZN(n5501) );
  OAI21_X1 U6638 ( .B1(n5502), .B2(n6086), .A(n5501), .ZN(U2988) );
  INV_X1 U6639 ( .A(n5503), .ZN(n5507) );
  AOI21_X1 U6640 ( .B1(n5505), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5504), 
        .ZN(n5506) );
  OAI21_X1 U6641 ( .B1(n5507), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5506), 
        .ZN(n5508) );
  AOI21_X1 U6642 ( .B1(n5509), .B2(n6097), .A(n5508), .ZN(n5510) );
  OAI21_X1 U6643 ( .B1(n5511), .B2(n6086), .A(n5510), .ZN(U2989) );
  NOR3_X1 U6644 ( .A1(n5525), .A2(n5513), .A3(n5512), .ZN(n5514) );
  AOI211_X1 U6645 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5523), .A(n5515), .B(n5514), .ZN(n5519) );
  INV_X1 U6646 ( .A(n5516), .ZN(n5517) );
  NAND2_X1 U6647 ( .A1(n5517), .A2(n6097), .ZN(n5518) );
  OAI211_X1 U6648 ( .C1(n5520), .C2(n6086), .A(n5519), .B(n5518), .ZN(U2990)
         );
  AOI21_X1 U6649 ( .B1(n5523), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5522), 
        .ZN(n5524) );
  OAI21_X1 U6650 ( .B1(n5525), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5524), 
        .ZN(n5526) );
  AOI21_X1 U6651 ( .B1(n3997), .B2(n6097), .A(n5526), .ZN(n5527) );
  OAI21_X1 U6652 ( .B1(n5528), .B2(n6086), .A(n5527), .ZN(U2991) );
  XNOR2_X1 U6653 ( .A(n5542), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5532)
         );
  NOR2_X1 U6654 ( .A1(n5546), .A2(n5529), .ZN(n5530) );
  AOI211_X1 U6655 ( .C1(n5543), .C2(n5532), .A(n5531), .B(n5530), .ZN(n5536)
         );
  INV_X1 U6656 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U6657 ( .A1(n5534), .A2(n6097), .ZN(n5535) );
  OAI211_X1 U6658 ( .C1(n5537), .C2(n6086), .A(n5536), .B(n5535), .ZN(U2992)
         );
  OAI21_X1 U6659 ( .B1(n5546), .B2(n5542), .A(n5538), .ZN(n5541) );
  NOR2_X1 U6660 ( .A1(n5539), .A2(n6079), .ZN(n5540) );
  AOI211_X1 U6661 ( .C1(n5543), .C2(n5542), .A(n5541), .B(n5540), .ZN(n5544)
         );
  OAI21_X1 U6662 ( .B1(n5545), .B2(n6086), .A(n5544), .ZN(U2993) );
  NAND3_X1 U6663 ( .A1(n5579), .A2(n5563), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5548) );
  AOI21_X1 U6664 ( .B1(n5548), .B2(n5547), .A(n5546), .ZN(n5549) );
  AOI211_X1 U6665 ( .C1(n5551), .C2(n6097), .A(n5550), .B(n5549), .ZN(n5552)
         );
  OAI21_X1 U6666 ( .B1(n5553), .B2(n6086), .A(n5552), .ZN(U2994) );
  INV_X1 U6667 ( .A(n5554), .ZN(n5556) );
  OAI21_X1 U6668 ( .B1(n5556), .B2(n5558), .A(n5555), .ZN(n5557) );
  AOI21_X1 U6669 ( .B1(n5640), .B2(n6097), .A(n5557), .ZN(n5560) );
  NAND3_X1 U6670 ( .A1(n5579), .A2(n5563), .A3(n5558), .ZN(n5559) );
  OAI211_X1 U6671 ( .C1(n5561), .C2(n6086), .A(n5560), .B(n5559), .ZN(U2995)
         );
  INV_X1 U6672 ( .A(n5579), .ZN(n5564) );
  NOR3_X1 U6673 ( .A1(n5564), .A2(n5563), .A3(n5562), .ZN(n5565) );
  AOI211_X1 U6674 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5574), .A(n5566), .B(n5565), .ZN(n5568) );
  NAND2_X1 U6675 ( .A1(n5647), .A2(n6097), .ZN(n5567) );
  OAI211_X1 U6676 ( .C1(n5569), .C2(n6086), .A(n5568), .B(n5567), .ZN(U2996)
         );
  OR2_X1 U6677 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  AND2_X1 U6678 ( .A1(n5573), .A2(n5572), .ZN(n5669) );
  NAND2_X1 U6679 ( .A1(n5574), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U6680 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  AOI21_X1 U6681 ( .B1(n5669), .B2(n6097), .A(n5577), .ZN(n5581) );
  INV_X1 U6682 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U6683 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  OAI211_X1 U6684 ( .C1(n5582), .C2(n6086), .A(n5581), .B(n5580), .ZN(U2997)
         );
  NOR2_X1 U6685 ( .A1(n5583), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5591)
         );
  INV_X1 U6686 ( .A(n5584), .ZN(n5585) );
  OR2_X1 U6687 ( .A1(n6030), .A2(n5585), .ZN(n5590) );
  NAND2_X1 U6688 ( .A1(n5586), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5588) );
  AOI21_X1 U6689 ( .B1(n6074), .B2(n5588), .A(n5587), .ZN(n5589) );
  NAND2_X1 U6690 ( .A1(n5590), .A2(n5589), .ZN(n5685) );
  OR2_X1 U6691 ( .A1(n5591), .A2(n5685), .ZN(n5613) );
  AND2_X1 U6692 ( .A1(n6031), .A2(n5615), .ZN(n5592) );
  NOR2_X1 U6693 ( .A1(n5613), .A2(n5592), .ZN(n5606) );
  NOR2_X1 U6694 ( .A1(n5690), .A2(n5593), .ZN(n5610) );
  NOR2_X1 U6695 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  NAND2_X1 U6696 ( .A1(n5610), .A2(n5596), .ZN(n5598) );
  OAI211_X1 U6697 ( .C1(n5606), .C2(n5599), .A(n5598), .B(n5597), .ZN(n5602)
         );
  NOR2_X1 U6698 ( .A1(n5600), .A2(n6086), .ZN(n5601) );
  AOI211_X1 U6699 ( .C1(n6097), .C2(n5603), .A(n5602), .B(n5601), .ZN(n5604)
         );
  INV_X1 U6700 ( .A(n5604), .ZN(U2998) );
  OAI21_X1 U6701 ( .B1(n5606), .B2(n5609), .A(n5605), .ZN(n5608) );
  NOR2_X1 U6702 ( .A1(n5668), .A2(n6079), .ZN(n5607) );
  AOI211_X1 U6703 ( .C1(n5610), .C2(n5609), .A(n5608), .B(n5607), .ZN(n5611)
         );
  OAI21_X1 U6704 ( .B1(n5612), .B2(n6086), .A(n5611), .ZN(U2999) );
  INV_X1 U6705 ( .A(n5613), .ZN(n5616) );
  OAI21_X1 U6706 ( .B1(n5616), .B2(n5615), .A(n5614), .ZN(n5619) );
  NOR3_X1 U6707 ( .A1(n5690), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5617), 
        .ZN(n5618) );
  AOI211_X1 U6708 ( .C1(n6097), .C2(n5759), .A(n5619), .B(n5618), .ZN(n5620)
         );
  OAI21_X1 U6709 ( .B1(n5621), .B2(n6086), .A(n5620), .ZN(U3000) );
  INV_X1 U6710 ( .A(n5630), .ZN(n6219) );
  OAI211_X1 U6711 ( .C1(n5622), .C2(STATEBS16_REG_SCAN_IN), .A(n6219), .B(
        n6218), .ZN(n5623) );
  OAI21_X1 U6712 ( .B1(n5626), .B2(n5624), .A(n5623), .ZN(n5625) );
  MUX2_X1 U6713 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5625), .S(n6108), 
        .Z(U3464) );
  OAI21_X1 U6714 ( .B1(n6219), .B2(n4518), .A(n6218), .ZN(n5633) );
  NOR2_X1 U6715 ( .A1(n5630), .A2(n6112), .ZN(n5627) );
  OAI22_X1 U6716 ( .A1(n5633), .A2(n5627), .B1(n4315), .B2(n5626), .ZN(n5628)
         );
  MUX2_X1 U6717 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5628), .S(n6108), 
        .Z(U3463) );
  NAND2_X1 U6718 ( .A1(n6146), .A2(n5629), .ZN(n5632) );
  NAND3_X1 U6719 ( .A1(n6217), .A2(n6218), .A3(n5630), .ZN(n5631) );
  OAI211_X1 U6720 ( .C1(n5633), .C2(n6110), .A(n5632), .B(n5631), .ZN(n5634)
         );
  MUX2_X1 U6721 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5634), .S(n6108), 
        .Z(U3462) );
  AOI22_X1 U6722 ( .A1(EBX_REG_23__SCAN_IN), .A2(n5848), .B1(n5635), .B2(n4892), .ZN(n5642) );
  AND2_X1 U6723 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5648), .ZN(n5645) );
  AOI21_X1 U6724 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5645), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5637) );
  OAI22_X1 U6725 ( .A1(n5638), .A2(n5810), .B1(n5637), .B2(n5636), .ZN(n5639)
         );
  AOI21_X1 U6726 ( .B1(n5640), .B2(n5825), .A(n5639), .ZN(n5641) );
  OAI211_X1 U6727 ( .C1(n5643), .C2(n5856), .A(n5642), .B(n5641), .ZN(U2804)
         );
  AOI22_X1 U6728 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5848), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5845), .ZN(n5653) );
  INV_X1 U6729 ( .A(n5644), .ZN(n5646) );
  INV_X1 U6730 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6484) );
  AOI22_X1 U6731 ( .A1(n5646), .A2(n4892), .B1(n5645), .B2(n6484), .ZN(n5652)
         );
  AOI22_X1 U6732 ( .A1(n5672), .A2(n4093), .B1(n5825), .B2(n5647), .ZN(n5651)
         );
  INV_X1 U6733 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U6734 ( .A1(n6480), .A2(n5648), .ZN(n5656) );
  INV_X1 U6735 ( .A(n5656), .ZN(n5649) );
  OAI21_X1 U6736 ( .B1(n5654), .B2(n5649), .A(REIP_REG_22__SCAN_IN), .ZN(n5650) );
  NAND4_X1 U6737 ( .A1(n5653), .A2(n5652), .A3(n5651), .A4(n5650), .ZN(U2805)
         );
  AOI22_X1 U6738 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5848), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5845), .ZN(n5659) );
  AOI22_X1 U6739 ( .A1(n5655), .A2(n4892), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5654), .ZN(n5658) );
  AOI22_X1 U6740 ( .A1(n5675), .A2(n4093), .B1(n5825), .B2(n5669), .ZN(n5657)
         );
  NAND4_X1 U6741 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(U2806)
         );
  AOI22_X1 U6742 ( .A1(n5660), .A2(n4892), .B1(REIP_REG_19__SCAN_IN), .B2(
        n5755), .ZN(n5661) );
  OAI211_X1 U6743 ( .C1(n5856), .C2(n3637), .A(n5661), .B(n5826), .ZN(n5666)
         );
  OAI21_X1 U6744 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5662), .ZN(n5663) );
  OAI22_X1 U6745 ( .A1(n5664), .A2(n5810), .B1(n5663), .B2(n5762), .ZN(n5665)
         );
  AOI211_X1 U6746 ( .C1(EBX_REG_19__SCAN_IN), .C2(n5848), .A(n5666), .B(n5665), 
        .ZN(n5667) );
  OAI21_X1 U6747 ( .B1(n5668), .B2(n5861), .A(n5667), .ZN(U2808) );
  AOI22_X1 U6748 ( .A1(n5675), .A2(n3900), .B1(n3996), .B2(n5669), .ZN(n5670)
         );
  OAI21_X1 U6749 ( .B1(n5878), .B2(n6644), .A(n5670), .ZN(U2838) );
  INV_X1 U6750 ( .A(n5671), .ZN(n5883) );
  AOI22_X1 U6751 ( .A1(n5672), .A2(n5883), .B1(n5882), .B2(DATAI_22_), .ZN(
        n5674) );
  AOI22_X1 U6752 ( .A1(n5886), .A2(DATAI_6_), .B1(n5885), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U6753 ( .A1(n5674), .A2(n5673), .ZN(U2869) );
  AOI22_X1 U6754 ( .A1(n5675), .A2(n5883), .B1(n5882), .B2(DATAI_21_), .ZN(
        n5677) );
  AOI22_X1 U6755 ( .A1(n5886), .A2(DATAI_5_), .B1(n5885), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U6756 ( .A1(n5677), .A2(n5676), .ZN(U2870) );
  AOI22_X1 U6757 ( .A1(n5678), .A2(n5883), .B1(n5882), .B2(DATAI_20_), .ZN(
        n5680) );
  AOI22_X1 U6758 ( .A1(n5886), .A2(DATAI_4_), .B1(n5885), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U6759 ( .A1(n5680), .A2(n5679), .ZN(U2871) );
  AOI22_X1 U6760 ( .A1(n6076), .A2(REIP_REG_13__SCAN_IN), .B1(n6006), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5684) );
  XNOR2_X1 U6761 ( .A(n5681), .B(n5682), .ZN(n5723) );
  AOI22_X1 U6762 ( .A1(n5723), .A2(n6011), .B1(n5446), .B2(n5795), .ZN(n5683)
         );
  OAI211_X1 U6763 ( .C1(n6015), .C2(n5792), .A(n5684), .B(n5683), .ZN(U2973)
         );
  AOI22_X1 U6764 ( .A1(n6076), .A2(REIP_REG_17__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5685), .ZN(n5689) );
  AOI22_X1 U6765 ( .A1(n5687), .A2(n6102), .B1(n6097), .B2(n5686), .ZN(n5688)
         );
  OAI211_X1 U6766 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5690), .A(n5689), .B(n5688), .ZN(U3001) );
  OAI21_X1 U6767 ( .B1(n5692), .B2(n5691), .A(n6024), .ZN(n5700) );
  OAI22_X1 U6768 ( .A1(n5693), .A2(n6086), .B1(n6079), .B2(n5774), .ZN(n5694)
         );
  AOI21_X1 U6769 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n5700), .A(n5694), 
        .ZN(n5696) );
  OAI221_X1 U6770 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5420), .C2(n6595), .A(n5701), 
        .ZN(n5695) );
  OAI211_X1 U6771 ( .C1(n6475), .C2(n6032), .A(n5696), .B(n5695), .ZN(U3002)
         );
  AOI22_X1 U6772 ( .A1(n5698), .A2(n6102), .B1(n6097), .B2(n5697), .ZN(n5703)
         );
  NOR2_X1 U6773 ( .A1(n6032), .A2(n5765), .ZN(n5699) );
  AOI221_X1 U6774 ( .B1(n5701), .B2(n5420), .C1(n5700), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5699), .ZN(n5702) );
  NAND2_X1 U6775 ( .A1(n5703), .A2(n5702), .ZN(U3003) );
  NOR2_X1 U6776 ( .A1(n6022), .A2(n5704), .ZN(n5709) );
  NOR3_X1 U6777 ( .A1(n4386), .A2(n5706), .A3(n5705), .ZN(n5707) );
  AND2_X1 U6778 ( .A1(n4234), .A2(n5709), .ZN(n5718) );
  OAI21_X1 U6779 ( .B1(n5708), .B2(n5707), .A(n5718), .ZN(n5725) );
  OAI211_X1 U6780 ( .C1(n5710), .C2(n5709), .A(n6024), .B(n5725), .ZN(n5711)
         );
  AOI21_X1 U6781 ( .B1(n5719), .B2(n5712), .A(n5711), .ZN(n5726) );
  NOR3_X1 U6782 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6016), .A3(n5712), 
        .ZN(n5715) );
  OAI22_X1 U6783 ( .A1(n5713), .A2(n6086), .B1(n6079), .B2(n5784), .ZN(n5714)
         );
  AOI211_X1 U6784 ( .C1(REIP_REG_14__SCAN_IN), .C2(n6076), .A(n5715), .B(n5714), .ZN(n5716) );
  OAI21_X1 U6785 ( .B1(n5726), .B2(n5458), .A(n5716), .ZN(U3004) );
  NAND2_X1 U6786 ( .A1(n6095), .A2(REIP_REG_13__SCAN_IN), .ZN(n5721) );
  NAND3_X1 U6787 ( .A1(n5719), .A2(n5718), .A3(n5717), .ZN(n5720) );
  OAI211_X1 U6788 ( .C1(n5793), .C2(n6079), .A(n5721), .B(n5720), .ZN(n5722)
         );
  AOI21_X1 U6789 ( .B1(n5723), .B2(n6102), .A(n5722), .ZN(n5724) );
  OAI211_X1 U6790 ( .C1(n5726), .C2(n4234), .A(n5725), .B(n5724), .ZN(U3005)
         );
  INV_X1 U6791 ( .A(n5852), .ZN(n5729) );
  NAND3_X1 U6792 ( .A1(n5729), .A2(n5728), .A3(n5727), .ZN(n5731) );
  OAI22_X1 U6793 ( .A1(n5732), .A2(n5731), .B1(n5730), .B2(n6521), .ZN(U3455)
         );
  INV_X1 U6794 ( .A(STATE_REG_1__SCAN_IN), .ZN(n5733) );
  OAI21_X1 U6795 ( .B1(n5733), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n5738) );
  NOR2_X2 U6796 ( .A1(STATE_REG_0__SCAN_IN), .A2(n5733), .ZN(n6547) );
  OAI21_X1 U6797 ( .B1(n5738), .B2(ADS_N_REG_SCAN_IN), .A(n6497), .ZN(n5734)
         );
  INV_X1 U6798 ( .A(n5734), .ZN(U2789) );
  INV_X1 U6799 ( .A(n6420), .ZN(n6426) );
  OAI21_X1 U6800 ( .B1(n5735), .B2(n6426), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5736) );
  OAI21_X1 U6801 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6425), .A(n5736), .ZN(
        U2790) );
  NOR2_X1 U6802 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5739) );
  OAI21_X1 U6803 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5739), .A(n6497), .ZN(n5737)
         );
  OAI21_X1 U6804 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6497), .A(n5737), .ZN(
        U2791) );
  NAND2_X1 U6805 ( .A1(n6497), .A2(n5738), .ZN(n6503) );
  INV_X1 U6806 ( .A(n6503), .ZN(n6507) );
  OAI21_X1 U6807 ( .B1(BS16_N), .B2(n5739), .A(n6507), .ZN(n6505) );
  OAI21_X1 U6808 ( .B1(n6507), .B2(n6322), .A(n6505), .ZN(U2792) );
  OAI21_X1 U6809 ( .B1(n5741), .B2(n5740), .A(n5992), .ZN(U2793) );
  INV_X1 U6810 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6506) );
  INV_X1 U6811 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6504) );
  NOR2_X1 U6812 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6692) );
  NOR4_X1 U6813 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6693) );
  OAI211_X1 U6814 ( .C1(n6506), .C2(n6504), .A(n6692), .B(n6693), .ZN(n5749)
         );
  OR4_X1 U6815 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5748) );
  OR4_X1 U6816 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(
        n5747) );
  NOR4_X1 U6817 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n5745) );
  NOR4_X1 U6818 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_14__SCAN_IN), .ZN(n5744)
         );
  NOR4_X1 U6819 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5743) );
  NOR4_X1 U6820 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5742) );
  NAND4_X1 U6821 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n5746)
         );
  NOR4_X2 U6822 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n6534)
         );
  INV_X1 U6823 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5751) );
  NOR3_X1 U6824 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5752) );
  OAI21_X1 U6825 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5752), .A(n6534), .ZN(n5750)
         );
  OAI21_X1 U6826 ( .B1(n6534), .B2(n5751), .A(n5750), .ZN(U2794) );
  AOI21_X1 U6827 ( .B1(n6527), .B2(n6506), .A(n5752), .ZN(n5754) );
  INV_X1 U6828 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5753) );
  INV_X1 U6829 ( .A(n6534), .ZN(n6529) );
  AOI22_X1 U6830 ( .A1(n6534), .A2(n5754), .B1(n5753), .B2(n6529), .ZN(U2795)
         );
  AOI22_X1 U6831 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5848), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5755), .ZN(n5756) );
  OAI21_X1 U6832 ( .B1(n5757), .B2(n5870), .A(n5756), .ZN(n5758) );
  AOI211_X1 U6833 ( .C1(n5845), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5854), 
        .B(n5758), .ZN(n5761) );
  AOI22_X1 U6834 ( .A1(n5879), .A2(n4093), .B1(n5825), .B2(n5759), .ZN(n5760)
         );
  OAI211_X1 U6835 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5762), .A(n5761), .B(n5760), .ZN(U2809) );
  AOI22_X1 U6836 ( .A1(n5766), .A2(n5765), .B1(n5764), .B2(n5763), .ZN(n5768)
         );
  AOI21_X1 U6837 ( .B1(n5845), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5854), 
        .ZN(n5767) );
  OAI221_X1 U6838 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5769), .C1(n6475), .C2(
        n5768), .A(n5767), .ZN(n5770) );
  AOI21_X1 U6839 ( .B1(EBX_REG_16__SCAN_IN), .B2(n5848), .A(n5770), .ZN(n5773)
         );
  AOI22_X1 U6840 ( .A1(n5884), .A2(n4093), .B1(n4892), .B2(n5771), .ZN(n5772)
         );
  OAI211_X1 U6841 ( .C1(n5861), .C2(n5774), .A(n5773), .B(n5772), .ZN(U2811)
         );
  AOI21_X1 U6842 ( .B1(n5845), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5854), 
        .ZN(n5775) );
  OAI221_X1 U6843 ( .B1(REIP_REG_14__SCAN_IN), .B2(n5777), .C1(n6473), .C2(
        n5776), .A(n5775), .ZN(n5778) );
  AOI21_X1 U6844 ( .B1(EBX_REG_14__SCAN_IN), .B2(n5848), .A(n5778), .ZN(n5783)
         );
  INV_X1 U6845 ( .A(n5779), .ZN(n5781) );
  AOI22_X1 U6846 ( .A1(n5781), .A2(n4093), .B1(n4892), .B2(n5780), .ZN(n5782)
         );
  OAI211_X1 U6847 ( .C1(n5861), .C2(n5784), .A(n5783), .B(n5782), .ZN(U2813)
         );
  INV_X1 U6848 ( .A(n5804), .ZN(n5786) );
  OAI211_X1 U6849 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5787), .A(n5786), .B(n5785), .ZN(n5790) );
  INV_X1 U6850 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5788) );
  OAI21_X1 U6851 ( .B1(n5856), .B2(n5788), .A(n5826), .ZN(n5789) );
  AOI221_X1 U6852 ( .B1(n5791), .B2(n6471), .C1(n5790), .C2(
        REIP_REG_13__SCAN_IN), .A(n5789), .ZN(n5797) );
  OAI22_X1 U6853 ( .A1(n5793), .A2(n5861), .B1(n5792), .B2(n5870), .ZN(n5794)
         );
  AOI21_X1 U6854 ( .B1(n5795), .B2(n4093), .A(n5794), .ZN(n5796) );
  OAI211_X1 U6855 ( .C1(n5798), .C2(n5858), .A(n5797), .B(n5796), .ZN(U2814)
         );
  AND2_X1 U6856 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  NOR2_X1 U6857 ( .A1(n5802), .A2(n5801), .ZN(n5871) );
  INV_X1 U6858 ( .A(n5803), .ZN(n5805) );
  AOI22_X1 U6859 ( .A1(n5825), .A2(n5871), .B1(n5805), .B2(n5804), .ZN(n5814)
         );
  OAI22_X1 U6860 ( .A1(n5807), .A2(n6467), .B1(n5806), .B2(n5856), .ZN(n5808)
         );
  AOI211_X1 U6861 ( .C1(n5848), .C2(EBX_REG_11__SCAN_IN), .A(n5854), .B(n5808), 
        .ZN(n5813) );
  INV_X1 U6862 ( .A(n5809), .ZN(n5986) );
  OAI22_X1 U6863 ( .A1(n5988), .A2(n5810), .B1(n5870), .B2(n5986), .ZN(n5811)
         );
  INV_X1 U6864 ( .A(n5811), .ZN(n5812) );
  NAND3_X1 U6865 ( .A1(n5814), .A2(n5813), .A3(n5812), .ZN(U2816) );
  INV_X1 U6866 ( .A(n5815), .ZN(n5876) );
  AOI22_X1 U6867 ( .A1(n5876), .A2(n4093), .B1(n4892), .B2(n5816), .ZN(n5832)
         );
  INV_X1 U6868 ( .A(n5817), .ZN(n5818) );
  NAND2_X1 U6869 ( .A1(n5819), .A2(n5818), .ZN(n5822) );
  INV_X1 U6870 ( .A(n5820), .ZN(n5821) );
  AOI21_X1 U6871 ( .B1(n5823), .B2(n5822), .A(n5821), .ZN(n6042) );
  AOI22_X1 U6872 ( .A1(n5825), .A2(n6042), .B1(REIP_REG_9__SCAN_IN), .B2(n5824), .ZN(n5827) );
  OAI211_X1 U6873 ( .C1(n5856), .C2(n5828), .A(n5827), .B(n5826), .ZN(n5829)
         );
  AOI211_X1 U6874 ( .C1(n5848), .C2(EBX_REG_9__SCAN_IN), .A(n5830), .B(n5829), 
        .ZN(n5831) );
  NAND2_X1 U6875 ( .A1(n5832), .A2(n5831), .ZN(U2818) );
  OAI22_X1 U6876 ( .A1(n5834), .A2(n5858), .B1(n5861), .B2(n5833), .ZN(n5835)
         );
  AOI211_X1 U6877 ( .C1(n5845), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5854), 
        .B(n5835), .ZN(n5839) );
  NAND2_X1 U6878 ( .A1(n5837), .A2(n5836), .ZN(n5838) );
  OAI211_X1 U6879 ( .C1(n5836), .C2(n5840), .A(n5839), .B(n5838), .ZN(n5841)
         );
  AOI21_X1 U6880 ( .B1(n4093), .B2(n5993), .A(n5841), .ZN(n5842) );
  OAI21_X1 U6881 ( .B1(n5997), .B2(n5870), .A(n5842), .ZN(U2821) );
  INV_X1 U6882 ( .A(n5843), .ZN(n5864) );
  OAI22_X1 U6883 ( .A1(n5844), .A2(n6456), .B1(n5861), .B2(n6078), .ZN(n5847)
         );
  AND2_X1 U6884 ( .A1(n5845), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5846)
         );
  AOI211_X1 U6885 ( .C1(EBX_REG_4__SCAN_IN), .C2(n5848), .A(n5847), .B(n5846), 
        .ZN(n5851) );
  NAND2_X1 U6886 ( .A1(n5849), .A2(n6456), .ZN(n5850) );
  OAI211_X1 U6887 ( .C1(n5859), .C2(n5852), .A(n5851), .B(n5850), .ZN(n5853)
         );
  AOI211_X1 U6888 ( .C1(n6002), .C2(n5864), .A(n5854), .B(n5853), .ZN(n5855)
         );
  OAI21_X1 U6889 ( .B1(n6005), .B2(n5870), .A(n5855), .ZN(U2823) );
  OAI22_X1 U6890 ( .A1(n5858), .A2(n5857), .B1(n3339), .B2(n5856), .ZN(n5863)
         );
  INV_X1 U6891 ( .A(n6096), .ZN(n5860) );
  OAI22_X1 U6892 ( .A1(n5861), .A2(n5860), .B1(n4315), .B2(n5859), .ZN(n5862)
         );
  AOI211_X1 U6893 ( .C1(n6010), .C2(n5864), .A(n5863), .B(n5862), .ZN(n5869)
         );
  AND2_X1 U6894 ( .A1(n5865), .A2(REIP_REG_1__SCAN_IN), .ZN(n5867) );
  OAI21_X1 U6895 ( .B1(n5867), .B2(REIP_REG_2__SCAN_IN), .A(n5866), .ZN(n5868)
         );
  OAI211_X1 U6896 ( .C1(n5870), .C2(n6014), .A(n5869), .B(n5868), .ZN(U2825)
         );
  INV_X1 U6897 ( .A(n5871), .ZN(n6017) );
  OAI22_X1 U6898 ( .A1(n5988), .A2(n5300), .B1(n5872), .B2(n6017), .ZN(n5873)
         );
  INV_X1 U6899 ( .A(n5873), .ZN(n5874) );
  OAI21_X1 U6900 ( .B1(n5878), .B2(n5875), .A(n5874), .ZN(U2848) );
  INV_X1 U6901 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U6902 ( .A1(n5876), .A2(n3900), .B1(n3996), .B2(n6042), .ZN(n5877)
         );
  OAI21_X1 U6903 ( .B1(n5878), .B2(n6655), .A(n5877), .ZN(U2850) );
  AOI22_X1 U6904 ( .A1(n5879), .A2(n5883), .B1(n5882), .B2(DATAI_18_), .ZN(
        n5881) );
  AOI22_X1 U6905 ( .A1(n5886), .A2(DATAI_2_), .B1(n5885), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U6906 ( .A1(n5881), .A2(n5880), .ZN(U2873) );
  AOI22_X1 U6907 ( .A1(n5884), .A2(n5883), .B1(n5882), .B2(DATAI_16_), .ZN(
        n5888) );
  AOI22_X1 U6908 ( .A1(n5886), .A2(DATAI_0_), .B1(n5885), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U6909 ( .A1(n5888), .A2(n5887), .ZN(U2875) );
  INV_X1 U6910 ( .A(n5889), .ZN(n5895) );
  AOI22_X1 U6911 ( .A1(n5895), .A2(EAX_REG_30__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5890) );
  OAI21_X1 U6912 ( .B1(n6610), .B2(n5915), .A(n5890), .ZN(U2893) );
  INV_X1 U6913 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n6694) );
  INV_X1 U6914 ( .A(n5917), .ZN(n5913) );
  AOI22_X1 U6915 ( .A1(n5895), .A2(EAX_REG_29__SCAN_IN), .B1(n6539), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U6916 ( .B1(n6694), .B2(n5913), .A(n5891), .ZN(U2894) );
  AOI22_X1 U6917 ( .A1(n5895), .A2(EAX_REG_27__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5892) );
  OAI21_X1 U6918 ( .B1(n6669), .B2(n5915), .A(n5892), .ZN(U2896) );
  AOI22_X1 U6919 ( .A1(n5895), .A2(EAX_REG_22__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5893) );
  OAI21_X1 U6920 ( .B1(n6571), .B2(n5915), .A(n5893), .ZN(U2901) );
  AOI22_X1 U6921 ( .A1(n5895), .A2(EAX_REG_21__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5894) );
  OAI21_X1 U6922 ( .B1(n6666), .B2(n5915), .A(n5894), .ZN(U2902) );
  AOI22_X1 U6923 ( .A1(n5895), .A2(EAX_REG_18__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5896) );
  OAI21_X1 U6924 ( .B1(n6582), .B2(n5915), .A(n5896), .ZN(U2905) );
  INV_X1 U6925 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5981) );
  AOI22_X1 U6926 ( .A1(n5898), .A2(LWORD_REG_15__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5897) );
  OAI21_X1 U6927 ( .B1(n5981), .B2(n5919), .A(n5897), .ZN(U2908) );
  INV_X1 U6928 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5976) );
  AOI22_X1 U6929 ( .A1(n5898), .A2(LWORD_REG_14__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5899) );
  OAI21_X1 U6930 ( .B1(n5976), .B2(n5919), .A(n5899), .ZN(U2909) );
  INV_X1 U6931 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n6589) );
  INV_X1 U6932 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5900) );
  INV_X1 U6933 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n6570) );
  OAI222_X1 U6934 ( .A1(n5915), .A2(n6589), .B1(n5919), .B2(n5900), .C1(n6570), 
        .C2(n5913), .ZN(U2910) );
  INV_X1 U6935 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5970) );
  AOI22_X1 U6936 ( .A1(n6539), .A2(LWORD_REG_12__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5901) );
  OAI21_X1 U6937 ( .B1(n5970), .B2(n5919), .A(n5901), .ZN(U2911) );
  INV_X1 U6938 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5967) );
  AOI22_X1 U6939 ( .A1(n6539), .A2(LWORD_REG_11__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5902) );
  OAI21_X1 U6940 ( .B1(n5967), .B2(n5919), .A(n5902), .ZN(U2912) );
  INV_X1 U6941 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5963) );
  AOI22_X1 U6942 ( .A1(n6539), .A2(LWORD_REG_10__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5903) );
  OAI21_X1 U6943 ( .B1(n5963), .B2(n5919), .A(n5903), .ZN(U2913) );
  INV_X1 U6944 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5960) );
  AOI22_X1 U6945 ( .A1(n6539), .A2(LWORD_REG_9__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5904) );
  OAI21_X1 U6946 ( .B1(n5960), .B2(n5919), .A(n5904), .ZN(U2914) );
  AOI22_X1 U6947 ( .A1(n6539), .A2(LWORD_REG_8__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5905) );
  OAI21_X1 U6948 ( .B1(n6641), .B2(n5919), .A(n5905), .ZN(U2915) );
  AOI22_X1 U6949 ( .A1(n6539), .A2(LWORD_REG_7__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5906) );
  OAI21_X1 U6950 ( .B1(n3456), .B2(n5919), .A(n5906), .ZN(U2916) );
  AOI22_X1 U6951 ( .A1(n6539), .A2(LWORD_REG_6__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5907) );
  OAI21_X1 U6952 ( .B1(n5953), .B2(n5919), .A(n5907), .ZN(U2917) );
  INV_X1 U6953 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6623) );
  OAI222_X1 U6954 ( .A1(n5909), .A2(n5915), .B1(n5919), .B2(n5908), .C1(n5913), 
        .C2(n6623), .ZN(U2918) );
  AOI22_X1 U6955 ( .A1(n6539), .A2(LWORD_REG_4__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5910) );
  OAI21_X1 U6956 ( .B1(n5950), .B2(n5919), .A(n5910), .ZN(U2919) );
  AOI22_X1 U6957 ( .A1(n6539), .A2(LWORD_REG_3__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5911) );
  OAI21_X1 U6958 ( .B1(n5947), .B2(n5919), .A(n5911), .ZN(U2920) );
  AOI22_X1 U6959 ( .A1(n6539), .A2(LWORD_REG_2__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5912) );
  OAI21_X1 U6960 ( .B1(n5944), .B2(n5919), .A(n5912), .ZN(U2921) );
  INV_X1 U6961 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5914) );
  INV_X1 U6962 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6596) );
  OAI222_X1 U6963 ( .A1(n5916), .A2(n5915), .B1(n5919), .B2(n5914), .C1(n5913), 
        .C2(n6596), .ZN(U2922) );
  AOI22_X1 U6964 ( .A1(n6539), .A2(LWORD_REG_0__SCAN_IN), .B1(n5917), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5918) );
  OAI21_X1 U6965 ( .B1(n5941), .B2(n5919), .A(n5918), .ZN(U2923) );
  AND2_X1 U6966 ( .A1(n5977), .A2(DATAI_0_), .ZN(n5939) );
  AOI21_X1 U6967 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n5965), .A(n5939), .ZN(n5920) );
  OAI21_X1 U6968 ( .B1(n5921), .B2(n5980), .A(n5920), .ZN(U2924) );
  AOI21_X1 U6969 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n5965), .A(n5922), .ZN(n5923) );
  OAI21_X1 U6970 ( .B1(n6626), .B2(n5980), .A(n5923), .ZN(U2925) );
  AND2_X1 U6971 ( .A1(n5977), .A2(DATAI_3_), .ZN(n5945) );
  AOI21_X1 U6972 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n5978), .A(n5945), .ZN(n5925) );
  OAI21_X1 U6973 ( .B1(n5926), .B2(n5980), .A(n5925), .ZN(U2927) );
  AND2_X1 U6974 ( .A1(n5977), .A2(DATAI_4_), .ZN(n5948) );
  AOI21_X1 U6975 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n5978), .A(n5948), .ZN(n5927) );
  OAI21_X1 U6976 ( .B1(n3668), .B2(n5980), .A(n5927), .ZN(U2928) );
  AND2_X1 U6977 ( .A1(n5977), .A2(DATAI_7_), .ZN(n5954) );
  AOI21_X1 U6978 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n5978), .A(n5954), .ZN(n5928) );
  OAI21_X1 U6979 ( .B1(n6670), .B2(n5980), .A(n5928), .ZN(U2931) );
  AND2_X1 U6980 ( .A1(n5977), .A2(DATAI_8_), .ZN(n5956) );
  AOI21_X1 U6981 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n5978), .A(n5956), .ZN(n5929) );
  OAI21_X1 U6982 ( .B1(n5930), .B2(n5980), .A(n5929), .ZN(U2932) );
  INV_X1 U6983 ( .A(DATAI_9_), .ZN(n5931) );
  NOR2_X1 U6984 ( .A1(n5936), .A2(n5931), .ZN(n5958) );
  AOI21_X1 U6985 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n5978), .A(n5958), .ZN(n5932) );
  OAI21_X1 U6986 ( .B1(n5933), .B2(n5980), .A(n5932), .ZN(U2933) );
  NOR2_X1 U6987 ( .A1(n5936), .A2(n6593), .ZN(n5961) );
  AOI21_X1 U6988 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n5978), .A(n5961), .ZN(
        n5934) );
  OAI21_X1 U6989 ( .B1(n3787), .B2(n5980), .A(n5934), .ZN(U2934) );
  INV_X1 U6990 ( .A(DATAI_12_), .ZN(n5935) );
  NOR2_X1 U6991 ( .A1(n5936), .A2(n5935), .ZN(n5968) );
  AOI21_X1 U6992 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n5978), .A(n5968), .ZN(
        n5937) );
  OAI21_X1 U6993 ( .B1(n4014), .B2(n5980), .A(n5937), .ZN(U2936) );
  AOI22_X1 U6994 ( .A1(n5978), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n5971), .ZN(n5938) );
  NAND2_X1 U6995 ( .A1(n5977), .A2(DATAI_13_), .ZN(n5972) );
  NAND2_X1 U6996 ( .A1(n5938), .A2(n5972), .ZN(U2937) );
  AOI21_X1 U6997 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n5978), .A(n5939), .ZN(n5940) );
  OAI21_X1 U6998 ( .B1(n5941), .B2(n5980), .A(n5940), .ZN(U2939) );
  AOI21_X1 U6999 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n5978), .A(n5942), .ZN(n5943) );
  OAI21_X1 U7000 ( .B1(n5944), .B2(n5980), .A(n5943), .ZN(U2941) );
  AOI21_X1 U7001 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n5978), .A(n5945), .ZN(n5946) );
  OAI21_X1 U7002 ( .B1(n5947), .B2(n5980), .A(n5946), .ZN(U2942) );
  AOI21_X1 U7003 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n5978), .A(n5948), .ZN(n5949) );
  OAI21_X1 U7004 ( .B1(n5950), .B2(n5980), .A(n5949), .ZN(U2943) );
  AOI21_X1 U7005 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n5965), .A(n5951), .ZN(n5952) );
  OAI21_X1 U7006 ( .B1(n5953), .B2(n5980), .A(n5952), .ZN(U2945) );
  AOI21_X1 U7007 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n5978), .A(n5954), .ZN(n5955) );
  OAI21_X1 U7008 ( .B1(n3456), .B2(n5980), .A(n5955), .ZN(U2946) );
  AOI21_X1 U7009 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n5978), .A(n5956), .ZN(n5957) );
  OAI21_X1 U7010 ( .B1(n6641), .B2(n5980), .A(n5957), .ZN(U2947) );
  AOI21_X1 U7011 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n5978), .A(n5958), .ZN(n5959) );
  OAI21_X1 U7012 ( .B1(n5960), .B2(n5980), .A(n5959), .ZN(U2948) );
  AOI21_X1 U7013 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n5978), .A(n5961), .ZN(
        n5962) );
  OAI21_X1 U7014 ( .B1(n5963), .B2(n5980), .A(n5962), .ZN(U2949) );
  AOI21_X1 U7015 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n5965), .A(n5964), .ZN(
        n5966) );
  OAI21_X1 U7016 ( .B1(n5967), .B2(n5980), .A(n5966), .ZN(U2950) );
  AOI21_X1 U7017 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n5978), .A(n5968), .ZN(
        n5969) );
  OAI21_X1 U7018 ( .B1(n5970), .B2(n5980), .A(n5969), .ZN(U2951) );
  AOI22_X1 U7019 ( .A1(n5978), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n5971), .ZN(n5973) );
  NAND2_X1 U7020 ( .A1(n5973), .A2(n5972), .ZN(U2952) );
  AOI21_X1 U7021 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n5978), .A(n5974), .ZN(
        n5975) );
  OAI21_X1 U7022 ( .B1(n5976), .B2(n5980), .A(n5975), .ZN(U2953) );
  AOI22_X1 U7023 ( .A1(n5978), .A2(LWORD_REG_15__SCAN_IN), .B1(n5977), .B2(
        DATAI_15_), .ZN(n5979) );
  OAI21_X1 U7024 ( .B1(n5981), .B2(n5980), .A(n5979), .ZN(U2954) );
  NAND2_X1 U7025 ( .A1(n5983), .A2(n5982), .ZN(n5985) );
  XNOR2_X1 U7026 ( .A(n4226), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5984)
         );
  XNOR2_X1 U7027 ( .A(n5985), .B(n5984), .ZN(n6018) );
  AOI22_X1 U7028 ( .A1(n6076), .A2(REIP_REG_11__SCAN_IN), .B1(n6006), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5991) );
  OAI22_X1 U7029 ( .A1(n5988), .A2(n5987), .B1(n6015), .B2(n5986), .ZN(n5989)
         );
  INV_X1 U7030 ( .A(n5989), .ZN(n5990) );
  OAI211_X1 U7031 ( .C1(n6018), .C2(n5992), .A(n5991), .B(n5990), .ZN(U2975)
         );
  AOI22_X1 U7032 ( .A1(n6076), .A2(REIP_REG_6__SCAN_IN), .B1(n6006), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5996) );
  AOI22_X1 U7033 ( .A1(n5994), .A2(n6011), .B1(n5446), .B2(n5993), .ZN(n5995)
         );
  OAI211_X1 U7034 ( .C1(n6015), .C2(n5997), .A(n5996), .B(n5995), .ZN(U2980)
         );
  AOI22_X1 U7035 ( .A1(n6076), .A2(REIP_REG_4__SCAN_IN), .B1(n6006), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6004) );
  OAI21_X1 U7036 ( .B1(n6000), .B2(n5999), .A(n5998), .ZN(n6001) );
  INV_X1 U7037 ( .A(n6001), .ZN(n6081) );
  AOI22_X1 U7038 ( .A1(n6081), .A2(n6011), .B1(n6002), .B2(n5446), .ZN(n6003)
         );
  OAI211_X1 U7039 ( .C1(n6015), .C2(n6005), .A(n6004), .B(n6003), .ZN(U2982)
         );
  AOI22_X1 U7040 ( .A1(n6076), .A2(REIP_REG_2__SCAN_IN), .B1(n6006), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6013) );
  XNOR2_X1 U7041 ( .A(n6007), .B(n6106), .ZN(n6008) );
  XNOR2_X1 U7042 ( .A(n6009), .B(n6008), .ZN(n6103) );
  AOI22_X1 U7043 ( .A1(n6103), .A2(n6011), .B1(n6010), .B2(n5446), .ZN(n6012)
         );
  OAI211_X1 U7044 ( .C1(n6015), .C2(n6014), .A(n6013), .B(n6012), .ZN(U2984)
         );
  INV_X1 U7045 ( .A(n6016), .ZN(n6021) );
  OAI22_X1 U7046 ( .A1(n6017), .A2(n6079), .B1(n6467), .B2(n6032), .ZN(n6020)
         );
  NOR2_X1 U7047 ( .A1(n6018), .A2(n6086), .ZN(n6019) );
  AOI211_X1 U7048 ( .C1(n6022), .C2(n6021), .A(n6020), .B(n6019), .ZN(n6023)
         );
  OAI21_X1 U7049 ( .B1(n6024), .B2(n6022), .A(n6023), .ZN(U3007) );
  OAI21_X1 U7050 ( .B1(n6099), .B2(n6026), .A(n6025), .ZN(n6027) );
  INV_X1 U7051 ( .A(n6027), .ZN(n6028) );
  OAI21_X1 U7052 ( .B1(n6030), .B2(n6029), .A(n6028), .ZN(n6061) );
  AOI21_X1 U7053 ( .B1(n6048), .B2(n6031), .A(n6061), .ZN(n6047) );
  OAI22_X1 U7054 ( .A1(n6033), .A2(n6079), .B1(n6465), .B2(n6032), .ZN(n6034)
         );
  AOI21_X1 U7055 ( .B1(n6035), .B2(n6102), .A(n6034), .ZN(n6039) );
  NAND2_X1 U7056 ( .A1(n6036), .A2(n6066), .ZN(n6065) );
  NOR2_X1 U7057 ( .A1(n6048), .A2(n6065), .ZN(n6043) );
  OAI211_X1 U7058 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6043), .B(n6037), .ZN(n6038) );
  OAI211_X1 U7059 ( .C1(n6047), .C2(n4230), .A(n6039), .B(n6038), .ZN(U3008)
         );
  INV_X1 U7060 ( .A(n6040), .ZN(n6041) );
  AOI21_X1 U7061 ( .B1(n6042), .B2(n6097), .A(n6041), .ZN(n6046) );
  AOI22_X1 U7062 ( .A1(n6044), .A2(n6102), .B1(n5047), .B2(n6043), .ZN(n6045)
         );
  OAI211_X1 U7063 ( .C1(n6047), .C2(n5047), .A(n6046), .B(n6045), .ZN(U3009)
         );
  OAI21_X1 U7064 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6048), .ZN(n6056) );
  INV_X1 U7065 ( .A(n6049), .ZN(n6050) );
  AOI21_X1 U7066 ( .B1(n6051), .B2(n6097), .A(n6050), .ZN(n6055) );
  INV_X1 U7067 ( .A(n6052), .ZN(n6053) );
  AOI22_X1 U7068 ( .A1(n6053), .A2(n6102), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6061), .ZN(n6054) );
  OAI211_X1 U7069 ( .C1(n6065), .C2(n6056), .A(n6055), .B(n6054), .ZN(U3010)
         );
  INV_X1 U7070 ( .A(n6057), .ZN(n6058) );
  AOI21_X1 U7071 ( .B1(n6059), .B2(n6097), .A(n6058), .ZN(n6064) );
  INV_X1 U7072 ( .A(n6060), .ZN(n6062) );
  AOI22_X1 U7073 ( .A1(n6062), .A2(n6102), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6061), .ZN(n6063) );
  OAI211_X1 U7074 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6065), .A(n6064), 
        .B(n6063), .ZN(U3011) );
  AOI21_X1 U7075 ( .B1(n6689), .B2(n6066), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6072) );
  INV_X1 U7076 ( .A(n6067), .ZN(n6069) );
  AOI22_X1 U7077 ( .A1(n6069), .A2(n6102), .B1(n6097), .B2(n6068), .ZN(n6071)
         );
  NAND2_X1 U7078 ( .A1(n6076), .A2(REIP_REG_5__SCAN_IN), .ZN(n6070) );
  OAI211_X1 U7079 ( .C1(n6073), .C2(n6072), .A(n6071), .B(n6070), .ZN(U3013)
         );
  AOI21_X1 U7080 ( .B1(n6074), .B2(n6093), .A(n6092), .ZN(n6091) );
  AOI211_X1 U7081 ( .C1(n6672), .C2(n6561), .A(n6689), .B(n6085), .ZN(n6075)
         );
  AOI21_X1 U7082 ( .B1(n6076), .B2(REIP_REG_4__SCAN_IN), .A(n6075), .ZN(n6077)
         );
  OAI21_X1 U7083 ( .B1(n6079), .B2(n6078), .A(n6077), .ZN(n6080) );
  AOI21_X1 U7084 ( .B1(n6081), .B2(n6102), .A(n6080), .ZN(n6082) );
  OAI21_X1 U7085 ( .B1(n6091), .B2(n6561), .A(n6082), .ZN(U3014) );
  AOI21_X1 U7086 ( .B1(n6097), .B2(n6084), .A(n6083), .ZN(n6090) );
  OAI22_X1 U7087 ( .A1(n6087), .A2(n6086), .B1(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n6085), .ZN(n6088) );
  INV_X1 U7088 ( .A(n6088), .ZN(n6089) );
  OAI211_X1 U7089 ( .C1(n6091), .C2(n6672), .A(n6090), .B(n6089), .ZN(U3015)
         );
  INV_X1 U7090 ( .A(n6092), .ZN(n6105) );
  AOI21_X1 U7091 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6094), .A(n6093), 
        .ZN(n6100) );
  AOI22_X1 U7092 ( .A1(n6097), .A2(n6096), .B1(n6095), .B2(REIP_REG_2__SCAN_IN), .ZN(n6098) );
  OAI21_X1 U7093 ( .B1(n6100), .B2(n6099), .A(n6098), .ZN(n6101) );
  AOI21_X1 U7094 ( .B1(n6103), .B2(n6102), .A(n6101), .ZN(n6104) );
  OAI221_X1 U7095 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6107), .C1(n6106), .C2(n6105), .A(n6104), .ZN(U3016) );
  NOR2_X1 U7096 ( .A1(n6398), .A2(n6108), .ZN(U3019) );
  NOR2_X1 U7097 ( .A1(n6111), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6138)
         );
  AOI22_X1 U7098 ( .A1(n6139), .A2(n6178), .B1(n6320), .B2(n6138), .ZN(n6124)
         );
  INV_X1 U7099 ( .A(n6120), .ZN(n6118) );
  NOR3_X1 U7100 ( .A1(n6219), .A2(n6113), .A3(n6112), .ZN(n6114) );
  NOR2_X1 U7101 ( .A1(n6114), .A2(n6325), .ZN(n6119) );
  AOI21_X1 U7102 ( .B1(n6115), .B2(n6382), .A(n6138), .ZN(n6121) );
  NAND2_X1 U7103 ( .A1(n6119), .A2(n6121), .ZN(n6117) );
  OAI211_X1 U7104 ( .C1(n6218), .C2(n6118), .A(n6117), .B(n6116), .ZN(n6141)
         );
  INV_X1 U7105 ( .A(n6119), .ZN(n6122) );
  OAI22_X1 U7106 ( .A1(n6122), .A2(n6121), .B1(n6120), .B2(n6414), .ZN(n6140)
         );
  AOI22_X1 U7107 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6141), .B1(n6321), 
        .B2(n6140), .ZN(n6123) );
  OAI211_X1 U7108 ( .C1(n6233), .C2(n6176), .A(n6124), .B(n6123), .ZN(U3044)
         );
  AOI22_X1 U7109 ( .A1(n6139), .A2(n6182), .B1(n6337), .B2(n6138), .ZN(n6126)
         );
  AOI22_X1 U7110 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6141), .B1(n6336), 
        .B2(n6140), .ZN(n6125) );
  OAI211_X1 U7111 ( .C1(n6280), .C2(n6176), .A(n6126), .B(n6125), .ZN(U3045)
         );
  AOI22_X1 U7112 ( .A1(n6139), .A2(n6187), .B1(n6342), .B2(n6138), .ZN(n6128)
         );
  AOI22_X1 U7113 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6141), .B1(n6343), 
        .B2(n6140), .ZN(n6127) );
  OAI211_X1 U7114 ( .C1(n6282), .C2(n6176), .A(n6128), .B(n6127), .ZN(U3046)
         );
  AOI22_X1 U7115 ( .A1(n6139), .A2(n6192), .B1(n6348), .B2(n6138), .ZN(n6130)
         );
  AOI22_X1 U7116 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6141), .B1(n6349), 
        .B2(n6140), .ZN(n6129) );
  OAI211_X1 U7117 ( .C1(n6290), .C2(n6176), .A(n6130), .B(n6129), .ZN(U3047)
         );
  AOI22_X1 U7118 ( .A1(n6139), .A2(n6131), .B1(n6354), .B2(n6138), .ZN(n6133)
         );
  AOI22_X1 U7119 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6141), .B1(n6355), 
        .B2(n6140), .ZN(n6132) );
  OAI211_X1 U7120 ( .C1(n6295), .C2(n6176), .A(n6133), .B(n6132), .ZN(U3048)
         );
  AOI22_X1 U7121 ( .A1(n6139), .A2(n6197), .B1(n6360), .B2(n6138), .ZN(n6135)
         );
  AOI22_X1 U7122 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6141), .B1(n6361), 
        .B2(n6140), .ZN(n6134) );
  OAI211_X1 U7123 ( .C1(n6297), .C2(n6176), .A(n6135), .B(n6134), .ZN(U3049)
         );
  AOI22_X1 U7124 ( .A1(n6139), .A2(n6202), .B1(n6366), .B2(n6138), .ZN(n6137)
         );
  AOI22_X1 U7125 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6141), .B1(n6367), 
        .B2(n6140), .ZN(n6136) );
  OAI211_X1 U7126 ( .C1(n6305), .C2(n6176), .A(n6137), .B(n6136), .ZN(U3050)
         );
  AOI22_X1 U7127 ( .A1(n6139), .A2(n6209), .B1(n6550), .B2(n6138), .ZN(n6143)
         );
  AOI22_X1 U7128 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6141), .B1(n6374), 
        .B2(n6140), .ZN(n6142) );
  OAI211_X1 U7129 ( .C1(n6314), .C2(n6176), .A(n6143), .B(n6142), .ZN(U3051)
         );
  NAND2_X1 U7130 ( .A1(n6327), .A2(n6218), .ZN(n6318) );
  INV_X1 U7131 ( .A(n6144), .ZN(n6145) );
  OAI22_X1 U7132 ( .A1(n6318), .A2(n6146), .B1(n6145), .B2(n6316), .ZN(n6172)
         );
  NOR2_X1 U7133 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6147), .ZN(n6171)
         );
  AOI22_X1 U7134 ( .A1(n6321), .A2(n6172), .B1(n6320), .B2(n6171), .ZN(n6158)
         );
  INV_X1 U7135 ( .A(n6148), .ZN(n6151) );
  OAI211_X1 U7136 ( .C1(n6176), .C2(n6151), .A(n6150), .B(n6149), .ZN(n6156)
         );
  INV_X1 U7137 ( .A(n6171), .ZN(n6154) );
  AOI211_X1 U7138 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6154), .A(n6153), .B(
        n6152), .ZN(n6155) );
  NAND2_X1 U7139 ( .A1(n6156), .A2(n6155), .ZN(n6173) );
  AOI22_X1 U7140 ( .A1(n6173), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6332), 
        .B2(n6208), .ZN(n6157) );
  OAI211_X1 U7141 ( .C1(n6335), .C2(n6176), .A(n6158), .B(n6157), .ZN(U3052)
         );
  AOI22_X1 U7142 ( .A1(n6337), .A2(n6171), .B1(n6336), .B2(n6172), .ZN(n6160)
         );
  AOI22_X1 U7143 ( .A1(n6173), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6338), 
        .B2(n6208), .ZN(n6159) );
  OAI211_X1 U7144 ( .C1(n6341), .C2(n6176), .A(n6160), .B(n6159), .ZN(U3053)
         );
  AOI22_X1 U7145 ( .A1(n6343), .A2(n6172), .B1(n6342), .B2(n6171), .ZN(n6162)
         );
  AOI22_X1 U7146 ( .A1(n6173), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6344), 
        .B2(n6208), .ZN(n6161) );
  OAI211_X1 U7147 ( .C1(n6347), .C2(n6176), .A(n6162), .B(n6161), .ZN(U3054)
         );
  AOI22_X1 U7148 ( .A1(n6349), .A2(n6172), .B1(n6348), .B2(n6171), .ZN(n6164)
         );
  AOI22_X1 U7149 ( .A1(n6173), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6350), 
        .B2(n6208), .ZN(n6163) );
  OAI211_X1 U7150 ( .C1(n6353), .C2(n6176), .A(n6164), .B(n6163), .ZN(U3055)
         );
  AOI22_X1 U7151 ( .A1(n6355), .A2(n6172), .B1(n6354), .B2(n6171), .ZN(n6166)
         );
  AOI22_X1 U7152 ( .A1(n6173), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6356), 
        .B2(n6208), .ZN(n6165) );
  OAI211_X1 U7153 ( .C1(n6359), .C2(n6176), .A(n6166), .B(n6165), .ZN(U3056)
         );
  AOI22_X1 U7154 ( .A1(n6361), .A2(n6172), .B1(n6360), .B2(n6171), .ZN(n6168)
         );
  AOI22_X1 U7155 ( .A1(n6173), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6362), 
        .B2(n6208), .ZN(n6167) );
  OAI211_X1 U7156 ( .C1(n6365), .C2(n6176), .A(n6168), .B(n6167), .ZN(U3057)
         );
  AOI22_X1 U7157 ( .A1(n6367), .A2(n6172), .B1(n6366), .B2(n6171), .ZN(n6170)
         );
  AOI22_X1 U7158 ( .A1(n6173), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6368), 
        .B2(n6208), .ZN(n6169) );
  OAI211_X1 U7159 ( .C1(n6371), .C2(n6176), .A(n6170), .B(n6169), .ZN(U3058)
         );
  AOI22_X1 U7160 ( .A1(n6374), .A2(n6172), .B1(n6550), .B2(n6171), .ZN(n6175)
         );
  AOI22_X1 U7161 ( .A1(n6173), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6556), 
        .B2(n6208), .ZN(n6174) );
  OAI211_X1 U7162 ( .C1(n6559), .C2(n6176), .A(n6175), .B(n6174), .ZN(U3059)
         );
  INV_X1 U7163 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6639) );
  OAI22_X1 U7164 ( .A1(n6558), .A2(n6233), .B1(n6215), .B2(n6206), .ZN(n6177)
         );
  INV_X1 U7165 ( .A(n6177), .ZN(n6180) );
  AOI22_X1 U7166 ( .A1(n6210), .A2(n6321), .B1(n6178), .B2(n6208), .ZN(n6179)
         );
  OAI211_X1 U7167 ( .C1(n6214), .C2(n6639), .A(n6180), .B(n6179), .ZN(U3060)
         );
  INV_X1 U7168 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6185) );
  OAI22_X1 U7169 ( .A1(n6558), .A2(n6280), .B1(n6275), .B2(n6206), .ZN(n6181)
         );
  INV_X1 U7170 ( .A(n6181), .ZN(n6184) );
  AOI22_X1 U7171 ( .A1(n6210), .A2(n6336), .B1(n6182), .B2(n6208), .ZN(n6183)
         );
  OAI211_X1 U7172 ( .C1(n6214), .C2(n6185), .A(n6184), .B(n6183), .ZN(U3061)
         );
  INV_X1 U7173 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6190) );
  OAI22_X1 U7174 ( .A1(n6558), .A2(n6282), .B1(n6281), .B2(n6206), .ZN(n6186)
         );
  INV_X1 U7175 ( .A(n6186), .ZN(n6189) );
  AOI22_X1 U7176 ( .A1(n6210), .A2(n6343), .B1(n6187), .B2(n6208), .ZN(n6188)
         );
  OAI211_X1 U7177 ( .C1(n6214), .C2(n6190), .A(n6189), .B(n6188), .ZN(U3062)
         );
  INV_X1 U7178 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n6195) );
  OAI22_X1 U7179 ( .A1(n6558), .A2(n6290), .B1(n6286), .B2(n6206), .ZN(n6191)
         );
  INV_X1 U7180 ( .A(n6191), .ZN(n6194) );
  AOI22_X1 U7181 ( .A1(n6210), .A2(n6349), .B1(n6192), .B2(n6208), .ZN(n6193)
         );
  OAI211_X1 U7182 ( .C1(n6214), .C2(n6195), .A(n6194), .B(n6193), .ZN(U3063)
         );
  INV_X1 U7183 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6200) );
  OAI22_X1 U7184 ( .A1(n6558), .A2(n6297), .B1(n6296), .B2(n6206), .ZN(n6196)
         );
  INV_X1 U7185 ( .A(n6196), .ZN(n6199) );
  AOI22_X1 U7186 ( .A1(n6210), .A2(n6361), .B1(n6197), .B2(n6208), .ZN(n6198)
         );
  OAI211_X1 U7187 ( .C1(n6214), .C2(n6200), .A(n6199), .B(n6198), .ZN(U3065)
         );
  INV_X1 U7188 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6205) );
  OAI22_X1 U7189 ( .A1(n6558), .A2(n6305), .B1(n6301), .B2(n6206), .ZN(n6201)
         );
  INV_X1 U7190 ( .A(n6201), .ZN(n6204) );
  AOI22_X1 U7191 ( .A1(n6210), .A2(n6367), .B1(n6202), .B2(n6208), .ZN(n6203)
         );
  OAI211_X1 U7192 ( .C1(n6214), .C2(n6205), .A(n6204), .B(n6203), .ZN(U3066)
         );
  INV_X1 U7193 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6213) );
  OAI22_X1 U7194 ( .A1(n6558), .A2(n6314), .B1(n6307), .B2(n6206), .ZN(n6207)
         );
  INV_X1 U7195 ( .A(n6207), .ZN(n6212) );
  AOI22_X1 U7196 ( .A1(n6210), .A2(n6374), .B1(n6209), .B2(n6208), .ZN(n6211)
         );
  OAI211_X1 U7197 ( .C1(n6214), .C2(n6213), .A(n6212), .B(n6211), .ZN(U3067)
         );
  OAI22_X1 U7198 ( .A1(n6253), .A2(n6335), .B1(n6252), .B2(n6215), .ZN(n6216)
         );
  INV_X1 U7199 ( .A(n6216), .ZN(n6232) );
  INV_X1 U7200 ( .A(n6217), .ZN(n6220) );
  OAI21_X1 U7201 ( .B1(n6220), .B2(n6219), .A(n6218), .ZN(n6230) );
  NOR2_X1 U7202 ( .A1(n2956), .A2(n6326), .ZN(n6223) );
  INV_X1 U7203 ( .A(n6252), .ZN(n6222) );
  AOI21_X1 U7204 ( .B1(n6224), .B2(n6223), .A(n6222), .ZN(n6229) );
  INV_X1 U7205 ( .A(n6229), .ZN(n6227) );
  AOI21_X1 U7206 ( .B1(n6228), .B2(n6325), .A(n6225), .ZN(n6226) );
  OAI21_X1 U7207 ( .B1(n6230), .B2(n6227), .A(n6226), .ZN(n6256) );
  OAI22_X1 U7208 ( .A1(n6230), .A2(n6229), .B1(n6228), .B2(n6414), .ZN(n6255)
         );
  AOI22_X1 U7209 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6256), .B1(n6321), 
        .B2(n6255), .ZN(n6231) );
  OAI211_X1 U7210 ( .C1(n6233), .C2(n6274), .A(n6232), .B(n6231), .ZN(U3076)
         );
  OAI22_X1 U7211 ( .A1(n6253), .A2(n6341), .B1(n6252), .B2(n6275), .ZN(n6234)
         );
  INV_X1 U7212 ( .A(n6234), .ZN(n6236) );
  AOI22_X1 U7213 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6256), .B1(n6336), 
        .B2(n6255), .ZN(n6235) );
  OAI211_X1 U7214 ( .C1(n6280), .C2(n6274), .A(n6236), .B(n6235), .ZN(U3077)
         );
  OAI22_X1 U7215 ( .A1(n6253), .A2(n6347), .B1(n6252), .B2(n6281), .ZN(n6237)
         );
  INV_X1 U7216 ( .A(n6237), .ZN(n6239) );
  AOI22_X1 U7217 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6256), .B1(n6343), 
        .B2(n6255), .ZN(n6238) );
  OAI211_X1 U7218 ( .C1(n6282), .C2(n6274), .A(n6239), .B(n6238), .ZN(U3078)
         );
  OAI22_X1 U7219 ( .A1(n6253), .A2(n6353), .B1(n6252), .B2(n6286), .ZN(n6240)
         );
  INV_X1 U7220 ( .A(n6240), .ZN(n6242) );
  AOI22_X1 U7221 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6256), .B1(n6349), 
        .B2(n6255), .ZN(n6241) );
  OAI211_X1 U7222 ( .C1(n6290), .C2(n6274), .A(n6242), .B(n6241), .ZN(U3079)
         );
  OAI22_X1 U7223 ( .A1(n6253), .A2(n6359), .B1(n6252), .B2(n6291), .ZN(n6243)
         );
  INV_X1 U7224 ( .A(n6243), .ZN(n6245) );
  AOI22_X1 U7225 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6256), .B1(n6355), 
        .B2(n6255), .ZN(n6244) );
  OAI211_X1 U7226 ( .C1(n6295), .C2(n6274), .A(n6245), .B(n6244), .ZN(U3080)
         );
  OAI22_X1 U7227 ( .A1(n6253), .A2(n6365), .B1(n6252), .B2(n6296), .ZN(n6246)
         );
  INV_X1 U7228 ( .A(n6246), .ZN(n6248) );
  AOI22_X1 U7229 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6256), .B1(n6361), 
        .B2(n6255), .ZN(n6247) );
  OAI211_X1 U7230 ( .C1(n6297), .C2(n6274), .A(n6248), .B(n6247), .ZN(U3081)
         );
  OAI22_X1 U7231 ( .A1(n6274), .A2(n6305), .B1(n6252), .B2(n6301), .ZN(n6249)
         );
  INV_X1 U7232 ( .A(n6249), .ZN(n6251) );
  AOI22_X1 U7233 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6256), .B1(n6367), 
        .B2(n6255), .ZN(n6250) );
  OAI211_X1 U7234 ( .C1(n6371), .C2(n6253), .A(n6251), .B(n6250), .ZN(U3082)
         );
  OAI22_X1 U7235 ( .A1(n6253), .A2(n6559), .B1(n6252), .B2(n6307), .ZN(n6254)
         );
  INV_X1 U7236 ( .A(n6254), .ZN(n6258) );
  AOI22_X1 U7237 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6256), .B1(n6374), 
        .B2(n6255), .ZN(n6257) );
  OAI211_X1 U7238 ( .C1(n6314), .C2(n6274), .A(n6258), .B(n6257), .ZN(U3083)
         );
  INV_X1 U7239 ( .A(n6259), .ZN(n6269) );
  AOI22_X1 U7240 ( .A1(n6269), .A2(n6336), .B1(n6337), .B2(n6268), .ZN(n6261)
         );
  AOI22_X1 U7241 ( .A1(n6271), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6338), 
        .B2(n6270), .ZN(n6260) );
  OAI211_X1 U7242 ( .C1(n6341), .C2(n6274), .A(n6261), .B(n6260), .ZN(U3085)
         );
  AOI22_X1 U7243 ( .A1(n6343), .A2(n6269), .B1(n6342), .B2(n6268), .ZN(n6263)
         );
  AOI22_X1 U7244 ( .A1(n6271), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6344), 
        .B2(n6270), .ZN(n6262) );
  OAI211_X1 U7245 ( .C1(n6347), .C2(n6274), .A(n6263), .B(n6262), .ZN(U3086)
         );
  AOI22_X1 U7246 ( .A1(n6355), .A2(n6269), .B1(n6354), .B2(n6268), .ZN(n6265)
         );
  AOI22_X1 U7247 ( .A1(n6271), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6356), 
        .B2(n6270), .ZN(n6264) );
  OAI211_X1 U7248 ( .C1(n6359), .C2(n6274), .A(n6265), .B(n6264), .ZN(U3088)
         );
  AOI22_X1 U7249 ( .A1(n6361), .A2(n6269), .B1(n6360), .B2(n6268), .ZN(n6267)
         );
  AOI22_X1 U7250 ( .A1(n6271), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6362), 
        .B2(n6270), .ZN(n6266) );
  OAI211_X1 U7251 ( .C1(n6365), .C2(n6274), .A(n6267), .B(n6266), .ZN(U3089)
         );
  AOI22_X1 U7252 ( .A1(n6374), .A2(n6269), .B1(n6550), .B2(n6268), .ZN(n6273)
         );
  AOI22_X1 U7253 ( .A1(n6271), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6556), 
        .B2(n6270), .ZN(n6272) );
  OAI211_X1 U7254 ( .C1(n6559), .C2(n6274), .A(n6273), .B(n6272), .ZN(U3091)
         );
  OAI22_X1 U7255 ( .A1(n6308), .A2(n6341), .B1(n6275), .B2(n6306), .ZN(n6276)
         );
  INV_X1 U7256 ( .A(n6276), .ZN(n6279) );
  INV_X1 U7257 ( .A(n6277), .ZN(n6311) );
  AOI22_X1 U7258 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6311), .B1(n6336), 
        .B2(n6310), .ZN(n6278) );
  OAI211_X1 U7259 ( .C1(n6280), .C2(n6379), .A(n6279), .B(n6278), .ZN(U3109)
         );
  OAI22_X1 U7260 ( .A1(n6379), .A2(n6282), .B1(n6281), .B2(n6306), .ZN(n6283)
         );
  INV_X1 U7261 ( .A(n6283), .ZN(n6285) );
  AOI22_X1 U7262 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6311), .B1(n6343), 
        .B2(n6310), .ZN(n6284) );
  OAI211_X1 U7263 ( .C1(n6347), .C2(n6308), .A(n6285), .B(n6284), .ZN(U3110)
         );
  OAI22_X1 U7264 ( .A1(n6308), .A2(n6353), .B1(n6286), .B2(n6306), .ZN(n6287)
         );
  INV_X1 U7265 ( .A(n6287), .ZN(n6289) );
  AOI22_X1 U7266 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6311), .B1(n6349), 
        .B2(n6310), .ZN(n6288) );
  OAI211_X1 U7267 ( .C1(n6290), .C2(n6379), .A(n6289), .B(n6288), .ZN(U3111)
         );
  OAI22_X1 U7268 ( .A1(n6308), .A2(n6359), .B1(n6291), .B2(n6306), .ZN(n6292)
         );
  INV_X1 U7269 ( .A(n6292), .ZN(n6294) );
  AOI22_X1 U7270 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6311), .B1(n6355), 
        .B2(n6310), .ZN(n6293) );
  OAI211_X1 U7271 ( .C1(n6295), .C2(n6379), .A(n6294), .B(n6293), .ZN(U3112)
         );
  OAI22_X1 U7272 ( .A1(n6379), .A2(n6297), .B1(n6296), .B2(n6306), .ZN(n6298)
         );
  INV_X1 U7273 ( .A(n6298), .ZN(n6300) );
  AOI22_X1 U7274 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6311), .B1(n6361), 
        .B2(n6310), .ZN(n6299) );
  OAI211_X1 U7275 ( .C1(n6365), .C2(n6308), .A(n6300), .B(n6299), .ZN(U3113)
         );
  OAI22_X1 U7276 ( .A1(n6308), .A2(n6371), .B1(n6301), .B2(n6306), .ZN(n6302)
         );
  INV_X1 U7277 ( .A(n6302), .ZN(n6304) );
  AOI22_X1 U7278 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6311), .B1(n6367), 
        .B2(n6310), .ZN(n6303) );
  OAI211_X1 U7279 ( .C1(n6305), .C2(n6379), .A(n6304), .B(n6303), .ZN(U3114)
         );
  OAI22_X1 U7280 ( .A1(n6308), .A2(n6559), .B1(n6307), .B2(n6306), .ZN(n6309)
         );
  INV_X1 U7281 ( .A(n6309), .ZN(n6313) );
  AOI22_X1 U7282 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6311), .B1(n6374), 
        .B2(n6310), .ZN(n6312) );
  OAI211_X1 U7283 ( .C1(n6314), .C2(n6379), .A(n6313), .B(n6312), .ZN(U3115)
         );
  OAI22_X1 U7284 ( .A1(n6318), .A2(n6317), .B1(n6316), .B2(n6315), .ZN(n6373)
         );
  NOR2_X1 U7285 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6319), .ZN(n6372)
         );
  AOI22_X1 U7286 ( .A1(n6321), .A2(n6373), .B1(n6320), .B2(n6372), .ZN(n6334)
         );
  INV_X1 U7287 ( .A(n6375), .ZN(n6323) );
  AOI21_X1 U7288 ( .B1(n6323), .B2(n6379), .A(n6322), .ZN(n6324) );
  AOI211_X1 U7289 ( .C1(n6327), .C2(n6326), .A(n6325), .B(n6324), .ZN(n6331)
         );
  OAI211_X1 U7290 ( .C1(n6512), .C2(n6372), .A(n6329), .B(n6328), .ZN(n6330)
         );
  AOI22_X1 U7291 ( .A1(n6376), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6332), 
        .B2(n6375), .ZN(n6333) );
  OAI211_X1 U7292 ( .C1(n6335), .C2(n6379), .A(n6334), .B(n6333), .ZN(U3116)
         );
  AOI22_X1 U7293 ( .A1(n6337), .A2(n6372), .B1(n6336), .B2(n6373), .ZN(n6340)
         );
  AOI22_X1 U7294 ( .A1(n6376), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6338), 
        .B2(n6375), .ZN(n6339) );
  OAI211_X1 U7295 ( .C1(n6341), .C2(n6379), .A(n6340), .B(n6339), .ZN(U3117)
         );
  AOI22_X1 U7296 ( .A1(n6343), .A2(n6373), .B1(n6342), .B2(n6372), .ZN(n6346)
         );
  AOI22_X1 U7297 ( .A1(n6376), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6344), 
        .B2(n6375), .ZN(n6345) );
  OAI211_X1 U7298 ( .C1(n6347), .C2(n6379), .A(n6346), .B(n6345), .ZN(U3118)
         );
  AOI22_X1 U7299 ( .A1(n6349), .A2(n6373), .B1(n6348), .B2(n6372), .ZN(n6352)
         );
  AOI22_X1 U7300 ( .A1(n6376), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6350), 
        .B2(n6375), .ZN(n6351) );
  OAI211_X1 U7301 ( .C1(n6353), .C2(n6379), .A(n6352), .B(n6351), .ZN(U3119)
         );
  AOI22_X1 U7302 ( .A1(n6355), .A2(n6373), .B1(n6354), .B2(n6372), .ZN(n6358)
         );
  AOI22_X1 U7303 ( .A1(n6376), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6356), 
        .B2(n6375), .ZN(n6357) );
  OAI211_X1 U7304 ( .C1(n6359), .C2(n6379), .A(n6358), .B(n6357), .ZN(U3120)
         );
  AOI22_X1 U7305 ( .A1(n6361), .A2(n6373), .B1(n6360), .B2(n6372), .ZN(n6364)
         );
  AOI22_X1 U7306 ( .A1(n6376), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6362), 
        .B2(n6375), .ZN(n6363) );
  OAI211_X1 U7307 ( .C1(n6365), .C2(n6379), .A(n6364), .B(n6363), .ZN(U3121)
         );
  AOI22_X1 U7308 ( .A1(n6367), .A2(n6373), .B1(n6366), .B2(n6372), .ZN(n6370)
         );
  AOI22_X1 U7309 ( .A1(n6376), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6368), 
        .B2(n6375), .ZN(n6369) );
  OAI211_X1 U7310 ( .C1(n6371), .C2(n6379), .A(n6370), .B(n6369), .ZN(U3122)
         );
  AOI22_X1 U7311 ( .A1(n6374), .A2(n6373), .B1(n6550), .B2(n6372), .ZN(n6378)
         );
  AOI22_X1 U7312 ( .A1(n6376), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6556), 
        .B2(n6375), .ZN(n6377) );
  OAI211_X1 U7313 ( .C1(n6559), .C2(n6379), .A(n6378), .B(n6377), .ZN(U3123)
         );
  AOI22_X1 U7314 ( .A1(n6382), .A2(n6381), .B1(n6380), .B2(n3041), .ZN(n6518)
         );
  NAND2_X1 U7315 ( .A1(n6383), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6526) );
  AND3_X1 U7316 ( .A1(n6518), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6526), 
        .ZN(n6389) );
  INV_X1 U7317 ( .A(n6389), .ZN(n6386) );
  OAI211_X1 U7318 ( .C1(n6387), .C2(n6386), .A(n6385), .B(n6384), .ZN(n6388)
         );
  OAI21_X1 U7319 ( .B1(n6389), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6388), 
        .ZN(n6392) );
  INV_X1 U7320 ( .A(n6392), .ZN(n6390) );
  NOR2_X1 U7321 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6390), .ZN(n6393)
         );
  OAI22_X1 U7322 ( .A1(n6394), .A2(n6393), .B1(n6392), .B2(n6391), .ZN(n6395)
         );
  OAI21_X1 U7323 ( .B1(n6396), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6395), 
        .ZN(n6399) );
  NAND2_X1 U7324 ( .A1(n6396), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6397) );
  NAND3_X1 U7325 ( .A1(n6399), .A2(n6398), .A3(n6397), .ZN(n6408) );
  NOR2_X1 U7326 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6402) );
  OAI211_X1 U7327 ( .C1(n6403), .C2(n6402), .A(n6401), .B(n6400), .ZN(n6404)
         );
  NOR2_X1 U7328 ( .A1(n6405), .A2(n6404), .ZN(n6407) );
  NAND3_X1 U7329 ( .A1(n6408), .A2(n6407), .A3(n6406), .ZN(n6419) );
  NAND2_X1 U7330 ( .A1(READY_N), .A2(n6539), .ZN(n6409) );
  OAI21_X1 U7331 ( .B1(n6419), .B2(n6426), .A(n6409), .ZN(n6413) );
  OR2_X1 U7332 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  AOI21_X1 U7333 ( .B1(READY_N), .B2(n6414), .A(n6508), .ZN(n6424) );
  NOR2_X1 U7334 ( .A1(n6512), .A2(n6430), .ZN(n6416) );
  AOI211_X1 U7335 ( .C1(n6416), .C2(n6415), .A(STATE2_REG_0__SCAN_IN), .B(
        n6508), .ZN(n6417) );
  AOI211_X1 U7336 ( .C1(n6420), .C2(n6419), .A(n6418), .B(n6417), .ZN(n6421)
         );
  OAI221_X1 U7337 ( .B1(n6423), .B2(n6424), .C1(n6423), .C2(n6422), .A(n6421), 
        .ZN(U3148) );
  NOR2_X1 U7338 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6433) );
  NOR3_X1 U7339 ( .A1(n6433), .A2(n6424), .A3(n6520), .ZN(n6428) );
  AOI221_X1 U7340 ( .B1(READY_N), .B2(n6426), .C1(n6425), .C2(n6426), .A(n6508), .ZN(n6427) );
  OR3_X1 U7341 ( .A1(n6429), .A2(n6428), .A3(n6427), .ZN(U3149) );
  OAI211_X1 U7342 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6538), .A(n6509), .B(
        n6430), .ZN(n6432) );
  OAI21_X1 U7343 ( .B1(n6433), .B2(n6432), .A(n6431), .ZN(U3150) );
  AND2_X1 U7344 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6503), .ZN(U3151) );
  INV_X1 U7345 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6568) );
  NOR2_X1 U7346 ( .A1(n6507), .A2(n6568), .ZN(U3152) );
  AND2_X1 U7347 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6503), .ZN(U3153) );
  AND2_X1 U7348 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6503), .ZN(U3154) );
  INV_X1 U7349 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6562) );
  NOR2_X1 U7350 ( .A1(n6507), .A2(n6562), .ZN(U3155) );
  INV_X1 U7351 ( .A(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6642) );
  NOR2_X1 U7352 ( .A1(n6507), .A2(n6642), .ZN(U3156) );
  AND2_X1 U7353 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6503), .ZN(U3157) );
  INV_X1 U7354 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6608) );
  NOR2_X1 U7355 ( .A1(n6507), .A2(n6608), .ZN(U3158) );
  AND2_X1 U7356 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6503), .ZN(U3159) );
  AND2_X1 U7357 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6503), .ZN(U3160) );
  INV_X1 U7358 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U7359 ( .A1(n6507), .A2(n6578), .ZN(U3161) );
  AND2_X1 U7360 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6503), .ZN(U3162) );
  AND2_X1 U7361 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6503), .ZN(U3163) );
  AND2_X1 U7362 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6503), .ZN(U3164) );
  INV_X1 U7363 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6632) );
  NOR2_X1 U7364 ( .A1(n6507), .A2(n6632), .ZN(U3165) );
  AND2_X1 U7365 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6503), .ZN(U3166) );
  INV_X1 U7366 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6657) );
  NOR2_X1 U7367 ( .A1(n6507), .A2(n6657), .ZN(U3167) );
  AND2_X1 U7368 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6503), .ZN(U3168) );
  AND2_X1 U7369 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6503), .ZN(U3169) );
  AND2_X1 U7370 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6503), .ZN(U3170) );
  AND2_X1 U7371 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6503), .ZN(U3171) );
  AND2_X1 U7372 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6503), .ZN(U3172) );
  AND2_X1 U7373 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6503), .ZN(U3173) );
  AND2_X1 U7374 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6503), .ZN(U3174) );
  AND2_X1 U7375 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6503), .ZN(U3175) );
  AND2_X1 U7376 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6503), .ZN(U3176) );
  AND2_X1 U7377 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6503), .ZN(U3177) );
  AND2_X1 U7378 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6503), .ZN(U3178) );
  AND2_X1 U7379 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6503), .ZN(U3179) );
  AND2_X1 U7380 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6503), .ZN(U3180) );
  NAND2_X1 U7381 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6437) );
  NAND2_X1 U7382 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6438) );
  NAND2_X1 U7383 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U7384 ( .A1(n6438), .A2(n6445), .ZN(n6444) );
  INV_X1 U7385 ( .A(NA_N), .ZN(n6446) );
  INV_X1 U7386 ( .A(n6435), .ZN(n6434) );
  AOI211_X1 U7387 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6446), .A(
        STATE_REG_0__SCAN_IN), .B(n6434), .ZN(n6450) );
  AOI21_X1 U7388 ( .B1(n6435), .B2(n6444), .A(n6450), .ZN(n6436) );
  OAI221_X1 U7389 ( .B1(n6547), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6547), 
        .C2(n6437), .A(n6436), .ZN(U3181) );
  AND2_X1 U7390 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6440) );
  INV_X1 U7391 ( .A(n6437), .ZN(n6439) );
  OAI21_X1 U7392 ( .B1(n6440), .B2(n6439), .A(n6438), .ZN(n6441) );
  NAND3_X1 U7393 ( .A1(n6442), .A2(n6445), .A3(n6441), .ZN(U3182) );
  AOI221_X1 U7394 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6538), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6443) );
  AOI22_X1 U7395 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6444), .B1(HOLD), .B2(n6443), .ZN(n6449) );
  INV_X1 U7396 ( .A(n6445), .ZN(n6447) );
  NAND4_X1 U7397 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6447), .A4(n6446), .ZN(n6448) );
  OAI221_X1 U7398 ( .B1(n6450), .B2(STATE_REG_0__SCAN_IN), .C1(n6450), .C2(
        n6449), .A(n6448), .ZN(U3183) );
  INV_X1 U7399 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U7400 ( .A1(n6547), .A2(n6451), .ZN(n6500) );
  INV_X1 U7401 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6452) );
  INV_X1 U7402 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U7403 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6547), .ZN(n6496) );
  OAI222_X1 U7404 ( .A1(n6500), .A2(n6452), .B1(n6629), .B2(n6547), .C1(n6527), 
        .C2(n6496), .ZN(U3184) );
  INV_X1 U7405 ( .A(n6496), .ZN(n6498) );
  AOI22_X1 U7406 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6497), .ZN(n6453) );
  OAI21_X1 U7407 ( .B1(n6454), .B2(n6500), .A(n6453), .ZN(U3185) );
  AOI22_X1 U7408 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6497), .ZN(n6455) );
  OAI21_X1 U7409 ( .B1(n6456), .B2(n6500), .A(n6455), .ZN(U3186) );
  AOI22_X1 U7410 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6497), .ZN(n6457) );
  OAI21_X1 U7411 ( .B1(n6458), .B2(n6500), .A(n6457), .ZN(U3187) );
  AOI22_X1 U7412 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6497), .ZN(n6459) );
  OAI21_X1 U7413 ( .B1(n5836), .B2(n6500), .A(n6459), .ZN(U3188) );
  AOI22_X1 U7414 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6497), .ZN(n6460) );
  OAI21_X1 U7415 ( .B1(n6461), .B2(n6500), .A(n6460), .ZN(U3189) );
  INV_X1 U7416 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6613) );
  OAI222_X1 U7417 ( .A1(n6496), .A2(n6461), .B1(n6613), .B2(n6547), .C1(n6463), 
        .C2(n6500), .ZN(U3190) );
  INV_X1 U7418 ( .A(n6500), .ZN(n6488) );
  AOI22_X1 U7419 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6497), .ZN(n6462) );
  OAI21_X1 U7420 ( .B1(n6463), .B2(n6496), .A(n6462), .ZN(U3191) );
  INV_X1 U7421 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6464) );
  INV_X1 U7422 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6647) );
  OAI222_X1 U7423 ( .A1(n6496), .A2(n6464), .B1(n6647), .B2(n6547), .C1(n6465), 
        .C2(n6500), .ZN(U3192) );
  INV_X1 U7424 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6604) );
  OAI222_X1 U7425 ( .A1(n6496), .A2(n6465), .B1(n6604), .B2(n6547), .C1(n6467), 
        .C2(n6500), .ZN(U3193) );
  AOI22_X1 U7426 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6497), .ZN(n6466) );
  OAI21_X1 U7427 ( .B1(n6467), .B2(n6496), .A(n6466), .ZN(U3194) );
  AOI22_X1 U7428 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6497), .ZN(n6468) );
  OAI21_X1 U7429 ( .B1(n6469), .B2(n6496), .A(n6468), .ZN(U3195) );
  AOI22_X1 U7430 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6497), .ZN(n6470) );
  OAI21_X1 U7431 ( .B1(n6471), .B2(n6496), .A(n6470), .ZN(U3196) );
  AOI22_X1 U7432 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6497), .ZN(n6472) );
  OAI21_X1 U7433 ( .B1(n6473), .B2(n6496), .A(n6472), .ZN(U3197) );
  AOI22_X1 U7434 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6497), .ZN(n6474) );
  OAI21_X1 U7435 ( .B1(n6475), .B2(n6500), .A(n6474), .ZN(U3198) );
  INV_X1 U7436 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6673) );
  OAI222_X1 U7437 ( .A1(n6496), .A2(n6475), .B1(n6673), .B2(n6547), .C1(n5434), 
        .C2(n6500), .ZN(U3199) );
  AOI22_X1 U7438 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6497), .ZN(n6476) );
  OAI21_X1 U7439 ( .B1(n5434), .B2(n6496), .A(n6476), .ZN(U3200) );
  INV_X1 U7440 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6478) );
  AOI22_X1 U7441 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6497), .ZN(n6477) );
  OAI21_X1 U7442 ( .B1(n6478), .B2(n6496), .A(n6477), .ZN(U3201) );
  AOI22_X1 U7443 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6497), .ZN(n6479) );
  OAI21_X1 U7444 ( .B1(n6481), .B2(n6500), .A(n6479), .ZN(U3202) );
  INV_X1 U7445 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6658) );
  OAI222_X1 U7446 ( .A1(n6496), .A2(n6481), .B1(n6658), .B2(n6547), .C1(n6480), 
        .C2(n6500), .ZN(U3203) );
  AOI22_X1 U7447 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6497), .ZN(n6482) );
  OAI21_X1 U7448 ( .B1(n6484), .B2(n6500), .A(n6482), .ZN(U3204) );
  AOI22_X1 U7449 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6497), .ZN(n6483) );
  OAI21_X1 U7450 ( .B1(n6484), .B2(n6496), .A(n6483), .ZN(U3205) );
  AOI22_X1 U7451 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6497), .ZN(n6485) );
  OAI21_X1 U7452 ( .B1(n6487), .B2(n6500), .A(n6485), .ZN(U3206) );
  AOI22_X1 U7453 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6497), .ZN(n6486) );
  OAI21_X1 U7454 ( .B1(n6487), .B2(n6496), .A(n6486), .ZN(U3207) );
  AOI22_X1 U7455 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6488), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6497), .ZN(n6489) );
  OAI21_X1 U7456 ( .B1(n6490), .B2(n6496), .A(n6489), .ZN(U3208) );
  AOI22_X1 U7457 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6497), .ZN(n6491) );
  OAI21_X1 U7458 ( .B1(n6611), .B2(n6500), .A(n6491), .ZN(U3209) );
  INV_X1 U7459 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6493) );
  AOI22_X1 U7460 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6497), .ZN(n6492) );
  OAI21_X1 U7461 ( .B1(n6493), .B2(n6500), .A(n6492), .ZN(U3210) );
  AOI22_X1 U7462 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6497), .ZN(n6494) );
  OAI21_X1 U7463 ( .B1(n6495), .B2(n6500), .A(n6494), .ZN(U3211) );
  INV_X1 U7464 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6580) );
  OAI222_X1 U7465 ( .A1(n6496), .A2(n6495), .B1(n6580), .B2(n6547), .C1(n4112), 
        .C2(n6500), .ZN(U3212) );
  INV_X1 U7466 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6501) );
  AOI22_X1 U7467 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6498), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6497), .ZN(n6499) );
  OAI21_X1 U7468 ( .B1(n6501), .B2(n6500), .A(n6499), .ZN(U3213) );
  MUX2_X1 U7469 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6547), .Z(U3445) );
  MUX2_X1 U7470 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6547), .Z(U3446) );
  MUX2_X1 U7471 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6547), .Z(U3447) );
  MUX2_X1 U7472 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6547), .Z(U3448) );
  INV_X1 U7473 ( .A(n6505), .ZN(n6502) );
  AOI21_X1 U7474 ( .B1(n6504), .B2(n6503), .A(n6502), .ZN(U3451) );
  OAI21_X1 U7475 ( .B1(n6507), .B2(n6506), .A(n6505), .ZN(U3452) );
  INV_X1 U7476 ( .A(n6508), .ZN(n6511) );
  OAI211_X1 U7477 ( .C1(n6512), .C2(n6511), .A(n6510), .B(n6509), .ZN(U3453)
         );
  INV_X1 U7478 ( .A(n6513), .ZN(n6516) );
  OAI22_X1 U7479 ( .A1(n6516), .A2(n6525), .B1(n6515), .B2(n6514), .ZN(n6517)
         );
  MUX2_X1 U7480 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6517), .S(n6521), 
        .Z(U3456) );
  OR2_X1 U7481 ( .A1(n6518), .A2(n6525), .ZN(n6519) );
  OAI21_X1 U7482 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6520), .A(n6519), 
        .ZN(n6523) );
  OAI22_X1 U7483 ( .A1(n6523), .A2(n6522), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6521), .ZN(n6524) );
  OAI21_X1 U7484 ( .B1(n6526), .B2(n6525), .A(n6524), .ZN(U3461) );
  AOI21_X1 U7485 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U7486 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6528), .B2(n6527), .ZN(n6531) );
  INV_X1 U7487 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6530) );
  AOI22_X1 U7488 ( .A1(n6534), .A2(n6531), .B1(n6530), .B2(n6529), .ZN(U3468)
         );
  INV_X1 U7489 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6533) );
  OAI21_X1 U7490 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6534), .ZN(n6532) );
  OAI21_X1 U7491 ( .B1(n6534), .B2(n6533), .A(n6532), .ZN(U3469) );
  NAND2_X1 U7492 ( .A1(n6497), .A2(W_R_N_REG_SCAN_IN), .ZN(n6535) );
  OAI21_X1 U7493 ( .B1(n6497), .B2(READREQUEST_REG_SCAN_IN), .A(n6535), .ZN(
        U3470) );
  AOI211_X1 U7494 ( .C1(n6539), .C2(n6538), .A(n6537), .B(n6536), .ZN(n6546)
         );
  OAI211_X1 U7495 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6541), .A(n6540), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6543) );
  AOI21_X1 U7496 ( .B1(n6543), .B2(STATE2_REG_0__SCAN_IN), .A(n6542), .ZN(
        n6545) );
  NAND2_X1 U7497 ( .A1(n6546), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6544) );
  OAI21_X1 U7498 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(U3472) );
  MUX2_X1 U7499 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6547), .Z(U3473) );
  AOI22_X1 U7500 ( .A1(n6550), .A2(n6549), .B1(INSTQUEUE_REG_6__7__SCAN_IN), 
        .B2(n6548), .ZN(n6551) );
  OAI21_X1 U7501 ( .B1(n6553), .B2(n6552), .A(n6551), .ZN(n6554) );
  AOI21_X1 U7502 ( .B1(n6556), .B2(n6555), .A(n6554), .ZN(n6557) );
  OAI21_X1 U7503 ( .B1(n6559), .B2(n6558), .A(n6557), .ZN(n6719) );
  INV_X1 U7504 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6703) );
  AOI22_X1 U7505 ( .A1(n6703), .A2(keyinput40), .B1(keyinput4), .B2(n6561), 
        .ZN(n6560) );
  OAI221_X1 U7506 ( .B1(n6703), .B2(keyinput40), .C1(n6561), .C2(keyinput4), 
        .A(n6560), .ZN(n6565) );
  XNOR2_X1 U7507 ( .A(n6562), .B(keyinput0), .ZN(n6564) );
  XOR2_X1 U7508 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput31), .Z(n6563)
         );
  OR3_X1 U7509 ( .A1(n6565), .A2(n6564), .A3(n6563), .ZN(n6574) );
  INV_X1 U7510 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6567) );
  AOI22_X1 U7511 ( .A1(n6568), .A2(keyinput21), .B1(n6567), .B2(keyinput8), 
        .ZN(n6566) );
  OAI221_X1 U7512 ( .B1(n6568), .B2(keyinput21), .C1(n6567), .C2(keyinput8), 
        .A(n6566), .ZN(n6573) );
  AOI22_X1 U7513 ( .A1(n6571), .A2(keyinput39), .B1(n6570), .B2(keyinput57), 
        .ZN(n6569) );
  OAI221_X1 U7514 ( .B1(n6571), .B2(keyinput39), .C1(n6570), .C2(keyinput57), 
        .A(n6569), .ZN(n6572) );
  NOR3_X1 U7515 ( .A1(n6574), .A2(n6573), .A3(n6572), .ZN(n6621) );
  INV_X1 U7516 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6576) );
  AOI22_X1 U7517 ( .A1(n6686), .A2(keyinput2), .B1(keyinput61), .B2(n6576), 
        .ZN(n6575) );
  OAI221_X1 U7518 ( .B1(n6686), .B2(keyinput2), .C1(n6576), .C2(keyinput61), 
        .A(n6575), .ZN(n6587) );
  AOI22_X1 U7519 ( .A1(n6578), .A2(keyinput24), .B1(keyinput44), .B2(n6694), 
        .ZN(n6577) );
  OAI221_X1 U7520 ( .B1(n6578), .B2(keyinput24), .C1(n6694), .C2(keyinput44), 
        .A(n6577), .ZN(n6586) );
  AOI22_X1 U7521 ( .A1(n6580), .A2(keyinput27), .B1(n3956), .B2(keyinput23), 
        .ZN(n6579) );
  OAI221_X1 U7522 ( .B1(n6580), .B2(keyinput27), .C1(n3956), .C2(keyinput23), 
        .A(n6579), .ZN(n6585) );
  INV_X1 U7523 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6583) );
  AOI22_X1 U7524 ( .A1(n6583), .A2(keyinput29), .B1(keyinput52), .B2(n6582), 
        .ZN(n6581) );
  OAI221_X1 U7525 ( .B1(n6583), .B2(keyinput29), .C1(n6582), .C2(keyinput52), 
        .A(n6581), .ZN(n6584) );
  NOR4_X1 U7526 ( .A1(n6587), .A2(n6586), .A3(n6585), .A4(n6584), .ZN(n6620)
         );
  AOI22_X1 U7527 ( .A1(n6590), .A2(keyinput56), .B1(keyinput45), .B2(n6589), 
        .ZN(n6588) );
  OAI221_X1 U7528 ( .B1(n6590), .B2(keyinput56), .C1(n6589), .C2(keyinput45), 
        .A(n6588), .ZN(n6602) );
  INV_X1 U7529 ( .A(DATAI_10_), .ZN(n6593) );
  AOI22_X1 U7530 ( .A1(n6593), .A2(keyinput14), .B1(keyinput50), .B2(n6592), 
        .ZN(n6591) );
  OAI221_X1 U7531 ( .B1(n6593), .B2(keyinput14), .C1(n6592), .C2(keyinput50), 
        .A(n6591), .ZN(n6601) );
  AOI22_X1 U7532 ( .A1(n6596), .A2(keyinput48), .B1(n6595), .B2(keyinput17), 
        .ZN(n6594) );
  OAI221_X1 U7533 ( .B1(n6596), .B2(keyinput48), .C1(n6595), .C2(keyinput17), 
        .A(n6594), .ZN(n6600) );
  XNOR2_X1 U7534 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .B(keyinput6), .ZN(
        n6598) );
  XNOR2_X1 U7535 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .B(keyinput9), .ZN(n6597)
         );
  NAND2_X1 U7536 ( .A1(n6598), .A2(n6597), .ZN(n6599) );
  NOR4_X1 U7537 ( .A1(n6602), .A2(n6601), .A3(n6600), .A4(n6599), .ZN(n6619)
         );
  AOI22_X1 U7538 ( .A1(n6605), .A2(keyinput54), .B1(n6604), .B2(keyinput59), 
        .ZN(n6603) );
  OAI221_X1 U7539 ( .B1(n6605), .B2(keyinput54), .C1(n6604), .C2(keyinput59), 
        .A(n6603), .ZN(n6617) );
  INV_X1 U7540 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6607) );
  AOI22_X1 U7541 ( .A1(n6608), .A2(keyinput15), .B1(n6607), .B2(keyinput19), 
        .ZN(n6606) );
  OAI221_X1 U7542 ( .B1(n6608), .B2(keyinput15), .C1(n6607), .C2(keyinput19), 
        .A(n6606), .ZN(n6616) );
  AOI22_X1 U7543 ( .A1(n6611), .A2(keyinput11), .B1(keyinput60), .B2(n6610), 
        .ZN(n6609) );
  OAI221_X1 U7544 ( .B1(n6611), .B2(keyinput11), .C1(n6610), .C2(keyinput60), 
        .A(n6609), .ZN(n6615) );
  AOI22_X1 U7545 ( .A1(n3339), .A2(keyinput18), .B1(keyinput33), .B2(n6613), 
        .ZN(n6612) );
  OAI221_X1 U7546 ( .B1(n3339), .B2(keyinput18), .C1(n6613), .C2(keyinput33), 
        .A(n6612), .ZN(n6614) );
  NOR4_X1 U7547 ( .A1(n6617), .A2(n6616), .A3(n6615), .A4(n6614), .ZN(n6618)
         );
  NAND4_X1 U7548 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n6685)
         );
  INV_X1 U7549 ( .A(DATAI_16_), .ZN(n6624) );
  AOI22_X1 U7550 ( .A1(n6624), .A2(keyinput47), .B1(keyinput62), .B2(n6623), 
        .ZN(n6622) );
  OAI221_X1 U7551 ( .B1(n6624), .B2(keyinput47), .C1(n6623), .C2(keyinput62), 
        .A(n6622), .ZN(n6636) );
  INV_X1 U7552 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U7553 ( .A1(n6627), .A2(keyinput35), .B1(keyinput7), .B2(n6626), 
        .ZN(n6625) );
  OAI221_X1 U7554 ( .B1(n6627), .B2(keyinput35), .C1(n6626), .C2(keyinput7), 
        .A(n6625), .ZN(n6635) );
  AOI22_X1 U7555 ( .A1(n6630), .A2(keyinput22), .B1(keyinput28), .B2(n6629), 
        .ZN(n6628) );
  OAI221_X1 U7556 ( .B1(n6630), .B2(keyinput22), .C1(n6629), .C2(keyinput28), 
        .A(n6628), .ZN(n6634) );
  AOI22_X1 U7557 ( .A1(n5836), .A2(keyinput58), .B1(keyinput3), .B2(n6632), 
        .ZN(n6631) );
  OAI221_X1 U7558 ( .B1(n5836), .B2(keyinput58), .C1(n6632), .C2(keyinput3), 
        .A(n6631), .ZN(n6633) );
  NOR4_X1 U7559 ( .A1(n6636), .A2(n6635), .A3(n6634), .A4(n6633), .ZN(n6683)
         );
  AOI22_X1 U7560 ( .A1(n6639), .A2(keyinput38), .B1(keyinput36), .B2(n6638), 
        .ZN(n6637) );
  OAI221_X1 U7561 ( .B1(n6639), .B2(keyinput38), .C1(n6638), .C2(keyinput36), 
        .A(n6637), .ZN(n6651) );
  AOI22_X1 U7562 ( .A1(n6642), .A2(keyinput16), .B1(n6641), .B2(keyinput49), 
        .ZN(n6640) );
  OAI221_X1 U7563 ( .B1(n6642), .B2(keyinput16), .C1(n6641), .C2(keyinput49), 
        .A(n6640), .ZN(n6650) );
  AOI22_X1 U7564 ( .A1(n5931), .A2(keyinput55), .B1(n6644), .B2(keyinput10), 
        .ZN(n6643) );
  OAI221_X1 U7565 ( .B1(n5931), .B2(keyinput55), .C1(n6644), .C2(keyinput10), 
        .A(n6643), .ZN(n6649) );
  AOI22_X1 U7566 ( .A1(n6647), .A2(keyinput5), .B1(n6646), .B2(keyinput42), 
        .ZN(n6645) );
  OAI221_X1 U7567 ( .B1(n6647), .B2(keyinput5), .C1(n6646), .C2(keyinput42), 
        .A(n6645), .ZN(n6648) );
  NOR4_X1 U7568 ( .A1(n6651), .A2(n6650), .A3(n6649), .A4(n6648), .ZN(n6682)
         );
  INV_X1 U7569 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6687) );
  AOI22_X1 U7570 ( .A1(n6687), .A2(keyinput53), .B1(keyinput37), .B2(n6653), 
        .ZN(n6652) );
  OAI221_X1 U7571 ( .B1(n6687), .B2(keyinput53), .C1(n6653), .C2(keyinput37), 
        .A(n6652), .ZN(n6664) );
  AOI22_X1 U7572 ( .A1(n6655), .A2(keyinput26), .B1(n6699), .B2(keyinput32), 
        .ZN(n6654) );
  OAI221_X1 U7573 ( .B1(n6655), .B2(keyinput26), .C1(n6699), .C2(keyinput32), 
        .A(n6654), .ZN(n6663) );
  AOI22_X1 U7574 ( .A1(n6658), .A2(keyinput1), .B1(n6657), .B2(keyinput12), 
        .ZN(n6656) );
  OAI221_X1 U7575 ( .B1(n6658), .B2(keyinput1), .C1(n6657), .C2(keyinput12), 
        .A(n6656), .ZN(n6662) );
  INV_X1 U7576 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6688) );
  AOI22_X1 U7577 ( .A1(n6660), .A2(keyinput30), .B1(n6688), .B2(keyinput46), 
        .ZN(n6659) );
  OAI221_X1 U7578 ( .B1(n6660), .B2(keyinput30), .C1(n6688), .C2(keyinput46), 
        .A(n6659), .ZN(n6661) );
  NOR4_X1 U7579 ( .A1(n6664), .A2(n6663), .A3(n6662), .A4(n6661), .ZN(n6681)
         );
  INV_X1 U7580 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6667) );
  AOI22_X1 U7581 ( .A1(n6667), .A2(keyinput41), .B1(keyinput34), .B2(n6666), 
        .ZN(n6665) );
  OAI221_X1 U7582 ( .B1(n6667), .B2(keyinput41), .C1(n6666), .C2(keyinput34), 
        .A(n6665), .ZN(n6679) );
  AOI22_X1 U7583 ( .A1(n6670), .A2(keyinput20), .B1(keyinput13), .B2(n6669), 
        .ZN(n6668) );
  OAI221_X1 U7584 ( .B1(n6670), .B2(keyinput20), .C1(n6669), .C2(keyinput13), 
        .A(n6668), .ZN(n6678) );
  AOI22_X1 U7585 ( .A1(n6673), .A2(keyinput63), .B1(n6672), .B2(keyinput25), 
        .ZN(n6671) );
  OAI221_X1 U7586 ( .B1(n6673), .B2(keyinput63), .C1(n6672), .C2(keyinput25), 
        .A(n6671), .ZN(n6677) );
  XNOR2_X1 U7587 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput43), .ZN(n6675)
         );
  XNOR2_X1 U7588 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .B(keyinput51), .ZN(n6674) );
  NAND2_X1 U7589 ( .A1(n6675), .A2(n6674), .ZN(n6676) );
  NOR4_X1 U7590 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6680)
         );
  NAND4_X1 U7591 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6684)
         );
  NOR2_X1 U7592 ( .A1(n6685), .A2(n6684), .ZN(n6717) );
  NAND4_X1 U7593 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n6688), .A3(n6687), 
        .A4(n6686), .ZN(n6715) );
  NAND2_X1 U7594 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n6689), .ZN(n6690) );
  NOR4_X1 U7595 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n6690), .A3(
        INSTQUEUE_REG_11__0__SCAN_IN), .A4(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n6691) );
  NAND3_X1 U7596 ( .A1(n6693), .A2(n6692), .A3(n6691), .ZN(n6714) );
  NOR4_X1 U7597 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(EBX_REG_9__SCAN_IN), 
        .A3(DATAO_REG_1__SCAN_IN), .A4(MORE_REG_SCAN_IN), .ZN(n6698) );
  NOR4_X1 U7598 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(EAX_REG_8__SCAN_IN), 
        .A3(DATAI_16_), .A4(LWORD_REG_13__SCAN_IN), .ZN(n6697) );
  NOR4_X1 U7599 ( .A1(EBX_REG_28__SCAN_IN), .A2(EBX_REG_23__SCAN_IN), .A3(
        EAX_REG_23__SCAN_IN), .A4(UWORD_REG_6__SCAN_IN), .ZN(n6696) );
  NOR4_X1 U7600 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(
        REIP_REG_23__SCAN_IN), .A3(DATAI_10_), .A4(n6694), .ZN(n6695) );
  NAND4_X1 U7601 ( .A1(n6698), .A2(n6697), .A3(n6696), .A4(n6695), .ZN(n6713)
         );
  NAND4_X1 U7602 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(DATAI_4_), .A4(n6699), .ZN(n6702) );
  NAND4_X1 U7603 ( .A1(EBX_REG_20__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        DATAI_9_), .A4(DATAI_8_), .ZN(n6701) );
  NAND4_X1 U7604 ( .A1(ADDRESS_REG_28__SCAN_IN), .A2(DATAO_REG_13__SCAN_IN), 
        .A3(DATAO_REG_5__SCAN_IN), .A4(ADDRESS_REG_0__SCAN_IN), .ZN(n6700) );
  NOR3_X1 U7605 ( .A1(n6702), .A2(n6701), .A3(n6700), .ZN(n6705) );
  NOR2_X1 U7606 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6703), .ZN(n6704) );
  AND4_X1 U7607 ( .A1(n6705), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .A3(n6704), 
        .A4(n6607), .ZN(n6711) );
  NAND4_X1 U7608 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(EAX_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(UWORD_REG_2__SCAN_IN), .ZN(n6708) );
  NAND4_X1 U7609 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(MEMORYFETCH_REG_SCAN_IN), 
        .A3(ADDRESS_REG_15__SCAN_IN), .A4(UWORD_REG_5__SCAN_IN), .ZN(n6707) );
  NAND3_X1 U7610 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        EBX_REG_21__SCAN_IN), .A3(REIP_REG_6__SCAN_IN), .ZN(n6706) );
  NOR4_X1 U7611 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6708), .A3(n6707), .A4(
        n6706), .ZN(n6710) );
  NOR4_X1 U7612 ( .A1(UWORD_REG_11__SCAN_IN), .A2(ADDRESS_REG_19__SCAN_IN), 
        .A3(ADDRESS_REG_9__SCAN_IN), .A4(ADDRESS_REG_8__SCAN_IN), .ZN(n6709)
         );
  NAND3_X1 U7613 ( .A1(n6711), .A2(n6710), .A3(n6709), .ZN(n6712) );
  NOR4_X1 U7614 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6716)
         );
  XNOR2_X1 U7615 ( .A(n6717), .B(n6716), .ZN(n6718) );
  XNOR2_X1 U7616 ( .A(n6719), .B(n6718), .ZN(U3075) );
  AND2_X2 U3937 ( .A1(n3053), .A2(n3047), .ZN(n3271) );
  AND4_X1 U3972 ( .A1(n3086), .A2(n3085), .A3(n3084), .A4(n3083), .ZN(n3092)
         );
  AND4_X1 U3959 ( .A1(n3074), .A2(n3073), .A3(n3072), .A4(n3071), .ZN(n3107)
         );
  XNOR2_X1 U3521 ( .A(n3292), .B(n3288), .ZN(n3300) );
  CLKBUF_X1 U3401 ( .A(n3265), .Z(n3363) );
  AND4_X1 U3423 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .ZN(n3091)
         );
  NOR2_X1 U3427 ( .A1(n3889), .A2(n4360), .ZN(n4373) );
  AOI21_X1 U3428 ( .B1(n3300), .B2(n3299), .A(n3293), .ZN(n3295) );
  CLKBUF_X1 U3502 ( .A(n3905), .Z(n5274) );
  AND2_X1 U3504 ( .A1(n3826), .A2(n3306), .ZN(n4890) );
  CLKBUF_X1 U3507 ( .A(n3186), .Z(n4337) );
  OAI21_X1 U3518 ( .B1(n4517), .B2(n4158), .A(n4176), .ZN(n4177) );
  INV_X1 U3561 ( .A(n4226), .ZN(n2953) );
  CLKBUF_X1 U3667 ( .A(n3188), .Z(n4487) );
  NOR2_X1 U3716 ( .A1(n5398), .A2(n5399), .ZN(n5397) );
  NAND2_X1 U3728 ( .A1(n5371), .A2(n4242), .ZN(n5412) );
  CLKBUF_X1 U3814 ( .A(n4459), .Z(n5624) );
  NAND2_X1 U3816 ( .A1(n3225), .A2(n3224), .ZN(n3250) );
  OAI21_X1 U4072 ( .B1(n3226), .B2(n3250), .A(n3225), .ZN(n3233) );
  NAND3_X1 U4079 ( .A1(n3219), .A2(n3220), .A3(n3218), .ZN(n3225) );
  NAND2_X1 U4082 ( .A1(n5441), .A2(n6720), .ZN(n5371) );
  AND2_X1 U4092 ( .A1(n4239), .A2(n4240), .ZN(n6720) );
  OR2_X1 U4112 ( .A1(n2953), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6721)
         );
  NAND2_X1 U5109 ( .A1(n6721), .A2(n5374), .ZN(n5393) );
  AND2_X1 U5182 ( .A1(n5441), .A2(n4239), .ZN(n5419) );
  CLKBUF_X1 U5185 ( .A(n3256), .Z(n3309) );
endmodule

