

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204;

  NOR3_X2 U7286 ( .A1(n14885), .A2(n10181), .A3(n8316), .ZN(n14845) );
  NAND2_X1 U7287 ( .A1(n7775), .A2(n14886), .ZN(n14885) );
  NAND2_X1 U7288 ( .A1(n16170), .A2(n14426), .ZN(n14432) );
  INV_X1 U7289 ( .A(n9352), .ZN(n9177) );
  INV_X4 U7290 ( .A(n13365), .ZN(n13340) );
  INV_X2 U7291 ( .A(n7191), .ZN(n13350) );
  CLKBUF_X1 U7292 ( .A(n14737), .Z(n7185) );
  OAI21_X1 U7293 ( .B1(n11562), .B2(n11559), .A(n15931), .ZN(n14737) );
  INV_X2 U7294 ( .A(n14585), .ZN(n14526) );
  OR2_X1 U7295 ( .A1(n13950), .A2(n7421), .ZN(n7420) );
  INV_X1 U7296 ( .A(n10835), .ZN(n10857) );
  CLKBUF_X2 U7297 ( .A(n11917), .Z(n14533) );
  OAI21_X1 U7298 ( .B1(n10995), .B2(n8937), .A(n8637), .ZN(n12437) );
  INV_X1 U7299 ( .A(n8421), .ZN(n8504) );
  INV_X1 U7301 ( .A(n11967), .ZN(n11878) );
  INV_X1 U7303 ( .A(n10551), .ZN(n13357) );
  OR2_X2 U7304 ( .A1(n14082), .A2(n14271), .ZN(n14075) );
  INV_X1 U7305 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n10415) );
  NOR2_X1 U7306 ( .A1(n14885), .A2(n15042), .ZN(n14872) );
  NAND2_X2 U7307 ( .A1(n11437), .A2(n8990), .ZN(n14589) );
  AND4_X1 U7308 ( .A1(n8570), .A2(n8569), .A3(n8568), .A4(n8567), .ZN(n15915)
         );
  INV_X2 U7309 ( .A(n8424), .ZN(n8421) );
  AND4_X1 U7310 ( .A1(n9107), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(n11418)
         );
  NAND2_X1 U7311 ( .A1(n9260), .A2(n9259), .ZN(n9277) );
  OAI21_X1 U7312 ( .B1(n11043), .B2(n7191), .A(n10465), .ZN(n13216) );
  NAND2_X1 U7313 ( .A1(n12559), .A2(n7425), .ZN(n12600) );
  NAND2_X1 U7314 ( .A1(n8709), .A2(n8708), .ZN(n14560) );
  INV_X1 U7315 ( .A(n8901), .ZN(n8977) );
  BUF_X1 U7316 ( .A(n15915), .Z(n7694) );
  NAND2_X1 U7317 ( .A1(n8632), .A2(n8631), .ZN(n8634) );
  INV_X2 U7318 ( .A(n16041), .ZN(n16156) );
  NAND2_X1 U7319 ( .A1(n10444), .A2(n10443), .ZN(n13399) );
  OR2_X1 U7320 ( .A1(n13285), .A2(n13284), .ZN(n7186) );
  AOI21_X2 U7321 ( .B1(n12976), .B2(n7988), .A(n7986), .ZN(n7985) );
  NAND2_X2 U7322 ( .A1(n9616), .A2(n12969), .ZN(n12976) );
  AOI21_X2 U7323 ( .B1(n13625), .B2(n9546), .A(n9545), .ZN(n9876) );
  NOR2_X2 U7324 ( .A1(n15838), .A2(n15839), .ZN(n15837) );
  NOR2_X2 U7325 ( .A1(n14919), .A2(n15055), .ZN(n7775) );
  NAND2_X2 U7326 ( .A1(n11638), .A2(n10618), .ZN(n11868) );
  INV_X1 U7327 ( .A(n8517), .ZN(n8512) );
  INV_X2 U7328 ( .A(n10109), .ZN(n10188) );
  OAI21_X2 U7329 ( .B1(n8634), .B2(n8433), .A(n7547), .ZN(n8666) );
  INV_X1 U7330 ( .A(n9140), .ZN(n9160) );
  INV_X1 U7331 ( .A(n11438), .ZN(n11437) );
  OAI21_X1 U7332 ( .B1(n11838), .B2(n8352), .A(n7278), .ZN(n7391) );
  OAI21_X2 U7333 ( .B1(n11836), .B2(n11835), .A(n14563), .ZN(n11838) );
  AOI21_X2 U7334 ( .B1(n10434), .B2(P2_IR_REG_22__SCAN_IN), .A(n10433), .ZN(
        n10435) );
  OAI211_X2 U7335 ( .C1(n7363), .C2(P2_IR_REG_31__SCAN_IN), .A(n7361), .B(
        n7360), .ZN(n10417) );
  INV_X4 U7337 ( .A(n7529), .ZN(n8972) );
  AOI21_X1 U7338 ( .B1(n7960), .B2(n7212), .A(n7195), .ZN(n7851) );
  NAND2_X1 U7339 ( .A1(n7282), .A2(n7212), .ZN(n7852) );
  OR2_X1 U7340 ( .A1(n10139), .A2(n10140), .ZN(n10141) );
  AOI21_X1 U7341 ( .B1(n13063), .B2(n14121), .A(n7488), .ZN(n14276) );
  AND2_X1 U7342 ( .A1(n7365), .A2(n8060), .ZN(n13063) );
  XNOR2_X1 U7343 ( .A(n8983), .B(n10227), .ZN(n14862) );
  OAI21_X1 U7344 ( .B1(n8041), .B2(n9859), .A(n11657), .ZN(n8040) );
  OR2_X1 U7345 ( .A1(n8041), .A2(n8039), .ZN(n8038) );
  NAND2_X1 U7346 ( .A1(n10853), .A2(n7222), .ZN(n13989) );
  NAND2_X1 U7347 ( .A1(n7487), .A2(n7486), .ZN(n14088) );
  NAND2_X1 U7348 ( .A1(n13919), .A2(n13920), .ZN(n10853) );
  NOR2_X1 U7349 ( .A1(n8317), .A2(n14878), .ZN(n14874) );
  NOR2_X1 U7350 ( .A1(n14896), .A2(n14898), .ZN(n14895) );
  AND2_X1 U7351 ( .A1(n10822), .A2(n10836), .ZN(n8215) );
  NAND2_X1 U7352 ( .A1(n7359), .A2(n8051), .ZN(n14133) );
  NAND2_X1 U7353 ( .A1(n7431), .A2(n7430), .ZN(n13904) );
  AOI21_X1 U7354 ( .B1(n12789), .B2(n9707), .A(n7319), .ZN(n12971) );
  AND2_X1 U7355 ( .A1(n8203), .A2(n7211), .ZN(n7430) );
  NAND2_X1 U7356 ( .A1(n7482), .A2(n7480), .ZN(n13000) );
  NAND2_X1 U7357 ( .A1(n10807), .A2(n10806), .ZN(n14295) );
  NAND2_X1 U7358 ( .A1(n8537), .A2(n8536), .ZN(n15073) );
  AND2_X1 U7359 ( .A1(n12952), .A2(n12829), .ZN(n12831) );
  OAI22_X1 U7360 ( .A1(n12445), .A2(n8167), .B1(n16108), .B2(n13578), .ZN(
        n12651) );
  OAI21_X1 U7361 ( .B1(n12600), .B2(n8219), .A(n8216), .ZN(n8228) );
  NAND2_X1 U7362 ( .A1(n8866), .A2(n8865), .ZN(n15105) );
  AND2_X1 U7363 ( .A1(n8206), .A2(n8205), .ZN(n8208) );
  AND2_X1 U7364 ( .A1(n8846), .A2(n8860), .ZN(n12384) );
  NOR2_X1 U7365 ( .A1(n12936), .A2(n14449), .ZN(n8324) );
  AND2_X1 U7366 ( .A1(n8841), .A2(n8859), .ZN(n8845) );
  OR2_X1 U7367 ( .A1(n8893), .A2(n8892), .ZN(n8895) );
  NAND2_X1 U7368 ( .A1(n10723), .A2(n10722), .ZN(n14332) );
  INV_X2 U7369 ( .A(n13637), .ZN(n13115) );
  OAI21_X1 U7370 ( .B1(n8826), .B2(n8825), .A(n8460), .ZN(n8839) );
  OAI21_X1 U7371 ( .B1(n9400), .B2(n8028), .A(n8025), .ZN(n9420) );
  NAND2_X1 U7372 ( .A1(n8457), .A2(n8456), .ZN(n8826) );
  NAND2_X1 U7373 ( .A1(n10476), .A2(n10475), .ZN(n13210) );
  OR2_X1 U7374 ( .A1(n8809), .A2(n8807), .ZN(n8457) );
  NAND2_X1 U7375 ( .A1(n8706), .A2(n8705), .ZN(n11043) );
  NAND2_X1 U7376 ( .A1(n8704), .A2(n8685), .ZN(n11041) );
  NAND2_X1 U7377 ( .A1(n8755), .A2(n8449), .ZN(n8772) );
  NAND2_X1 U7378 ( .A1(n7805), .A2(n7803), .ZN(n8720) );
  NAND2_X1 U7379 ( .A1(n9760), .A2(n9763), .ZN(n9713) );
  AND2_X1 U7380 ( .A1(n9768), .A2(n9765), .ZN(n11957) );
  INV_X1 U7381 ( .A(n13588), .ZN(n11228) );
  NAND2_X1 U7382 ( .A1(n10511), .A2(n10510), .ZN(n13168) );
  INV_X2 U7383 ( .A(n13715), .ZN(n7188) );
  NAND2_X1 U7384 ( .A1(n8595), .A2(n8594), .ZN(n14566) );
  NAND2_X1 U7385 ( .A1(n13590), .A2(n11669), .ZN(n11494) );
  INV_X1 U7386 ( .A(n12281), .ZN(n8581) );
  NOR2_X1 U7387 ( .A1(P2_U3088), .A2(n11057), .ZN(P2_U3947) );
  NAND2_X1 U7388 ( .A1(n8280), .A2(n8580), .ZN(n12281) );
  NAND4_X1 U7389 ( .A1(n9094), .A2(n9093), .A3(n9092), .A4(n9091), .ZN(n13590)
         );
  AND4_X1 U7390 ( .A1(n9121), .A2(n9120), .A3(n9119), .A4(n9118), .ZN(n15961)
         );
  INV_X1 U7391 ( .A(n11669), .ZN(n11592) );
  NAND2_X1 U7392 ( .A1(n9115), .A2(n9114), .ZN(n15970) );
  NAND2_X1 U7393 ( .A1(n10549), .A2(n10548), .ZN(n14248) );
  NOR2_X2 U7394 ( .A1(n9961), .A2(n9966), .ZN(n15844) );
  INV_X1 U7395 ( .A(n15934), .ZN(n15917) );
  INV_X1 U7396 ( .A(n7694), .ZN(n14768) );
  AND2_X1 U7397 ( .A1(n7696), .A2(n7532), .ZN(n15934) );
  INV_X1 U7398 ( .A(n9080), .ZN(n13881) );
  BUF_X2 U7399 ( .A(n10109), .Z(n10182) );
  NAND2_X1 U7400 ( .A1(n10517), .A2(n7224), .ZN(n14026) );
  NAND4_X1 U7401 ( .A1(n10557), .A2(n10556), .A3(n10555), .A4(n10554), .ZN(
        n14027) );
  NAND2_X2 U7402 ( .A1(n10941), .A2(n13024), .ZN(n10938) );
  INV_X8 U7403 ( .A(n13393), .ZN(n13365) );
  XNOR2_X1 U7404 ( .A(n9074), .B(n13872), .ZN(n9078) );
  INV_X2 U7405 ( .A(n10519), .ZN(n10552) );
  OAI21_X1 U7406 ( .B1(n11054), .B2(P2_IR_REG_0__SCAN_IN), .A(n10528), .ZN(
        n15895) );
  INV_X2 U7407 ( .A(n8937), .ZN(n10171) );
  OAI211_X1 U7408 ( .C1(P3_IR_REG_31__SCAN_IN), .C2(P3_IR_REG_28__SCAN_IN), 
        .A(n9088), .B(n8148), .ZN(n9598) );
  NAND2_X1 U7409 ( .A1(n9076), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9074) );
  NAND2_X2 U7410 ( .A1(n8563), .A2(n8421), .ZN(n8937) );
  NAND2_X2 U7411 ( .A1(n8512), .A2(n15156), .ZN(n8976) );
  AND2_X1 U7412 ( .A1(n10042), .A2(n12389), .ZN(n11438) );
  NAND2_X2 U7413 ( .A1(n13464), .A2(n10425), .ZN(n10553) );
  CLKBUF_X3 U7414 ( .A(n9969), .Z(n13132) );
  AND2_X2 U7415 ( .A1(n8517), .A2(n8518), .ZN(n8951) );
  INV_X1 U7416 ( .A(n8518), .ZN(n15156) );
  XNOR2_X1 U7417 ( .A(n8348), .B(P1_IR_REG_22__SCAN_IN), .ZN(n10040) );
  INV_X1 U7418 ( .A(n10425), .ZN(n14372) );
  NAND2_X1 U7419 ( .A1(n7406), .A2(n7404), .ZN(n13455) );
  XNOR2_X1 U7420 ( .A(n7364), .B(P2_IR_REG_29__SCAN_IN), .ZN(n10425) );
  XNOR2_X1 U7421 ( .A(n9424), .B(n9423), .ZN(n11505) );
  NAND2_X1 U7422 ( .A1(n8509), .A2(n8502), .ZN(n15161) );
  NAND2_X1 U7423 ( .A1(n7217), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8348) );
  OR2_X1 U7424 ( .A1(n14365), .A2(n7362), .ZN(n7361) );
  NAND2_X2 U7425 ( .A1(n10986), .A2(P1_U3086), .ZN(n15157) );
  XNOR2_X1 U7426 ( .A(n10442), .B(P2_IR_REG_21__SCAN_IN), .ZN(n13445) );
  MUX2_X1 U7427 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8501), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n8502) );
  NAND2_X2 U7428 ( .A1(n10986), .A2(P2_U3088), .ZN(n14378) );
  XNOR2_X1 U7429 ( .A(n8864), .B(P1_IR_REG_19__SCAN_IN), .ZN(n14835) );
  NAND2_X1 U7430 ( .A1(n10447), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7364) );
  INV_X1 U7431 ( .A(n13024), .ZN(n10458) );
  NOR2_X1 U7432 ( .A1(n7407), .A2(n7265), .ZN(n7406) );
  NAND2_X2 U7433 ( .A1(n10986), .A2(P3_U3151), .ZN(n13880) );
  NAND2_X1 U7434 ( .A1(n7405), .A2(n7257), .ZN(n7404) );
  NOR2_X1 U7435 ( .A1(n10436), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n10431) );
  NAND2_X1 U7436 ( .A1(n8421), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8141) );
  NAND4_X1 U7437 ( .A1(n7197), .A2(n8792), .A3(n8394), .A4(n8491), .ZN(n8863)
         );
  NAND2_X1 U7438 ( .A1(n7732), .A2(n7731), .ZN(n10446) );
  AND2_X2 U7439 ( .A1(n7506), .A2(n8578), .ZN(n8792) );
  NAND2_X1 U7440 ( .A1(n7932), .A2(n7933), .ZN(n8424) );
  AND2_X1 U7441 ( .A1(n8171), .A2(n8170), .ZN(n8169) );
  AND2_X1 U7442 ( .A1(n10438), .A2(n10412), .ZN(n8411) );
  AND2_X1 U7443 ( .A1(n7403), .A2(n7402), .ZN(n10438) );
  AND4_X1 U7444 ( .A1(n10706), .A2(n10410), .A3(n10449), .A4(n10705), .ZN(
        n10411) );
  AND3_X1 U7445 ( .A1(n10407), .A2(n10460), .A3(n8043), .ZN(n8042) );
  AND4_X1 U7446 ( .A1(n8498), .A2(n8497), .A3(n8496), .A4(n8400), .ZN(n8412)
         );
  AND2_X1 U7447 ( .A1(n8491), .A2(n8490), .ZN(n7505) );
  AND2_X1 U7448 ( .A1(n8554), .A2(n8495), .ZN(n8578) );
  AND2_X1 U7449 ( .A1(n9084), .A2(n7543), .ZN(n9108) );
  AND2_X1 U7450 ( .A1(n9063), .A2(n9070), .ZN(n8171) );
  NOR2_X1 U7451 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n8487) );
  NOR2_X1 U7452 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8488) );
  INV_X1 U7453 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8813) );
  INV_X1 U7454 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9645) );
  NOR2_X1 U7455 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n8346) );
  NOR2_X1 U7456 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8345) );
  INV_X4 U7457 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7458 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n10430) );
  INV_X1 U7459 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10705) );
  NOR2_X1 U7460 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n10706) );
  INV_X1 U7461 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8043) );
  INV_X1 U7462 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10915) );
  INV_X4 U7463 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7464 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10926) );
  INV_X1 U7465 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n10919) );
  NOR2_X1 U7466 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n10412) );
  INV_X1 U7467 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n10449) );
  NOR2_X1 U7468 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n10408) );
  NOR2_X1 U7469 ( .A1(n14955), .A2(n14954), .ZN(n14953) );
  NOR2_X2 U7470 ( .A1(n12463), .A2(n14387), .ZN(n8323) );
  NOR2_X4 U7471 ( .A1(n12963), .A2(n16148), .ZN(n12962) );
  INV_X1 U7472 ( .A(n10854), .ZN(n7189) );
  INV_X1 U7473 ( .A(n7189), .ZN(n7190) );
  INV_X1 U7474 ( .A(n7189), .ZN(n7191) );
  NAND2_X1 U7475 ( .A1(n13464), .A2(n10425), .ZN(n7192) );
  INV_X1 U7476 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U7477 ( .A1(n7935), .A2(n10050), .ZN(n10053) );
  MUX2_X1 U7478 ( .A(n10049), .B(n10048), .S(n12281), .Z(n10050) );
  OAI211_X1 U7479 ( .C1(n10043), .C2(n10109), .A(n10047), .B(n7936), .ZN(n7935) );
  NAND2_X1 U7480 ( .A1(n7724), .A2(n13246), .ZN(n7723) );
  NAND2_X1 U7481 ( .A1(n7726), .A2(n8190), .ZN(n7724) );
  NOR2_X1 U7482 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n9067) );
  NOR2_X1 U7483 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n9065) );
  NOR2_X1 U7484 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n9066) );
  INV_X1 U7485 ( .A(n7646), .ZN(n7645) );
  OAI21_X1 U7486 ( .B1(n9165), .B2(n7647), .A(n9185), .ZN(n7646) );
  INV_X1 U7487 ( .A(n7824), .ZN(n7823) );
  OAI21_X1 U7488 ( .B1(n7825), .B2(n8092), .A(n7200), .ZN(n7824) );
  NAND2_X1 U7489 ( .A1(n8936), .A2(n8483), .ZN(n8962) );
  INV_X1 U7490 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7543) );
  INV_X1 U7491 ( .A(n8010), .ZN(n9087) );
  XNOR2_X1 U7492 ( .A(n9090), .B(n9089), .ZN(n9969) );
  OAI21_X1 U7493 ( .B1(n9630), .B2(P3_IR_REG_26__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9090) );
  XNOR2_X1 U7494 ( .A(n9631), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U7495 ( .A1(n7367), .A2(n8061), .ZN(n8060) );
  AND2_X1 U7496 ( .A1(n7303), .A2(n13433), .ZN(n8061) );
  NOR2_X1 U7497 ( .A1(n7817), .A2(n13051), .ZN(n7816) );
  INV_X1 U7498 ( .A(n13050), .ZN(n7817) );
  INV_X1 U7499 ( .A(n11054), .ZN(n10740) );
  NAND2_X1 U7500 ( .A1(n11054), .A2(n8421), .ZN(n10546) );
  NAND2_X1 U7501 ( .A1(n11054), .A2(n10986), .ZN(n10854) );
  NAND2_X2 U7502 ( .A1(n10950), .A2(n13455), .ZN(n11054) );
  NAND2_X1 U7503 ( .A1(n13074), .A2(n13073), .ZN(n13072) );
  AND2_X1 U7504 ( .A1(n8344), .A2(n8343), .ZN(n8342) );
  INV_X1 U7505 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8343) );
  INV_X1 U7506 ( .A(n8494), .ZN(n7506) );
  OR2_X1 U7507 ( .A1(n10044), .A2(n10188), .ZN(n7936) );
  NAND2_X1 U7508 ( .A1(n10053), .A2(n10054), .ZN(n10052) );
  NAND2_X1 U7509 ( .A1(n10063), .A2(n10062), .ZN(n7846) );
  NAND2_X1 U7510 ( .A1(n10067), .A2(n10066), .ZN(n7845) );
  OAI22_X1 U7511 ( .A1(n7944), .A2(n7254), .B1(n10079), .B2(n7946), .ZN(n10081) );
  NAND2_X1 U7512 ( .A1(n10077), .A2(n7945), .ZN(n7944) );
  NAND2_X1 U7513 ( .A1(n10079), .A2(n7946), .ZN(n7945) );
  OR2_X1 U7514 ( .A1(n13213), .A2(n7203), .ZN(n8184) );
  OAI22_X1 U7515 ( .A1(n7949), .A2(n7253), .B1(n10094), .B2(n7951), .ZN(n10096) );
  NAND2_X1 U7516 ( .A1(n10092), .A2(n7950), .ZN(n7949) );
  NAND2_X1 U7517 ( .A1(n10094), .A2(n7951), .ZN(n7950) );
  INV_X1 U7518 ( .A(n7722), .ZN(n7721) );
  OAI21_X1 U7519 ( .B1(n7723), .B2(n7726), .A(n7725), .ZN(n7722) );
  OAI21_X1 U7520 ( .B1(n7276), .B2(n7957), .A(n7956), .ZN(n10121) );
  OR2_X1 U7521 ( .A1(n7959), .A2(n10119), .ZN(n7956) );
  NAND2_X1 U7522 ( .A1(n10117), .A2(n7958), .ZN(n7957) );
  OR2_X1 U7523 ( .A1(n9735), .A2(n9734), .ZN(n9737) );
  OR2_X1 U7524 ( .A1(n9877), .A2(n9722), .ZN(n9740) );
  AND3_X1 U7525 ( .A1(n10165), .A2(n10235), .A3(n10164), .ZN(n10233) );
  INV_X1 U7526 ( .A(n8718), .ZN(n8331) );
  NOR2_X1 U7527 ( .A1(n8111), .A2(n10169), .ZN(n8110) );
  INV_X1 U7528 ( .A(n8113), .ZN(n8111) );
  NAND2_X1 U7529 ( .A1(n11226), .A2(n11225), .ZN(n11350) );
  AND3_X1 U7530 ( .A1(n7997), .A2(n9697), .A3(n9865), .ZN(n7996) );
  INV_X1 U7531 ( .A(n8005), .ZN(n7998) );
  NAND2_X1 U7532 ( .A1(n9862), .A2(n9694), .ZN(n9724) );
  NAND2_X1 U7533 ( .A1(n7627), .A2(n7625), .ZN(n9862) );
  NOR2_X1 U7534 ( .A1(n13593), .A2(n7626), .ZN(n7625) );
  INV_X1 U7535 ( .A(n9682), .ZN(n7626) );
  NAND2_X1 U7536 ( .A1(n15731), .A2(n7538), .ZN(n9949) );
  NAND2_X1 U7537 ( .A1(n15737), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7538) );
  OR2_X1 U7538 ( .A1(n9669), .A2(n13610), .ZN(n9861) );
  OR2_X1 U7539 ( .A1(n13123), .A2(n13470), .ZN(n9858) );
  NAND2_X1 U7540 ( .A1(n13123), .A2(n13470), .ZN(n9860) );
  NAND2_X1 U7541 ( .A1(n9875), .A2(n9558), .ZN(n8177) );
  OR2_X1 U7542 ( .A1(n13560), .A2(n13115), .ZN(n9732) );
  OR2_X1 U7543 ( .A1(n13522), .A2(n13504), .ZN(n9742) );
  OR2_X1 U7544 ( .A1(n13474), .A2(n13676), .ZN(n9748) );
  OR2_X1 U7545 ( .A1(n13539), .A2(n13496), .ZN(n9750) );
  AND2_X1 U7546 ( .A1(n12793), .A2(n7886), .ZN(n7885) );
  NAND2_X1 U7547 ( .A1(n12748), .A2(n9752), .ZN(n7886) );
  AOI21_X1 U7548 ( .B1(n7215), .B2(n7632), .A(n7347), .ZN(n7629) );
  INV_X1 U7549 ( .A(n9208), .ZN(n7687) );
  NAND2_X1 U7550 ( .A1(n7826), .A2(n13059), .ZN(n7825) );
  NAND2_X1 U7551 ( .A1(n8092), .A2(n8094), .ZN(n7826) );
  OR2_X1 U7552 ( .A1(n14285), .A2(n14090), .ZN(n13402) );
  OR2_X1 U7553 ( .A1(n12624), .A2(n13024), .ZN(n13354) );
  NAND2_X1 U7554 ( .A1(n8360), .A2(n7400), .ZN(n8358) );
  NOR2_X1 U7555 ( .A1(n13073), .A2(n7579), .ZN(n7578) );
  INV_X1 U7556 ( .A(n7581), .ZN(n7579) );
  INV_X1 U7557 ( .A(n14746), .ZN(n14531) );
  AND2_X1 U7558 ( .A1(n15099), .A2(n14750), .ZN(n8891) );
  AND2_X1 U7559 ( .A1(n8248), .A2(n15004), .ZN(n7684) );
  NOR2_X1 U7560 ( .A1(n8245), .A2(n8250), .ZN(n8248) );
  NAND2_X1 U7561 ( .A1(n8564), .A2(n15934), .ZN(n10035) );
  NAND2_X1 U7562 ( .A1(n8967), .A2(n8966), .ZN(n8971) );
  AND2_X1 U7563 ( .A1(n8813), .A2(n8486), .ZN(n7498) );
  AOI21_X1 U7564 ( .B1(n7553), .B2(n7552), .A(n7327), .ZN(n7551) );
  NAND2_X1 U7565 ( .A1(n8909), .A2(n8908), .ZN(n8911) );
  NAND2_X1 U7566 ( .A1(n8403), .A2(n8985), .ZN(n8402) );
  INV_X1 U7567 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8985) );
  INV_X1 U7568 ( .A(n8404), .ZN(n8403) );
  NAND2_X1 U7569 ( .A1(n8448), .A2(SI_13_), .ZN(n8449) );
  INV_X1 U7570 ( .A(n8737), .ZN(n8131) );
  AOI21_X1 U7571 ( .B1(n7806), .B2(n7808), .A(n7804), .ZN(n7803) );
  NAND2_X1 U7572 ( .A1(n8666), .A2(n7806), .ZN(n7805) );
  INV_X1 U7573 ( .A(n8442), .ZN(n7804) );
  OR2_X1 U7574 ( .A1(n8421), .A2(n10980), .ZN(n8142) );
  XNOR2_X1 U7575 ( .A(n10298), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n10342) );
  AND2_X1 U7576 ( .A1(n7604), .A2(n7287), .ZN(n10337) );
  NAND2_X1 U7577 ( .A1(n7605), .A2(n7913), .ZN(n7604) );
  INV_X1 U7578 ( .A(n10339), .ZN(n7605) );
  AOI21_X1 U7579 ( .B1(n12614), .B2(n12613), .A(n7305), .ZN(n12615) );
  NAND2_X1 U7580 ( .A1(n13088), .A2(n13734), .ZN(n8296) );
  INV_X1 U7581 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U7582 ( .A1(n11756), .A2(n7542), .ZN(n9943) );
  OR2_X1 U7583 ( .A1(n10005), .A2(n16073), .ZN(n7542) );
  XNOR2_X1 U7584 ( .A(n9949), .B(n15745), .ZN(n15747) );
  NAND2_X1 U7585 ( .A1(n15747), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n15746) );
  OR2_X1 U7586 ( .A1(n15764), .A2(n15763), .ZN(n15761) );
  AOI21_X1 U7587 ( .B1(n7741), .B2(n7740), .A(n7328), .ZN(n7739) );
  INV_X1 U7588 ( .A(n15729), .ZN(n7740) );
  OR2_X1 U7589 ( .A1(n15730), .A2(n7742), .ZN(n7738) );
  NOR2_X1 U7590 ( .A1(n8177), .A2(n13608), .ZN(n13609) );
  NAND2_X1 U7591 ( .A1(n7872), .A2(n9748), .ZN(n13650) );
  NAND2_X1 U7592 ( .A1(n13662), .A2(n13663), .ZN(n7872) );
  AOI21_X1 U7593 ( .B1(n7904), .B2(n7906), .A(n7903), .ZN(n7902) );
  NAND2_X1 U7594 ( .A1(n7987), .A2(n13750), .ZN(n7986) );
  NAND2_X1 U7595 ( .A1(n7988), .A2(n9719), .ZN(n7987) );
  OR2_X1 U7596 ( .A1(n11236), .A2(n11657), .ZN(n15960) );
  BUF_X1 U7597 ( .A(n9262), .Z(n9691) );
  INV_X1 U7598 ( .A(n9148), .ZN(n9690) );
  AND2_X1 U7599 ( .A1(n9637), .A2(n9648), .ZN(n9649) );
  AND2_X1 U7600 ( .A1(n9077), .A2(n9076), .ZN(n9080) );
  MUX2_X1 U7601 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9075), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n9077) );
  NAND2_X1 U7602 ( .A1(n9567), .A2(n9566), .ZN(n9580) );
  AND2_X1 U7603 ( .A1(n7436), .A2(n9071), .ZN(n7435) );
  AND2_X1 U7604 ( .A1(n8169), .A2(n9072), .ZN(n7436) );
  INV_X1 U7605 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9072) );
  AND2_X1 U7606 ( .A1(n9071), .A2(n8169), .ZN(n8168) );
  NAND2_X1 U7607 ( .A1(n9467), .A2(n9466), .ZN(n9471) );
  INV_X1 U7608 ( .A(n8023), .ZN(n8022) );
  OAI21_X1 U7609 ( .B1(n9345), .B2(n8024), .A(n9364), .ZN(n8023) );
  OR2_X1 U7610 ( .A1(n9309), .A2(n9308), .ZN(n9310) );
  AOI21_X1 U7611 ( .B1(n7651), .B2(n7649), .A(n7648), .ZN(n9327) );
  AND2_X1 U7612 ( .A1(n9279), .A2(n7650), .ZN(n7649) );
  NOR2_X1 U7613 ( .A1(n7652), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7648) );
  NOR2_X1 U7614 ( .A1(n7654), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7650) );
  AND2_X1 U7615 ( .A1(n9238), .A2(n9224), .ZN(n9225) );
  AND2_X1 U7616 ( .A1(n9187), .A2(n9168), .ZN(n9185) );
  OR2_X1 U7617 ( .A1(n14267), .A2(n13889), .ZN(n14045) );
  NAND3_X1 U7618 ( .A1(n7401), .A2(n10566), .A3(n8200), .ZN(n11599) );
  AND2_X1 U7619 ( .A1(n10565), .A2(n10562), .ZN(n8200) );
  AOI21_X1 U7620 ( .B1(n13904), .B2(n13903), .A(n7429), .ZN(n13960) );
  AND2_X1 U7621 ( .A1(n10755), .A2(n10756), .ZN(n7429) );
  NOR2_X1 U7622 ( .A1(n11695), .A2(n15408), .ZN(n10954) );
  INV_X1 U7623 ( .A(n10943), .ZN(n10879) );
  NAND2_X1 U7624 ( .A1(n7810), .A2(n7235), .ZN(n14147) );
  AOI21_X1 U7625 ( .B1(n7816), .B2(n13048), .A(n7259), .ZN(n7815) );
  AND2_X1 U7626 ( .A1(n7371), .A2(n8044), .ZN(n14226) );
  NAND2_X1 U7627 ( .A1(n12898), .A2(n7370), .ZN(n7371) );
  AND2_X1 U7628 ( .A1(n12527), .A2(n12529), .ZN(n8064) );
  INV_X1 U7629 ( .A(n13417), .ZN(n12529) );
  AND2_X1 U7630 ( .A1(n11465), .A2(n10950), .ZN(n14091) );
  NAND2_X1 U7631 ( .A1(n10446), .A2(n10445), .ZN(n10440) );
  INV_X1 U7632 ( .A(n14744), .ZN(n14587) );
  AND2_X1 U7633 ( .A1(n14584), .A2(n8382), .ZN(n8381) );
  NAND2_X1 U7634 ( .A1(n8383), .A2(n14723), .ZN(n8382) );
  INV_X1 U7635 ( .A(n14720), .ZN(n8383) );
  NOR2_X1 U7636 ( .A1(n14684), .A2(n8387), .ZN(n8386) );
  INV_X1 U7637 ( .A(n14489), .ZN(n8387) );
  AOI21_X1 U7638 ( .B1(n8365), .B2(n8368), .A(n8364), .ZN(n8363) );
  INV_X1 U7639 ( .A(n14465), .ZN(n8364) );
  NAND2_X1 U7640 ( .A1(n7384), .A2(n7383), .ZN(n7382) );
  NAND2_X1 U7641 ( .A1(n14412), .A2(n14413), .ZN(n7383) );
  NAND2_X1 U7642 ( .A1(n15036), .A2(n14383), .ZN(n8316) );
  XNOR2_X1 U7643 ( .A(n15063), .B(n14747), .ZN(n14916) );
  NOR2_X1 U7644 ( .A1(n14945), .A2(n14932), .ZN(n8272) );
  AOI21_X1 U7645 ( .B1(n14961), .B2(n14963), .A(n8408), .ZN(n14955) );
  OR2_X1 U7646 ( .A1(n15099), .A2(n9015), .ZN(n9016) );
  OAI21_X1 U7647 ( .B1(n12857), .B2(n7521), .A(n7207), .ZN(n15007) );
  NAND2_X1 U7648 ( .A1(n7520), .A2(n7519), .ZN(n7518) );
  AND2_X1 U7649 ( .A1(n8256), .A2(n9013), .ZN(n7598) );
  NAND2_X1 U7650 ( .A1(n8563), .A2(n10986), .ZN(n7529) );
  NAND2_X1 U7651 ( .A1(n15927), .A2(n15881), .ZN(n16139) );
  AND2_X1 U7652 ( .A1(n11845), .A2(n9055), .ZN(n11557) );
  AND2_X1 U7653 ( .A1(n11844), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9055) );
  AND2_X1 U7654 ( .A1(n8511), .A2(n7575), .ZN(n8518) );
  MUX2_X1 U7655 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8510), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8511) );
  NOR2_X1 U7656 ( .A1(n7504), .A2(n7503), .ZN(n8499) );
  INV_X1 U7657 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8496) );
  NOR2_X1 U7658 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8497) );
  NAND2_X1 U7659 ( .A1(n8126), .A2(n8124), .ZN(n8755) );
  NOR2_X1 U7660 ( .A1(n8125), .A2(n8752), .ZN(n8124) );
  INV_X1 U7661 ( .A(n8128), .ZN(n8125) );
  INV_X1 U7662 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U7663 ( .A1(n15603), .A2(n7615), .ZN(n7614) );
  OR2_X1 U7664 ( .A1(n15603), .A2(n7615), .ZN(n7613) );
  NOR2_X1 U7665 ( .A1(n15711), .A2(n15712), .ZN(n15710) );
  OR2_X1 U7666 ( .A1(n15728), .A2(n15727), .ZN(n7969) );
  NAND2_X1 U7667 ( .A1(n10874), .A2(n10873), .ZN(n14271) );
  AOI21_X1 U7668 ( .B1(n11868), .B2(n10621), .A(n11867), .ZN(n11980) );
  AND2_X1 U7669 ( .A1(n12550), .A2(n10645), .ZN(n8234) );
  NAND2_X1 U7670 ( .A1(n8235), .A2(n12145), .ZN(n8233) );
  NAND2_X1 U7671 ( .A1(n10628), .A2(n8235), .ZN(n7426) );
  NAND2_X1 U7672 ( .A1(n10457), .A2(n10456), .ZN(n13237) );
  NAND2_X1 U7673 ( .A1(n7366), .A2(n14042), .ZN(n7365) );
  NAND2_X1 U7674 ( .A1(n7367), .A2(n7303), .ZN(n7366) );
  XNOR2_X1 U7675 ( .A(n12665), .B(n15535), .ZN(n15531) );
  AND2_X1 U7676 ( .A1(n8394), .A2(n7293), .ZN(n7862) );
  NAND2_X1 U7677 ( .A1(n13072), .A2(n7236), .ZN(n15041) );
  NAND2_X1 U7678 ( .A1(n15578), .A2(n15577), .ZN(n15576) );
  OAI21_X1 U7679 ( .B1(n13135), .B2(n13136), .A(n13134), .ZN(n13141) );
  OR2_X1 U7680 ( .A1(n10059), .A2(n10061), .ZN(n7965) );
  AOI22_X1 U7681 ( .A1(n14027), .A2(n13393), .B1(n13365), .B2(n14248), .ZN(
        n13161) );
  NAND2_X1 U7682 ( .A1(n10069), .A2(n7941), .ZN(n7940) );
  NAND2_X1 U7683 ( .A1(n7273), .A2(n13179), .ZN(n7704) );
  NOR2_X1 U7684 ( .A1(n7273), .A2(n13179), .ZN(n8178) );
  NAND2_X1 U7685 ( .A1(n7842), .A2(n10080), .ZN(n7841) );
  NAND2_X1 U7686 ( .A1(n10081), .A2(n10082), .ZN(n7842) );
  OR2_X1 U7687 ( .A1(n10081), .A2(n10082), .ZN(n7840) );
  NAND2_X1 U7688 ( .A1(n10084), .A2(n7948), .ZN(n7947) );
  AND2_X1 U7689 ( .A1(n8182), .A2(n8180), .ZN(n13219) );
  INV_X1 U7690 ( .A(n8183), .ZN(n8181) );
  NAND2_X1 U7691 ( .A1(n13213), .A2(n7203), .ZN(n8183) );
  NAND2_X1 U7692 ( .A1(n7837), .A2(n10095), .ZN(n7836) );
  NAND2_X1 U7693 ( .A1(n10096), .A2(n10097), .ZN(n7837) );
  OR2_X1 U7694 ( .A1(n10096), .A2(n10097), .ZN(n7835) );
  NAND2_X1 U7695 ( .A1(n10099), .A2(n7943), .ZN(n7942) );
  AOI21_X1 U7696 ( .B1(n7721), .B2(n7723), .A(n7715), .ZN(n7714) );
  NAND2_X1 U7697 ( .A1(n7256), .A2(n7716), .ZN(n7715) );
  NAND2_X1 U7698 ( .A1(n7726), .A2(n7717), .ZN(n7716) );
  NOR2_X1 U7699 ( .A1(n7721), .A2(n7720), .ZN(n7719) );
  NOR2_X1 U7700 ( .A1(n13246), .A2(n7727), .ZN(n7720) );
  NAND2_X1 U7701 ( .A1(n10111), .A2(n7953), .ZN(n7952) );
  AOI21_X1 U7702 ( .B1(n7201), .B2(n7736), .A(n7279), .ZN(n7733) );
  AND2_X1 U7703 ( .A1(n13257), .A2(n13258), .ZN(n7736) );
  NAND2_X1 U7704 ( .A1(n7707), .A2(n7706), .ZN(n7705) );
  INV_X1 U7705 ( .A(n13276), .ZN(n8188) );
  NAND2_X1 U7706 ( .A1(n7832), .A2(n10120), .ZN(n7831) );
  NAND2_X1 U7707 ( .A1(n10121), .A2(n10122), .ZN(n7832) );
  OR2_X1 U7708 ( .A1(n10121), .A2(n10122), .ZN(n7830) );
  NAND2_X1 U7709 ( .A1(n10124), .A2(n7939), .ZN(n7938) );
  NAND2_X1 U7710 ( .A1(n8196), .A2(n8197), .ZN(n13295) );
  NAND2_X1 U7711 ( .A1(n13290), .A2(n7310), .ZN(n8197) );
  INV_X1 U7712 ( .A(n9466), .ZN(n7631) );
  NAND2_X1 U7713 ( .A1(n7861), .A2(n10041), .ZN(n7857) );
  INV_X1 U7714 ( .A(n7859), .ZN(n7856) );
  INV_X1 U7715 ( .A(n9740), .ZN(n9743) );
  NOR2_X1 U7716 ( .A1(n8003), .A2(n9698), .ZN(n8000) );
  NAND2_X1 U7717 ( .A1(n13342), .A2(n13339), .ZN(n13385) );
  NAND2_X1 U7718 ( .A1(n7850), .A2(n7849), .ZN(n10139) );
  NAND2_X1 U7719 ( .A1(n10134), .A2(n10136), .ZN(n7849) );
  AOI21_X1 U7720 ( .B1(n8771), .B2(n8452), .A(n8147), .ZN(n8146) );
  INV_X1 U7721 ( .A(n8790), .ZN(n8147) );
  INV_X1 U7722 ( .A(n8452), .ZN(n8144) );
  NOR2_X1 U7723 ( .A1(n10299), .A2(n7914), .ZN(n10301) );
  AND2_X1 U7724 ( .A1(n10300), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7914) );
  AND2_X1 U7725 ( .A1(n13556), .A2(n8286), .ZN(n8285) );
  OR2_X1 U7726 ( .A1(n13502), .A2(n8287), .ZN(n8286) );
  INV_X1 U7727 ( .A(n13114), .ZN(n8287) );
  NOR2_X1 U7728 ( .A1(n13529), .A2(n8312), .ZN(n8311) );
  INV_X1 U7729 ( .A(n13092), .ZN(n8312) );
  INV_X1 U7730 ( .A(n13492), .ZN(n8310) );
  INV_X1 U7731 ( .A(n8000), .ZN(n7999) );
  CLKBUF_X1 U7732 ( .A(n9084), .Z(n9930) );
  AOI21_X1 U7733 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10999), .A(n15638), .ZN(
        n9899) );
  OR2_X1 U7734 ( .A1(n9902), .A2(n11620), .ZN(n7973) );
  NAND2_X1 U7735 ( .A1(n15765), .A2(n7345), .ZN(n9953) );
  AND2_X1 U7736 ( .A1(n7751), .A2(n7750), .ZN(n10030) );
  NAND2_X1 U7737 ( .A1(n10029), .A2(n15821), .ZN(n7750) );
  NAND2_X1 U7738 ( .A1(n15802), .A2(n7540), .ZN(n9957) );
  OR2_X1 U7739 ( .A1(n15798), .A2(n9955), .ZN(n7540) );
  INV_X1 U7740 ( .A(n13608), .ZN(n9623) );
  INV_X1 U7741 ( .A(n9578), .ZN(n7442) );
  AND2_X1 U7742 ( .A1(n13123), .A2(n9881), .ZN(n9578) );
  AND2_X1 U7743 ( .A1(n7196), .A2(n7454), .ZN(n7453) );
  NAND2_X1 U7744 ( .A1(n7457), .A2(n9498), .ZN(n7454) );
  INV_X1 U7745 ( .A(n9498), .ZN(n7455) );
  INV_X1 U7746 ( .A(n13639), .ZN(n13635) );
  NOR2_X1 U7747 ( .A1(n13096), .A2(n8162), .ZN(n8161) );
  INV_X1 U7748 ( .A(n9452), .ZN(n8162) );
  NOR2_X1 U7749 ( .A1(n9840), .A2(n7908), .ZN(n7907) );
  NOR2_X1 U7750 ( .A1(n13704), .A2(n8164), .ZN(n8163) );
  INV_X1 U7751 ( .A(n9437), .ZN(n8164) );
  NOR2_X1 U7752 ( .A1(n8155), .A2(n7452), .ZN(n7451) );
  INV_X1 U7753 ( .A(n13012), .ZN(n7452) );
  INV_X1 U7754 ( .A(n8156), .ZN(n8155) );
  INV_X1 U7755 ( .A(n7451), .ZN(n7450) );
  NOR2_X1 U7756 ( .A1(n13750), .A2(n8157), .ZN(n8156) );
  INV_X1 U7757 ( .A(n9380), .ZN(n8157) );
  INV_X1 U7758 ( .A(n9760), .ZN(n7876) );
  NAND2_X1 U7759 ( .A1(n9756), .A2(n9608), .ZN(n9758) );
  NOR2_X1 U7760 ( .A1(n7660), .A2(n12626), .ZN(n7659) );
  OR2_X1 U7761 ( .A1(n9515), .A2(n7660), .ZN(n7657) );
  INV_X1 U7762 ( .A(n9399), .ZN(n8027) );
  AND2_X1 U7763 ( .A1(n9367), .A2(n9387), .ZN(n8315) );
  INV_X1 U7764 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9063) );
  NOR2_X1 U7765 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n9060) );
  NOR2_X1 U7766 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7865) );
  AND2_X1 U7767 ( .A1(n9062), .A2(n9061), .ZN(n7866) );
  INV_X1 U7768 ( .A(n9167), .ZN(n7647) );
  OR2_X1 U7769 ( .A1(n13886), .A2(n8242), .ZN(n8241) );
  INV_X1 U7770 ( .A(n10872), .ZN(n8242) );
  NAND2_X1 U7771 ( .A1(n14027), .A2(n10938), .ZN(n10560) );
  INV_X1 U7772 ( .A(n10852), .ZN(n8243) );
  NAND2_X1 U7773 ( .A1(n13399), .A2(n13024), .ZN(n13356) );
  NOR2_X1 U7774 ( .A1(n7825), .A2(n7822), .ZN(n7821) );
  INV_X1 U7775 ( .A(n13054), .ZN(n7822) );
  OR2_X1 U7776 ( .A1(n14087), .A2(n8091), .ZN(n8090) );
  INV_X1 U7777 ( .A(n13060), .ZN(n8091) );
  INV_X1 U7778 ( .A(n8093), .ZN(n8092) );
  OAI21_X1 U7779 ( .B1(n8095), .B2(n8094), .A(n13058), .ZN(n8093) );
  NAND2_X1 U7780 ( .A1(n14128), .A2(n13054), .ZN(n13056) );
  NOR2_X1 U7781 ( .A1(n8054), .A2(n7358), .ZN(n7357) );
  INV_X1 U7782 ( .A(n13032), .ZN(n7358) );
  OR3_X1 U7783 ( .A1(n10810), .A2(n10809), .A3(n10808), .ZN(n10825) );
  NOR2_X1 U7784 ( .A1(n13035), .A2(n8057), .ZN(n8056) );
  INV_X1 U7785 ( .A(n13033), .ZN(n8057) );
  NOR2_X1 U7786 ( .A1(n13249), .A2(n14342), .ZN(n7763) );
  AOI21_X1 U7787 ( .B1(n12536), .B2(n8074), .A(n8072), .ZN(n8071) );
  INV_X1 U7788 ( .A(n12699), .ZN(n8072) );
  NAND2_X1 U7789 ( .A1(n7492), .A2(n14019), .ZN(n8078) );
  INV_X1 U7790 ( .A(n11698), .ZN(n13136) );
  AND2_X1 U7791 ( .A1(n13399), .A2(n13445), .ZN(n11698) );
  NOR2_X1 U7792 ( .A1(n15896), .A2(n13442), .ZN(n10941) );
  NAND2_X1 U7793 ( .A1(n10437), .A2(n8411), .ZN(n10436) );
  INV_X1 U7794 ( .A(n14633), .ZN(n8373) );
  AND2_X1 U7795 ( .A1(n7399), .A2(n8365), .ZN(n7396) );
  NAND2_X1 U7796 ( .A1(n7249), .A2(n7199), .ZN(n7581) );
  NAND2_X1 U7797 ( .A1(n7199), .A2(n7583), .ZN(n7582) );
  INV_X1 U7798 ( .A(n8279), .ZN(n7583) );
  INV_X1 U7799 ( .A(n14913), .ZN(n14516) );
  NOR2_X1 U7800 ( .A1(n15077), .A2(n14748), .ZN(n7667) );
  NOR2_X1 U7801 ( .A1(n14932), .A2(n8274), .ZN(n8271) );
  NOR2_X1 U7802 ( .A1(n14738), .A2(n7773), .ZN(n7771) );
  INV_X1 U7803 ( .A(n12263), .ZN(n7779) );
  INV_X1 U7804 ( .A(n7587), .ZN(n7586) );
  OAI21_X1 U7805 ( .B1(n11803), .B2(n7588), .A(n9002), .ZN(n7587) );
  INV_X1 U7806 ( .A(n9001), .ZN(n7588) );
  INV_X1 U7807 ( .A(n8995), .ZN(n7563) );
  NAND2_X1 U7808 ( .A1(n10206), .A2(n8993), .ZN(n10037) );
  NAND2_X1 U7809 ( .A1(n15917), .A2(n8555), .ZN(n8993) );
  NAND2_X1 U7810 ( .A1(n15924), .A2(n15914), .ZN(n15912) );
  INV_X1 U7811 ( .A(n15073), .ZN(n14939) );
  AOI21_X1 U7812 ( .B1(n8110), .B2(n8115), .A(n7216), .ZN(n8108) );
  NOR2_X1 U7813 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n8492) );
  INV_X1 U7814 ( .A(n8478), .ZN(n8140) );
  INV_X1 U7815 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8490) );
  INV_X1 U7816 ( .A(SI_22_), .ZN(n15295) );
  NAND2_X1 U7817 ( .A1(n8895), .A2(n8469), .ZN(n8530) );
  AOI21_X1 U7818 ( .B1(n8119), .B2(n8122), .A(n7325), .ZN(n8117) );
  AOI21_X1 U7819 ( .B1(n8462), .B2(n8463), .A(n7324), .ZN(n8123) );
  INV_X1 U7820 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U7821 ( .A1(n7493), .A2(SI_5_), .ZN(n8428) );
  NAND2_X1 U7822 ( .A1(n7828), .A2(SI_4_), .ZN(n8426) );
  NAND2_X1 U7823 ( .A1(n7546), .A2(SI_3_), .ZN(n8425) );
  AND2_X1 U7824 ( .A1(n8141), .A2(n7377), .ZN(n7375) );
  XNOR2_X1 U7825 ( .A(n10301), .B(n10302), .ZN(n10339) );
  OAI22_X1 U7826 ( .A1(n10320), .A2(n10371), .B1(P3_ADDR_REG_11__SCAN_IN), 
        .B2(n10319), .ZN(n10374) );
  INV_X1 U7827 ( .A(n11350), .ZN(n12498) );
  AOI21_X1 U7828 ( .B1(n13537), .B2(n13496), .A(n13104), .ZN(n13107) );
  AND2_X1 U7829 ( .A1(n12780), .A2(n12781), .ZN(n12778) );
  NAND2_X1 U7830 ( .A1(n15374), .A2(n9475), .ZN(n9492) );
  NAND2_X1 U7831 ( .A1(n11227), .A2(n11228), .ZN(n11347) );
  INV_X1 U7832 ( .A(n8296), .ZN(n8293) );
  NAND2_X1 U7833 ( .A1(n8295), .A2(n8294), .ZN(n13510) );
  INV_X1 U7834 ( .A(n13512), .ZN(n8295) );
  NAND2_X1 U7835 ( .A1(n12814), .A2(n12813), .ZN(n12888) );
  NAND2_X1 U7836 ( .A1(n9860), .A2(n9926), .ZN(n8039) );
  NOR2_X1 U7837 ( .A1(n9724), .A2(n9696), .ZN(n9865) );
  NOR2_X1 U7838 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9084) );
  NAND2_X1 U7839 ( .A1(n11371), .A2(n7240), .ZN(n9897) );
  NAND2_X1 U7840 ( .A1(n15663), .A2(n15662), .ZN(n15661) );
  NOR2_X1 U7841 ( .A1(n7974), .A2(n9903), .ZN(n11763) );
  NOR2_X1 U7842 ( .A1(n11614), .A2(n11908), .ZN(n7974) );
  OR2_X1 U7843 ( .A1(n11763), .A2(n11762), .ZN(n7470) );
  AND2_X1 U7844 ( .A1(n12059), .A2(n10010), .ZN(n15704) );
  NAND2_X1 U7845 ( .A1(n15704), .A2(n15703), .ZN(n15702) );
  NAND2_X1 U7846 ( .A1(n15730), .A2(n15729), .ZN(n7743) );
  NAND2_X1 U7847 ( .A1(n7743), .A2(n7741), .ZN(n15748) );
  NAND2_X1 U7848 ( .A1(n7969), .A2(n7968), .ZN(n7468) );
  NAND2_X1 U7849 ( .A1(n15737), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7968) );
  AND2_X1 U7850 ( .A1(n7738), .A2(n7331), .ZN(n15774) );
  INV_X1 U7851 ( .A(n15775), .ZN(n7737) );
  NAND2_X1 U7852 ( .A1(n15746), .A2(n9950), .ZN(n15766) );
  NAND2_X1 U7853 ( .A1(n15761), .A2(n9917), .ZN(n7975) );
  XNOR2_X1 U7854 ( .A(n10025), .B(n10024), .ZN(n15792) );
  NOR2_X1 U7855 ( .A1(n15792), .A2(n15791), .ZN(n15790) );
  XNOR2_X1 U7856 ( .A(n9953), .B(n10024), .ZN(n15786) );
  NAND2_X1 U7857 ( .A1(n15786), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n15785) );
  NAND2_X1 U7858 ( .A1(n15801), .A2(n15800), .ZN(n15799) );
  INV_X1 U7859 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9367) );
  AND2_X1 U7860 ( .A1(n9590), .A2(n9348), .ZN(n9368) );
  OR2_X1 U7861 ( .A1(n15824), .A2(n15825), .ZN(n7751) );
  XNOR2_X1 U7862 ( .A(n9957), .B(n9956), .ZN(n15818) );
  NAND2_X1 U7863 ( .A1(n15818), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n15817) );
  XNOR2_X1 U7864 ( .A(n10030), .B(n15833), .ZN(n15838) );
  NOR2_X1 U7865 ( .A1(n9623), .A2(n9877), .ZN(n8005) );
  OAI21_X1 U7866 ( .B1(n9623), .B2(n8004), .A(n9858), .ZN(n8003) );
  AND2_X2 U7867 ( .A1(n9858), .A2(n9860), .ZN(n13608) );
  INV_X1 U7868 ( .A(n13628), .ZN(n7881) );
  INV_X1 U7869 ( .A(n7880), .ZN(n7879) );
  OAI21_X1 U7870 ( .B1(n7881), .B2(n9621), .A(n9732), .ZN(n7880) );
  AND2_X1 U7871 ( .A1(n13651), .A2(n9513), .ZN(n13640) );
  AND2_X1 U7872 ( .A1(n9742), .A2(n9739), .ZN(n13654) );
  AND4_X1 U7873 ( .A1(n9528), .A2(n9527), .A3(n9526), .A4(n9525), .ZN(n13656)
         );
  NAND2_X1 U7874 ( .A1(n13664), .A2(n9498), .ZN(n13653) );
  OR2_X1 U7875 ( .A1(n13653), .A2(n13654), .ZN(n13651) );
  NAND2_X1 U7876 ( .A1(n7873), .A2(n7991), .ZN(n13662) );
  NOR2_X1 U7877 ( .A1(n7243), .A2(n7993), .ZN(n7991) );
  NAND2_X1 U7878 ( .A1(n13684), .A2(n7261), .ZN(n7873) );
  OR2_X1 U7879 ( .A1(n13697), .A2(n13675), .ZN(n13097) );
  AND2_X1 U7880 ( .A1(n9750), .A2(n9751), .ZN(n13678) );
  NAND2_X1 U7881 ( .A1(n13684), .A2(n13689), .ZN(n13686) );
  AND2_X1 U7882 ( .A1(n13097), .A2(n13099), .ZN(n13689) );
  AOI21_X1 U7883 ( .B1(n13730), .B2(n7907), .A(n7905), .ZN(n7904) );
  INV_X1 U7884 ( .A(n7907), .ZN(n7906) );
  NAND2_X1 U7885 ( .A1(n13738), .A2(n13737), .ZN(n13736) );
  AOI21_X1 U7886 ( .B1(n13017), .B2(n7990), .A(n7989), .ZN(n7988) );
  INV_X1 U7887 ( .A(n9817), .ZN(n7990) );
  INV_X1 U7888 ( .A(n9821), .ZN(n7989) );
  AND4_X1 U7889 ( .A1(n9414), .A2(n9413), .A3(n9412), .A4(n9411), .ZN(n13745)
         );
  AND2_X1 U7890 ( .A1(n9826), .A2(n9833), .ZN(n13750) );
  NAND2_X1 U7891 ( .A1(n9379), .A2(n9719), .ZN(n13014) );
  NAND2_X1 U7892 ( .A1(n12970), .A2(n13012), .ZN(n9379) );
  AOI21_X1 U7893 ( .B1(n7885), .B2(n7887), .A(n7884), .ZN(n7883) );
  OAI21_X1 U7894 ( .B1(n12747), .B2(n7887), .A(n7885), .ZN(n12974) );
  NAND2_X1 U7895 ( .A1(n12749), .A2(n12748), .ZN(n9326) );
  NAND2_X1 U7896 ( .A1(n12747), .A2(n12746), .ZN(n12745) );
  AOI21_X1 U7897 ( .B1(n7891), .B2(n7893), .A(n7890), .ZN(n7889) );
  INV_X1 U7898 ( .A(n12449), .ZN(n7890) );
  AND2_X1 U7899 ( .A1(n9802), .A2(n9803), .ZN(n12449) );
  NAND2_X1 U7900 ( .A1(n7432), .A2(n9269), .ZN(n12445) );
  NAND2_X1 U7901 ( .A1(n7433), .A2(n8165), .ZN(n7432) );
  AOI21_X1 U7902 ( .B1(n7227), .B2(n9249), .A(n8166), .ZN(n8165) );
  INV_X1 U7903 ( .A(n12229), .ZN(n7896) );
  AND4_X1 U7904 ( .A1(n9255), .A2(n9254), .A3(n9253), .A4(n9252), .ZN(n12497)
         );
  NOR2_X1 U7905 ( .A1(n12212), .A2(n8152), .ZN(n8151) );
  INV_X1 U7906 ( .A(n9213), .ZN(n8152) );
  NAND2_X1 U7907 ( .A1(n11904), .A2(n11903), .ZN(n11902) );
  AND4_X1 U7908 ( .A1(n9183), .A2(n9182), .A3(n9181), .A4(n9180), .ZN(n12025)
         );
  AND2_X1 U7909 ( .A1(n9176), .A2(n9156), .ZN(n8150) );
  NAND2_X1 U7910 ( .A1(n9610), .A2(n9769), .ZN(n11880) );
  AND2_X1 U7911 ( .A1(n9776), .A2(n9775), .ZN(n11884) );
  NAND2_X1 U7912 ( .A1(n11960), .A2(n9137), .ZN(n11894) );
  NAND2_X1 U7913 ( .A1(n11894), .A2(n11893), .ZN(n11892) );
  AND2_X1 U7914 ( .A1(n15904), .A2(n9758), .ZN(n15955) );
  NAND2_X1 U7915 ( .A1(n15955), .A2(n15957), .ZN(n15954) );
  OAI211_X1 U7916 ( .C1(n11663), .C2(n11662), .A(n11661), .B(n11660), .ZN(
        n11667) );
  INV_X1 U7917 ( .A(n12000), .ZN(n9755) );
  NAND2_X1 U7918 ( .A1(n9693), .A2(n9692), .ZN(n13596) );
  NAND2_X1 U7919 ( .A1(n9551), .A2(n9550), .ZN(n13117) );
  NAND2_X1 U7920 ( .A1(n9536), .A2(n9535), .ZN(n13560) );
  NOR2_X1 U7921 ( .A1(n9148), .A2(n8032), .ZN(n8031) );
  OR2_X1 U7922 ( .A1(n12564), .A2(n9148), .ZN(n9522) );
  NAND2_X1 U7923 ( .A1(n9505), .A2(n9504), .ZN(n13522) );
  NAND2_X1 U7924 ( .A1(n9490), .A2(n9489), .ZN(n13474) );
  NAND2_X1 U7925 ( .A1(n9446), .A2(n9445), .ZN(n13532) );
  OR2_X1 U7926 ( .A1(n11733), .A2(n9148), .ZN(n9446) );
  NAND2_X1 U7927 ( .A1(n9391), .A2(n9390), .ZN(n13807) );
  NAND2_X1 U7928 ( .A1(n9580), .A2(n9579), .ZN(n9677) );
  NAND2_X1 U7929 ( .A1(n7434), .A2(n8008), .ZN(n8010) );
  AND2_X1 U7930 ( .A1(n9073), .A2(n9089), .ZN(n8008) );
  INV_X1 U7931 ( .A(n9630), .ZN(n7434) );
  NAND2_X1 U7932 ( .A1(n9563), .A2(n9562), .ZN(n9567) );
  NAND2_X1 U7933 ( .A1(n9515), .A2(n7661), .ZN(n9519) );
  NAND2_X1 U7934 ( .A1(n9519), .A2(n9518), .ZN(n9530) );
  OR2_X1 U7935 ( .A1(n9502), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9515) );
  INV_X1 U7936 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9068) );
  NAND2_X1 U7937 ( .A1(n9471), .A2(n9470), .ZN(n9488) );
  NAND2_X1 U7938 ( .A1(n9594), .A2(n9592), .ZN(n9644) );
  AOI21_X1 U7939 ( .B1(n9453), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n8014), .ZN(
        n8012) );
  INV_X1 U7940 ( .A(n9456), .ZN(n8014) );
  NAND2_X1 U7941 ( .A1(n9590), .A2(n9589), .ZN(n9595) );
  INV_X1 U7942 ( .A(n9588), .ZN(n9589) );
  INV_X1 U7943 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9596) );
  OR2_X1 U7944 ( .A1(n9441), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U7945 ( .A1(n9368), .A2(n8313), .ZN(n9422) );
  AND2_X1 U7946 ( .A1(n8315), .A2(n8314), .ZN(n8313) );
  INV_X1 U7947 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8314) );
  AOI21_X1 U7948 ( .B1(n8022), .B2(n8024), .A(n8021), .ZN(n8020) );
  INV_X1 U7949 ( .A(n9381), .ZN(n8021) );
  AND2_X1 U7950 ( .A1(n9399), .A2(n9383), .ZN(n9384) );
  AND2_X1 U7951 ( .A1(n9381), .A2(n9363), .ZN(n9364) );
  INV_X1 U7952 ( .A(n9361), .ZN(n8024) );
  AND2_X1 U7953 ( .A1(n9361), .A2(n9344), .ZN(n9345) );
  NAND2_X1 U7954 ( .A1(n9346), .A2(n9345), .ZN(n9362) );
  INV_X1 U7955 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9348) );
  AND2_X1 U7956 ( .A1(n9327), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8037) );
  NOR2_X1 U7957 ( .A1(n9302), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n9590) );
  AOI21_X1 U7958 ( .B1(n9279), .B2(n8018), .A(n8017), .ZN(n8016) );
  INV_X1 U7959 ( .A(n9294), .ZN(n8017) );
  INV_X1 U7960 ( .A(n9276), .ZN(n8018) );
  NAND2_X1 U7961 ( .A1(n7651), .A2(n9279), .ZN(n7655) );
  AND3_X1 U7962 ( .A1(n9108), .A2(n7198), .A3(n7866), .ZN(n9064) );
  XNOR2_X1 U7963 ( .A(n9221), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10005) );
  INV_X1 U7964 ( .A(n7622), .ZN(n7621) );
  OAI21_X1 U7965 ( .B1(n7687), .B2(n7623), .A(n9225), .ZN(n7622) );
  NAND2_X1 U7966 ( .A1(n7624), .A2(n7687), .ZN(n9223) );
  INV_X1 U7967 ( .A(n9209), .ZN(n7624) );
  NAND2_X1 U7968 ( .A1(n9152), .A2(n9151), .ZN(n9166) );
  AND2_X1 U7969 ( .A1(n9167), .A2(n9153), .ZN(n9165) );
  NAND2_X1 U7970 ( .A1(n14026), .A2(n10938), .ZN(n10563) );
  INV_X1 U7971 ( .A(n8208), .ZN(n8202) );
  NAND2_X1 U7972 ( .A1(n8208), .A2(n8209), .ZN(n8204) );
  INV_X1 U7973 ( .A(n14054), .ZN(n13889) );
  NAND2_X1 U7974 ( .A1(n10819), .A2(n10821), .ZN(n10822) );
  XNOR2_X1 U7975 ( .A(n13210), .B(n10835), .ZN(n10624) );
  NAND2_X1 U7976 ( .A1(n8214), .A2(n10772), .ZN(n8213) );
  INV_X1 U7977 ( .A(n8211), .ZN(n8210) );
  INV_X1 U7978 ( .A(n13911), .ZN(n8214) );
  NAND2_X1 U7979 ( .A1(n13144), .A2(n10938), .ZN(n10541) );
  NOR2_X1 U7980 ( .A1(n7417), .A2(n7416), .ZN(n7414) );
  INV_X1 U7981 ( .A(n10570), .ZN(n7417) );
  OR2_X1 U7982 ( .A1(n12739), .A2(n8226), .ZN(n8225) );
  INV_X1 U7983 ( .A(n12597), .ZN(n8226) );
  AND2_X1 U7984 ( .A1(n8222), .A2(n10677), .ZN(n8221) );
  OR2_X1 U7985 ( .A1(n12739), .A2(n8223), .ZN(n8222) );
  AND4_X1 U7986 ( .A1(n13436), .A2(n13435), .A3(n13434), .A4(n14056), .ZN(
        n13439) );
  AND2_X1 U7987 ( .A1(n10435), .A2(n13445), .ZN(n11465) );
  NAND2_X1 U7988 ( .A1(n13318), .A2(n13317), .ZN(n14032) );
  AND2_X1 U7989 ( .A1(n10875), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n10892) );
  NAND2_X1 U7990 ( .A1(n8060), .A2(n7306), .ZN(n14071) );
  OR2_X1 U7991 ( .A1(n14066), .A2(n14072), .ZN(n14069) );
  NAND2_X1 U7992 ( .A1(n14081), .A2(n13039), .ZN(n7367) );
  NAND2_X1 U7993 ( .A1(n8089), .A2(n13060), .ZN(n14043) );
  NAND2_X1 U7994 ( .A1(n14088), .A2(n14087), .ZN(n8089) );
  NAND2_X1 U7995 ( .A1(n14131), .A2(n13036), .ZN(n14111) );
  NAND2_X1 U7996 ( .A1(n14111), .A2(n14114), .ZN(n14113) );
  NAND2_X1 U7997 ( .A1(n14133), .A2(n14132), .ZN(n14131) );
  NAND2_X1 U7998 ( .A1(n14172), .A2(n14144), .ZN(n8059) );
  NAND2_X1 U7999 ( .A1(n13034), .A2(n8056), .ZN(n8055) );
  NAND2_X1 U8000 ( .A1(n13047), .A2(n7494), .ZN(n7810) );
  AND2_X1 U8001 ( .A1(n7286), .A2(n13046), .ZN(n7494) );
  INV_X1 U8002 ( .A(n13052), .ZN(n7814) );
  AOI21_X1 U8003 ( .B1(n7815), .B2(n7813), .A(n7277), .ZN(n7812) );
  NOR2_X1 U8004 ( .A1(n7816), .A2(n13052), .ZN(n7813) );
  NAND2_X1 U8005 ( .A1(n14175), .A2(n13032), .ZN(n13034) );
  NOR2_X1 U8006 ( .A1(n14194), .A2(n8049), .ZN(n8048) );
  INV_X1 U8007 ( .A(n13029), .ZN(n8049) );
  INV_X1 U8008 ( .A(n10938), .ZN(n11781) );
  NAND2_X1 U8009 ( .A1(n13047), .A2(n13046), .ZN(n14188) );
  INV_X1 U8010 ( .A(n12993), .ZN(n8046) );
  AOI21_X1 U8011 ( .B1(n12899), .B2(n7485), .A(n7250), .ZN(n7484) );
  INV_X1 U8012 ( .A(n12823), .ZN(n7485) );
  NAND2_X1 U8013 ( .A1(n7483), .A2(n12899), .ZN(n7482) );
  NAND2_X1 U8014 ( .A1(n12898), .A2(n12897), .ZN(n12992) );
  NAND2_X1 U8015 ( .A1(n12831), .A2(n12830), .ZN(n12898) );
  NAND2_X1 U8016 ( .A1(n12704), .A2(n7368), .ZN(n8062) );
  NOR2_X1 U8017 ( .A1(n12827), .A2(n7369), .ZN(n7368) );
  INV_X1 U8018 ( .A(n12703), .ZN(n7369) );
  AND2_X1 U8019 ( .A1(n12528), .A2(n12699), .ZN(n13417) );
  NAND2_X1 U8020 ( .A1(n12526), .A2(n12525), .ZN(n12582) );
  NAND2_X1 U8021 ( .A1(n12533), .A2(n12532), .ZN(n12535) );
  OAI211_X1 U8022 ( .C1(n12077), .C2(n7356), .A(n8063), .B(n7354), .ZN(n12166)
         );
  AND2_X1 U8023 ( .A1(n13413), .A2(n12078), .ZN(n8063) );
  NAND2_X1 U8024 ( .A1(n13412), .A2(n7355), .ZN(n7354) );
  INV_X1 U8025 ( .A(n13412), .ZN(n7356) );
  NAND2_X1 U8026 ( .A1(n10489), .A2(n10488), .ZN(n13202) );
  OR2_X1 U8027 ( .A1(n10483), .A2(n7191), .ZN(n10489) );
  NOR2_X1 U8028 ( .A1(n13413), .A2(n8083), .ZN(n8082) );
  INV_X1 U8029 ( .A(n12072), .ZN(n8083) );
  NAND2_X1 U8030 ( .A1(n8085), .A2(n8086), .ZN(n8084) );
  INV_X1 U8031 ( .A(n12188), .ZN(n8085) );
  NAND2_X1 U8032 ( .A1(n10608), .A2(n10607), .ZN(n13195) );
  NAND2_X1 U8033 ( .A1(n12077), .A2(n12076), .ZN(n12181) );
  NAND2_X1 U8034 ( .A1(n12181), .A2(n13412), .ZN(n12180) );
  NAND2_X1 U8035 ( .A1(n11770), .A2(n13407), .ZN(n7352) );
  NAND2_X1 U8036 ( .A1(n15948), .A2(n15895), .ZN(n11701) );
  INV_X1 U8037 ( .A(n7190), .ZN(n7428) );
  INV_X1 U8038 ( .A(n14089), .ZN(n14189) );
  INV_X1 U8039 ( .A(n14091), .ZN(n14191) );
  OR2_X1 U8040 ( .A1(n12623), .A2(n7191), .ZN(n10795) );
  NAND2_X1 U8041 ( .A1(n10912), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10920) );
  OR2_X1 U8042 ( .A1(n10911), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n10912) );
  XNOR2_X1 U8043 ( .A(n10927), .B(n10926), .ZN(n12734) );
  NAND2_X1 U8044 ( .A1(n10436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10442) );
  INV_X1 U8045 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n10441) );
  NOR2_X1 U8046 ( .A1(n7244), .A2(n10415), .ZN(n7731) );
  INV_X1 U8047 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n10445) );
  OR2_X1 U8048 ( .A1(n10484), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U8049 ( .A1(n7373), .A2(SI_2_), .ZN(n8423) );
  NAND2_X1 U8050 ( .A1(n8142), .A2(n8141), .ZN(n7373) );
  INV_X1 U8051 ( .A(n7545), .ZN(n8588) );
  OAI21_X1 U8052 ( .B1(n7546), .B2(SI_3_), .A(n8425), .ZN(n7545) );
  NAND2_X1 U8053 ( .A1(n8401), .A2(n8400), .ZN(n8399) );
  INV_X1 U8054 ( .A(n8402), .ZN(n8401) );
  NOR2_X1 U8055 ( .A1(n8358), .A2(n11912), .ZN(n8356) );
  NAND2_X1 U8056 ( .A1(n8361), .A2(n8351), .ZN(n8350) );
  INV_X1 U8057 ( .A(n8358), .ZN(n8359) );
  INV_X1 U8058 ( .A(n11837), .ZN(n8351) );
  INV_X1 U8059 ( .A(n8361), .ZN(n8352) );
  OAI21_X1 U8060 ( .B1(n8358), .B2(n8354), .A(n12090), .ZN(n8353) );
  INV_X1 U8061 ( .A(n11912), .ZN(n8355) );
  INV_X1 U8062 ( .A(n12349), .ZN(n8390) );
  NAND2_X1 U8063 ( .A1(n14400), .A2(n14652), .ZN(n8391) );
  AOI21_X1 U8064 ( .B1(n8381), .B2(n8384), .A(n7326), .ZN(n8380) );
  INV_X1 U8065 ( .A(n14723), .ZN(n8384) );
  NAND2_X1 U8066 ( .A1(n8373), .A2(n14444), .ZN(n8370) );
  OR2_X1 U8067 ( .A1(n14488), .A2(n14487), .ZN(n14489) );
  NAND2_X1 U8068 ( .A1(n7228), .A2(n8361), .ZN(n8360) );
  NAND2_X1 U8069 ( .A1(n12004), .A2(n12003), .ZN(n8361) );
  NAND2_X1 U8070 ( .A1(n11838), .A2(n11837), .ZN(n11911) );
  OR2_X1 U8071 ( .A1(n11913), .A2(n11912), .ZN(n8362) );
  NOR2_X1 U8072 ( .A1(n10281), .A2(n7559), .ZN(n7558) );
  OR2_X1 U8073 ( .A1(n7560), .A2(n10282), .ZN(n7559) );
  NAND2_X1 U8074 ( .A1(n10155), .A2(n10154), .ZN(n10245) );
  INV_X1 U8075 ( .A(n14872), .ZN(n8317) );
  AND2_X1 U8076 ( .A1(n15055), .A2(n14516), .ZN(n8279) );
  INV_X1 U8077 ( .A(n7528), .ZN(n14933) );
  NAND2_X1 U8078 ( .A1(n14933), .A2(n14932), .ZN(n14931) );
  INV_X1 U8079 ( .A(n8271), .ZN(n8270) );
  OAI211_X1 U8080 ( .C1(n7569), .C2(n15010), .A(n7568), .B(n7566), .ZN(n7565)
         );
  AND2_X1 U8081 ( .A1(n7567), .A2(n7291), .ZN(n7566) );
  NAND2_X1 U8082 ( .A1(n7684), .A2(n14960), .ZN(n7569) );
  NAND2_X1 U8083 ( .A1(n10222), .A2(n8254), .ZN(n8246) );
  NAND2_X1 U8084 ( .A1(n8246), .A2(n8244), .ZN(n8249) );
  NOR2_X1 U8085 ( .A1(n8250), .A2(n8245), .ZN(n8244) );
  NAND2_X1 U8086 ( .A1(n14991), .A2(n14990), .ZN(n14989) );
  NAND2_X1 U8087 ( .A1(n8831), .A2(n8830), .ZN(n14449) );
  AOI21_X1 U8088 ( .B1(n7590), .B2(n7598), .A(n8837), .ZN(n7589) );
  NAND2_X1 U8089 ( .A1(n12480), .A2(n7592), .ZN(n7591) );
  INV_X1 U8090 ( .A(n7595), .ZN(n7590) );
  NOR2_X1 U8091 ( .A1(n8257), .A2(n7596), .ZN(n7595) );
  INV_X1 U8092 ( .A(n9010), .ZN(n7596) );
  OR2_X1 U8093 ( .A1(n12856), .A2(n8258), .ZN(n8257) );
  NAND2_X1 U8094 ( .A1(n12633), .A2(n9012), .ZN(n8258) );
  NAND2_X1 U8095 ( .A1(n12855), .A2(n7520), .ZN(n12932) );
  NAND2_X1 U8096 ( .A1(n12857), .A2(n12856), .ZN(n12855) );
  NAND2_X1 U8097 ( .A1(n7597), .A2(n9010), .ZN(n12629) );
  NAND2_X1 U8098 ( .A1(n7517), .A2(n8329), .ZN(n12400) );
  NAND2_X1 U8099 ( .A1(n12315), .A2(n12314), .ZN(n12313) );
  INV_X1 U8100 ( .A(n10214), .ZN(n12314) );
  INV_X1 U8101 ( .A(n12200), .ZN(n12196) );
  AOI21_X1 U8102 ( .B1(n12255), .B2(n12254), .A(n9003), .ZN(n12199) );
  NAND2_X1 U8103 ( .A1(n11804), .A2(n11803), .ZN(n11802) );
  NAND2_X1 U8104 ( .A1(n12289), .A2(n12290), .ZN(n8999) );
  INV_X1 U8105 ( .A(n15916), .ZN(n14914) );
  OAI21_X1 U8106 ( .B1(n8563), .B2(n14773), .A(n7530), .ZN(n7532) );
  NAND2_X1 U8107 ( .A1(n7698), .A2(n7697), .ZN(n7696) );
  NAND2_X1 U8108 ( .A1(n8563), .A2(n7531), .ZN(n7530) );
  INV_X1 U8109 ( .A(n14848), .ZN(n15035) );
  NAND2_X1 U8110 ( .A1(n8897), .A2(n8896), .ZN(n15086) );
  NAND2_X1 U8111 ( .A1(n7861), .A2(n8347), .ZN(n15880) );
  INV_X1 U8112 ( .A(n10040), .ZN(n8347) );
  XNOR2_X1 U8113 ( .A(n10168), .B(n10170), .ZN(n13351) );
  NAND2_X1 U8114 ( .A1(n8112), .A2(n8113), .ZN(n10168) );
  XNOR2_X1 U8115 ( .A(n10148), .B(n10147), .ZN(n14369) );
  NAND2_X1 U8116 ( .A1(n8932), .A2(n8482), .ZN(n8936) );
  NAND2_X1 U8117 ( .A1(n8911), .A2(n8478), .ZN(n8922) );
  NAND2_X1 U8118 ( .A1(n8490), .A2(n9031), .ZN(n9035) );
  INV_X1 U8119 ( .A(n9033), .ZN(n9031) );
  OAI21_X1 U8120 ( .B1(n8772), .B2(n8771), .A(n8452), .ZN(n8791) );
  AOI21_X1 U8121 ( .B1(n8130), .B2(n8129), .A(n7275), .ZN(n8128) );
  INV_X1 U8122 ( .A(n8445), .ZN(n8129) );
  NAND2_X1 U8123 ( .A1(n8127), .A2(n8130), .ZN(n8126) );
  AOI21_X1 U8124 ( .B1(n7807), .B2(n8436), .A(n7263), .ZN(n7806) );
  NAND2_X1 U8125 ( .A1(n7478), .A2(n8439), .ZN(n8704) );
  INV_X1 U8126 ( .A(n8684), .ZN(n7478) );
  AOI21_X1 U8127 ( .B1(n8648), .B2(n7549), .A(n7548), .ZN(n7547) );
  INV_X1 U8128 ( .A(n8434), .ZN(n7548) );
  INV_X1 U8129 ( .A(n8431), .ZN(n7549) );
  INV_X1 U8130 ( .A(n8425), .ZN(n8105) );
  INV_X1 U8131 ( .A(n8426), .ZN(n8104) );
  NAND2_X1 U8132 ( .A1(n8589), .A2(n8588), .ZN(n7379) );
  XNOR2_X1 U8133 ( .A(n10343), .B(n10346), .ZN(n10345) );
  XNOR2_X1 U8134 ( .A(n10339), .B(n7913), .ZN(n10350) );
  OAI22_X1 U8135 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n10306), .B1(n10305), .B2(
        n10354), .ZN(n10358) );
  INV_X1 U8136 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10306) );
  NAND2_X1 U8137 ( .A1(n7911), .A2(n7252), .ZN(n7910) );
  AOI21_X1 U8138 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n10316), .A(n10315), .ZN(
        n10336) );
  NOR2_X1 U8139 ( .A1(n10369), .A2(n10368), .ZN(n10315) );
  AND2_X1 U8140 ( .A1(n7923), .A2(n7924), .ZN(n10377) );
  NAND2_X1 U8141 ( .A1(n10373), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U8142 ( .A1(n15574), .A2(n15573), .ZN(n10373) );
  NAND2_X1 U8143 ( .A1(n12372), .A2(n7525), .ZN(n12495) );
  AND2_X1 U8144 ( .A1(n12363), .A2(n12364), .ZN(n7525) );
  NOR2_X1 U8145 ( .A1(n8300), .A2(n7264), .ZN(n8299) );
  OAI21_X1 U8146 ( .B1(n11227), .B2(n11228), .A(n11347), .ZN(n11230) );
  NOR2_X1 U8147 ( .A1(n11230), .A2(n11229), .ZN(n11349) );
  AND4_X1 U8148 ( .A1(n9512), .A2(n9511), .A3(n9510), .A4(n9509), .ZN(n13504)
         );
  NAND2_X1 U8149 ( .A1(n12373), .A2(n12374), .ZN(n12372) );
  AND4_X1 U8150 ( .A1(n9378), .A2(n9377), .A3(n9376), .A4(n9375), .ZN(n13746)
         );
  INV_X1 U8151 ( .A(n13504), .ZN(n13665) );
  INV_X1 U8152 ( .A(n13746), .ZN(n13573) );
  AND2_X1 U8153 ( .A1(n9147), .A2(n9169), .ZN(n15650) );
  NOR2_X1 U8154 ( .A1(n15710), .A2(n9909), .ZN(n15728) );
  XNOR2_X1 U8155 ( .A(n7468), .B(n11030), .ZN(n15754) );
  NOR2_X1 U8156 ( .A1(n15754), .A2(n15755), .ZN(n15756) );
  NAND2_X1 U8157 ( .A1(n7475), .A2(n7474), .ZN(n7477) );
  AOI21_X1 U8158 ( .B1(n9922), .B2(n7476), .A(n7346), .ZN(n7474) );
  NAND2_X1 U8159 ( .A1(n7535), .A2(n7753), .ZN(n7534) );
  INV_X1 U8160 ( .A(n10033), .ZN(n7753) );
  NAND2_X1 U8161 ( .A1(n7443), .A2(n9606), .ZN(n13600) );
  NAND2_X1 U8162 ( .A1(n7439), .A2(n7438), .ZN(n7443) );
  AND3_X1 U8163 ( .A1(n9175), .A2(n9174), .A3(n9173), .ZN(n16022) );
  NOR2_X1 U8164 ( .A1(n8405), .A2(n7226), .ZN(n9115) );
  NAND2_X1 U8165 ( .A1(n9100), .A2(n8006), .ZN(n11669) );
  OAI22_X1 U8166 ( .A1(n9262), .A2(n15267), .B1(n11016), .B2(n9928), .ZN(n8007) );
  NOR2_X1 U8167 ( .A1(n13600), .A2(n9627), .ZN(n10405) );
  AND2_X1 U8168 ( .A1(n13599), .A2(n16160), .ZN(n9627) );
  NAND2_X1 U8169 ( .A1(n9428), .A2(n9427), .ZN(n13860) );
  NAND2_X1 U8170 ( .A1(n16169), .A2(n16107), .ZN(n13864) );
  AND2_X1 U8171 ( .A1(n9925), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13870) );
  AND2_X1 U8172 ( .A1(n9643), .A2(n9642), .ZN(n13871) );
  INV_X1 U8173 ( .A(n14005), .ZN(n14101) );
  INV_X1 U8174 ( .A(n14007), .ZN(n14145) );
  NOR2_X1 U8175 ( .A1(n10628), .A2(n12145), .ZN(n12138) );
  NAND2_X1 U8176 ( .A1(n10743), .A2(n10742), .ZN(n14317) );
  AND2_X1 U8177 ( .A1(n11736), .A2(n10617), .ZN(n10618) );
  INV_X1 U8178 ( .A(n14108), .ZN(n14285) );
  NAND2_X1 U8179 ( .A1(n11484), .A2(n10570), .ZN(n7415) );
  NAND2_X1 U8180 ( .A1(n10768), .A2(n10767), .ZN(n14314) );
  OR2_X1 U8181 ( .A1(n10646), .A2(n10647), .ZN(n7425) );
  INV_X1 U8182 ( .A(n13144), .ZN(n12036) );
  NAND2_X1 U8183 ( .A1(n10942), .A2(n16038), .ZN(n13999) );
  NAND2_X1 U8184 ( .A1(n13441), .A2(n13440), .ZN(n13453) );
  NAND2_X1 U8185 ( .A1(n13439), .A2(n13024), .ZN(n13440) );
  NAND2_X1 U8186 ( .A1(n13438), .A2(n13437), .ZN(n13441) );
  NOR2_X1 U8187 ( .A1(n13439), .A2(n13024), .ZN(n13437) );
  AOI21_X1 U8188 ( .B1(n10448), .B2(n7239), .A(n7409), .ZN(n7408) );
  NAND2_X1 U8189 ( .A1(n10885), .A2(n10884), .ZN(n14092) );
  NAND4_X1 U8190 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(
        n14025) );
  NAND2_X1 U8191 ( .A1(n10652), .A2(n10651), .ZN(n16148) );
  NAND2_X1 U8192 ( .A1(n15409), .A2(n11474), .ZN(n16038) );
  INV_X1 U8193 ( .A(n13063), .ZN(n14277) );
  NAND2_X1 U8194 ( .A1(n12095), .A2(n12094), .ZN(n12346) );
  NAND2_X1 U8195 ( .A1(n14718), .A2(n14723), .ZN(n7686) );
  INV_X1 U8196 ( .A(n14584), .ZN(n7685) );
  NAND2_X1 U8197 ( .A1(n8778), .A2(n8777), .ZN(n16177) );
  NAND2_X1 U8198 ( .A1(n7380), .A2(n8397), .ZN(n16172) );
  NAND2_X1 U8199 ( .A1(n14417), .A2(n8398), .ZN(n8397) );
  NAND2_X1 U8200 ( .A1(n7382), .A2(n7381), .ZN(n7380) );
  OR2_X1 U8201 ( .A1(n11043), .A2(n8937), .ZN(n8709) );
  NAND2_X1 U8202 ( .A1(n8816), .A2(n8815), .ZN(n16199) );
  NAND2_X1 U8203 ( .A1(n7557), .A2(n8912), .ZN(n15063) );
  NAND2_X1 U8204 ( .A1(n12607), .A2(n10171), .ZN(n7557) );
  NAND2_X1 U8205 ( .A1(n14571), .A2(n14476), .ZN(n14601) );
  NAND2_X1 U8206 ( .A1(n11555), .A2(n11554), .ZN(n14740) );
  NAND4_X1 U8207 ( .A1(n8587), .A2(n8586), .A3(n8585), .A4(n8584), .ZN(n14767)
         );
  NAND2_X1 U8208 ( .A1(n15530), .A2(n12667), .ZN(n12669) );
  INV_X1 U8209 ( .A(n12665), .ZN(n12666) );
  OAI21_X1 U8210 ( .B1(n14833), .B2(n15859), .A(n7799), .ZN(n7798) );
  AOI21_X1 U8211 ( .B1(n14834), .B2(n15869), .A(n15862), .ZN(n7799) );
  NAND2_X1 U8212 ( .A1(n13076), .A2(n7683), .ZN(n7682) );
  INV_X1 U8213 ( .A(n13075), .ZN(n7683) );
  OR2_X1 U8214 ( .A1(n13071), .A2(n16134), .ZN(n13076) );
  NAND2_X1 U8215 ( .A1(n8883), .A2(n8882), .ZN(n15099) );
  NAND2_X1 U8216 ( .A1(n8621), .A2(n8620), .ZN(n12159) );
  OR2_X2 U8217 ( .A1(n11560), .A2(n11558), .ZN(n15931) );
  NAND2_X1 U8218 ( .A1(n8278), .A2(n16019), .ZN(n8277) );
  AND2_X1 U8219 ( .A1(n8412), .A2(n7574), .ZN(n7573) );
  INV_X1 U8220 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7574) );
  OR2_X1 U8221 ( .A1(n7919), .A2(n15552), .ZN(n7916) );
  INV_X1 U8222 ( .A(n10353), .ZN(n7920) );
  OR2_X1 U8223 ( .A1(n15559), .A2(n15560), .ZN(n7911) );
  XNOR2_X1 U8224 ( .A(n7910), .B(n7909), .ZN(n15563) );
  INV_X1 U8225 ( .A(n10366), .ZN(n7909) );
  AND2_X1 U8226 ( .A1(n7611), .A2(n7610), .ZN(n15569) );
  INV_X1 U8227 ( .A(n15564), .ZN(n7611) );
  NAND2_X1 U8228 ( .A1(n10370), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7610) );
  XNOR2_X1 U8229 ( .A(n10377), .B(n7922), .ZN(n15578) );
  INV_X1 U8230 ( .A(n10376), .ZN(n7922) );
  OAI21_X1 U8231 ( .B1(n15581), .B2(n15580), .A(n7693), .ZN(n7692) );
  INV_X1 U8232 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7693) );
  NOR2_X1 U8233 ( .A1(n10389), .A2(n15597), .ZN(n15601) );
  NAND2_X1 U8234 ( .A1(n7618), .A2(n7617), .ZN(n7927) );
  INV_X1 U8235 ( .A(n15600), .ZN(n7617) );
  INV_X1 U8236 ( .A(n15601), .ZN(n7618) );
  NAND2_X1 U8237 ( .A1(n7929), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U8238 ( .A1(n15601), .A2(n15600), .ZN(n7929) );
  XNOR2_X1 U8239 ( .A(n10399), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n10400) );
  NAND2_X1 U8240 ( .A1(n7964), .A2(n7963), .ZN(n10064) );
  NOR2_X1 U8241 ( .A1(n13173), .A2(n13170), .ZN(n7703) );
  NAND2_X1 U8242 ( .A1(n7844), .A2(n7843), .ZN(n10073) );
  NAND2_X1 U8243 ( .A1(n10068), .A2(n10070), .ZN(n7843) );
  NAND2_X1 U8244 ( .A1(n10073), .A2(n10074), .ZN(n10072) );
  NAND2_X1 U8245 ( .A1(n13187), .A2(n7223), .ZN(n13192) );
  INV_X1 U8246 ( .A(n7283), .ZN(n7713) );
  INV_X1 U8247 ( .A(n13198), .ZN(n7712) );
  NAND2_X1 U8248 ( .A1(n13198), .A2(n7283), .ZN(n7711) );
  AOI21_X1 U8249 ( .B1(n7194), .B2(n7711), .A(n7204), .ZN(n7709) );
  NAND2_X1 U8250 ( .A1(n7839), .A2(n7838), .ZN(n10088) );
  NAND2_X1 U8251 ( .A1(n10083), .A2(n10085), .ZN(n7838) );
  NAND2_X1 U8252 ( .A1(n13221), .A2(n7729), .ZN(n13229) );
  INV_X1 U8253 ( .A(n13220), .ZN(n7730) );
  NOR2_X1 U8254 ( .A1(n13239), .A2(n13241), .ZN(n8190) );
  NAND2_X1 U8255 ( .A1(n13229), .A2(n13230), .ZN(n13228) );
  AND2_X1 U8256 ( .A1(n8190), .A2(n7718), .ZN(n7717) );
  INV_X1 U8257 ( .A(n13246), .ZN(n7718) );
  NAND2_X1 U8258 ( .A1(n7834), .A2(n7833), .ZN(n10103) );
  NAND2_X1 U8259 ( .A1(n10098), .A2(n10100), .ZN(n7833) );
  INV_X1 U8260 ( .A(n13252), .ZN(n8192) );
  NOR2_X1 U8261 ( .A1(n13258), .A2(n13257), .ZN(n7735) );
  NOR2_X1 U8262 ( .A1(n13264), .A2(n7272), .ZN(n8185) );
  NAND2_X1 U8263 ( .A1(n7848), .A2(n7847), .ZN(n10115) );
  NAND2_X1 U8264 ( .A1(n10110), .A2(n10112), .ZN(n7847) );
  NOR2_X1 U8265 ( .A1(n13272), .A2(n8189), .ZN(n7706) );
  NOR2_X1 U8266 ( .A1(n13276), .A2(n13278), .ZN(n8189) );
  NAND2_X1 U8267 ( .A1(n13269), .A2(n13268), .ZN(n7707) );
  NAND2_X1 U8268 ( .A1(n10119), .A2(n7959), .ZN(n7958) );
  NAND2_X1 U8269 ( .A1(n13285), .A2(n13284), .ZN(n13283) );
  NAND2_X1 U8270 ( .A1(n7829), .A2(n7937), .ZN(n10128) );
  NAND2_X1 U8271 ( .A1(n10123), .A2(n10125), .ZN(n7937) );
  OAI22_X1 U8272 ( .A1(n13296), .A2(n7728), .B1(n13301), .B2(n13299), .ZN(
        n13308) );
  OAI21_X1 U8273 ( .B1(n13295), .B2(n13294), .A(n7270), .ZN(n7728) );
  AND2_X1 U8274 ( .A1(n10222), .A2(n14979), .ZN(n7556) );
  NAND2_X1 U8275 ( .A1(n10135), .A2(n7955), .ZN(n7954) );
  MUX2_X1 U8276 ( .A(n9745), .B(n9744), .S(n11657), .Z(n9746) );
  INV_X1 U8277 ( .A(n9518), .ZN(n7660) );
  NOR2_X1 U8278 ( .A1(n9499), .A2(n7634), .ZN(n7633) );
  NAND2_X1 U8279 ( .A1(n9470), .A2(n7631), .ZN(n7630) );
  INV_X1 U8280 ( .A(n9487), .ZN(n7634) );
  INV_X1 U8281 ( .A(n9470), .ZN(n7632) );
  NOR2_X1 U8282 ( .A1(n13343), .A2(n13344), .ZN(n8133) );
  INV_X1 U8283 ( .A(n13384), .ZN(n8137) );
  INV_X1 U8284 ( .A(n13383), .ZN(n8136) );
  INV_X1 U8285 ( .A(n13057), .ZN(n8094) );
  NOR2_X1 U8286 ( .A1(n14301), .A2(n14295), .ZN(n7766) );
  NOR2_X1 U8287 ( .A1(n8852), .A2(n8851), .ZN(n8850) );
  NAND2_X1 U8288 ( .A1(n8892), .A2(n8469), .ZN(n7555) );
  INV_X1 U8289 ( .A(n8469), .ZN(n7552) );
  AOI21_X1 U8290 ( .B1(n8121), .B2(n8123), .A(n8120), .ZN(n8119) );
  INV_X1 U8291 ( .A(n8880), .ZN(n8120) );
  INV_X1 U8292 ( .A(n8462), .ZN(n8121) );
  INV_X1 U8293 ( .A(n8123), .ZN(n8122) );
  NAND2_X1 U8294 ( .A1(n8455), .A2(SI_16_), .ZN(n8456) );
  INV_X1 U8295 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7801) );
  INV_X1 U8296 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8106) );
  INV_X1 U8297 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n10302) );
  OR2_X1 U8298 ( .A1(n15654), .A2(n7541), .ZN(n9939) );
  NOR2_X1 U8299 ( .A1(n15650), .A2(n9985), .ZN(n7541) );
  NAND2_X1 U8300 ( .A1(n15696), .A2(n7539), .ZN(n9945) );
  OR2_X1 U8301 ( .A1(n15705), .A2(n16104), .ZN(n7539) );
  NAND2_X1 U8302 ( .A1(n11258), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7979) );
  INV_X1 U8303 ( .A(n13097), .ZN(n7992) );
  INV_X1 U8304 ( .A(n12973), .ZN(n7884) );
  OR2_X1 U8305 ( .A1(n13577), .A2(n12853), .ZN(n9807) );
  INV_X1 U8306 ( .A(n12509), .ZN(n8166) );
  NAND2_X1 U8307 ( .A1(n12231), .A2(n9249), .ZN(n7433) );
  NAND2_X1 U8308 ( .A1(n9232), .A2(n9231), .ZN(n9250) );
  INV_X1 U8309 ( .A(n8036), .ZN(n8032) );
  NOR2_X1 U8310 ( .A1(n10990), .A2(n9660), .ZN(n9888) );
  INV_X1 U8311 ( .A(n9678), .ZN(n7640) );
  INV_X1 U8312 ( .A(n7639), .ZN(n7638) );
  OAI21_X1 U8313 ( .B1(n9676), .B2(n7640), .A(n9687), .ZN(n7639) );
  INV_X1 U8314 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8170) );
  INV_X1 U8315 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9501) );
  INV_X1 U8316 ( .A(n7653), .ZN(n7652) );
  OAI21_X1 U8317 ( .B1(n8016), .B2(n7654), .A(n9306), .ZN(n7653) );
  OR2_X1 U8318 ( .A1(n9220), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9244) );
  NOR2_X1 U8319 ( .A1(n8241), .A2(n7423), .ZN(n7422) );
  INV_X1 U8320 ( .A(n13920), .ZN(n7423) );
  OAI21_X1 U8321 ( .B1(n8218), .B2(n8230), .A(n8229), .ZN(n8217) );
  NAND2_X1 U8322 ( .A1(n8221), .A2(n8225), .ZN(n8218) );
  OAI22_X1 U8323 ( .A1(n13911), .A2(n8212), .B1(n10786), .B2(n10787), .ZN(
        n8211) );
  OR2_X1 U8324 ( .A1(n13959), .A2(n10771), .ZN(n8212) );
  NAND2_X1 U8325 ( .A1(n8186), .A2(n8187), .ZN(n13388) );
  NAND2_X1 U8326 ( .A1(n13316), .A2(n7309), .ZN(n8187) );
  OAI211_X1 U8327 ( .C1(n13385), .C2(n8135), .A(n8134), .B(n8132), .ZN(n13386)
         );
  NAND2_X1 U8328 ( .A1(n8137), .A2(n8136), .ZN(n8135) );
  NAND2_X1 U8329 ( .A1(n13342), .A2(n8133), .ZN(n8132) );
  INV_X1 U8330 ( .A(n13382), .ZN(n8134) );
  NOR2_X1 U8331 ( .A1(n13385), .A2(n13341), .ZN(n13387) );
  NAND2_X1 U8332 ( .A1(n14061), .A2(n7758), .ZN(n7757) );
  AND2_X1 U8333 ( .A1(n13428), .A2(n13055), .ZN(n8095) );
  INV_X1 U8334 ( .A(n10775), .ZN(n10773) );
  NAND2_X1 U8335 ( .A1(n10757), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n10775) );
  INV_X1 U8336 ( .A(n10759), .ZN(n10757) );
  NAND2_X1 U8337 ( .A1(n10731), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n10745) );
  INV_X1 U8338 ( .A(n10733), .ZN(n10731) );
  AND2_X1 U8339 ( .A1(n8045), .A2(n12897), .ZN(n7370) );
  NAND2_X1 U8340 ( .A1(n8077), .A2(n8076), .ZN(n8075) );
  INV_X1 U8341 ( .A(n12076), .ZN(n7355) );
  NOR2_X1 U8342 ( .A1(n11717), .A2(n13168), .ZN(n11687) );
  AND2_X1 U8343 ( .A1(n14167), .A2(n7206), .ZN(n14122) );
  NAND2_X1 U8344 ( .A1(n14167), .A2(n7766), .ZN(n14134) );
  AND2_X1 U8345 ( .A1(n14201), .A2(n14185), .ZN(n14180) );
  NAND2_X1 U8346 ( .A1(n11775), .A2(n11774), .ZN(n11943) );
  INV_X1 U8347 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7363) );
  INV_X1 U8348 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7403) );
  INV_X1 U8349 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8639) );
  INV_X1 U8350 ( .A(n14589), .ZN(n14529) );
  NOR2_X1 U8351 ( .A1(n8801), .A2(n8800), .ZN(n8799) );
  AOI21_X1 U8352 ( .B1(n10253), .B2(n10252), .A(n10251), .ZN(n10257) );
  NOR2_X1 U8353 ( .A1(n10287), .A2(n10283), .ZN(n7560) );
  NAND2_X1 U8354 ( .A1(n10145), .A2(n7854), .ZN(n7853) );
  NAND2_X1 U8355 ( .A1(n10141), .A2(n7961), .ZN(n7960) );
  NAND2_X1 U8356 ( .A1(n10143), .A2(n7962), .ZN(n7961) );
  NOR2_X1 U8357 ( .A1(n12114), .A2(n7794), .ZN(n12664) );
  AND2_X1 U8358 ( .A1(n12115), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7794) );
  AND2_X1 U8359 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n8941), .ZN(n8514) );
  OR2_X1 U8360 ( .A1(n14963), .A2(n9016), .ZN(n7567) );
  OR2_X1 U8361 ( .A1(n8249), .A2(n14963), .ZN(n7568) );
  AND2_X1 U8362 ( .A1(n8850), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8884) );
  INV_X1 U8363 ( .A(n12856), .ZN(n7519) );
  INV_X1 U8364 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8851) );
  AND2_X1 U8365 ( .A1(n7598), .A2(n12481), .ZN(n7592) );
  INV_X1 U8366 ( .A(n8263), .ZN(n8259) );
  INV_X1 U8367 ( .A(n8700), .ZN(n7516) );
  AND2_X1 U8368 ( .A1(n8710), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8727) );
  NOR2_X1 U8369 ( .A1(n8711), .A2(n11332), .ZN(n8710) );
  XNOR2_X1 U8370 ( .A(n14560), .B(n14760), .ZN(n10214) );
  NOR2_X1 U8371 ( .A1(n11632), .A2(n12437), .ZN(n11800) );
  AND2_X1 U8372 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8608) );
  OR2_X1 U8373 ( .A1(n8976), .A2(n11151), .ZN(n8567) );
  OR2_X1 U8374 ( .A1(n8953), .A2(n8566), .ZN(n8569) );
  NAND2_X1 U8375 ( .A1(n10986), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7531) );
  INV_X1 U8376 ( .A(n8937), .ZN(n7698) );
  NAND2_X1 U8377 ( .A1(n14992), .A2(n14984), .ZN(n14964) );
  NOR2_X1 U8378 ( .A1(n12293), .A2(n16008), .ZN(n12295) );
  AOI21_X1 U8379 ( .B1(n8114), .B2(n10147), .A(n7340), .ZN(n8113) );
  INV_X1 U8380 ( .A(n8970), .ZN(n8114) );
  INV_X1 U8381 ( .A(n10147), .ZN(n8115) );
  AND2_X1 U8382 ( .A1(n8500), .A2(n8503), .ZN(n8344) );
  OAI21_X1 U8383 ( .B1(n8962), .B2(n8961), .A(n8960), .ZN(n8967) );
  OAI21_X1 U8384 ( .B1(n8772), .B2(n8145), .A(n8143), .ZN(n8809) );
  AOI21_X1 U8385 ( .B1(n8146), .B2(n8144), .A(n7321), .ZN(n8143) );
  INV_X1 U8386 ( .A(n8146), .ZN(n8145) );
  OR2_X1 U8387 ( .A1(n8635), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n8652) );
  NOR2_X1 U8388 ( .A1(n8105), .A2(n8104), .ZN(n8103) );
  OAI21_X1 U8389 ( .B1(n8424), .B2(n7665), .A(n7664), .ZN(n8417) );
  NAND2_X1 U8390 ( .A1(n8424), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7664) );
  INV_X1 U8391 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10300) );
  OAI22_X1 U8392 ( .A1(n10337), .A2(n10304), .B1(P1_ADDR_REG_4__SCAN_IN), .B2(
        n10303), .ZN(n10354) );
  AOI22_X1 U8393 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10308), .B1(n10307), .B2(
        n10358), .ZN(n10309) );
  OR2_X1 U8394 ( .A1(n10308), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10307) );
  INV_X1 U8395 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10308) );
  OAI21_X1 U8396 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n10326), .A(n10325), .ZN(
        n10333) );
  OR2_X1 U8397 ( .A1(n10332), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U8398 ( .A1(n12023), .A2(n13583), .ZN(n8301) );
  NAND2_X1 U8399 ( .A1(n8283), .A2(n8282), .ZN(n13467) );
  AOI21_X1 U8400 ( .B1(n8285), .B2(n8287), .A(n7308), .ZN(n8282) );
  AND2_X1 U8401 ( .A1(n8305), .A2(n8303), .ZN(n8298) );
  NOR2_X1 U8402 ( .A1(n8301), .A2(n12103), .ZN(n8300) );
  INV_X1 U8403 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15346) );
  INV_X1 U8404 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15348) );
  AOI21_X1 U8405 ( .B1(n8288), .B2(n7512), .A(n7269), .ZN(n7511) );
  INV_X1 U8406 ( .A(n12813), .ZN(n7512) );
  NAND2_X1 U8407 ( .A1(n11649), .A2(n11648), .ZN(n11650) );
  AOI21_X1 U8408 ( .B1(n7511), .B2(n8289), .A(n7510), .ZN(n7509) );
  INV_X1 U8409 ( .A(n13082), .ZN(n7510) );
  NAND2_X1 U8410 ( .A1(n13093), .A2(n8311), .ZN(n13527) );
  INV_X1 U8411 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15369) );
  AND2_X1 U8412 ( .A1(n9447), .A2(n15369), .ZN(n9461) );
  NOR2_X1 U8413 ( .A1(n9288), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9319) );
  NOR2_X1 U8414 ( .A1(n8310), .A2(n8309), .ZN(n8308) );
  OAI21_X1 U8415 ( .B1(n8310), .B2(n13095), .A(n8307), .ZN(n8306) );
  INV_X1 U8416 ( .A(n8311), .ZN(n8309) );
  AND2_X1 U8417 ( .A1(n9461), .A2(n15348), .ZN(n9475) );
  OR2_X1 U8418 ( .A1(n9409), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U8419 ( .A1(n11988), .A2(n11994), .ZN(n11989) );
  OR2_X1 U8420 ( .A1(n9523), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9539) );
  NOR4_X1 U8421 ( .A1(n9724), .A2(n9863), .A3(n9723), .A4(n9747), .ZN(n9726)
         );
  INV_X1 U8422 ( .A(n9700), .ZN(n7995) );
  NAND2_X1 U8423 ( .A1(n9139), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U8424 ( .A1(n9103), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U8425 ( .A1(n9930), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7461) );
  NAND3_X1 U8426 ( .A1(n7462), .A2(n9085), .A3(n7460), .ZN(n7459) );
  OR2_X1 U8427 ( .A1(n11398), .A2(n11397), .ZN(n11400) );
  NAND2_X1 U8428 ( .A1(n7749), .A2(n7748), .ZN(n9971) );
  OR2_X1 U8429 ( .A1(n13132), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U8430 ( .A1(n13132), .A2(n9970), .ZN(n7748) );
  NAND2_X1 U8431 ( .A1(n11372), .A2(n11373), .ZN(n11371) );
  OR2_X1 U8432 ( .A1(n15621), .A2(n15622), .ZN(n7467) );
  XNOR2_X1 U8433 ( .A(n9939), .B(n15664), .ZN(n15670) );
  INV_X1 U8434 ( .A(n9900), .ZN(n7981) );
  NAND2_X1 U8435 ( .A1(n7982), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7980) );
  NAND3_X1 U8436 ( .A1(n7971), .A2(n7970), .A3(n7972), .ZN(n11614) );
  NAND2_X1 U8437 ( .A1(n9902), .A2(n11620), .ZN(n7972) );
  NAND2_X1 U8438 ( .A1(n15661), .A2(n9994), .ZN(n15682) );
  AND2_X1 U8439 ( .A1(n7470), .A2(n7469), .ZN(n9905) );
  NAND2_X1 U8440 ( .A1(n11760), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7469) );
  NAND2_X1 U8441 ( .A1(n7745), .A2(n7744), .ZN(n12059) );
  INV_X1 U8442 ( .A(n12062), .ZN(n7744) );
  INV_X1 U8443 ( .A(n12061), .ZN(n7745) );
  NAND2_X1 U8444 ( .A1(n12055), .A2(n9944), .ZN(n15698) );
  NAND2_X1 U8445 ( .A1(n15698), .A2(n15697), .ZN(n15696) );
  NOR2_X1 U8446 ( .A1(n9905), .A2(n9904), .ZN(n9906) );
  XNOR2_X1 U8447 ( .A(n9945), .B(n10015), .ZN(n15716) );
  NAND2_X1 U8448 ( .A1(n15702), .A2(n10013), .ZN(n15714) );
  NOR2_X1 U8449 ( .A1(n15694), .A2(n7691), .ZN(n9908) );
  NOR2_X1 U8450 ( .A1(n15705), .A2(n9907), .ZN(n7691) );
  INV_X1 U8451 ( .A(n7975), .ZN(n9918) );
  NOR2_X1 U8452 ( .A1(n15790), .A2(n7752), .ZN(n15801) );
  AND2_X1 U8453 ( .A1(n10027), .A2(n15789), .ZN(n7752) );
  NAND2_X1 U8454 ( .A1(n15785), .A2(n9954), .ZN(n15803) );
  OAI21_X1 U8455 ( .B1(n7472), .B2(n15782), .A(n7471), .ZN(n9921) );
  NAND2_X1 U8456 ( .A1(n15808), .A2(n7979), .ZN(n7471) );
  OR2_X1 U8457 ( .A1(n9919), .A2(n7473), .ZN(n7472) );
  INV_X1 U8458 ( .A(n7979), .ZN(n7473) );
  INV_X1 U8459 ( .A(n15846), .ZN(n7476) );
  XNOR2_X1 U8460 ( .A(n10031), .B(n10032), .ZN(n7754) );
  NAND2_X1 U8461 ( .A1(n15817), .A2(n9958), .ZN(n15836) );
  OAI21_X1 U8462 ( .B1(n13609), .B2(n7441), .A(n7440), .ZN(n7437) );
  AOI21_X1 U8463 ( .B1(n9706), .B2(n9578), .A(n15959), .ZN(n7440) );
  NAND2_X1 U8464 ( .A1(n9587), .A2(n7442), .ZN(n7441) );
  NAND2_X1 U8465 ( .A1(n13609), .A2(n9706), .ZN(n7438) );
  NAND2_X1 U8466 ( .A1(n8174), .A2(n8173), .ZN(n13625) );
  AOI21_X1 U8467 ( .B1(n7196), .B2(n13654), .A(n7271), .ZN(n8173) );
  OAI21_X1 U8468 ( .B1(n9486), .B2(n7455), .A(n7453), .ZN(n8174) );
  NAND2_X1 U8469 ( .A1(n9486), .A2(n7456), .ZN(n13664) );
  AOI21_X1 U8470 ( .B1(n8161), .B2(n8159), .A(n7208), .ZN(n8158) );
  INV_X1 U8471 ( .A(n8161), .ZN(n8160) );
  INV_X1 U8472 ( .A(n8163), .ZN(n8159) );
  NAND2_X1 U8473 ( .A1(n13706), .A2(n9452), .ZN(n13690) );
  NAND2_X1 U8474 ( .A1(n9438), .A2(n8163), .ZN(n13706) );
  NAND2_X1 U8475 ( .A1(n7447), .A2(n7446), .ZN(n13719) );
  AOI21_X1 U8476 ( .B1(n7448), .B2(n7450), .A(n7320), .ZN(n7446) );
  NAND2_X1 U8477 ( .A1(n12971), .A2(n7448), .ZN(n7447) );
  AND2_X1 U8478 ( .A1(n8153), .A2(n7449), .ZN(n7448) );
  NAND2_X1 U8479 ( .A1(n7451), .A2(n12969), .ZN(n7449) );
  AND2_X1 U8480 ( .A1(n9415), .A2(n8154), .ZN(n8153) );
  NAND2_X1 U8481 ( .A1(n8156), .A2(n13017), .ZN(n8154) );
  OR2_X1 U8482 ( .A1(n12971), .A2(n7450), .ZN(n7445) );
  NOR2_X1 U8483 ( .A1(n9353), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9373) );
  OR2_X1 U8484 ( .A1(n9336), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9353) );
  OAI21_X1 U8485 ( .B1(n12651), .B2(n7322), .A(n7444), .ZN(n12749) );
  OR2_X1 U8486 ( .A1(n12853), .A2(n12776), .ZN(n7444) );
  NOR2_X1 U8487 ( .A1(n9615), .A2(n12499), .ZN(n8167) );
  OR2_X1 U8488 ( .A1(n9270), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9288) );
  OR2_X1 U8489 ( .A1(n9250), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9270) );
  OAI21_X1 U8490 ( .B1(n12231), .B2(n7227), .A(n9249), .ZN(n12508) );
  INV_X1 U8491 ( .A(n11002), .ZN(n15664) );
  OAI21_X1 U8492 ( .B1(n15955), .B2(n7876), .A(n7874), .ZN(n9609) );
  INV_X1 U8493 ( .A(n7875), .ZN(n7874) );
  OAI21_X1 U8494 ( .B1(n15957), .B2(n7876), .A(n11957), .ZN(n7875) );
  NAND2_X1 U8495 ( .A1(n9136), .A2(n9135), .ZN(n11960) );
  NOR2_X1 U8496 ( .A1(n13590), .A2(n11592), .ZN(n11496) );
  AND2_X1 U8497 ( .A1(n9629), .A2(n11500), .ZN(n11659) );
  NAND2_X1 U8498 ( .A1(n7627), .A2(n9682), .ZN(n13591) );
  NAND2_X1 U8499 ( .A1(n9474), .A2(n9473), .ZN(n13539) );
  OR2_X1 U8500 ( .A1(n12002), .A2(n9148), .ZN(n9474) );
  INV_X1 U8501 ( .A(n9691), .ZN(n9426) );
  OR2_X1 U8502 ( .A1(n16057), .A2(n16103), .ZN(n16160) );
  NOR2_X1 U8503 ( .A1(n9889), .A2(n9888), .ZN(n11251) );
  OR2_X1 U8504 ( .A1(n9628), .A2(n11657), .ZN(n11500) );
  NAND2_X1 U8505 ( .A1(n9755), .A2(n11967), .ZN(n16157) );
  AOI21_X1 U8506 ( .B1(n7638), .B2(n7640), .A(n7348), .ZN(n7635) );
  AND2_X1 U8507 ( .A1(n9579), .A2(n9565), .ZN(n9566) );
  AOI21_X1 U8508 ( .B1(n9503), .B2(n7659), .A(n7658), .ZN(n7656) );
  XNOR2_X1 U8509 ( .A(n9646), .B(n9645), .ZN(n9925) );
  OAI21_X1 U8510 ( .B1(n9644), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9646) );
  AOI21_X1 U8511 ( .B1(n9402), .B2(n8027), .A(n8026), .ZN(n8025) );
  INV_X1 U8512 ( .A(n9402), .ZN(n8028) );
  INV_X1 U8513 ( .A(n9416), .ZN(n8026) );
  AND2_X1 U8514 ( .A1(n9439), .A2(n9418), .ZN(n9419) );
  NAND2_X1 U8515 ( .A1(n9368), .A2(n8315), .ZN(n9405) );
  AND2_X1 U8516 ( .A1(n9276), .A2(n9258), .ZN(n9259) );
  NOR2_X1 U8517 ( .A1(n9244), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9264) );
  INV_X1 U8518 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9263) );
  AND2_X1 U8519 ( .A1(n9256), .A2(n9240), .ZN(n9241) );
  AOI21_X1 U8520 ( .B1(n7645), .B2(n7647), .A(n7643), .ZN(n7642) );
  INV_X1 U8521 ( .A(n9187), .ZN(n7643) );
  OR2_X1 U8522 ( .A1(n9146), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9169) );
  NOR2_X1 U8523 ( .A1(n9169), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9200) );
  NOR2_X1 U8524 ( .A1(n9130), .A2(n9129), .ZN(n9980) );
  NAND2_X1 U8525 ( .A1(n9110), .A2(n9109), .ZN(n7619) );
  XNOR2_X1 U8526 ( .A(n13195), .B(n10835), .ZN(n10619) );
  NOR2_X1 U8527 ( .A1(n12600), .A2(n12596), .ZN(n8227) );
  INV_X1 U8528 ( .A(n7422), .ZN(n7421) );
  NAND2_X1 U8529 ( .A1(n7422), .A2(n7419), .ZN(n7418) );
  INV_X1 U8530 ( .A(n10840), .ZN(n7419) );
  INV_X1 U8531 ( .A(n8240), .ZN(n8239) );
  OAI22_X1 U8532 ( .A1(n7222), .A2(n8241), .B1(n10888), .B2(n10889), .ZN(n8240) );
  INV_X1 U8533 ( .A(n8236), .ZN(n8235) );
  NAND2_X1 U8534 ( .A1(n13960), .A2(n13959), .ZN(n13958) );
  NAND2_X1 U8535 ( .A1(n8238), .A2(n12472), .ZN(n8236) );
  INV_X1 U8536 ( .A(n10726), .ZN(n8205) );
  OR2_X1 U8537 ( .A1(n10649), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n10678) );
  OR2_X1 U8538 ( .A1(n10571), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n10708) );
  NAND2_X1 U8539 ( .A1(n13353), .A2(n13352), .ZN(n14035) );
  NOR3_X1 U8540 ( .A1(n14075), .A2(n7757), .A3(n14035), .ZN(n14036) );
  OR2_X1 U8541 ( .A1(n14075), .A2(n7757), .ZN(n14060) );
  AOI21_X1 U8542 ( .B1(n7200), .B2(n8091), .A(n7237), .ZN(n8088) );
  INV_X1 U8543 ( .A(n7825), .ZN(n7486) );
  NAND2_X1 U8544 ( .A1(n13056), .A2(n8092), .ZN(n7487) );
  XNOR2_X1 U8545 ( .A(n14098), .B(n14099), .ZN(n7672) );
  NAND2_X1 U8546 ( .A1(n14117), .A2(n13057), .ZN(n14098) );
  NAND2_X1 U8547 ( .A1(n13056), .A2(n13055), .ZN(n14115) );
  NAND2_X1 U8548 ( .A1(n13056), .A2(n8095), .ZN(n14117) );
  AOI21_X1 U8549 ( .B1(n8053), .B2(n8052), .A(n7242), .ZN(n8051) );
  NAND2_X1 U8550 ( .A1(n14175), .A2(n7357), .ZN(n7359) );
  INV_X1 U8551 ( .A(n8056), .ZN(n8052) );
  AND2_X1 U8552 ( .A1(n14180), .A2(n14172), .ZN(n14167) );
  NAND2_X1 U8553 ( .A1(n14167), .A2(n14152), .ZN(n14154) );
  NOR2_X1 U8554 ( .A1(n14317), .A2(n14216), .ZN(n14201) );
  NOR2_X1 U8555 ( .A1(n14332), .A2(n7761), .ZN(n7759) );
  OR2_X1 U8556 ( .A1(n10683), .A2(n10682), .ZN(n10700) );
  NAND2_X1 U8557 ( .A1(n10698), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10717) );
  INV_X1 U8558 ( .A(n10700), .ZN(n10698) );
  NAND2_X1 U8559 ( .A1(n12962), .A2(n7763), .ZN(n12994) );
  NOR2_X1 U8560 ( .A1(n12991), .A2(n7481), .ZN(n7480) );
  INV_X1 U8561 ( .A(n7484), .ZN(n7481) );
  NAND2_X1 U8562 ( .A1(n12962), .A2(n16183), .ZN(n12903) );
  INV_X1 U8563 ( .A(n10655), .ZN(n10654) );
  OR2_X1 U8564 ( .A1(n10637), .A2(n10423), .ZN(n10655) );
  NAND2_X1 U8565 ( .A1(n7491), .A2(n7490), .ZN(n12957) );
  NAND2_X1 U8566 ( .A1(n8070), .A2(n8071), .ZN(n12701) );
  NAND2_X1 U8567 ( .A1(n12581), .A2(n8074), .ZN(n8070) );
  OR2_X1 U8568 ( .A1(n10635), .A2(n12473), .ZN(n10637) );
  NAND2_X1 U8569 ( .A1(n8075), .A2(n8074), .ZN(n12700) );
  NOR2_X1 U8570 ( .A1(n12589), .A2(n13216), .ZN(n12588) );
  NAND2_X1 U8571 ( .A1(n7756), .A2(n7755), .ZN(n12589) );
  AOI21_X1 U8572 ( .B1(n8082), .B2(n12073), .A(n8081), .ZN(n8080) );
  INV_X1 U8573 ( .A(n12167), .ZN(n8081) );
  AND2_X1 U8574 ( .A1(n12184), .A2(n16063), .ZN(n12182) );
  NOR2_X1 U8575 ( .A1(n11949), .A2(n16043), .ZN(n12184) );
  AOI21_X1 U8576 ( .B1(n11942), .B2(n8068), .A(n7229), .ZN(n8067) );
  INV_X1 U8577 ( .A(n11774), .ZN(n8068) );
  INV_X1 U8578 ( .A(n11942), .ZN(n8069) );
  INV_X1 U8579 ( .A(n13410), .ZN(n11945) );
  NAND2_X1 U8580 ( .A1(n11716), .A2(n11676), .ZN(n11677) );
  XNOR2_X1 U8581 ( .A(n15995), .B(n14026), .ZN(n13405) );
  CLKBUF_X1 U8582 ( .A(n10941), .Z(n14302) );
  INV_X1 U8583 ( .A(n16182), .ZN(n14343) );
  AND2_X1 U8584 ( .A1(n10968), .A2(n12734), .ZN(n10959) );
  NAND2_X1 U8585 ( .A1(n8410), .A2(n8096), .ZN(n10416) );
  AND2_X1 U8586 ( .A1(n8098), .A2(n8232), .ZN(n8097) );
  INV_X1 U8587 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U8588 ( .A1(n10916), .A2(n10915), .ZN(n10918) );
  OR2_X1 U8589 ( .A1(n10486), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n10631) );
  AND2_X1 U8590 ( .A1(n10487), .A2(n10486), .ZN(n11070) );
  INV_X1 U8591 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8779) );
  INV_X1 U8592 ( .A(n14672), .ZN(n7381) );
  INV_X1 U8593 ( .A(n16173), .ZN(n8395) );
  OR2_X1 U8594 ( .A1(n8833), .A2(n8832), .ZN(n8852) );
  INV_X1 U8595 ( .A(n14766), .ZN(n11840) );
  OR2_X1 U8596 ( .A1(n12348), .A2(n12349), .ZN(n8393) );
  OR2_X1 U8597 ( .A1(n8762), .A2(n8761), .ZN(n8780) );
  NAND2_X1 U8598 ( .A1(n8898), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8899) );
  AND2_X1 U8599 ( .A1(n14707), .A2(n8366), .ZN(n8365) );
  NAND2_X1 U8600 ( .A1(n8372), .A2(n8367), .ZN(n8366) );
  OR2_X1 U8601 ( .A1(n8780), .A2(n8779), .ZN(n8801) );
  INV_X1 U8602 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U8603 ( .A1(n15162), .A2(n10042), .ZN(n11552) );
  AND4_X1 U8604 ( .A1(n8982), .A2(n8981), .A3(n8980), .A4(n8979), .ZN(n14594)
         );
  INV_X1 U8605 ( .A(n8976), .ZN(n10156) );
  INV_X1 U8606 ( .A(n8953), .ZN(n10157) );
  OR2_X1 U8607 ( .A1(n8953), .A2(n8556), .ZN(n8560) );
  OR2_X1 U8608 ( .A1(n11330), .A2(n11331), .ZN(n7783) );
  AND2_X1 U8609 ( .A1(n7783), .A2(n7782), .ZN(n14795) );
  NAND2_X1 U8610 ( .A1(n11528), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U8611 ( .A1(n14795), .A2(n14794), .ZN(n14793) );
  NAND2_X1 U8612 ( .A1(n14793), .A2(n7781), .ZN(n11525) );
  OR2_X1 U8613 ( .A1(n14805), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7781) );
  XNOR2_X1 U8614 ( .A(n12664), .B(n7793), .ZN(n12116) );
  OR2_X1 U8615 ( .A1(n11818), .A2(n11817), .ZN(n12112) );
  OR2_X1 U8616 ( .A1(n12873), .A2(n12872), .ZN(n7789) );
  NAND2_X1 U8617 ( .A1(n7789), .A2(n7788), .ZN(n7787) );
  NAND2_X1 U8618 ( .A1(n14814), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7788) );
  AND2_X1 U8619 ( .A1(n7787), .A2(n14826), .ZN(n14823) );
  AND2_X1 U8620 ( .A1(n8810), .A2(n8813), .ZN(n8394) );
  AOI21_X1 U8621 ( .B1(n8339), .B2(n13069), .A(n8965), .ZN(n8337) );
  AND2_X1 U8622 ( .A1(n14878), .A2(n14744), .ZN(n8965) );
  NAND2_X1 U8623 ( .A1(n7577), .A2(n7576), .ZN(n14867) );
  AOI21_X1 U8624 ( .B1(n7578), .B2(n7582), .A(n7205), .ZN(n7576) );
  NAND2_X1 U8625 ( .A1(n14895), .A2(n7578), .ZN(n7577) );
  NAND2_X1 U8626 ( .A1(n14383), .A2(n14595), .ZN(n8341) );
  AOI21_X1 U8627 ( .B1(n14587), .B2(n14878), .A(n9018), .ZN(n14871) );
  NOR2_X1 U8628 ( .A1(n14871), .A2(n8340), .ZN(n8339) );
  INV_X1 U8629 ( .A(n8341), .ZN(n8340) );
  AOI21_X2 U8630 ( .B1(n14883), .B2(n14884), .A(n7300), .ZN(n13074) );
  NAND2_X1 U8631 ( .A1(n7580), .A2(n7581), .ZN(n13070) );
  OR2_X1 U8632 ( .A1(n14895), .A2(n7582), .ZN(n7580) );
  INV_X1 U8633 ( .A(n8332), .ZN(n7666) );
  AOI21_X1 U8634 ( .B1(n8333), .B2(n10225), .A(n8920), .ZN(n8332) );
  INV_X1 U8635 ( .A(n8524), .ZN(n8914) );
  INV_X1 U8636 ( .A(n9017), .ZN(n8265) );
  NOR2_X1 U8637 ( .A1(n8271), .A2(n8267), .ZN(n8266) );
  OR2_X1 U8638 ( .A1(n9017), .A2(n8268), .ZN(n8267) );
  INV_X1 U8639 ( .A(n14916), .ZN(n8268) );
  NOR2_X1 U8640 ( .A1(n7225), .A2(n15077), .ZN(n14947) );
  AOI21_X1 U8641 ( .B1(n8326), .B2(n8328), .A(n8325), .ZN(n14961) );
  INV_X1 U8642 ( .A(n8327), .ZN(n8325) );
  AOI21_X1 U8643 ( .B1(n10222), .B2(n8328), .A(n8891), .ZN(n8327) );
  NAND2_X1 U8644 ( .A1(n8324), .A2(n8857), .ZN(n15022) );
  NOR2_X1 U8645 ( .A1(n15022), .A2(n15105), .ZN(n14992) );
  NOR2_X1 U8646 ( .A1(n15010), .A2(n15009), .ZN(n15008) );
  NAND2_X1 U8647 ( .A1(n8323), .A2(n7238), .ZN(n12936) );
  INV_X1 U8648 ( .A(n16199), .ZN(n7770) );
  NAND2_X1 U8649 ( .A1(n8323), .A2(n7771), .ZN(n12858) );
  INV_X1 U8650 ( .A(n16177), .ZN(n7774) );
  NAND2_X1 U8651 ( .A1(n8323), .A2(n8322), .ZN(n12634) );
  NOR2_X1 U8652 ( .A1(n14661), .A2(n14703), .ZN(n7776) );
  NOR2_X1 U8653 ( .A1(n12316), .A2(n14560), .ZN(n12394) );
  AND2_X1 U8654 ( .A1(n9004), .A2(n8699), .ZN(n12200) );
  NAND2_X1 U8655 ( .A1(n8319), .A2(n8318), .ZN(n12263) );
  NAND2_X1 U8656 ( .A1(n7779), .A2(n7778), .ZN(n12316) );
  NAND2_X1 U8657 ( .A1(n7585), .A2(n7584), .ZN(n12255) );
  AOI21_X1 U8658 ( .B1(n7586), .B2(n7588), .A(n7258), .ZN(n7585) );
  NAND2_X1 U8659 ( .A1(n7496), .A2(n8596), .ZN(n12288) );
  XNOR2_X1 U8660 ( .A(n12299), .B(n11840), .ZN(n12290) );
  INV_X1 U8661 ( .A(n8996), .ZN(n7564) );
  AND2_X1 U8662 ( .A1(n7562), .A2(n8997), .ZN(n7561) );
  INV_X1 U8663 ( .A(n14566), .ZN(n11825) );
  NAND2_X1 U8664 ( .A1(n12280), .A2(n11825), .ZN(n12293) );
  NAND2_X1 U8665 ( .A1(n7497), .A2(n8565), .ZN(n12269) );
  NAND2_X1 U8666 ( .A1(n15912), .A2(n10207), .ZN(n7497) );
  AND2_X1 U8667 ( .A1(n15978), .A2(n7780), .ZN(n12280) );
  NOR2_X1 U8668 ( .A1(n15914), .A2(n15917), .ZN(n7780) );
  NOR2_X1 U8669 ( .A1(n10037), .A2(n10036), .ZN(n15921) );
  OR2_X1 U8670 ( .A1(n12318), .A2(n14835), .ZN(n15927) );
  AOI21_X1 U8671 ( .B1(n9052), .B2(n9051), .A(n11029), .ZN(n11579) );
  INV_X1 U8672 ( .A(n14865), .ZN(n8278) );
  AND2_X1 U8673 ( .A1(n14939), .A2(n14947), .ZN(n15069) );
  NAND2_X1 U8674 ( .A1(n8742), .A2(n8741), .ZN(n14387) );
  INV_X1 U8675 ( .A(n16139), .ZN(n16015) );
  NOR2_X1 U8676 ( .A1(n11580), .A2(n11579), .ZN(n12152) );
  OR2_X1 U8677 ( .A1(n8992), .A2(n15162), .ZN(n15881) );
  NAND2_X1 U8678 ( .A1(n8109), .A2(n8108), .ZN(n10153) );
  AND2_X1 U8679 ( .A1(n8578), .A2(n8344), .ZN(n7500) );
  INV_X1 U8680 ( .A(n7504), .ZN(n7502) );
  XNOR2_X1 U8681 ( .A(n8967), .B(n8966), .ZN(n14374) );
  XNOR2_X1 U8682 ( .A(n8962), .B(n8485), .ZN(n13007) );
  NAND2_X1 U8683 ( .A1(n8139), .A2(n8138), .ZN(n8932) );
  NAND2_X1 U8684 ( .A1(n7214), .A2(n7299), .ZN(n8138) );
  AND2_X1 U8685 ( .A1(n8911), .A2(n8910), .ZN(n12607) );
  XNOR2_X1 U8686 ( .A(n8535), .B(n8534), .ZN(n12731) );
  XNOR2_X1 U8687 ( .A(n8530), .B(n15295), .ZN(n10788) );
  AND2_X1 U8688 ( .A1(n8895), .A2(n8894), .ZN(n12478) );
  NAND2_X1 U8689 ( .A1(n8984), .A2(n7863), .ZN(n8404) );
  NAND2_X1 U8690 ( .A1(n8118), .A2(n8123), .ZN(n8881) );
  NAND2_X1 U8691 ( .A1(n8839), .A2(n8462), .ZN(n8118) );
  INV_X1 U8692 ( .A(n8437), .ZN(n7809) );
  NAND2_X1 U8693 ( .A1(n8681), .A2(SI_9_), .ZN(n8702) );
  NAND2_X1 U8694 ( .A1(n8702), .A2(n7479), .ZN(n8684) );
  OR2_X1 U8695 ( .A1(n8681), .A2(SI_9_), .ZN(n7479) );
  AND2_X1 U8696 ( .A1(n8688), .A2(n8721), .ZN(n11334) );
  NAND2_X1 U8697 ( .A1(n8598), .A2(n8597), .ZN(n8600) );
  OR2_X1 U8698 ( .A1(n8592), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8602) );
  OAI211_X1 U8699 ( .C1(n8142), .C2(n7377), .A(n7376), .B(n7374), .ZN(n8572)
         );
  NAND2_X1 U8700 ( .A1(n8142), .A2(n7375), .ZN(n7374) );
  OAI21_X1 U8701 ( .B1(SI_1_), .B2(n8417), .A(n8420), .ZN(n8551) );
  OAI21_X1 U8702 ( .B1(n10342), .B2(n10346), .A(n7931), .ZN(n7930) );
  NAND2_X1 U8703 ( .A1(n10298), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7931) );
  XNOR2_X1 U8704 ( .A(n10337), .B(n7304), .ZN(n10338) );
  AOI21_X1 U8705 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n10314), .A(n10313), .ZN(
        n10369) );
  INV_X1 U8706 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7609) );
  OAI21_X1 U8707 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n10318), .A(n10317), .ZN(
        n10371) );
  AOI21_X1 U8708 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n10322), .A(n10321), .ZN(
        n10379) );
  NOR2_X1 U8709 ( .A1(n10375), .A2(n10374), .ZN(n10321) );
  NAND2_X1 U8710 ( .A1(n15584), .A2(n7603), .ZN(n7601) );
  OR2_X1 U8711 ( .A1(n15584), .A2(n7603), .ZN(n7602) );
  AND2_X1 U8712 ( .A1(n15587), .A2(n15589), .ZN(n10385) );
  OR2_X1 U8713 ( .A1(n11414), .A2(n11415), .ZN(n7676) );
  AOI21_X1 U8714 ( .B1(n8292), .B2(n13513), .A(n7274), .ZN(n8291) );
  NAND2_X1 U8715 ( .A1(n13527), .A2(n13095), .ZN(n13494) );
  NAND2_X1 U8716 ( .A1(n7508), .A2(n7511), .ZN(n13083) );
  OR2_X1 U8717 ( .A1(n12814), .A2(n8289), .ZN(n7508) );
  AND2_X1 U8718 ( .A1(n12358), .A2(n13581), .ZN(n7526) );
  AND3_X1 U8719 ( .A1(n9248), .A2(n9247), .A3(n9246), .ZN(n12379) );
  INV_X1 U8720 ( .A(n13566), .ZN(n13476) );
  NAND2_X1 U8721 ( .A1(n13093), .A2(n13092), .ZN(n13530) );
  AND4_X1 U8722 ( .A1(n9497), .A2(n9496), .A3(n9495), .A4(n9494), .ZN(n13676)
         );
  NAND2_X1 U8723 ( .A1(n12495), .A2(n7311), .ZN(n12614) );
  NOR2_X1 U8724 ( .A1(n11349), .A2(n11348), .ZN(n11353) );
  AND3_X1 U8725 ( .A1(n9435), .A2(n9434), .A3(n9433), .ZN(n13735) );
  NAND2_X1 U8726 ( .A1(n13510), .A2(n8296), .ZN(n13546) );
  NAND2_X1 U8727 ( .A1(n13510), .A2(n8292), .ZN(n13547) );
  NAND2_X1 U8728 ( .A1(n8284), .A2(n13114), .ZN(n13555) );
  NAND2_X1 U8729 ( .A1(n13501), .A2(n13502), .ZN(n8284) );
  NAND2_X1 U8730 ( .A1(n11242), .A2(n11241), .ZN(n13561) );
  OR2_X1 U8731 ( .A1(n11239), .A2(n11238), .ZN(n13551) );
  NAND2_X1 U8732 ( .A1(n12888), .A2(n12887), .ZN(n12889) );
  NAND2_X1 U8733 ( .A1(n12888), .A2(n8288), .ZN(n12985) );
  NAND2_X1 U8734 ( .A1(n11411), .A2(n12136), .ZN(n13564) );
  NAND2_X1 U8735 ( .A1(n9866), .A2(n11245), .ZN(n9867) );
  OR2_X1 U8736 ( .A1(n9866), .A2(n11664), .ZN(n8406) );
  AOI21_X1 U8737 ( .B1(n9865), .B2(n7681), .A(n9864), .ZN(n9866) );
  AND4_X1 U8738 ( .A1(n9686), .A2(n9685), .A3(n9684), .A4(n9683), .ZN(n13593)
         );
  AND4_X1 U8739 ( .A1(n9686), .A2(n9604), .A3(n9603), .A4(n9602), .ZN(n12033)
         );
  INV_X1 U8740 ( .A(n13627), .ZN(n13568) );
  INV_X1 U8741 ( .A(n13656), .ZN(n13569) );
  NAND2_X1 U8742 ( .A1(n9483), .A2(n9482), .ZN(n13688) );
  INV_X1 U8743 ( .A(n13735), .ZN(n13707) );
  INV_X1 U8744 ( .A(n12025), .ZN(n13583) );
  NAND2_X1 U8745 ( .A1(n7462), .A2(n9085), .ZN(n11410) );
  AND2_X1 U8746 ( .A1(n11386), .A2(n7746), .ZN(n11396) );
  NAND2_X1 U8747 ( .A1(n11410), .A2(n7747), .ZN(n7746) );
  INV_X1 U8748 ( .A(n9971), .ZN(n7747) );
  NOR2_X1 U8749 ( .A1(n7544), .A2(n9108), .ZN(n11391) );
  OAI22_X1 U8750 ( .A1(n9084), .A2(n7983), .B1(P3_IR_REG_2__SCAN_IN), .B2(
        P3_IR_REG_31__SCAN_IN), .ZN(n7544) );
  NAND2_X1 U8751 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7983) );
  NOR2_X1 U8752 ( .A1(n15652), .A2(n15651), .ZN(n15654) );
  OAI21_X1 U8753 ( .B1(n15621), .B2(n7464), .A(n7463), .ZN(n15638) );
  NAND2_X1 U8754 ( .A1(n7465), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7464) );
  INV_X1 U8755 ( .A(n9898), .ZN(n7466) );
  NOR2_X1 U8756 ( .A1(n9900), .A2(n7980), .ZN(n15658) );
  NAND2_X1 U8757 ( .A1(n7981), .A2(n7982), .ZN(n15659) );
  NOR2_X1 U8758 ( .A1(n15677), .A2(n15676), .ZN(n15675) );
  AND2_X1 U8759 ( .A1(n7981), .A2(n7980), .ZN(n15677) );
  OAI21_X1 U8760 ( .B1(n15682), .B2(n15678), .A(n15679), .ZN(n11612) );
  NAND2_X1 U8761 ( .A1(n11615), .A2(n9942), .ZN(n11757) );
  NAND2_X1 U8762 ( .A1(n11757), .A2(n11758), .ZN(n11756) );
  INV_X1 U8763 ( .A(n7470), .ZN(n11761) );
  XNOR2_X1 U8764 ( .A(n9905), .B(n9904), .ZN(n12054) );
  XNOR2_X1 U8765 ( .A(n9943), .B(n9904), .ZN(n12056) );
  NOR2_X1 U8766 ( .A1(n12054), .A2(n12053), .ZN(n12052) );
  OAI21_X1 U8767 ( .B1(n12054), .B2(n7977), .A(n7976), .ZN(n15694) );
  NAND2_X1 U8768 ( .A1(n7978), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U8769 ( .A1(n9906), .A2(n7978), .ZN(n7976) );
  INV_X1 U8770 ( .A(n15695), .ZN(n7978) );
  XNOR2_X1 U8771 ( .A(n9908), .B(n10015), .ZN(n15711) );
  AND2_X1 U8772 ( .A1(n7743), .A2(n7302), .ZN(n15750) );
  INV_X1 U8773 ( .A(n7468), .ZN(n9913) );
  NAND2_X1 U8774 ( .A1(n7738), .A2(n7739), .ZN(n15776) );
  XNOR2_X1 U8775 ( .A(n7975), .B(n15789), .ZN(n15783) );
  NOR2_X1 U8776 ( .A1(n15784), .A2(n15783), .ZN(n15782) );
  NOR2_X1 U8777 ( .A1(n9919), .A2(n15782), .ZN(n15809) );
  AND2_X1 U8778 ( .A1(n9368), .A2(n9367), .ZN(n9388) );
  XNOR2_X1 U8779 ( .A(n9921), .B(n9956), .ZN(n15815) );
  INV_X1 U8780 ( .A(n7751), .ZN(n15823) );
  INV_X1 U8781 ( .A(n9967), .ZN(n7967) );
  NAND2_X1 U8782 ( .A1(n8001), .A2(n8002), .ZN(n9699) );
  INV_X1 U8783 ( .A(n8003), .ZN(n8002) );
  OAI21_X1 U8784 ( .B1(n9877), .B2(n7879), .A(n8004), .ZN(n7878) );
  NOR3_X1 U8785 ( .A1(n9622), .A2(n7881), .A3(n9877), .ZN(n7877) );
  OAI21_X1 U8786 ( .B1(n13609), .B2(n8175), .A(n13612), .ZN(n13763) );
  OAI21_X1 U8787 ( .B1(n9883), .B2(n15959), .A(n9882), .ZN(n13622) );
  AOI21_X1 U8788 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(n9882) );
  NOR2_X1 U8789 ( .A1(n13115), .A2(n15960), .ZN(n9879) );
  NAND2_X1 U8790 ( .A1(n9622), .A2(n9621), .ZN(n13629) );
  NAND2_X1 U8791 ( .A1(n13651), .A2(n7196), .ZN(n13638) );
  NAND2_X1 U8792 ( .A1(n13686), .A2(n13097), .ZN(n13677) );
  NAND2_X1 U8793 ( .A1(n9460), .A2(n9459), .ZN(n13697) );
  OAI21_X1 U8794 ( .B1(n13738), .B2(n7906), .A(n7904), .ZN(n13703) );
  NAND2_X1 U8795 ( .A1(n13736), .A2(n9830), .ZN(n13723) );
  OAI21_X1 U8796 ( .B1(n12976), .B2(n9719), .A(n7988), .ZN(n13751) );
  NAND2_X1 U8797 ( .A1(n13014), .A2(n9380), .ZN(n13744) );
  NAND2_X1 U8798 ( .A1(n13018), .A2(n13017), .ZN(n13016) );
  NAND2_X1 U8799 ( .A1(n12976), .A2(n9817), .ZN(n13018) );
  NAND2_X1 U8800 ( .A1(n12745), .A2(n9752), .ZN(n12794) );
  NAND2_X1 U8801 ( .A1(n7888), .A2(n7891), .ZN(n12450) );
  NAND2_X1 U8802 ( .A1(n12229), .A2(n7894), .ZN(n7888) );
  NAND2_X1 U8803 ( .A1(n7895), .A2(n9711), .ZN(n12507) );
  NAND2_X1 U8804 ( .A1(n7896), .A2(n7897), .ZN(n7895) );
  AND3_X1 U8805 ( .A1(n9268), .A2(n9267), .A3(n9266), .ZN(n12516) );
  NAND2_X1 U8806 ( .A1(n11668), .A2(n15966), .ZN(n13754) );
  NAND2_X1 U8807 ( .A1(n11902), .A2(n9213), .ZN(n12211) );
  NAND2_X1 U8808 ( .A1(n11892), .A2(n9156), .ZN(n11883) );
  NAND2_X1 U8809 ( .A1(n15954), .A2(n9760), .ZN(n11956) );
  OR2_X1 U8810 ( .A1(n11665), .A2(n11664), .ZN(n15967) );
  INV_X1 U8811 ( .A(n13596), .ZN(n13824) );
  AOI21_X1 U8812 ( .B1(n13762), .B2(n16160), .A(n13763), .ZN(n13825) );
  INV_X1 U8813 ( .A(n13505), .ZN(n13836) );
  INV_X1 U8814 ( .A(n13522), .ZN(n13840) );
  INV_X1 U8815 ( .A(n13474), .ZN(n13844) );
  INV_X1 U8816 ( .A(n13539), .ZN(n13848) );
  INV_X1 U8817 ( .A(n13532), .ZN(n13856) );
  INV_X1 U8818 ( .A(n15908), .ZN(n11538) );
  AND2_X1 U8819 ( .A1(n9640), .A2(n9639), .ZN(n13869) );
  NAND2_X1 U8820 ( .A1(n7636), .A2(n7635), .ZN(n9681) );
  INV_X1 U8821 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13872) );
  NOR2_X1 U8822 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), .ZN(
        n7871) );
  NAND2_X1 U8823 ( .A1(n7637), .A2(n9678), .ZN(n9689) );
  XNOR2_X1 U8824 ( .A(n9677), .B(n9675), .ZN(n13879) );
  INV_X1 U8825 ( .A(SI_28_), .ZN(n15177) );
  NAND2_X1 U8826 ( .A1(n8010), .A2(n8009), .ZN(n8148) );
  NOR2_X1 U8827 ( .A1(n9369), .A2(n8149), .ZN(n8009) );
  NAND2_X1 U8828 ( .A1(n7663), .A2(n7662), .ZN(n9568) );
  INV_X1 U8829 ( .A(n9566), .ZN(n7662) );
  INV_X1 U8830 ( .A(SI_27_), .ZN(n15283) );
  NAND2_X1 U8831 ( .A1(n9534), .A2(n7658), .ZN(n8036) );
  NOR2_X1 U8832 ( .A1(n9534), .A2(n7658), .ZN(n8035) );
  NAND2_X1 U8833 ( .A1(n8029), .A2(n9534), .ZN(n8033) );
  OR2_X1 U8834 ( .A1(n9519), .A2(n9518), .ZN(n9520) );
  NAND2_X1 U8835 ( .A1(n9515), .A2(n9503), .ZN(n9514) );
  NAND2_X1 U8836 ( .A1(n9633), .A2(n7220), .ZN(n12562) );
  NAND2_X1 U8837 ( .A1(n9488), .A2(n9487), .ZN(n9500) );
  XNOR2_X1 U8838 ( .A(n9593), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12000) );
  OAI211_X1 U8839 ( .C1(n9594), .C2(n7523), .A(n9644), .B(n7522), .ZN(n11967)
         );
  NAND2_X1 U8840 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n7523) );
  NAND2_X1 U8841 ( .A1(n9592), .A2(n9369), .ZN(n7522) );
  INV_X1 U8842 ( .A(SI_20_), .ZN(n11731) );
  XNOR2_X1 U8843 ( .A(n9597), .B(n9596), .ZN(n11732) );
  NAND2_X1 U8844 ( .A1(n9453), .A2(n9442), .ZN(n9443) );
  INV_X1 U8845 ( .A(SI_19_), .ZN(n15192) );
  INV_X1 U8846 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9423) );
  OAI21_X1 U8847 ( .B1(n9422), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9424) );
  INV_X1 U8848 ( .A(SI_18_), .ZN(n11424) );
  NAND2_X1 U8849 ( .A1(n9403), .A2(n9402), .ZN(n9417) );
  NAND2_X1 U8850 ( .A1(n9400), .A2(n9399), .ZN(n9403) );
  INV_X1 U8851 ( .A(SI_17_), .ZN(n15275) );
  OAI21_X1 U8852 ( .B1(n9346), .B2(n8024), .A(n8022), .ZN(n9382) );
  NAND2_X1 U8853 ( .A1(n9362), .A2(n9361), .ZN(n9365) );
  INV_X1 U8854 ( .A(SI_14_), .ZN(n11037) );
  NAND2_X1 U8855 ( .A1(n9327), .A2(n9310), .ZN(n9311) );
  NAND2_X1 U8856 ( .A1(n9302), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9313) );
  INV_X1 U8857 ( .A(SI_12_), .ZN(n15307) );
  NAND2_X1 U8858 ( .A1(n9298), .A2(n9297), .ZN(n9307) );
  NAND2_X1 U8859 ( .A1(n7655), .A2(n8016), .ZN(n9298) );
  INV_X1 U8860 ( .A(n9064), .ZN(n9300) );
  INV_X1 U8861 ( .A(SI_11_), .ZN(n15313) );
  NAND2_X1 U8862 ( .A1(n9280), .A2(n9279), .ZN(n9295) );
  NAND2_X1 U8863 ( .A1(n9277), .A2(n9276), .ZN(n9280) );
  INV_X1 U8864 ( .A(n10005), .ZN(n11760) );
  NAND2_X1 U8865 ( .A1(n9223), .A2(n9222), .ZN(n9226) );
  NAND2_X1 U8866 ( .A1(n7644), .A2(n9167), .ZN(n9186) );
  NAND2_X1 U8867 ( .A1(n9166), .A2(n9165), .ZN(n7644) );
  INV_X1 U8868 ( .A(n9980), .ZN(n15630) );
  OR2_X1 U8869 ( .A1(n10968), .A2(n10967), .ZN(n11057) );
  NAND2_X1 U8870 ( .A1(n13989), .A2(n10872), .ZN(n13885) );
  NOR2_X1 U8871 ( .A1(n8227), .A2(n8225), .ZN(n12737) );
  NAND2_X1 U8872 ( .A1(n8224), .A2(n12597), .ZN(n12738) );
  INV_X1 U8873 ( .A(n8227), .ZN(n8224) );
  INV_X1 U8874 ( .A(n10563), .ZN(n10518) );
  NAND2_X1 U8875 ( .A1(n13926), .A2(n8201), .ZN(n7431) );
  NAND2_X1 U8876 ( .A1(n13958), .A2(n10772), .ZN(n13912) );
  XNOR2_X1 U8877 ( .A(n10849), .B(n10850), .ZN(n13920) );
  NAND2_X1 U8878 ( .A1(n13902), .A2(n10822), .ZN(n13949) );
  INV_X1 U8879 ( .A(n14021), .ZN(n12169) );
  NAND2_X1 U8880 ( .A1(n11054), .A2(n14379), .ZN(n10528) );
  OR2_X1 U8881 ( .A1(n12138), .A2(n8236), .ZN(n12549) );
  INV_X1 U8882 ( .A(n8238), .ZN(n8237) );
  NAND2_X1 U8883 ( .A1(n8207), .A2(n8208), .ZN(n13980) );
  OR2_X1 U8884 ( .A1(n13926), .A2(n8209), .ZN(n8207) );
  NAND2_X1 U8885 ( .A1(n10604), .A2(n10603), .ZN(n11638) );
  OAI21_X1 U8886 ( .B1(n11484), .B2(n7411), .A(n7413), .ZN(n11637) );
  AOI21_X1 U8887 ( .B1(n7417), .B2(n11483), .A(n7416), .ZN(n7413) );
  AND2_X1 U8888 ( .A1(n10848), .A2(n10847), .ZN(n14118) );
  NAND2_X1 U8889 ( .A1(n10856), .A2(n10855), .ZN(n14278) );
  OAI21_X1 U8890 ( .B1(n8220), .B2(n8225), .A(n8221), .ZN(n8231) );
  INV_X1 U8891 ( .A(n12600), .ZN(n8220) );
  NAND2_X1 U8892 ( .A1(n10415), .A2(n10430), .ZN(n10432) );
  INV_X1 U8893 ( .A(n14118), .ZN(n14090) );
  NAND2_X1 U8894 ( .A1(n10552), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10555) );
  NAND2_X1 U8895 ( .A1(n10552), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10533) );
  CLKBUF_X2 U8896 ( .A(P2_U3947), .Z(n15405) );
  INV_X1 U8897 ( .A(n14035), .ZN(n14258) );
  AOI21_X1 U8898 ( .B1(n14053), .B2(n14236), .A(n14052), .ZN(n14263) );
  OR2_X1 U8899 ( .A1(n14267), .A2(n14054), .ZN(n14055) );
  NAND2_X1 U8900 ( .A1(n13323), .A2(n13322), .ZN(n14260) );
  AND2_X1 U8901 ( .A1(n8060), .A2(n7301), .ZN(n14073) );
  AND2_X1 U8902 ( .A1(n10894), .A2(n10878), .ZN(n13887) );
  OAI21_X1 U8903 ( .B1(n7489), .B2(n14214), .A(n13062), .ZN(n7488) );
  XNOR2_X1 U8904 ( .A(n14043), .B(n13433), .ZN(n7489) );
  AND2_X1 U8905 ( .A1(n10842), .A2(n10841), .ZN(n14108) );
  NAND2_X1 U8906 ( .A1(n7671), .A2(n7669), .ZN(n14283) );
  INV_X1 U8907 ( .A(n7670), .ZN(n7669) );
  NAND2_X1 U8908 ( .A1(n7672), .A2(n14236), .ZN(n7671) );
  OAI22_X1 U8909 ( .A1(n14101), .A2(n14191), .B1(n14189), .B2(n14100), .ZN(
        n7670) );
  NAND2_X1 U8910 ( .A1(n14113), .A2(n13037), .ZN(n14097) );
  AND2_X1 U8911 ( .A1(n14113), .A2(n14112), .ZN(n14288) );
  NAND2_X1 U8912 ( .A1(n8055), .A2(n8059), .ZN(n14150) );
  NAND2_X1 U8913 ( .A1(n8055), .A2(n8053), .ZN(n14300) );
  NAND2_X1 U8914 ( .A1(n7810), .A2(n7812), .ZN(n14143) );
  NAND2_X1 U8915 ( .A1(n7811), .A2(n7815), .ZN(n14164) );
  NAND2_X1 U8916 ( .A1(n14188), .A2(n7816), .ZN(n7811) );
  NAND2_X1 U8917 ( .A1(n13034), .A2(n13033), .ZN(n14162) );
  NAND2_X1 U8918 ( .A1(n7818), .A2(n13050), .ZN(n14176) );
  OR2_X1 U8919 ( .A1(n14188), .A2(n13048), .ZN(n7818) );
  NAND2_X1 U8920 ( .A1(n8050), .A2(n13029), .ZN(n14193) );
  NAND2_X1 U8921 ( .A1(n12992), .A2(n12991), .ZN(n8047) );
  NAND2_X1 U8922 ( .A1(n10681), .A2(n10680), .ZN(n14342) );
  NAND2_X1 U8923 ( .A1(n12959), .A2(n12823), .ZN(n12900) );
  NAND2_X1 U8924 ( .A1(n8062), .A2(n12828), .ZN(n12954) );
  NAND2_X1 U8925 ( .A1(n12704), .A2(n12703), .ZN(n12826) );
  NAND2_X1 U8926 ( .A1(n12582), .A2(n12527), .ZN(n12530) );
  NAND2_X1 U8927 ( .A1(n10634), .A2(n10633), .ZN(n13224) );
  OR2_X1 U8928 ( .A1(n11041), .A2(n7191), .ZN(n10476) );
  NAND2_X1 U8929 ( .A1(n12180), .A2(n12078), .ZN(n12080) );
  NAND2_X1 U8930 ( .A1(n8084), .A2(n8082), .ZN(n12168) );
  AND2_X1 U8931 ( .A1(n16041), .A2(n12082), .ZN(n14151) );
  NAND2_X1 U8932 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  INV_X1 U8933 ( .A(n16045), .ZN(n16150) );
  INV_X1 U8934 ( .A(n10547), .ZN(n10549) );
  OR2_X1 U8935 ( .A1(n7191), .A2(n11022), .ZN(n10548) );
  OR2_X1 U8936 ( .A1(n11700), .A2(n10458), .ZN(n16045) );
  NAND2_X2 U8937 ( .A1(n7219), .A2(n7427), .ZN(n13143) );
  OR2_X1 U8938 ( .A1(n11054), .A2(n11059), .ZN(n7767) );
  AND2_X1 U8939 ( .A1(n16041), .A2(n11699), .ZN(n16147) );
  AND2_X1 U8940 ( .A1(n10959), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15409) );
  NAND2_X1 U8941 ( .A1(n10934), .A2(n10933), .ZN(n15408) );
  XNOR2_X1 U8942 ( .A(n10914), .B(P2_IR_REG_26__SCAN_IN), .ZN(n12802) );
  NAND2_X1 U8943 ( .A1(n10918), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10914) );
  INV_X1 U8944 ( .A(n13445), .ZN(n13452) );
  NAND2_X1 U8945 ( .A1(n10440), .A2(n10439), .ZN(n10444) );
  NOR2_X1 U8946 ( .A1(n10415), .A2(n10441), .ZN(n10439) );
  INV_X1 U8947 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11521) );
  INV_X1 U8948 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n11187) );
  INV_X1 U8949 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n11042) );
  INV_X1 U8950 ( .A(n11193), .ZN(n11277) );
  INV_X1 U8951 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n11039) );
  INV_X1 U8952 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n11025) );
  INV_X1 U8953 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n11017) );
  INV_X1 U8954 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10993) );
  INV_X1 U8955 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10983) );
  INV_X1 U8956 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10982) );
  INV_X1 U8957 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10989) );
  INV_X1 U8958 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9053) );
  OAI21_X1 U8959 ( .B1(n7217), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9054) );
  INV_X1 U8960 ( .A(n8353), .ZN(n7392) );
  NAND2_X1 U8961 ( .A1(n8356), .A2(n11838), .ZN(n7390) );
  NAND2_X1 U8962 ( .A1(n14546), .A2(n14504), .ZN(n14549) );
  OAI22_X1 U8963 ( .A1(n12348), .A2(n8389), .B1(n8388), .B2(n7262), .ZN(n14555) );
  INV_X1 U8964 ( .A(n8391), .ZN(n8388) );
  NAND2_X1 U8965 ( .A1(n8391), .A2(n8390), .ZN(n8389) );
  NAND2_X1 U8966 ( .A1(n14621), .A2(n14525), .ZN(n14719) );
  NAND2_X1 U8967 ( .A1(n14593), .A2(n8378), .ZN(n8377) );
  INV_X1 U8968 ( .A(n8381), .ZN(n8378) );
  NAND2_X1 U8969 ( .A1(n8380), .A2(n14593), .ZN(n8379) );
  NAND2_X1 U8970 ( .A1(n12346), .A2(n7388), .ZN(n12348) );
  NAND2_X1 U8971 ( .A1(n12345), .A2(n7389), .ZN(n7388) );
  INV_X1 U8972 ( .A(n12347), .ZN(n7389) );
  INV_X1 U8973 ( .A(n15086), .ZN(n14967) );
  NAND2_X1 U8974 ( .A1(n7387), .A2(n7386), .ZN(n7385) );
  INV_X1 U8975 ( .A(n14610), .ZN(n7387) );
  INV_X1 U8976 ( .A(n14611), .ZN(n7386) );
  NAND2_X1 U8977 ( .A1(n16193), .A2(n16194), .ZN(n14632) );
  NAND2_X1 U8978 ( .A1(n8362), .A2(n11911), .ZN(n12005) );
  NAND2_X1 U8979 ( .A1(n8369), .A2(n8370), .ZN(n14631) );
  NAND2_X1 U8980 ( .A1(n16193), .A2(n8371), .ZN(n8369) );
  INV_X1 U8981 ( .A(n7394), .ZN(n7393) );
  OAI21_X1 U8982 ( .B1(n14504), .B2(n7395), .A(n14644), .ZN(n7394) );
  INV_X1 U8983 ( .A(n14646), .ZN(n7395) );
  INV_X1 U8984 ( .A(n7382), .ZN(n14673) );
  NAND2_X1 U8985 ( .A1(n14600), .A2(n14489), .ZN(n14683) );
  OAI22_X1 U8986 ( .A1(n14555), .A2(n14554), .B1(n14405), .B2(n14404), .ZN(
        n14694) );
  INV_X1 U8987 ( .A(n14740), .ZN(n16195) );
  NAND2_X1 U8988 ( .A1(n8357), .A2(n8360), .ZN(n12091) );
  NAND2_X1 U8989 ( .A1(n7341), .A2(n8362), .ZN(n8357) );
  AND2_X1 U8990 ( .A1(n11557), .A2(n11846), .ZN(n11561) );
  AND3_X1 U8991 ( .A1(n7558), .A2(n10267), .A3(n7288), .ZN(n10284) );
  NAND4_X1 U8992 ( .A1(n8629), .A2(n8628), .A3(n8627), .A4(n8626), .ZN(n14765)
         );
  NOR2_X1 U8993 ( .A1(n11290), .A2(n7785), .ZN(n11312) );
  AND2_X1 U8994 ( .A1(n11295), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U8995 ( .A1(n11312), .A2(n11311), .ZN(n11310) );
  NAND2_X1 U8996 ( .A1(n11310), .A2(n7784), .ZN(n11292) );
  NAND2_X1 U8997 ( .A1(n11321), .A2(n11291), .ZN(n7784) );
  NAND2_X1 U8998 ( .A1(n11292), .A2(n11293), .ZN(n11329) );
  INV_X1 U8999 ( .A(n7783), .ZN(n11523) );
  NOR2_X1 U9000 ( .A1(n11812), .A2(n11813), .ZN(n12114) );
  NAND2_X1 U9001 ( .A1(n11811), .A2(n7795), .ZN(n11812) );
  OR2_X1 U9002 ( .A1(n11815), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7795) );
  OR2_X1 U9003 ( .A1(n12116), .A2(n12773), .ZN(n12663) );
  NAND2_X1 U9004 ( .A1(n15531), .A2(n8798), .ZN(n15530) );
  INV_X1 U9005 ( .A(n7789), .ZN(n14813) );
  NOR2_X1 U9006 ( .A1(n14823), .A2(n7786), .ZN(n14817) );
  NOR2_X1 U9007 ( .A1(n7787), .A2(n14826), .ZN(n7786) );
  NAND2_X1 U9008 ( .A1(n10173), .A2(n10172), .ZN(n14848) );
  AOI211_X1 U9009 ( .C1(n9026), .C2(n10181), .A(n14845), .B(n16077), .ZN(
        n14861) );
  OR2_X1 U9010 ( .A1(n14874), .A2(n14873), .ZN(n15038) );
  AOI22_X1 U9011 ( .A1(n7524), .A2(n14871), .B1(n13072), .B2(n8339), .ZN(
        n15040) );
  NAND2_X1 U9012 ( .A1(n13072), .A2(n8341), .ZN(n7524) );
  NAND2_X1 U9013 ( .A1(n8924), .A2(n8923), .ZN(n15055) );
  NAND2_X1 U9014 ( .A1(n14931), .A2(n8334), .ZN(n14911) );
  AOI21_X1 U9015 ( .B1(n14944), .B2(n14954), .A(n8273), .ZN(n14930) );
  NAND2_X1 U9016 ( .A1(n8269), .A2(n8270), .ZN(n14929) );
  NAND2_X1 U9017 ( .A1(n7571), .A2(n7570), .ZN(n14962) );
  AND2_X1 U9018 ( .A1(n8249), .A2(n9016), .ZN(n7570) );
  NAND2_X1 U9019 ( .A1(n14989), .A2(n8879), .ZN(n14978) );
  AND2_X1 U9020 ( .A1(n14989), .A2(n8328), .ZN(n14977) );
  NAND2_X1 U9021 ( .A1(n8251), .A2(n8247), .ZN(n14976) );
  AND2_X1 U9022 ( .A1(n7571), .A2(n8249), .ZN(n14975) );
  NAND2_X1 U9023 ( .A1(n8246), .A2(n8252), .ZN(n8251) );
  NAND2_X1 U9024 ( .A1(n12932), .A2(n8838), .ZN(n15005) );
  INV_X1 U9025 ( .A(n8324), .ZN(n15118) );
  INV_X1 U9026 ( .A(n7593), .ZN(n12935) );
  AOI21_X1 U9027 ( .B1(n7597), .B2(n7595), .A(n7594), .ZN(n7593) );
  INV_X1 U9028 ( .A(n7598), .ZN(n7594) );
  NAND2_X1 U9029 ( .A1(n8263), .A2(n8788), .ZN(n8260) );
  NAND2_X1 U9030 ( .A1(n12629), .A2(n8263), .ZN(n8261) );
  NAND2_X1 U9031 ( .A1(n8264), .A2(n9011), .ZN(n12687) );
  OR2_X1 U9032 ( .A1(n12629), .A2(n8788), .ZN(n8264) );
  NAND2_X1 U9033 ( .A1(n12482), .A2(n8770), .ZN(n12632) );
  NAND2_X1 U9034 ( .A1(n12400), .A2(n8736), .ZN(n12456) );
  NAND2_X1 U9035 ( .A1(n12313), .A2(n8718), .ZN(n12402) );
  INV_X1 U9036 ( .A(n14974), .ZN(n15001) );
  NAND2_X1 U9037 ( .A1(n11802), .A2(n9001), .ZN(n12126) );
  NAND2_X1 U9038 ( .A1(n12274), .A2(n8995), .ZN(n11585) );
  INV_X1 U9039 ( .A(n15933), .ZN(n15026) );
  INV_X1 U9040 ( .A(n12281), .ZN(n15978) );
  OR2_X1 U9041 ( .A1(n15894), .A2(n12154), .ZN(n15933) );
  INV_X1 U9042 ( .A(n14958), .ZN(n15936) );
  AOI21_X1 U9043 ( .B1(n15041), .B2(n7680), .A(n7679), .ZN(n7695) );
  INV_X1 U9044 ( .A(n15044), .ZN(n7679) );
  INV_X1 U9045 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U9046 ( .A1(n7575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8508) );
  NOR2_X1 U9047 ( .A1(n8493), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n8321) );
  XNOR2_X1 U9048 ( .A(n9039), .B(P1_IR_REG_26__SCAN_IN), .ZN(n12804) );
  XNOR2_X1 U9049 ( .A(n9032), .B(P1_IR_REG_25__SCAN_IN), .ZN(n12649) );
  NAND2_X1 U9050 ( .A1(n9035), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9032) );
  AND2_X1 U9051 ( .A1(n9036), .A2(n9035), .ZN(n12608) );
  INV_X1 U9053 ( .A(n14835), .ZN(n12471) );
  INV_X1 U9054 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11861) );
  INV_X1 U9055 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U9056 ( .A1(n8792), .A2(n7197), .ZN(n8811) );
  INV_X1 U9057 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11519) );
  NAND2_X1 U9058 ( .A1(n8126), .A2(n8128), .ZN(n8753) );
  INV_X1 U9059 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n11188) );
  INV_X1 U9060 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n11044) );
  INV_X1 U9061 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n11040) );
  INV_X1 U9062 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n11026) );
  OR2_X1 U9063 ( .A1(n8666), .A2(n8665), .ZN(n8667) );
  INV_X1 U9064 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U9065 ( .A1(n8649), .A2(n8648), .ZN(n8650) );
  NAND2_X1 U9066 ( .A1(n8634), .A2(n8431), .ZN(n8649) );
  INV_X1 U9067 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10994) );
  NAND2_X1 U9068 ( .A1(n8633), .A2(n8634), .ZN(n10995) );
  AOI21_X1 U9069 ( .B1(n8597), .B2(n8105), .A(n8104), .ZN(n8102) );
  NAND2_X1 U9070 ( .A1(n8576), .A2(n7790), .ZN(n11147) );
  AOI22_X1 U9071 ( .A1(n7281), .A2(n15398), .B1(n7792), .B2(n7791), .ZN(n7790)
         );
  INV_X1 U9072 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7792) );
  CLKBUF_X1 U9073 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n15398) );
  NOR2_X1 U9074 ( .A1(n10348), .A2(n15606), .ZN(n15546) );
  INV_X1 U9075 ( .A(n10350), .ZN(n7912) );
  NOR2_X1 U9076 ( .A1(n15561), .A2(n10367), .ZN(n15566) );
  INV_X1 U9077 ( .A(n7910), .ZN(n10365) );
  NOR2_X1 U9078 ( .A1(n15566), .A2(n15565), .ZN(n15564) );
  NAND2_X1 U9079 ( .A1(n7607), .A2(n7606), .ZN(n15574) );
  NAND2_X1 U9080 ( .A1(n15570), .A2(n7609), .ZN(n7606) );
  NAND2_X1 U9081 ( .A1(n15569), .A2(n7608), .ZN(n7607) );
  OR2_X1 U9082 ( .A1(n15570), .A2(n7609), .ZN(n7608) );
  NOR2_X1 U9083 ( .A1(n15574), .A2(n15573), .ZN(n15572) );
  NAND2_X1 U9084 ( .A1(n15576), .A2(n10378), .ZN(n15581) );
  NAND2_X1 U9085 ( .A1(n7600), .A2(n7599), .ZN(n15590) );
  AND2_X1 U9086 ( .A1(n10384), .A2(n7601), .ZN(n7599) );
  NOR2_X1 U9087 ( .A1(n10385), .A2(n10386), .ZN(n15593) );
  NAND2_X1 U9088 ( .A1(n10385), .A2(n10386), .ZN(n15595) );
  NAND2_X1 U9089 ( .A1(n15595), .A2(n15596), .ZN(n15592) );
  AND2_X1 U9090 ( .A1(n13870), .A2(n9895), .ZN(P3_U3897) );
  INV_X1 U9091 ( .A(n7969), .ZN(n15726) );
  AOI21_X1 U9092 ( .B1(n10034), .B2(n15844), .A(n7534), .ZN(n7533) );
  OAI21_X1 U9093 ( .B1(n13825), .B2(n9674), .A(n7898), .ZN(P3_U3487) );
  AOI21_X1 U9094 ( .B1(n13123), .B2(n7900), .A(n7899), .ZN(n7898) );
  NOR2_X1 U9095 ( .A1(n16165), .A2(n13764), .ZN(n7899) );
  INV_X1 U9096 ( .A(n13806), .ZN(n7900) );
  OAI21_X1 U9097 ( .B1(n13601), .B2(n13864), .A(n10402), .ZN(n10403) );
  NAND2_X1 U9098 ( .A1(n7415), .A2(n11483), .ZN(n11488) );
  XNOR2_X1 U9099 ( .A(n7686), .B(n7685), .ZN(n14542) );
  OAI21_X1 U9100 ( .B1(n14836), .B2(n14835), .A(n7796), .ZN(P1_U3262) );
  AOI21_X1 U9101 ( .B1(n7798), .B2(n14835), .A(n7797), .ZN(n7796) );
  OAI21_X1 U9102 ( .B1(n15876), .B2(n8107), .A(n14837), .ZN(n7797) );
  INV_X1 U9103 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8275) );
  NOR2_X1 U9104 ( .A1(n15604), .A2(n15603), .ZN(n15602) );
  AND2_X1 U9105 ( .A1(n7230), .A2(n7915), .ZN(n15604) );
  INV_X1 U9106 ( .A(n7911), .ZN(n15558) );
  NOR2_X1 U9107 ( .A1(n15569), .A2(n15570), .ZN(n15568) );
  NAND2_X1 U9108 ( .A1(n15585), .A2(n15584), .ZN(n15583) );
  NAND2_X1 U9109 ( .A1(n7927), .A2(n7616), .ZN(n7668) );
  NAND2_X1 U9110 ( .A1(n15601), .A2(n15600), .ZN(n7616) );
  XNOR2_X1 U9111 ( .A(n7926), .B(n7925), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9112 ( .A(n10400), .B(n7350), .ZN(n7925) );
  NAND2_X1 U9113 ( .A1(n7928), .A2(n7927), .ZN(n7926) );
  AND2_X1 U9114 ( .A1(n7713), .A2(n7712), .ZN(n7194) );
  AND2_X1 U9115 ( .A1(n10144), .A2(n10146), .ZN(n7195) );
  AND2_X1 U9116 ( .A1(n7398), .A2(n7399), .ZN(n16193) );
  AND2_X1 U9117 ( .A1(n13639), .A2(n9513), .ZN(n7196) );
  INV_X1 U9118 ( .A(n14979), .ZN(n8250) );
  AND4_X1 U9119 ( .A1(n8489), .A2(n8486), .A3(n8488), .A4(n8487), .ZN(n7197)
         );
  AND3_X1 U9120 ( .A1(n9060), .A2(n7865), .A3(n7864), .ZN(n7198) );
  INV_X1 U9121 ( .A(n15639), .ZN(n7465) );
  NAND2_X1 U9122 ( .A1(n15047), .A2(n14531), .ZN(n7199) );
  AND2_X1 U9123 ( .A1(n14042), .A2(n8090), .ZN(n7200) );
  NOR2_X1 U9124 ( .A1(n8185), .A2(n7735), .ZN(n7201) );
  NAND2_X1 U9125 ( .A1(n10784), .A2(n10783), .ZN(n14309) );
  INV_X1 U9126 ( .A(n10225), .ZN(n14932) );
  INV_X1 U9127 ( .A(n13513), .ZN(n8294) );
  AND2_X1 U9128 ( .A1(n15163), .A2(n8563), .ZN(n15077) );
  OR2_X1 U9129 ( .A1(n11629), .A2(n7677), .ZN(n7202) );
  NAND2_X1 U9130 ( .A1(n8796), .A2(n8795), .ZN(n14738) );
  NOR2_X1 U9131 ( .A1(n14916), .A2(n8335), .ZN(n8333) );
  AND2_X1 U9132 ( .A1(n13209), .A2(n13208), .ZN(n7203) );
  AND2_X1 U9133 ( .A1(n9617), .A2(n13735), .ZN(n9840) );
  AND2_X1 U9134 ( .A1(n13201), .A2(n13200), .ZN(n7204) );
  AND2_X1 U9135 ( .A1(n15042), .A2(n14595), .ZN(n7205) );
  INV_X1 U9136 ( .A(n14383), .ZN(n15042) );
  AND2_X1 U9137 ( .A1(n8506), .A2(n8505), .ZN(n14383) );
  AND2_X1 U9138 ( .A1(n7766), .A2(n7765), .ZN(n7206) );
  AND2_X1 U9139 ( .A1(n7280), .A2(n7518), .ZN(n7207) );
  NOR2_X1 U9140 ( .A1(n13697), .A2(n13709), .ZN(n7208) );
  AND2_X1 U9141 ( .A1(n7515), .A2(n8736), .ZN(n7209) );
  INV_X1 U9142 ( .A(n13582), .ZN(n12214) );
  AND2_X1 U9143 ( .A1(n9294), .A2(n9278), .ZN(n9279) );
  INV_X1 U9144 ( .A(n7827), .ZN(n8597) );
  OAI21_X1 U9145 ( .B1(n7828), .B2(SI_4_), .A(n8426), .ZN(n7827) );
  AND2_X1 U9146 ( .A1(n8788), .A2(n8770), .ZN(n7210) );
  NAND2_X1 U9147 ( .A1(n10738), .A2(n10739), .ZN(n7211) );
  INV_X1 U9148 ( .A(n13704), .ZN(n7903) );
  INV_X1 U9149 ( .A(n14149), .ZN(n8058) );
  AND2_X1 U9150 ( .A1(n7329), .A2(n7853), .ZN(n7212) );
  AND2_X1 U9151 ( .A1(n9305), .A2(n9304), .ZN(n12610) );
  INV_X1 U9152 ( .A(n12610), .ZN(n12853) );
  NAND2_X1 U9153 ( .A1(n8964), .A2(n8963), .ZN(n14878) );
  AND2_X1 U9154 ( .A1(n8047), .A2(n12993), .ZN(n7213) );
  OR2_X1 U9155 ( .A1(n8921), .A2(n8140), .ZN(n7214) );
  INV_X1 U9156 ( .A(n13210), .ZN(n7756) );
  INV_X1 U9157 ( .A(n12073), .ZN(n8086) );
  AND2_X1 U9158 ( .A1(n7633), .A2(n7630), .ZN(n7215) );
  NAND2_X1 U9159 ( .A1(n12240), .A2(n11800), .ZN(n12261) );
  INV_X1 U9160 ( .A(n12261), .ZN(n8319) );
  NAND2_X1 U9161 ( .A1(n9303), .A2(n9302), .ZN(n15737) );
  AND2_X1 U9162 ( .A1(n10150), .A2(SI_30_), .ZN(n7216) );
  INV_X1 U9163 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7791) );
  OR2_X1 U9164 ( .A1(n8863), .A2(n8399), .ZN(n7217) );
  INV_X2 U9165 ( .A(n8901), .ZN(n8609) );
  INV_X2 U9166 ( .A(n9160), .ZN(n9477) );
  NAND3_X1 U9167 ( .A1(n10525), .A2(n10524), .A3(n10523), .ZN(n13138) );
  AND4_X1 U9168 ( .A1(n8198), .A2(n8199), .A3(n10545), .A4(n10406), .ZN(n7218)
         );
  NAND2_X1 U9169 ( .A1(n9928), .A2(n10986), .ZN(n9262) );
  AND2_X1 U9170 ( .A1(n7767), .A2(n7768), .ZN(n7219) );
  NAND2_X1 U9171 ( .A1(n8168), .A2(n9064), .ZN(n7220) );
  NOR2_X1 U9172 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8554) );
  NAND2_X1 U9173 ( .A1(n9522), .A2(n9521), .ZN(n13505) );
  AND2_X1 U9174 ( .A1(n10458), .A2(n11698), .ZN(n7221) );
  NAND2_X1 U9175 ( .A1(n9087), .A2(n7871), .ZN(n9076) );
  NAND2_X1 U9176 ( .A1(n13014), .A2(n8156), .ZN(n13729) );
  INV_X1 U9177 ( .A(n9138), .ZN(n9480) );
  INV_X1 U9178 ( .A(n9719), .ZN(n13017) );
  INV_X1 U9179 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8491) );
  NOR2_X1 U9180 ( .A1(n13991), .A2(n8243), .ZN(n7222) );
  OR2_X1 U9181 ( .A1(n13186), .A2(n13185), .ZN(n7223) );
  AND3_X1 U9182 ( .A1(n10516), .A2(n10515), .A3(n10514), .ZN(n7224) );
  OR2_X1 U9183 ( .A1(n14964), .A2(n15086), .ZN(n7225) );
  NOR2_X1 U9184 ( .A1(n9928), .A2(n11391), .ZN(n7226) );
  INV_X1 U9185 ( .A(n14593), .ZN(n8385) );
  NOR2_X1 U9186 ( .A1(n13580), .A2(n12379), .ZN(n7227) );
  NOR2_X1 U9187 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n10537) );
  INV_X1 U9188 ( .A(n12536), .ZN(n8076) );
  AND2_X1 U9189 ( .A1(n8974), .A2(n8973), .ZN(n14858) );
  INV_X1 U9190 ( .A(n14858), .ZN(n10181) );
  NOR2_X1 U9191 ( .A1(n12004), .A2(n12003), .ZN(n7228) );
  AND4_X1 U9192 ( .A1(n8561), .A2(n8560), .A3(n8559), .A4(n8558), .ZN(n11441)
         );
  XNOR2_X1 U9193 ( .A(n8508), .B(n8507), .ZN(n8517) );
  CLKBUF_X1 U9194 ( .A(n8564), .Z(n14769) );
  INV_X1 U9195 ( .A(n8289), .ZN(n8288) );
  NAND2_X1 U9196 ( .A1(n12891), .A2(n12887), .ZN(n8289) );
  NAND2_X1 U9197 ( .A1(n8607), .A2(n8606), .ZN(n16008) );
  INV_X1 U9198 ( .A(n8368), .ZN(n8367) );
  NAND2_X1 U9199 ( .A1(n8370), .A2(n14455), .ZN(n8368) );
  INV_X1 U9200 ( .A(n7808), .ZN(n7807) );
  OR2_X1 U9201 ( .A1(n8441), .A2(n7809), .ZN(n7808) );
  INV_X1 U9202 ( .A(n13123), .ZN(n13828) );
  OAI21_X1 U9203 ( .B1(n12801), .B2(n9148), .A(n9569), .ZN(n13123) );
  NAND2_X1 U9204 ( .A1(n13950), .A2(n10840), .ZN(n13919) );
  NAND2_X1 U9205 ( .A1(n8849), .A2(n8848), .ZN(n15025) );
  INV_X1 U9206 ( .A(n15004), .ZN(n15009) );
  AND2_X1 U9207 ( .A1(n13182), .A2(n11944), .ZN(n7229) );
  NAND2_X1 U9208 ( .A1(n15105), .A2(n8877), .ZN(n8252) );
  INV_X1 U9209 ( .A(n8252), .ZN(n8245) );
  XNOR2_X1 U9210 ( .A(n13143), .B(n10835), .ZN(n10540) );
  NAND2_X1 U9211 ( .A1(n10853), .A2(n10852), .ZN(n13988) );
  OR2_X1 U9212 ( .A1(n10356), .A2(n10357), .ZN(n7230) );
  NOR2_X1 U9213 ( .A1(n13117), .A2(n13627), .ZN(n9735) );
  INV_X1 U9214 ( .A(n9735), .ZN(n8004) );
  NAND2_X2 U9215 ( .A1(n9928), .A2(n8421), .ZN(n9148) );
  AND4_X1 U9216 ( .A1(n10704), .A2(n10411), .A3(n7218), .A4(n8232), .ZN(n7231)
         );
  NOR2_X1 U9217 ( .A1(n15809), .A2(n15808), .ZN(n7232) );
  NOR2_X1 U9218 ( .A1(n15847), .A2(n15846), .ZN(n7233) );
  NAND2_X1 U9219 ( .A1(n10665), .A2(n10664), .ZN(n13249) );
  AND2_X1 U9220 ( .A1(n8065), .A2(n13410), .ZN(n7234) );
  AND2_X1 U9221 ( .A1(n7812), .A2(n14149), .ZN(n7235) );
  INV_X1 U9222 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8810) );
  OR2_X1 U9223 ( .A1(n13074), .A2(n13073), .ZN(n7236) );
  AND2_X1 U9224 ( .A1(n14271), .A2(n14044), .ZN(n7237) );
  INV_X1 U9225 ( .A(n14301), .ZN(n14152) );
  NAND2_X1 U9226 ( .A1(n10795), .A2(n10794), .ZN(n14301) );
  AND2_X1 U9227 ( .A1(n7771), .A2(n7770), .ZN(n7238) );
  INV_X1 U9228 ( .A(n7775), .ZN(n14902) );
  AND2_X1 U9229 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n7239) );
  AND2_X1 U9230 ( .A1(n9818), .A2(n9817), .ZN(n12969) );
  OR2_X1 U9231 ( .A1(n11391), .A2(n9974), .ZN(n7240) );
  INV_X1 U9232 ( .A(n11994), .ZN(n13584) );
  AND4_X1 U9233 ( .A1(n9164), .A2(n9163), .A3(n9162), .A4(n9161), .ZN(n11994)
         );
  NOR2_X1 U9234 ( .A1(n15675), .A2(n9902), .ZN(n7241) );
  AND2_X1 U9235 ( .A1(n14301), .A2(n14008), .ZN(n7242) );
  AND2_X1 U9236 ( .A1(n13678), .A2(n7992), .ZN(n7243) );
  INV_X1 U9237 ( .A(n7727), .ZN(n7726) );
  AND2_X1 U9238 ( .A1(n10438), .A2(n10415), .ZN(n7244) );
  AND2_X1 U9239 ( .A1(n13234), .A2(n13233), .ZN(n7245) );
  AND2_X1 U9240 ( .A1(n9486), .A2(n9485), .ZN(n7246) );
  AND2_X1 U9241 ( .A1(n8879), .A2(n8250), .ZN(n8328) );
  AND2_X1 U9242 ( .A1(n14931), .A2(n8333), .ZN(n7247) );
  AND2_X1 U9243 ( .A1(n12956), .A2(n12828), .ZN(n7248) );
  AND2_X1 U9244 ( .A1(n14886), .A2(n14746), .ZN(n7249) );
  AND2_X1 U9245 ( .A1(n13249), .A2(n13251), .ZN(n7250) );
  OR2_X1 U9246 ( .A1(n8188), .A2(n13277), .ZN(n7251) );
  OR2_X1 U9247 ( .A1(n10362), .A2(n10360), .ZN(n7252) );
  INV_X1 U9248 ( .A(n8335), .ZN(n8334) );
  INV_X1 U9249 ( .A(n8254), .ZN(n8253) );
  AND2_X1 U9250 ( .A1(n10087), .A2(n10086), .ZN(n7253) );
  AND2_X1 U9251 ( .A1(n10072), .A2(n10071), .ZN(n7254) );
  INV_X1 U9252 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7863) );
  INV_X1 U9253 ( .A(n12909), .ZN(n8230) );
  AND2_X1 U9254 ( .A1(n8239), .A2(n7418), .ZN(n7255) );
  OR2_X1 U9255 ( .A1(n13252), .A2(n13254), .ZN(n7256) );
  AND2_X1 U9256 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7257) );
  NOR2_X1 U9257 ( .A1(n12129), .A2(n12256), .ZN(n7258) );
  INV_X1 U9258 ( .A(n8054), .ZN(n8053) );
  NAND2_X1 U9259 ( .A1(n8058), .A2(n8059), .ZN(n8054) );
  NOR2_X1 U9260 ( .A1(n14314), .A2(n14192), .ZN(n7259) );
  OR2_X1 U9261 ( .A1(n8863), .A2(n8404), .ZN(n7260) );
  AND2_X1 U9262 ( .A1(n13678), .A2(n13689), .ZN(n7261) );
  AND2_X1 U9263 ( .A1(n14401), .A2(n8392), .ZN(n7262) );
  INV_X1 U9264 ( .A(n7892), .ZN(n7891) );
  OAI21_X1 U9265 ( .B1(n7897), .B2(n7893), .A(n9796), .ZN(n7892) );
  INV_X1 U9266 ( .A(n8274), .ZN(n8273) );
  OR2_X1 U9267 ( .A1(n8701), .A2(n8440), .ZN(n7263) );
  AND2_X1 U9268 ( .A1(n12102), .A2(n13582), .ZN(n7264) );
  AND2_X1 U9269 ( .A1(n8232), .A2(n10415), .ZN(n7265) );
  NAND3_X1 U9270 ( .A1(n7197), .A2(n8792), .A3(n7862), .ZN(n7266) );
  NAND3_X1 U9271 ( .A1(n8499), .A2(n8412), .A3(n8792), .ZN(n7267) );
  AND2_X1 U9272 ( .A1(n7708), .A2(n7711), .ZN(n7268) );
  AND2_X1 U9273 ( .A1(n12984), .A2(n13574), .ZN(n7269) );
  INV_X1 U9274 ( .A(n11020), .ZN(n7697) );
  INV_X1 U9275 ( .A(n7761), .ZN(n7760) );
  NAND2_X1 U9276 ( .A1(n7763), .A2(n7762), .ZN(n7761) );
  INV_X1 U9277 ( .A(n7773), .ZN(n7772) );
  NAND2_X1 U9278 ( .A1(n8322), .A2(n7774), .ZN(n7773) );
  OR2_X1 U9279 ( .A1(n13300), .A2(n13302), .ZN(n7270) );
  AND2_X1 U9280 ( .A1(n13505), .A2(n13569), .ZN(n7271) );
  AND2_X1 U9281 ( .A1(n13261), .A2(n13260), .ZN(n7272) );
  AND2_X1 U9282 ( .A1(n13175), .A2(n13174), .ZN(n7273) );
  AND2_X1 U9283 ( .A1(n13090), .A2(n13571), .ZN(n7274) );
  AND2_X1 U9284 ( .A1(n8447), .A2(n15307), .ZN(n7275) );
  AND2_X1 U9285 ( .A1(n10114), .A2(n10113), .ZN(n7276) );
  INV_X1 U9286 ( .A(n7521), .ZN(n7520) );
  NAND2_X1 U9287 ( .A1(n8837), .A2(n8824), .ZN(n7521) );
  NOR2_X1 U9288 ( .A1(n14172), .A2(n14009), .ZN(n7277) );
  AND2_X1 U9289 ( .A1(n8359), .A2(n8350), .ZN(n7278) );
  NAND2_X1 U9290 ( .A1(n7435), .A2(n9064), .ZN(n9630) );
  AND2_X1 U9291 ( .A1(n7272), .A2(n13264), .ZN(n7279) );
  AND2_X1 U9292 ( .A1(n15009), .A2(n8838), .ZN(n7280) );
  INV_X1 U9293 ( .A(n12389), .ZN(n7860) );
  NAND2_X1 U9294 ( .A1(n8989), .A2(n8988), .ZN(n12389) );
  AND2_X1 U9295 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7281) );
  AND2_X1 U9296 ( .A1(n13138), .A2(n13135), .ZN(n11452) );
  AND2_X1 U9297 ( .A1(n10138), .A2(n10137), .ZN(n7282) );
  AND2_X1 U9298 ( .A1(n13194), .A2(n13193), .ZN(n7283) );
  INV_X1 U9299 ( .A(n14878), .ZN(n15036) );
  AND2_X1 U9300 ( .A1(n8270), .A2(n8265), .ZN(n7284) );
  AND2_X1 U9301 ( .A1(n14922), .A2(n14508), .ZN(n8920) );
  INV_X1 U9302 ( .A(n9706), .ZN(n9587) );
  INV_X1 U9303 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8232) );
  INV_X1 U9304 ( .A(n8372), .ZN(n8371) );
  NAND2_X1 U9305 ( .A1(n8373), .A2(n16194), .ZN(n8372) );
  INV_X1 U9306 ( .A(n7457), .ZN(n7456) );
  NAND2_X1 U9307 ( .A1(n7458), .A2(n9485), .ZN(n7457) );
  AND2_X1 U9308 ( .A1(n9591), .A2(n9596), .ZN(n9594) );
  NOR2_X1 U9309 ( .A1(n14895), .A2(n8279), .ZN(n7285) );
  AND2_X1 U9310 ( .A1(n7815), .A2(n7814), .ZN(n7286) );
  OR2_X1 U9311 ( .A1(n10301), .A2(n10302), .ZN(n7287) );
  OR2_X1 U9312 ( .A1(n10271), .A2(n10286), .ZN(n7288) );
  INV_X1 U9313 ( .A(n13428), .ZN(n14114) );
  OR2_X1 U9314 ( .A1(n13290), .A2(n7310), .ZN(n7289) );
  NOR2_X1 U9315 ( .A1(n13545), .A2(n8293), .ZN(n8292) );
  INV_X1 U9316 ( .A(n9222), .ZN(n7623) );
  AND2_X1 U9317 ( .A1(n8184), .A2(n13220), .ZN(n7290) );
  NAND2_X1 U9318 ( .A1(n14967), .A2(n14749), .ZN(n7291) );
  AOI21_X1 U9319 ( .B1(n8045), .B2(n13423), .A(n8413), .ZN(n8044) );
  AND2_X1 U9320 ( .A1(n7206), .A2(n14108), .ZN(n7292) );
  OAI21_X1 U9321 ( .B1(n7493), .B2(SI_5_), .A(n8428), .ZN(n8427) );
  AND2_X1 U9322 ( .A1(n8491), .A2(n7863), .ZN(n7293) );
  INV_X1 U9323 ( .A(n8736), .ZN(n7514) );
  AND2_X1 U9324 ( .A1(n8385), .A2(n8381), .ZN(n7294) );
  OR2_X1 U9325 ( .A1(n8192), .A2(n13253), .ZN(n7295) );
  AND2_X1 U9326 ( .A1(n7284), .A2(n8269), .ZN(n7296) );
  AND2_X1 U9327 ( .A1(n9453), .A2(n8015), .ZN(n7297) );
  INV_X1 U9328 ( .A(n10587), .ZN(n7416) );
  INV_X1 U9329 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9089) );
  INV_X1 U9330 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8503) );
  INV_X1 U9331 ( .A(n12103), .ZN(n8305) );
  INV_X1 U9332 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10526) );
  INV_X1 U9333 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10980) );
  INV_X1 U9334 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8400) );
  INV_X1 U9335 ( .A(n11628), .ZN(n7677) );
  NOR2_X1 U9336 ( .A1(n13001), .A2(n8046), .ZN(n8045) );
  INV_X1 U9337 ( .A(n7675), .ZN(n7674) );
  NAND2_X1 U9338 ( .A1(n11568), .A2(n13586), .ZN(n7675) );
  INV_X1 U9339 ( .A(n9793), .ZN(n7897) );
  INV_X1 U9340 ( .A(n9103), .ZN(n9352) );
  AND2_X1 U9341 ( .A1(n10218), .A2(n9011), .ZN(n8263) );
  NAND2_X1 U9342 ( .A1(n12480), .A2(n12481), .ZN(n7597) );
  AND2_X1 U9343 ( .A1(n8323), .A2(n7772), .ZN(n7298) );
  INV_X1 U9344 ( .A(n12671), .ZN(n7793) );
  NAND2_X1 U9345 ( .A1(n12195), .A2(n8700), .ZN(n12315) );
  INV_X1 U9346 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7864) );
  OR2_X1 U9347 ( .A1(n10437), .A2(n10415), .ZN(n10721) );
  NAND2_X1 U9348 ( .A1(n12971), .A2(n9360), .ZN(n12970) );
  INV_X1 U9349 ( .A(n8074), .ZN(n8073) );
  AND2_X1 U9350 ( .A1(n8078), .A2(n13417), .ZN(n8074) );
  NAND2_X1 U9351 ( .A1(n8480), .A2(n15290), .ZN(n7299) );
  INV_X1 U9352 ( .A(n9829), .ZN(n7905) );
  AND2_X1 U9353 ( .A1(n15047), .A2(n14746), .ZN(n7300) );
  INV_X1 U9354 ( .A(n13663), .ZN(n7458) );
  NAND2_X1 U9355 ( .A1(n14271), .A2(n14092), .ZN(n7301) );
  NAND2_X1 U9356 ( .A1(n10019), .A2(n15737), .ZN(n7302) );
  OR2_X1 U9357 ( .A1(n14278), .A2(n14005), .ZN(n7303) );
  NAND2_X1 U9358 ( .A1(n9326), .A2(n9325), .ZN(n12789) );
  NAND2_X1 U9359 ( .A1(n9607), .A2(n9608), .ZN(n9708) );
  INV_X1 U9360 ( .A(n9830), .ZN(n7908) );
  NAND2_X1 U9361 ( .A1(n8939), .A2(n8938), .ZN(n15047) );
  XOR2_X1 U9362 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P3_ADDR_REG_4__SCAN_IN), .Z(
        n7304) );
  NAND2_X1 U9363 ( .A1(n10891), .A2(n10890), .ZN(n14267) );
  INV_X1 U9364 ( .A(n14267), .ZN(n7758) );
  INV_X1 U9365 ( .A(n9752), .ZN(n7887) );
  AND4_X1 U9366 ( .A1(n9293), .A2(n9292), .A3(n9291), .A4(n9290), .ZN(n12776)
         );
  INV_X1 U9367 ( .A(n15010), .ZN(n7572) );
  XNOR2_X1 U9368 ( .A(n9265), .B(P3_IR_REG_10__SCAN_IN), .ZN(n15705) );
  NAND2_X1 U9369 ( .A1(n8062), .A2(n7248), .ZN(n12952) );
  AND2_X1 U9370 ( .A1(n12612), .A2(n13578), .ZN(n7305) );
  AND2_X1 U9371 ( .A1(n14072), .A2(n7301), .ZN(n7306) );
  INV_X1 U9372 ( .A(n13491), .ZN(n8307) );
  AND2_X1 U9373 ( .A1(n7445), .A2(n7448), .ZN(n7307) );
  AND2_X1 U9374 ( .A1(n13116), .A2(n13115), .ZN(n7308) );
  AND3_X1 U9375 ( .A1(n8042), .A2(n10409), .A3(n10408), .ZN(n10704) );
  AND2_X1 U9376 ( .A1(n13314), .A2(n13313), .ZN(n7309) );
  AND2_X1 U9377 ( .A1(n13288), .A2(n13287), .ZN(n7310) );
  INV_X1 U9378 ( .A(n13734), .ZN(n13572) );
  AND4_X1 U9379 ( .A1(n9398), .A2(n9397), .A3(n9396), .A4(n9395), .ZN(n13734)
         );
  NAND2_X1 U9380 ( .A1(n12962), .A2(n7760), .ZN(n7764) );
  OR2_X1 U9381 ( .A1(n12496), .A2(n12497), .ZN(n7311) );
  AND2_X1 U9382 ( .A1(n9438), .A2(n9437), .ZN(n7312) );
  AND2_X1 U9383 ( .A1(n8075), .A2(n8078), .ZN(n7313) );
  OR2_X1 U9384 ( .A1(n14517), .A2(n14516), .ZN(n7314) );
  NAND2_X1 U9385 ( .A1(n8047), .A2(n8045), .ZN(n7315) );
  AND2_X1 U9386 ( .A1(n8264), .A2(n8263), .ZN(n7316) );
  AND2_X1 U9387 ( .A1(n7895), .A2(n7894), .ZN(n7317) );
  AND2_X1 U9388 ( .A1(n7482), .A2(n7484), .ZN(n7318) );
  INV_X1 U9389 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9369) );
  INV_X1 U9390 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7913) );
  NOR2_X1 U9391 ( .A1(n16158), .A2(n12784), .ZN(n7319) );
  NOR2_X1 U9392 ( .A1(n13544), .A2(n13571), .ZN(n7320) );
  AND2_X1 U9393 ( .A1(n8454), .A2(n15305), .ZN(n7321) );
  AND2_X1 U9394 ( .A1(n12853), .A2(n12776), .ZN(n7322) );
  NAND3_X1 U9395 ( .A1(n8792), .A2(n7197), .A3(n8810), .ZN(n7323) );
  AND2_X1 U9396 ( .A1(n8465), .A2(n15192), .ZN(n7324) );
  AND2_X1 U9397 ( .A1(n8467), .A2(n11731), .ZN(n7325) );
  AND2_X1 U9398 ( .A1(n14583), .A2(n14582), .ZN(n7326) );
  OR2_X1 U9399 ( .A1(n14693), .A2(n7385), .ZN(n7384) );
  NAND2_X1 U9400 ( .A1(n8475), .A2(n8532), .ZN(n7327) );
  NOR2_X1 U9401 ( .A1(n10020), .A2(n11030), .ZN(n7328) );
  INV_X1 U9402 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9592) );
  OR2_X1 U9403 ( .A1(n10143), .A2(n7962), .ZN(n7329) );
  NOR2_X1 U9404 ( .A1(n15008), .A2(n8253), .ZN(n7330) );
  AND2_X1 U9405 ( .A1(n7739), .A2(n7737), .ZN(n7331) );
  AND2_X1 U9406 ( .A1(n13401), .A2(n13037), .ZN(n7332) );
  AND2_X1 U9407 ( .A1(n12855), .A2(n8824), .ZN(n7333) );
  INV_X1 U9408 ( .A(n9297), .ZN(n7654) );
  AND2_X1 U9409 ( .A1(n9306), .A2(n9296), .ZN(n9297) );
  AND2_X1 U9410 ( .A1(n7299), .A2(n8908), .ZN(n7334) );
  OR2_X1 U9411 ( .A1(n13316), .A2(n7309), .ZN(n7335) );
  INV_X1 U9412 ( .A(n7742), .ZN(n7741) );
  NAND2_X1 U9413 ( .A1(n15749), .A2(n7302), .ZN(n7742) );
  INV_X1 U9414 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11393) );
  NAND2_X1 U9415 ( .A1(n9279), .A2(n9297), .ZN(n7336) );
  INV_X1 U9416 ( .A(n7554), .ZN(n7553) );
  NAND2_X1 U9417 ( .A1(n7555), .A2(n8472), .ZN(n7554) );
  INV_X1 U9418 ( .A(n15942), .ZN(n15894) );
  AND2_X1 U9419 ( .A1(n14853), .A2(n15931), .ZN(n14997) );
  INV_X1 U9420 ( .A(n10435), .ZN(n12624) );
  INV_X1 U9421 ( .A(n13216), .ZN(n7492) );
  AND2_X1 U9422 ( .A1(n7217), .A2(n8349), .ZN(n10042) );
  INV_X1 U9423 ( .A(n10042), .ZN(n7861) );
  NAND2_X1 U9424 ( .A1(n10711), .A2(n10710), .ZN(n14337) );
  INV_X1 U9425 ( .A(n14337), .ZN(n7762) );
  NAND2_X1 U9426 ( .A1(n8760), .A2(n8759), .ZN(n14679) );
  INV_X1 U9427 ( .A(n14679), .ZN(n8322) );
  NAND2_X1 U9428 ( .A1(n8150), .A2(n11892), .ZN(n11881) );
  NAND2_X1 U9429 ( .A1(n10834), .A2(n10833), .ZN(n14290) );
  INV_X1 U9430 ( .A(n14290), .ZN(n7765) );
  OAI21_X2 U9431 ( .B1(n11041), .B2(n8937), .A(n8689), .ZN(n14661) );
  INV_X1 U9432 ( .A(n14661), .ZN(n7778) );
  NAND2_X1 U9433 ( .A1(n12209), .A2(n9230), .ZN(n12231) );
  NAND2_X1 U9434 ( .A1(n12166), .A2(n12165), .ZN(n12522) );
  AND2_X1 U9435 ( .A1(n8302), .A2(n8301), .ZN(n7337) );
  NAND2_X1 U9436 ( .A1(n10040), .A2(n14835), .ZN(n10041) );
  NOR2_X1 U9437 ( .A1(n14694), .A2(n14695), .ZN(n14693) );
  INV_X1 U9438 ( .A(n14560), .ZN(n7777) );
  INV_X1 U9439 ( .A(n8323), .ZN(n12485) );
  INV_X1 U9440 ( .A(n7894), .ZN(n7893) );
  NOR2_X1 U9441 ( .A1(n9794), .A2(n12509), .ZN(n7894) );
  NOR2_X1 U9442 ( .A1(n12052), .A2(n9906), .ZN(n7338) );
  INV_X1 U9443 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7402) );
  AND2_X1 U9444 ( .A1(n8084), .A2(n12072), .ZN(n7339) );
  NAND2_X1 U9445 ( .A1(n11902), .A2(n8151), .ZN(n12209) );
  AND2_X1 U9446 ( .A1(n10149), .A2(n15277), .ZN(n7340) );
  NAND2_X1 U9447 ( .A1(n12182), .A2(n12305), .ZN(n12175) );
  INV_X1 U9448 ( .A(n12175), .ZN(n7755) );
  AND2_X1 U9449 ( .A1(n11911), .A2(n8361), .ZN(n7341) );
  AND2_X1 U9450 ( .A1(n8393), .A2(n8392), .ZN(n7342) );
  NOR2_X1 U9451 ( .A1(n12138), .A2(n8237), .ZN(n7343) );
  INV_X1 U9452 ( .A(n9012), .ZN(n8262) );
  AND2_X1 U9453 ( .A1(n12000), .A2(n11878), .ZN(n9926) );
  INV_X1 U9454 ( .A(n9926), .ZN(n11657) );
  INV_X1 U9455 ( .A(n16133), .ZN(n16009) );
  INV_X1 U9456 ( .A(n16076), .ZN(n8318) );
  INV_X1 U9457 ( .A(n15881), .ZN(n7680) );
  NAND2_X1 U9458 ( .A1(n13354), .A2(n11459), .ZN(n14236) );
  NAND2_X1 U9459 ( .A1(n8582), .A2(n10038), .ZN(n11582) );
  OR2_X1 U9460 ( .A1(n15984), .A2(n8275), .ZN(n7344) );
  INV_X1 U9461 ( .A(n9529), .ZN(n7658) );
  OR2_X1 U9462 ( .A1(n15768), .A2(n16164), .ZN(n7345) );
  AND2_X1 U9463 ( .A1(n9887), .A2(n9728), .ZN(n15959) );
  AND2_X1 U9464 ( .A1(n11423), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7346) );
  OR2_X1 U9465 ( .A1(n12012), .A2(n12011), .ZN(n7400) );
  AND2_X1 U9466 ( .A1(n9501), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7347) );
  INV_X1 U9467 ( .A(n7527), .ZN(n11567) );
  OR2_X1 U9468 ( .A1(n11416), .A2(n7676), .ZN(n7527) );
  NOR2_X1 U9469 ( .A1(n10416), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n14365) );
  INV_X1 U9470 ( .A(n7378), .ZN(n15395) );
  AND2_X1 U9471 ( .A1(n13128), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7348) );
  AND2_X1 U9472 ( .A1(n7467), .A2(n7466), .ZN(n7349) );
  INV_X1 U9473 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8107) );
  XOR2_X1 U9474 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n7350) );
  INV_X1 U9475 ( .A(SI_2_), .ZN(n7377) );
  INV_X1 U9476 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7665) );
  INV_X1 U9477 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7802) );
  INV_X1 U9478 ( .A(n15126), .ZN(n16133) );
  INV_X1 U9479 ( .A(n14376), .ZN(n14370) );
  NOR2_X1 U9480 ( .A1(n10986), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14376) );
  NAND3_X1 U9481 ( .A1(n8198), .A2(n8199), .A3(n10545), .ZN(n7351) );
  AND2_X1 U9482 ( .A1(n7351), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10508) );
  NAND3_X1 U9483 ( .A1(n7353), .A2(n7352), .A3(n11776), .ZN(n11939) );
  NAND3_X1 U9484 ( .A1(n11770), .A2(n11716), .A3(n11676), .ZN(n7353) );
  NAND2_X1 U9485 ( .A1(n11677), .A2(n11683), .ZN(n11771) );
  INV_X2 U9486 ( .A(n10417), .ZN(n13464) );
  NAND2_X1 U9487 ( .A1(n14365), .A2(P2_IR_REG_30__SCAN_IN), .ZN(n7360) );
  NAND2_X1 U9488 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n7363), .ZN(n7362) );
  NAND2_X2 U9489 ( .A1(n10417), .A2(n10425), .ZN(n10943) );
  NAND2_X1 U9490 ( .A1(n14226), .A2(n14225), .ZN(n14224) );
  INV_X1 U9491 ( .A(n8141), .ZN(n7372) );
  NAND2_X1 U9492 ( .A1(n7372), .A2(SI_2_), .ZN(n7376) );
  NAND2_X1 U9493 ( .A1(n7379), .A2(n8103), .ZN(n8101) );
  NAND2_X1 U9494 ( .A1(n7379), .A2(n8425), .ZN(n8598) );
  OAI211_X1 U9495 ( .C1(n7379), .C2(n7827), .A(n8102), .B(n8427), .ZN(n8617)
         );
  NAND2_X1 U9496 ( .A1(n8590), .A2(n7379), .ZN(n7378) );
  NAND3_X1 U9497 ( .A1(n7392), .A2(n7391), .A3(n7390), .ZN(n12095) );
  OAI21_X2 U9498 ( .B1(n14546), .B2(n7395), .A(n7393), .ZN(n14648) );
  NAND2_X1 U9499 ( .A1(n14648), .A2(n14515), .ZN(n14622) );
  NAND2_X1 U9500 ( .A1(n14732), .A2(n14731), .ZN(n7398) );
  NAND2_X1 U9501 ( .A1(n7398), .A2(n7396), .ZN(n7397) );
  NAND2_X1 U9502 ( .A1(n7397), .A2(n8363), .ZN(n14572) );
  NAND2_X2 U9503 ( .A1(n14572), .A2(n14573), .ZN(n14571) );
  NAND2_X1 U9504 ( .A1(n14433), .A2(n14434), .ZN(n7399) );
  NAND2_X1 U9505 ( .A1(n7401), .A2(n10562), .ZN(n11515) );
  NOR2_X1 U9506 ( .A1(n14001), .A2(n7401), .ZN(n10976) );
  NAND2_X1 U9507 ( .A1(n10558), .A2(n10971), .ZN(n7401) );
  NAND2_X1 U9508 ( .A1(n10437), .A2(n8410), .ZN(n7405) );
  INV_X1 U9509 ( .A(n10448), .ZN(n7407) );
  NAND2_X1 U9510 ( .A1(n10447), .A2(n7408), .ZN(n10950) );
  NOR2_X1 U9511 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n7409) );
  NAND2_X1 U9512 ( .A1(n7412), .A2(n7410), .ZN(n10604) );
  NAND2_X1 U9513 ( .A1(n10587), .A2(n7411), .ZN(n7410) );
  INV_X1 U9514 ( .A(n11483), .ZN(n7411) );
  NAND2_X1 U9515 ( .A1(n11484), .A2(n7414), .ZN(n7412) );
  NAND2_X2 U9516 ( .A1(n7420), .A2(n7255), .ZN(n7424) );
  XNOR2_X2 U9517 ( .A(n7424), .B(n10835), .ZN(n10937) );
  NAND3_X1 U9518 ( .A1(n7426), .A2(n8233), .A3(n8234), .ZN(n12559) );
  XNOR2_X1 U9519 ( .A(n10540), .B(n10541), .ZN(n11365) );
  NAND2_X1 U9520 ( .A1(n7428), .A2(n7697), .ZN(n7427) );
  NAND2_X2 U9521 ( .A1(n13927), .A2(n13928), .ZN(n13926) );
  AND2_X2 U9522 ( .A1(n9080), .A2(n9078), .ZN(n9103) );
  NAND2_X1 U9523 ( .A1(n13588), .A2(n11538), .ZN(n9607) );
  NAND2_X1 U9524 ( .A1(n7868), .A2(n7867), .ZN(n13588) );
  NAND2_X1 U9525 ( .A1(n9708), .A2(n11494), .ZN(n9102) );
  INV_X1 U9526 ( .A(n7437), .ZN(n7439) );
  NOR2_X1 U9527 ( .A1(n15756), .A2(n9914), .ZN(n15764) );
  INV_X1 U9528 ( .A(n9930), .ZN(n7462) );
  NAND2_X1 U9529 ( .A1(n7459), .A2(n7461), .ZN(n11398) );
  INV_X1 U9530 ( .A(n15609), .ZN(n7460) );
  NAND2_X1 U9531 ( .A1(n9898), .A2(n7465), .ZN(n7463) );
  XNOR2_X1 U9532 ( .A(n9897), .B(n15630), .ZN(n15621) );
  INV_X1 U9533 ( .A(n7467), .ZN(n15620) );
  NAND2_X1 U9534 ( .A1(n15814), .A2(n7476), .ZN(n7475) );
  NOR2_X1 U9535 ( .A1(n15814), .A2(n9922), .ZN(n15847) );
  XNOR2_X1 U9536 ( .A(n7477), .B(n7967), .ZN(n7537) );
  INV_X1 U9537 ( .A(n12959), .ZN(n7483) );
  NAND2_X1 U9538 ( .A1(n12957), .A2(n12955), .ZN(n7819) );
  NAND2_X1 U9539 ( .A1(n8077), .A2(n8071), .ZN(n7490) );
  AOI21_X1 U9540 ( .B1(n8071), .B2(n8073), .A(n13419), .ZN(n7491) );
  MUX2_X1 U9541 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8421), .Z(n7493) );
  OAI21_X1 U9542 ( .B1(n12288), .B2(n8615), .A(n7495), .ZN(n11627) );
  OR2_X1 U9543 ( .A1(n12299), .A2(n11840), .ZN(n7495) );
  NAND2_X1 U9544 ( .A1(n11582), .A2(n11583), .ZN(n7496) );
  NAND2_X1 U9545 ( .A1(n8993), .A2(n10035), .ZN(n10207) );
  NAND4_X1 U9546 ( .A1(n7505), .A2(n7498), .A3(n8488), .A4(n8487), .ZN(n7504)
         );
  NAND2_X1 U9547 ( .A1(n7499), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8501) );
  NAND4_X1 U9548 ( .A1(n7502), .A2(n7501), .A3(n7500), .A4(n8412), .ZN(n7499)
         );
  NOR2_X1 U9549 ( .A1(n7503), .A2(n8494), .ZN(n7501) );
  NAND3_X1 U9550 ( .A1(n7505), .A2(n8492), .A3(n8813), .ZN(n8493) );
  NAND2_X1 U9551 ( .A1(n8489), .A2(n8492), .ZN(n7503) );
  NAND2_X1 U9552 ( .A1(n7507), .A2(n7509), .ZN(n13087) );
  NAND2_X1 U9553 ( .A1(n12814), .A2(n7511), .ZN(n7507) );
  NAND2_X1 U9554 ( .A1(n12195), .A2(n7209), .ZN(n7513) );
  NOR2_X1 U9555 ( .A1(n8331), .A2(n7516), .ZN(n7515) );
  OAI211_X1 U9556 ( .C1(n7514), .C2(n8329), .A(n7513), .B(n12455), .ZN(n12454)
         );
  NAND2_X1 U9557 ( .A1(n12195), .A2(n7515), .ZN(n7517) );
  NAND2_X1 U9558 ( .A1(n9702), .A2(n11967), .ZN(n11223) );
  AOI21_X2 U9559 ( .B1(n12360), .B2(n12359), .A(n7526), .ZN(n12373) );
  NAND3_X1 U9560 ( .A1(n7527), .A2(n7675), .A3(n11571), .ZN(n11649) );
  NOR2_X1 U9561 ( .A1(n11567), .A2(n7674), .ZN(n11572) );
  AOI21_X2 U9562 ( .B1(n7528), .B2(n8333), .A(n7666), .ZN(n14899) );
  OR2_X2 U9563 ( .A1(n14953), .A2(n7667), .ZN(n7528) );
  INV_X2 U9564 ( .A(n8563), .ZN(n11032) );
  NAND4_X1 U9565 ( .A1(n9108), .A2(n7198), .A3(n7866), .A4(n9063), .ZN(n9302)
         );
  NAND2_X1 U9566 ( .A1(n7536), .A2(n7533), .ZN(P3_U3201) );
  NAND2_X1 U9567 ( .A1(n7754), .A2(n15806), .ZN(n7535) );
  NAND2_X1 U9568 ( .A1(n7537), .A2(n15845), .ZN(n7536) );
  INV_X2 U9569 ( .A(n8421), .ZN(n10986) );
  MUX2_X1 U9570 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n8421), .Z(n7546) );
  OR2_X1 U9571 ( .A1(n8893), .A2(n7554), .ZN(n7550) );
  NAND2_X1 U9572 ( .A1(n7550), .A2(n7551), .ZN(n8909) );
  NAND3_X1 U9573 ( .A1(n10223), .A2(n14916), .A3(n7556), .ZN(n10224) );
  INV_X1 U9574 ( .A(n12270), .ZN(n12271) );
  OAI21_X2 U9575 ( .B1(n8581), .B2(n15915), .A(n10038), .ZN(n12270) );
  NAND2_X1 U9576 ( .A1(n8581), .A2(n15915), .ZN(n10038) );
  OAI21_X1 U9577 ( .B1(n12274), .B2(n7564), .A(n7561), .ZN(n12289) );
  NAND2_X1 U9578 ( .A1(n7563), .A2(n8996), .ZN(n7562) );
  INV_X1 U9579 ( .A(n12290), .ZN(n10208) );
  INV_X1 U9580 ( .A(n7565), .ZN(n14944) );
  NAND2_X1 U9581 ( .A1(n7572), .A2(n7684), .ZN(n7571) );
  NAND4_X1 U9582 ( .A1(n8499), .A2(n8792), .A3(n8342), .A4(n8412), .ZN(n8509)
         );
  NAND4_X1 U9583 ( .A1(n8499), .A2(n8792), .A3(n8342), .A4(n7573), .ZN(n7575)
         );
  NOR2_X1 U9584 ( .A1(n14867), .A2(n14868), .ZN(n14866) );
  NAND2_X1 U9585 ( .A1(n11804), .A2(n7586), .ZN(n7584) );
  NAND2_X1 U9586 ( .A1(n7591), .A2(n7589), .ZN(n12933) );
  NOR2_X1 U9587 ( .A1(n15563), .A2(n15562), .ZN(n15561) );
  NAND2_X1 U9588 ( .A1(n15585), .A2(n7602), .ZN(n7600) );
  NAND2_X1 U9589 ( .A1(n7600), .A2(n7601), .ZN(n10383) );
  NAND2_X1 U9590 ( .A1(n15590), .A2(n15591), .ZN(n15587) );
  INV_X1 U9591 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9592 ( .A1(n7612), .A2(n7614), .ZN(n10362) );
  NAND3_X1 U9593 ( .A1(n7230), .A2(n7915), .A3(n7613), .ZN(n7612) );
  INV_X1 U9594 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U9595 ( .A1(n7619), .A2(n9112), .ZN(n9123) );
  AND2_X1 U9596 ( .A1(n10526), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9109) );
  XNOR2_X1 U9597 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9110) );
  NAND2_X1 U9598 ( .A1(n9209), .A2(n9222), .ZN(n7620) );
  NAND2_X1 U9599 ( .A1(n7620), .A2(n7621), .ZN(n9239) );
  NAND2_X1 U9600 ( .A1(n13877), .A2(n9690), .ZN(n7627) );
  NAND2_X1 U9601 ( .A1(n7628), .A2(n7629), .ZN(n9502) );
  NAND2_X1 U9602 ( .A1(n9467), .A2(n7215), .ZN(n7628) );
  NAND2_X1 U9603 ( .A1(n9677), .A2(n7638), .ZN(n7636) );
  NAND2_X1 U9604 ( .A1(n9677), .A2(n9676), .ZN(n7637) );
  NAND2_X1 U9605 ( .A1(n9166), .A2(n7645), .ZN(n7641) );
  NAND2_X1 U9606 ( .A1(n7641), .A2(n7642), .ZN(n9204) );
  INV_X1 U9607 ( .A(n9277), .ZN(n7651) );
  OAI21_X1 U9608 ( .B1(n9277), .B2(n7336), .A(n7652), .ZN(n9309) );
  NAND2_X1 U9609 ( .A1(n9503), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U9610 ( .A1(n7657), .A2(n7656), .ZN(n8034) );
  OAI21_X1 U9611 ( .B1(n9442), .B2(n8013), .A(n8012), .ZN(n9467) );
  NAND2_X1 U9612 ( .A1(n9206), .A2(n9205), .ZN(n9209) );
  NAND2_X1 U9613 ( .A1(n8011), .A2(n9124), .ZN(n9150) );
  NAND2_X1 U9614 ( .A1(n9441), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U9615 ( .A1(n9343), .A2(n9342), .ZN(n9346) );
  NAND2_X1 U9616 ( .A1(n9331), .A2(n9330), .ZN(n9343) );
  NAND2_X1 U9617 ( .A1(n9239), .A2(n9238), .ZN(n9242) );
  INV_X1 U9618 ( .A(n9567), .ZN(n7663) );
  NAND2_X1 U9619 ( .A1(n9440), .A2(n9439), .ZN(n9441) );
  NAND2_X1 U9620 ( .A1(n7996), .A2(n9874), .ZN(n7994) );
  OAI21_X1 U9621 ( .B1(n12686), .B2(n10218), .A(n8806), .ZN(n12857) );
  NAND2_X1 U9622 ( .A1(n14897), .A2(n7314), .ZN(n14883) );
  NAND2_X1 U9623 ( .A1(n12124), .A2(n12125), .ZN(n12123) );
  NAND2_X1 U9624 ( .A1(n12197), .A2(n12196), .ZN(n12195) );
  NAND2_X1 U9625 ( .A1(n12251), .A2(n8680), .ZN(n12197) );
  AOI21_X2 U9626 ( .B1(n15041), .B2(n15877), .A(n7682), .ZN(n15045) );
  NAND2_X1 U9627 ( .A1(n11799), .A2(n11798), .ZN(n11797) );
  NAND2_X1 U9628 ( .A1(n11625), .A2(n8630), .ZN(n11799) );
  NAND2_X1 U9629 ( .A1(n12630), .A2(n8789), .ZN(n12686) );
  NAND2_X1 U9630 ( .A1(n14899), .A2(n14898), .ZN(n14897) );
  AOI22_X1 U9631 ( .A1(n8951), .A2(P1_REG1_REG_1__SCAN_IN), .B1(n8901), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7673) );
  AND2_X2 U9632 ( .A1(n8512), .A2(n8518), .ZN(n8901) );
  NAND2_X1 U9633 ( .A1(n12454), .A2(n8751), .ZN(n12484) );
  NAND2_X1 U9634 ( .A1(n12123), .A2(n8664), .ZN(n12253) );
  XNOR2_X1 U9635 ( .A(n7668), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  XNOR2_X1 U9636 ( .A(n10362), .B(n10360), .ZN(n15559) );
  NAND2_X1 U9637 ( .A1(n7692), .A2(n15579), .ZN(n15585) );
  INV_X1 U9638 ( .A(n7930), .ZN(n10341) );
  AOI21_X1 U9639 ( .B1(n9743), .B2(n9742), .A(n9741), .ZN(n9744) );
  NAND2_X1 U9640 ( .A1(n7920), .A2(n10357), .ZN(n7919) );
  OAI21_X1 U9641 ( .B1(n12314), .B2(n8331), .A(n12401), .ZN(n8330) );
  NAND2_X1 U9642 ( .A1(n7819), .A2(n13420), .ZN(n12959) );
  INV_X1 U9643 ( .A(n8100), .ZN(n8099) );
  INV_X1 U9644 ( .A(n12581), .ZN(n8077) );
  OR2_X1 U9645 ( .A1(n8953), .A2(n8546), .ZN(n8548) );
  NAND2_X2 U9646 ( .A1(n8517), .A2(n15156), .ZN(n8953) );
  NAND3_X1 U9647 ( .A1(n7673), .A2(n8548), .A3(n8547), .ZN(n8564) );
  NAND2_X1 U9648 ( .A1(n9649), .A2(n9641), .ZN(n9643) );
  NAND2_X1 U9649 ( .A1(n8290), .A2(n8291), .ZN(n13484) );
  NAND2_X1 U9650 ( .A1(n13038), .A2(n13402), .ZN(n14081) );
  INV_X1 U9651 ( .A(n13143), .ZN(n15948) );
  NAND2_X1 U9652 ( .A1(n14210), .A2(n13028), .ZN(n8050) );
  NAND2_X1 U9653 ( .A1(n7231), .A2(n8410), .ZN(n10448) );
  NAND2_X1 U9654 ( .A1(n7678), .A2(n7677), .ZN(n11625) );
  NAND2_X1 U9655 ( .A1(n15135), .A2(n15984), .ZN(n8276) );
  INV_X1 U9656 ( .A(n11627), .ZN(n7678) );
  NAND2_X1 U9657 ( .A1(n9548), .A2(n9547), .ZN(n9561) );
  NAND3_X1 U9658 ( .A1(n8038), .A2(n8040), .A3(n9861), .ZN(n7681) );
  NAND2_X1 U9659 ( .A1(n15007), .A2(n8858), .ZN(n14991) );
  NAND2_X1 U9660 ( .A1(n8276), .A2(n7344), .ZN(P1_U3525) );
  AOI21_X1 U9661 ( .B1(n7996), .B2(n7999), .A(n7995), .ZN(n7699) );
  OAI21_X1 U9662 ( .B1(n12312), .B2(n12314), .A(n9005), .ZN(n12392) );
  NAND2_X1 U9663 ( .A1(n8272), .A2(n14944), .ZN(n8269) );
  NOR2_X1 U9664 ( .A1(n7689), .A2(n15039), .ZN(n7688) );
  NOR2_X1 U9665 ( .A1(n14870), .A2(n14869), .ZN(n8416) );
  NAND2_X1 U9666 ( .A1(n8266), .A2(n8269), .ZN(n14915) );
  OR2_X1 U9667 ( .A1(n9727), .A2(n11223), .ZN(n7700) );
  NAND2_X1 U9668 ( .A1(n9310), .A2(n8037), .ZN(n9328) );
  NAND2_X1 U9669 ( .A1(n9257), .A2(n9256), .ZN(n9260) );
  NAND2_X1 U9670 ( .A1(n8396), .A2(n8395), .ZN(n16170) );
  NAND2_X1 U9671 ( .A1(n9857), .A2(n9856), .ZN(n8041) );
  NAND2_X1 U9672 ( .A1(n7690), .A2(n7688), .ZN(n15136) );
  INV_X1 U9673 ( .A(n8416), .ZN(n7689) );
  NAND2_X1 U9674 ( .A1(n15040), .A2(n16139), .ZN(n7690) );
  NAND2_X1 U9675 ( .A1(n12269), .A2(n12271), .ZN(n8582) );
  NAND2_X1 U9676 ( .A1(n8509), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U9677 ( .A1(n8034), .A2(n9534), .ZN(n9548) );
  NAND2_X1 U9678 ( .A1(n9385), .A2(n9384), .ZN(n9400) );
  NAND2_X1 U9679 ( .A1(n15045), .A2(n7695), .ZN(n15137) );
  NAND2_X1 U9680 ( .A1(n11797), .A2(n8647), .ZN(n12124) );
  INV_X1 U9681 ( .A(n15572), .ZN(n7924) );
  XNOR2_X1 U9682 ( .A(n10351), .B(n7912), .ZN(n15551) );
  NAND2_X1 U9683 ( .A1(n12482), .A2(n7210), .ZN(n12630) );
  NAND2_X2 U9684 ( .A1(n15161), .A2(n13009), .ZN(n8563) );
  NAND2_X1 U9685 ( .A1(n12484), .A2(n12483), .ZN(n12482) );
  NAND2_X1 U9686 ( .A1(n8704), .A2(n8703), .ZN(n8706) );
  NAND2_X1 U9687 ( .A1(n9420), .A2(n9419), .ZN(n9440) );
  INV_X1 U9688 ( .A(n8330), .ZN(n8329) );
  NAND2_X1 U9689 ( .A1(n8019), .A2(n8020), .ZN(n9385) );
  OAI21_X1 U9690 ( .B1(n9729), .B2(n9728), .A(n7700), .ZN(n9870) );
  NAND2_X1 U9691 ( .A1(n7699), .A2(n7994), .ZN(n9701) );
  NAND2_X1 U9692 ( .A1(n8000), .A2(n7998), .ZN(n7997) );
  NAND2_X1 U9693 ( .A1(n7934), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7933) );
  NAND2_X1 U9694 ( .A1(n8668), .A2(n8437), .ZN(n8681) );
  NAND2_X1 U9695 ( .A1(n8320), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7769) );
  NOR2_X1 U9696 ( .A1(n11022), .A2(n8937), .ZN(n8281) );
  NAND2_X1 U9697 ( .A1(n7701), .A2(n7704), .ZN(n13186) );
  OR2_X1 U9698 ( .A1(n8178), .A2(n7702), .ZN(n7701) );
  OAI22_X1 U9699 ( .A1(n7703), .A2(n13171), .B1(n13172), .B2(n13169), .ZN(
        n7702) );
  NAND2_X1 U9700 ( .A1(n7705), .A2(n7251), .ZN(n13285) );
  OR2_X1 U9701 ( .A1(n13199), .A2(n7194), .ZN(n7708) );
  NAND2_X1 U9702 ( .A1(n13199), .A2(n7711), .ZN(n7710) );
  NAND2_X1 U9703 ( .A1(n7710), .A2(n7709), .ZN(n13205) );
  OAI21_X1 U9704 ( .B1(n7245), .B2(n7719), .A(n7714), .ZN(n8191) );
  INV_X1 U9705 ( .A(n13245), .ZN(n7725) );
  NOR2_X1 U9706 ( .A1(n13238), .A2(n13240), .ZN(n7727) );
  NAND3_X1 U9707 ( .A1(n8179), .A2(n8183), .A3(n7730), .ZN(n7729) );
  AND3_X1 U9708 ( .A1(n10704), .A2(n7218), .A3(n10411), .ZN(n10437) );
  NAND4_X1 U9709 ( .A1(n10438), .A2(n10704), .A3(n7218), .A4(n10411), .ZN(
        n7732) );
  NAND2_X1 U9710 ( .A1(n13259), .A2(n7201), .ZN(n7734) );
  NAND2_X1 U9711 ( .A1(n7734), .A2(n7733), .ZN(n13271) );
  INV_X1 U9712 ( .A(n14036), .ZN(n14037) );
  NOR2_X1 U9713 ( .A1(n14075), .A2(n14267), .ZN(n14074) );
  NAND2_X1 U9714 ( .A1(n12962), .A2(n7759), .ZN(n14229) );
  INV_X1 U9715 ( .A(n7764), .ZN(n14228) );
  NAND2_X1 U9716 ( .A1(n14167), .A2(n7292), .ZN(n14102) );
  NAND2_X1 U9717 ( .A1(n10535), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7768) );
  XNOR2_X2 U9718 ( .A(n7769), .B(n8503), .ZN(n13009) );
  NAND3_X1 U9719 ( .A1(n7777), .A2(n7776), .A3(n7779), .ZN(n12463) );
  NAND3_X1 U9720 ( .A1(n9028), .A2(n9029), .A3(n8277), .ZN(n15135) );
  MUX2_X1 U9721 ( .A(n11140), .B(P1_REG1_REG_1__SCAN_IN), .S(n11147), .Z(
        n14772) );
  NAND2_X1 U9722 ( .A1(n7800), .A2(n8107), .ZN(n7932) );
  NAND3_X1 U9723 ( .A1(n7802), .A2(n7801), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7800) );
  NAND2_X1 U9724 ( .A1(n8666), .A2(n8665), .ZN(n8668) );
  OAI21_X1 U9725 ( .B1(n8666), .B2(n7808), .A(n7806), .ZN(n8705) );
  NAND2_X1 U9726 ( .A1(n7820), .A2(n7823), .ZN(n8087) );
  NAND2_X1 U9727 ( .A1(n14128), .A2(n7821), .ZN(n7820) );
  MUX2_X1 U9728 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n8421), .Z(n7828) );
  NAND3_X1 U9729 ( .A1(n7831), .A2(n7938), .A3(n7830), .ZN(n7829) );
  NAND3_X1 U9730 ( .A1(n7836), .A2(n7942), .A3(n7835), .ZN(n7834) );
  NAND3_X1 U9731 ( .A1(n7841), .A2(n7947), .A3(n7840), .ZN(n7839) );
  NAND3_X1 U9732 ( .A1(n7846), .A2(n7845), .A3(n7940), .ZN(n7844) );
  OR2_X1 U9733 ( .A1(n10115), .A2(n10116), .ZN(n10117) );
  NAND3_X1 U9734 ( .A1(n10108), .A2(n7952), .A3(n10107), .ZN(n7848) );
  NAND3_X1 U9735 ( .A1(n10133), .A2(n7954), .A3(n10132), .ZN(n7850) );
  NAND2_X1 U9736 ( .A1(n7852), .A2(n7851), .ZN(n10289) );
  INV_X1 U9737 ( .A(n10144), .ZN(n7854) );
  OR2_X1 U9738 ( .A1(n10040), .A2(n14835), .ZN(n7859) );
  OAI211_X2 U9739 ( .C1(n7857), .C2(n7856), .A(n7858), .B(n7855), .ZN(n10109)
         );
  OR2_X1 U9740 ( .A1(n12389), .A2(n10041), .ZN(n7855) );
  NAND2_X1 U9741 ( .A1(n7859), .A2(n10041), .ZN(n10175) );
  OR2_X1 U9742 ( .A1(n7859), .A2(n12389), .ZN(n7858) );
  NAND3_X1 U9743 ( .A1(n7197), .A2(n8792), .A3(n8394), .ZN(n8828) );
  NAND3_X1 U9744 ( .A1(n7868), .A2(n7867), .A3(n15908), .ZN(n9608) );
  AND2_X1 U9745 ( .A1(n9081), .A2(n9082), .ZN(n7867) );
  AND2_X1 U9746 ( .A1(n7870), .A2(n7869), .ZN(n7868) );
  NAND2_X1 U9747 ( .A1(n9087), .A2(n8149), .ZN(n9088) );
  NOR2_X1 U9748 ( .A1(n7877), .A2(n7878), .ZN(n13607) );
  OAI21_X2 U9749 ( .B1(n9622), .B2(n7881), .A(n7879), .ZN(n9874) );
  NAND2_X1 U9750 ( .A1(n12747), .A2(n7885), .ZN(n7882) );
  NAND2_X1 U9751 ( .A1(n7882), .A2(n7883), .ZN(n9616) );
  OAI21_X2 U9752 ( .B1(n12229), .B2(n7892), .A(n7889), .ZN(n12448) );
  NAND2_X1 U9753 ( .A1(n13738), .A2(n7904), .ZN(n7901) );
  NAND2_X1 U9754 ( .A1(n7901), .A2(n7902), .ZN(n9619) );
  NAND3_X1 U9755 ( .A1(n7917), .A2(P2_ADDR_REG_5__SCAN_IN), .A3(n7916), .ZN(
        n7915) );
  NAND2_X1 U9756 ( .A1(n7917), .A2(n7916), .ZN(n15557) );
  INV_X1 U9757 ( .A(n7915), .ZN(n15555) );
  NOR2_X1 U9758 ( .A1(n15552), .A2(n10353), .ZN(n10356) );
  OAI21_X1 U9759 ( .B1(n15552), .B2(n10353), .A(n7918), .ZN(n7917) );
  INV_X1 U9760 ( .A(n10357), .ZN(n7918) );
  INV_X1 U9761 ( .A(n15589), .ZN(n15588) );
  NAND2_X1 U9762 ( .A1(n10383), .A2(n7921), .ZN(n15589) );
  INV_X1 U9763 ( .A(n10384), .ZN(n7921) );
  NAND3_X1 U9764 ( .A1(n8106), .A2(n15853), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7934) );
  INV_X1 U9765 ( .A(n10123), .ZN(n7939) );
  INV_X1 U9766 ( .A(n10068), .ZN(n7941) );
  INV_X1 U9767 ( .A(n10098), .ZN(n7943) );
  INV_X1 U9768 ( .A(n10078), .ZN(n7946) );
  INV_X1 U9769 ( .A(n10083), .ZN(n7948) );
  INV_X1 U9770 ( .A(n10093), .ZN(n7951) );
  INV_X1 U9771 ( .A(n10110), .ZN(n7953) );
  INV_X1 U9772 ( .A(n10134), .ZN(n7955) );
  INV_X1 U9773 ( .A(n10118), .ZN(n7959) );
  INV_X1 U9774 ( .A(n10142), .ZN(n7962) );
  OR2_X1 U9775 ( .A1(n10060), .A2(n7966), .ZN(n7963) );
  NAND3_X1 U9776 ( .A1(n10058), .A2(n10057), .A3(n7965), .ZN(n7964) );
  INV_X1 U9777 ( .A(n10059), .ZN(n7966) );
  NAND2_X1 U9778 ( .A1(n15675), .A2(n11620), .ZN(n7970) );
  OR2_X1 U9779 ( .A1(n15675), .A2(n7973), .ZN(n7971) );
  NAND2_X1 U9780 ( .A1(n9899), .A2(n15664), .ZN(n7982) );
  NAND2_X1 U9781 ( .A1(n11927), .A2(n9778), .ZN(n9611) );
  NAND2_X1 U9782 ( .A1(n7984), .A2(n9776), .ZN(n11927) );
  NAND2_X1 U9783 ( .A1(n11880), .A2(n11884), .ZN(n7984) );
  INV_X1 U9784 ( .A(n7985), .ZN(n13749) );
  OR2_X1 U9785 ( .A1(n9708), .A2(n11496), .ZN(n15904) );
  INV_X1 U9786 ( .A(n9750), .ZN(n7993) );
  NAND2_X1 U9787 ( .A1(n9874), .A2(n8005), .ZN(n8001) );
  INV_X1 U9788 ( .A(n8007), .ZN(n8006) );
  NAND2_X4 U9789 ( .A1(n7187), .A2(n9969), .ZN(n9928) );
  NAND2_X2 U9790 ( .A1(n9614), .A2(n9613), .ZN(n12229) );
  NAND2_X1 U9791 ( .A1(n9123), .A2(n9122), .ZN(n8011) );
  INV_X1 U9792 ( .A(n9453), .ZN(n8013) );
  NAND2_X1 U9793 ( .A1(n9454), .A2(n9453), .ZN(n9457) );
  NAND2_X1 U9794 ( .A1(n7297), .A2(n9442), .ZN(n9454) );
  INV_X1 U9795 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U9796 ( .A1(n9346), .A2(n8022), .ZN(n8019) );
  NAND3_X1 U9797 ( .A1(n8033), .A2(n8031), .A3(n8030), .ZN(n9536) );
  NAND2_X1 U9798 ( .A1(n9530), .A2(n8035), .ZN(n8030) );
  INV_X1 U9799 ( .A(n9530), .ZN(n8029) );
  NAND3_X1 U9800 ( .A1(n8033), .A2(n8036), .A3(n8030), .ZN(n12646) );
  NAND2_X1 U9801 ( .A1(n9328), .A2(n9327), .ZN(n9331) );
  NAND4_X1 U9802 ( .A1(n10409), .A2(n10407), .A3(n10460), .A4(n10408), .ZN(
        n10450) );
  NAND2_X1 U9803 ( .A1(n8050), .A2(n8048), .ZN(n14196) );
  NAND2_X1 U9804 ( .A1(n14113), .A2(n7332), .ZN(n13038) );
  NAND2_X1 U9805 ( .A1(n12582), .A2(n8064), .ZN(n12704) );
  NAND2_X1 U9806 ( .A1(n8406), .A2(n9867), .ZN(n9869) );
  OAI21_X1 U9807 ( .B1(n11775), .B2(n8069), .A(n8067), .ZN(n12068) );
  NAND2_X1 U9808 ( .A1(n8066), .A2(n7234), .ZN(n12071) );
  NAND2_X1 U9809 ( .A1(n8067), .A2(n8069), .ZN(n8065) );
  NAND2_X1 U9810 ( .A1(n11775), .A2(n8067), .ZN(n8066) );
  NAND2_X1 U9811 ( .A1(n8082), .A2(n12188), .ZN(n8079) );
  NAND2_X1 U9812 ( .A1(n8079), .A2(n8080), .ZN(n12533) );
  NAND2_X1 U9813 ( .A1(n8087), .A2(n8088), .ZN(n14066) );
  AND4_X2 U9814 ( .A1(n10704), .A2(n10411), .A3(n7218), .A4(n8097), .ZN(n8096)
         );
  OAI21_X1 U9815 ( .B1(n8597), .B2(n8104), .A(n8616), .ZN(n8100) );
  NAND2_X1 U9816 ( .A1(n8101), .A2(n8099), .ZN(n8618) );
  OR2_X1 U9817 ( .A1(n8971), .A2(n8115), .ZN(n8112) );
  NAND2_X1 U9818 ( .A1(n8971), .A2(n8110), .ZN(n8109) );
  NAND2_X1 U9819 ( .A1(n8971), .A2(n8970), .ZN(n10148) );
  NAND2_X1 U9820 ( .A1(n8839), .A2(n8119), .ZN(n8116) );
  NAND2_X1 U9821 ( .A1(n8116), .A2(n8117), .ZN(n8893) );
  INV_X1 U9822 ( .A(n8720), .ZN(n8127) );
  OAI21_X1 U9823 ( .B1(n8720), .B2(n8719), .A(n8445), .ZN(n8738) );
  AOI21_X1 U9824 ( .B1(n8719), .B2(n8445), .A(n8131), .ZN(n8130) );
  NAND2_X1 U9825 ( .A1(n8909), .A2(n7334), .ZN(n8139) );
  INV_X1 U9826 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U9827 ( .A1(n11881), .A2(n9192), .ZN(n11928) );
  OAI21_X2 U9828 ( .B1(n9438), .B2(n8160), .A(n8158), .ZN(n13673) );
  NAND3_X1 U9829 ( .A1(n9064), .A2(n9071), .A3(n8171), .ZN(n8172) );
  NAND2_X1 U9830 ( .A1(n8176), .A2(n13705), .ZN(n8175) );
  NAND2_X1 U9831 ( .A1(n8177), .A2(n13608), .ZN(n8176) );
  NAND2_X4 U9832 ( .A1(n13354), .A2(n7221), .ZN(n13393) );
  NAND2_X1 U9833 ( .A1(n16041), .A2(n7221), .ZN(n12713) );
  NAND3_X1 U9834 ( .A1(n13207), .A2(n13206), .A3(n8184), .ZN(n8179) );
  NAND2_X1 U9835 ( .A1(n8181), .A2(n13220), .ZN(n8180) );
  NAND3_X1 U9836 ( .A1(n13207), .A2(n13206), .A3(n7290), .ZN(n8182) );
  NOR2_X1 U9837 ( .A1(n13271), .A2(n13270), .ZN(n13272) );
  NAND3_X1 U9838 ( .A1(n13312), .A2(n13311), .A3(n7335), .ZN(n8186) );
  NAND2_X1 U9839 ( .A1(n8191), .A2(n7295), .ZN(n13259) );
  OAI22_X1 U9840 ( .A1(n13192), .A2(n8193), .B1(n13191), .B2(n13190), .ZN(
        n13199) );
  NOR2_X1 U9841 ( .A1(n8194), .A2(n8195), .ZN(n8193) );
  INV_X1 U9842 ( .A(n13190), .ZN(n8194) );
  INV_X1 U9843 ( .A(n13191), .ZN(n8195) );
  NAND3_X1 U9844 ( .A1(n7186), .A2(n13286), .A3(n7289), .ZN(n8196) );
  INV_X1 U9845 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8199) );
  INV_X1 U9846 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8198) );
  INV_X2 U9847 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U9848 ( .A1(n10567), .A2(n11599), .ZN(n11484) );
  NAND2_X1 U9849 ( .A1(n10566), .A2(n10565), .ZN(n11514) );
  NOR2_X1 U9850 ( .A1(n13979), .A2(n8202), .ZN(n8201) );
  OR2_X1 U9851 ( .A1(n13979), .A2(n8204), .ZN(n8203) );
  NAND2_X1 U9852 ( .A1(n13939), .A2(n10714), .ZN(n8206) );
  INV_X1 U9853 ( .A(n13939), .ZN(n8209) );
  NAND2_X1 U9854 ( .A1(n13938), .A2(n13939), .ZN(n13937) );
  NAND2_X1 U9855 ( .A1(n13926), .A2(n10715), .ZN(n13938) );
  OAI21_X1 U9856 ( .B1(n13960), .B2(n8213), .A(n8210), .ZN(n10804) );
  XNOR2_X1 U9857 ( .A(n10804), .B(n10796), .ZN(n13970) );
  NAND2_X1 U9858 ( .A1(n13902), .A2(n8215), .ZN(n13950) );
  NAND2_X1 U9859 ( .A1(n12596), .A2(n12597), .ZN(n8223) );
  INV_X1 U9860 ( .A(n8217), .ZN(n8216) );
  NAND2_X1 U9861 ( .A1(n12909), .A2(n8221), .ZN(n8219) );
  INV_X1 U9862 ( .A(n8231), .ZN(n12910) );
  INV_X1 U9863 ( .A(n8228), .ZN(n13927) );
  NAND2_X1 U9864 ( .A1(n10693), .A2(n10694), .ZN(n8229) );
  NAND2_X1 U9865 ( .A1(n10630), .A2(n10629), .ZN(n8238) );
  NAND3_X1 U9866 ( .A1(n7572), .A2(n15004), .A3(n8252), .ZN(n8247) );
  NAND2_X1 U9867 ( .A1(n8857), .A2(n14752), .ZN(n8254) );
  NOR2_X1 U9868 ( .A1(n12856), .A2(n8262), .ZN(n8255) );
  NAND2_X1 U9869 ( .A1(n8259), .A2(n8255), .ZN(n8256) );
  NAND3_X1 U9870 ( .A1(n8261), .A2(n8260), .A3(n9012), .ZN(n12854) );
  NAND2_X1 U9871 ( .A1(n15077), .A2(n14490), .ZN(n8274) );
  AOI21_X1 U9872 ( .B1(n8972), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n8281), .ZN(
        n8280) );
  NAND2_X1 U9873 ( .A1(n13501), .A2(n8285), .ZN(n8283) );
  NAND2_X1 U9874 ( .A1(n13512), .A2(n8292), .ZN(n8290) );
  NAND2_X1 U9875 ( .A1(n11990), .A2(n8298), .ZN(n8297) );
  NAND2_X1 U9876 ( .A1(n11990), .A2(n8303), .ZN(n8302) );
  NAND2_X1 U9877 ( .A1(n8297), .A2(n8299), .ZN(n12360) );
  NAND2_X1 U9878 ( .A1(n11990), .A2(n11989), .ZN(n11991) );
  INV_X1 U9879 ( .A(n8302), .ZN(n12022) );
  NOR2_X1 U9880 ( .A1(n11992), .A2(n8304), .ZN(n8303) );
  INV_X1 U9881 ( .A(n11989), .ZN(n8304) );
  AOI21_X1 U9882 ( .B1(n13093), .B2(n8308), .A(n8306), .ZN(n13103) );
  NAND4_X1 U9883 ( .A1(n8792), .A2(n8321), .A3(n8412), .A4(n7197), .ZN(n8320)
         );
  INV_X1 U9884 ( .A(n14991), .ZN(n8326) );
  NOR2_X1 U9885 ( .A1(n14939), .A2(n14686), .ZN(n8335) );
  OAI21_X1 U9886 ( .B1(n13074), .B2(n8338), .A(n8337), .ZN(n8336) );
  INV_X1 U9887 ( .A(n8336), .ZN(n8983) );
  INV_X1 U9888 ( .A(n8339), .ZN(n8338) );
  NAND3_X1 U9889 ( .A1(n8346), .A2(n8345), .A3(n8603), .ZN(n8494) );
  NOR2_X4 U9890 ( .A1(n15880), .A2(n7860), .ZN(n16012) );
  MUX2_X1 U9891 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8986), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8349) );
  NAND2_X1 U9892 ( .A1(n8355), .A2(n11837), .ZN(n8354) );
  NOR2_X1 U9893 ( .A1(n11838), .A2(n11837), .ZN(n11913) );
  OAI21_X1 U9894 ( .B1(n16193), .B2(n8368), .A(n8365), .ZN(n14706) );
  NAND2_X1 U9895 ( .A1(n14719), .A2(n14720), .ZN(n14718) );
  OAI211_X1 U9896 ( .C1(n14719), .C2(n8379), .A(n8375), .B(n8374), .ZN(n14599)
         );
  NAND2_X1 U9897 ( .A1(n14719), .A2(n7294), .ZN(n8374) );
  OAI21_X1 U9898 ( .B1(n8385), .B2(n8380), .A(n8376), .ZN(n8375) );
  NAND2_X1 U9899 ( .A1(n8380), .A2(n8377), .ZN(n8376) );
  NAND2_X2 U9900 ( .A1(n14600), .A2(n8386), .ZN(n14546) );
  NAND2_X2 U9901 ( .A1(n14601), .A2(n14485), .ZN(n14600) );
  INV_X1 U9902 ( .A(n8393), .ZN(n14391) );
  NAND2_X1 U9903 ( .A1(n14392), .A2(n14393), .ZN(n8392) );
  INV_X1 U9904 ( .A(n16172), .ZN(n8396) );
  INV_X1 U9905 ( .A(n14418), .ZN(n8398) );
  OR2_X1 U9906 ( .A1(n8863), .A2(n8402), .ZN(n8988) );
  OR2_X1 U9907 ( .A1(n10943), .A2(n14245), .ZN(n10557) );
  OR2_X1 U9908 ( .A1(n10943), .A2(n11133), .ZN(n10523) );
  OAI21_X1 U9909 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9873) );
  NAND4_X2 U9910 ( .A1(n10534), .A2(n10533), .A3(n10532), .A4(n10531), .ZN(
        n13144) );
  INV_X1 U9911 ( .A(n8951), .ZN(n10161) );
  OAI21_X1 U9912 ( .B1(n13398), .B2(n13397), .A(n13396), .ZN(n13447) );
  AOI21_X1 U9913 ( .B1(n13970), .B2(n13969), .A(n10805), .ZN(n10819) );
  INV_X1 U9914 ( .A(n11505), .ZN(n9725) );
  MUX2_X2 U9915 ( .A(n13826), .B(n13825), .S(n16169), .Z(n13827) );
  OAI21_X1 U9916 ( .B1(n15880), .B2(n12471), .A(n12154), .ZN(n15126) );
  NAND2_X1 U9917 ( .A1(n13464), .A2(n14372), .ZN(n10551) );
  OAI22_X1 U9918 ( .A1(n11605), .A2(n11606), .B1(n11547), .B2(n11546), .ZN(
        n11832) );
  NAND2_X1 U9919 ( .A1(n16012), .A2(n14835), .ZN(n11560) );
  AND2_X4 U9920 ( .A1(n9079), .A2(n9080), .ZN(n9139) );
  INV_X1 U9921 ( .A(n8839), .ZN(n8840) );
  INV_X1 U9922 ( .A(n15105), .ZN(n8878) );
  NOR2_X1 U9923 ( .A1(n9961), .A2(n9929), .ZN(n15845) );
  AND3_X2 U9924 ( .A1(n9668), .A2(n11660), .A3(n9667), .ZN(n16165) );
  INV_X1 U9925 ( .A(n16165), .ZN(n9674) );
  NOR2_X1 U9926 ( .A1(n13601), .A2(n13806), .ZN(n9670) );
  NAND2_X2 U9927 ( .A1(n11667), .A2(n15967), .ZN(n13715) );
  NOR2_X1 U9928 ( .A1(n9262), .A2(SI_2_), .ZN(n8405) );
  INV_X1 U9929 ( .A(n15025), .ZN(n8857) );
  OR2_X1 U9930 ( .A1(n13768), .A2(n13864), .ZN(n8407) );
  AND2_X1 U9931 ( .A1(n14967), .A2(n14666), .ZN(n8408) );
  AND4_X1 U9932 ( .A1(n10430), .A2(n10414), .A3(n10926), .A4(n10413), .ZN(
        n8409) );
  AND4_X1 U9933 ( .A1(n8411), .A2(n8409), .A3(n10915), .A4(n10919), .ZN(n8410)
         );
  INV_X1 U9934 ( .A(n9969), .ZN(n9966) );
  INV_X1 U9935 ( .A(n14751), .ZN(n8877) );
  INV_X1 U9936 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10303) );
  AND4_X1 U9937 ( .A1(n9359), .A2(n9358), .A3(n9357), .A4(n9356), .ZN(n12983)
         );
  NAND2_X1 U9938 ( .A1(n11236), .A2(n9926), .ZN(n15962) );
  INV_X1 U9939 ( .A(n15962), .ZN(n9880) );
  INV_X1 U9940 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9308) );
  INV_X1 U9941 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9158) );
  INV_X1 U9942 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9318) );
  INV_X1 U9943 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U9944 ( .A1(n11507), .A2(n15408), .ZN(n16190) );
  NAND2_X1 U9945 ( .A1(n11507), .A2(n11477), .ZN(n16188) );
  INV_X2 U9946 ( .A(n16188), .ZN(n16189) );
  AND2_X2 U9947 ( .A1(n9892), .A2(n11234), .ZN(n16169) );
  NAND2_X1 U9948 ( .A1(n12152), .A2(n11581), .ZN(n16142) );
  INV_X1 U9949 ( .A(n16141), .ZN(n16140) );
  AND2_X2 U9950 ( .A1(n11581), .A2(n9057), .ZN(n16141) );
  INV_X1 U9951 ( .A(n12969), .ZN(n9360) );
  AND2_X1 U9952 ( .A1(n14337), .A2(n14014), .ZN(n8413) );
  AND2_X1 U9953 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8414) );
  AND3_X1 U9954 ( .A1(n14263), .A2(n14262), .A3(n14261), .ZN(n8415) );
  NAND2_X2 U9955 ( .A1(n11700), .A2(n16038), .ZN(n16041) );
  AND2_X1 U9956 ( .A1(n10954), .A2(n10936), .ZN(n13940) );
  OAI21_X1 U9957 ( .B1(n15895), .B2(n13136), .A(n13393), .ZN(n13137) );
  INV_X1 U9958 ( .A(n13137), .ZN(n13139) );
  NAND2_X1 U9959 ( .A1(n13365), .A2(n13143), .ZN(n13146) );
  NAND2_X1 U9960 ( .A1(n14027), .A2(n13365), .ZN(n13152) );
  INV_X1 U9961 ( .A(n13154), .ZN(n13155) );
  OAI21_X1 U9962 ( .B1(n13226), .B2(n13393), .A(n13225), .ZN(n13227) );
  INV_X1 U9963 ( .A(n13253), .ZN(n13254) );
  INV_X1 U9964 ( .A(n13267), .ZN(n13268) );
  INV_X1 U9965 ( .A(n13277), .ZN(n13278) );
  INV_X1 U9966 ( .A(n13281), .ZN(n13282) );
  INV_X1 U9967 ( .A(n11884), .ZN(n9176) );
  INV_X1 U9968 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n10407) );
  NAND2_X1 U9969 ( .A1(n9117), .A2(n9116), .ZN(n11958) );
  INV_X1 U9970 ( .A(n10035), .ZN(n10036) );
  OAI21_X1 U9971 ( .B1(n11505), .B2(n11878), .A(n11732), .ZN(n11226) );
  INV_X1 U9972 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9387) );
  NAND2_X1 U9973 ( .A1(n10837), .A2(n10839), .ZN(n10840) );
  INV_X1 U9974 ( .A(n10825), .ZN(n10823) );
  INV_X1 U9975 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10423) );
  AND2_X1 U9976 ( .A1(n10862), .A2(n10861), .ZN(n10875) );
  INV_X1 U9977 ( .A(n13414), .ZN(n12525) );
  AND2_X1 U9978 ( .A1(n14665), .A2(n14664), .ZN(n14476) );
  AND2_X1 U9979 ( .A1(n8514), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8947) );
  AND2_X1 U9980 ( .A1(n15073), .A2(n14686), .ZN(n9017) );
  NAND2_X1 U9981 ( .A1(n15038), .A2(n15037), .ZN(n15039) );
  INV_X1 U9982 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15357) );
  INV_X1 U9983 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9231) );
  OR2_X1 U9984 ( .A1(n12886), .A2(n13575), .ZN(n12887) );
  AND2_X1 U9985 ( .A1(n9897), .A2(n15630), .ZN(n9898) );
  INV_X1 U9986 ( .A(n15721), .ZN(n10015) );
  INV_X1 U9987 ( .A(n13470), .ZN(n9881) );
  AND2_X1 U9988 ( .A1(n11658), .A2(n11657), .ZN(n11663) );
  AND2_X1 U9989 ( .A1(n10804), .A2(n10803), .ZN(n10805) );
  INV_X1 U9990 ( .A(n13948), .ZN(n10836) );
  NAND2_X1 U9991 ( .A1(n13400), .A2(n13399), .ZN(n13438) );
  NAND2_X1 U9992 ( .A1(n10823), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n10860) );
  NAND2_X1 U9993 ( .A1(n10773), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n10810) );
  OR2_X1 U9994 ( .A1(n10745), .A2(n10744), .ZN(n10759) );
  OR2_X1 U9995 ( .A1(n10943), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10515) );
  INV_X1 U9996 ( .A(n13399), .ZN(n13442) );
  NAND2_X1 U9997 ( .A1(n10654), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10669) );
  NOR2_X1 U9998 ( .A1(n14319), .A2(n13024), .ZN(n11474) );
  INV_X1 U9999 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n10406) );
  INV_X1 U10000 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8761) );
  AND2_X1 U10001 ( .A1(n14602), .A2(n14603), .ZN(n14485) );
  INV_X1 U10002 ( .A(n14586), .ZN(n14480) );
  INV_X1 U10003 ( .A(n8925), .ZN(n8941) );
  INV_X1 U10004 ( .A(n8913), .ZN(n8926) );
  INV_X1 U10005 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U10006 ( .A1(n8857), .A2(n8856), .ZN(n8858) );
  INV_X1 U10007 ( .A(n12633), .ZN(n8788) );
  NAND2_X1 U10008 ( .A1(n8727), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8762) );
  OR2_X1 U10009 ( .A1(n8692), .A2(n8513), .ZN(n8711) );
  INV_X1 U10010 ( .A(n10207), .ZN(n15920) );
  INV_X1 U10011 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8500) );
  INV_X1 U10012 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8984) );
  OR2_X1 U10013 ( .A1(n8739), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8740) );
  INV_X1 U10014 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10322) );
  NOR2_X1 U10015 ( .A1(n9194), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9214) );
  OR2_X1 U10016 ( .A1(n9552), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9572) );
  NOR2_X1 U10017 ( .A1(n9429), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9447) );
  AND2_X1 U10018 ( .A1(n9214), .A2(n15346), .ZN(n9232) );
  INV_X1 U10019 ( .A(n13688), .ZN(n13496) );
  AND2_X1 U10020 ( .A1(n9373), .A2(n15357), .ZN(n9393) );
  NAND2_X1 U10021 ( .A1(n9393), .A2(n9392), .ZN(n9409) );
  XNOR2_X1 U10022 ( .A(n11351), .B(n11350), .ZN(n11412) );
  INV_X1 U10023 ( .A(n13549), .ZN(n13559) );
  OR2_X1 U10024 ( .A1(n11240), .A2(n16157), .ZN(n11665) );
  AND2_X1 U10025 ( .A1(n9748), .A2(n9749), .ZN(n13663) );
  AND2_X1 U10026 ( .A1(n9807), .A2(n9806), .ZN(n12653) );
  OR2_X1 U10027 ( .A1(n9178), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U10028 ( .A1(n13586), .A2(n9134), .ZN(n9765) );
  INV_X1 U10029 ( .A(n13869), .ZN(n11662) );
  INV_X1 U10030 ( .A(n9605), .ZN(n9606) );
  INV_X1 U10031 ( .A(n9928), .ZN(n9425) );
  INV_X1 U10032 ( .A(n12379), .ZN(n16084) );
  NAND2_X1 U10033 ( .A1(n13870), .A2(n11244), .ZN(n11240) );
  AND2_X1 U10034 ( .A1(n9416), .A2(n9401), .ZN(n9402) );
  AND2_X1 U10035 ( .A1(n9342), .A2(n9329), .ZN(n9330) );
  AND2_X1 U10036 ( .A1(n9151), .A2(n9126), .ZN(n9149) );
  INV_X1 U10037 ( .A(n11636), .ZN(n10603) );
  NAND2_X1 U10038 ( .A1(n10564), .A2(n10563), .ZN(n10565) );
  OR2_X1 U10039 ( .A1(n10974), .A2(n10960), .ZN(n10961) );
  XNOR2_X1 U10040 ( .A(n13202), .B(n10857), .ZN(n11981) );
  INV_X1 U10041 ( .A(n10803), .ZN(n10796) );
  INV_X1 U10042 ( .A(n14092), .ZN(n14044) );
  OR2_X1 U10043 ( .A1(n10717), .A2(n10716), .ZN(n10733) );
  INV_X1 U10044 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n12473) );
  AND2_X1 U10045 ( .A1(n11074), .A2(n14375), .ZN(n11073) );
  INV_X1 U10046 ( .A(n14302), .ZN(n14319) );
  INV_X1 U10047 ( .A(n14018), .ZN(n13226) );
  INV_X1 U10048 ( .A(n16147), .ZN(n14231) );
  INV_X1 U10049 ( .A(n13430), .ZN(n14132) );
  INV_X1 U10050 ( .A(n13421), .ZN(n12830) );
  INV_X1 U10051 ( .A(n14236), .ZN(n14214) );
  NAND2_X1 U10052 ( .A1(n11466), .A2(n10835), .ZN(n14197) );
  AND2_X1 U10053 ( .A1(n10930), .A2(n10929), .ZN(n11471) );
  NAND2_X1 U10054 ( .A1(n10913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10916) );
  NOR2_X1 U10055 ( .A1(n8899), .A2(n14688), .ZN(n8538) );
  OR2_X1 U10056 ( .A1(n12150), .A2(n11551), .ZN(n11562) );
  AND2_X1 U10057 ( .A1(n8884), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8898) );
  INV_X1 U10058 ( .A(n13069), .ZN(n13073) );
  INV_X1 U10059 ( .A(n15925), .ZN(n15012) );
  INV_X1 U10060 ( .A(n11552), .ZN(n11033) );
  OR2_X1 U10061 ( .A1(n11552), .A2(n11449), .ZN(n15916) );
  INV_X1 U10062 ( .A(n16012), .ZN(n16077) );
  OR2_X1 U10063 ( .A1(n8687), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n8721) );
  INV_X1 U10064 ( .A(n8571), .ZN(n8573) );
  OAI21_X1 U10065 ( .B1(P3_ADDR_REG_13__SCAN_IN), .B2(n10324), .A(n10323), 
        .ZN(n10382) );
  AND2_X1 U10066 ( .A1(n11237), .A2(n11238), .ZN(n13549) );
  XNOR2_X1 U10067 ( .A(n13103), .B(n13101), .ZN(n13537) );
  NOR2_X1 U10068 ( .A1(n11353), .A2(n11352), .ZN(n11416) );
  INV_X1 U10069 ( .A(n13561), .ZN(n12504) );
  INV_X1 U10070 ( .A(n12136), .ZN(n9868) );
  AND4_X1 U10071 ( .A1(n9577), .A2(n9576), .A3(n9575), .A4(n9574), .ZN(n13470)
         );
  OR2_X1 U10072 ( .A1(n9962), .A2(n9963), .ZN(n9961) );
  INV_X1 U10073 ( .A(n15822), .ZN(n15834) );
  INV_X1 U10074 ( .A(n13717), .ZN(n13757) );
  INV_X1 U10075 ( .A(n15959), .ZN(n13705) );
  INV_X1 U10076 ( .A(n15967), .ZN(n15909) );
  AND3_X1 U10077 ( .A1(n9884), .A2(n9662), .A3(n9889), .ZN(n11660) );
  AND2_X1 U10078 ( .A1(n11879), .A2(n9755), .ZN(n16103) );
  NAND2_X1 U10079 ( .A1(n11658), .A2(n9626), .ZN(n16057) );
  INV_X1 U10080 ( .A(n9649), .ZN(n10990) );
  NAND2_X1 U10081 ( .A1(n14045), .A2(n10902), .ZN(n14072) );
  AND2_X1 U10082 ( .A1(n10961), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13994) );
  OR2_X1 U10083 ( .A1(n10955), .A2(n10943), .ZN(n10901) );
  INV_X1 U10084 ( .A(n15494), .ZN(n15508) );
  AND2_X1 U10085 ( .A1(n11073), .A2(n13455), .ZN(n15494) );
  AND2_X1 U10086 ( .A1(n15452), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15504) );
  AND2_X1 U10087 ( .A1(n11465), .A2(n10951), .ZN(n14089) );
  INV_X1 U10088 ( .A(n14197), .ZN(n14121) );
  INV_X1 U10089 ( .A(n15408), .ZN(n11477) );
  OR2_X1 U10090 ( .A1(n10435), .A2(n13443), .ZN(n16182) );
  INV_X1 U10091 ( .A(n16186), .ZN(n14346) );
  AND3_X1 U10092 ( .A1(n11476), .A2(n15401), .A3(n11475), .ZN(n11507) );
  AND2_X1 U10093 ( .A1(n12802), .A2(n10922), .ZN(n15403) );
  AND2_X1 U10094 ( .A1(n10650), .A2(n10678), .ZN(n15489) );
  AND4_X1 U10095 ( .A1(n8523), .A2(n8522), .A3(n8521), .A4(n8520), .ZN(n14595)
         );
  OR2_X1 U10096 ( .A1(n12732), .A2(n11557), .ZN(n11137) );
  NOR2_X1 U10097 ( .A1(n15529), .A2(n11449), .ZN(n15862) );
  INV_X1 U10098 ( .A(n10222), .ZN(n14990) );
  AND2_X1 U10099 ( .A1(n14860), .A2(n16012), .ZN(n14958) );
  INV_X1 U10100 ( .A(n14997), .ZN(n15942) );
  AND2_X1 U10101 ( .A1(n10041), .A2(n10166), .ZN(n16134) );
  INV_X1 U10102 ( .A(n16134), .ZN(n16019) );
  AND3_X1 U10103 ( .A1(n11560), .A2(n11549), .A3(n11548), .ZN(n11581) );
  AND2_X1 U10104 ( .A1(n9964), .A2(n9963), .ZN(n15832) );
  INV_X1 U10105 ( .A(n13564), .ZN(n12382) );
  NAND2_X1 U10106 ( .A1(n11235), .A2(n11234), .ZN(n13566) );
  AND4_X1 U10107 ( .A1(n9686), .A2(n9586), .A3(n9585), .A4(n9584), .ZN(n13610)
         );
  OAI211_X1 U10108 ( .C1(n9160), .C2(n9451), .A(n9450), .B(n9449), .ZN(n13687)
         );
  INV_X1 U10109 ( .A(n12776), .ZN(n13577) );
  INV_X1 U10110 ( .A(n15845), .ZN(n15830) );
  NAND2_X1 U10111 ( .A1(n13715), .A2(n15974), .ZN(n13717) );
  INV_X1 U10112 ( .A(n13117), .ZN(n13768) );
  NAND2_X1 U10113 ( .A1(n16165), .A2(n16107), .ZN(n13806) );
  INV_X1 U10114 ( .A(n13591), .ZN(n13821) );
  INV_X1 U10115 ( .A(n13560), .ZN(n13832) );
  INV_X1 U10116 ( .A(n16169), .ZN(n16166) );
  NAND2_X1 U10117 ( .A1(n10990), .A2(n13870), .ZN(n10991) );
  INV_X1 U10118 ( .A(SI_25_), .ZN(n15290) );
  INV_X1 U10119 ( .A(SI_15_), .ZN(n15305) );
  OR2_X1 U10120 ( .A1(n14001), .A2(n11781), .ZN(n13897) );
  OR2_X1 U10121 ( .A1(n13984), .A2(n14189), .ZN(n13992) );
  OR2_X1 U10122 ( .A1(n13984), .A2(n14191), .ZN(n13996) );
  INV_X1 U10123 ( .A(n13999), .ZN(n13978) );
  NAND2_X1 U10124 ( .A1(n10869), .A2(n10868), .ZN(n14005) );
  INV_X1 U10125 ( .A(n15504), .ZN(n15468) );
  INV_X1 U10126 ( .A(n15512), .ZN(n15412) );
  INV_X1 U10127 ( .A(n14151), .ZN(n14244) );
  AND2_X1 U10128 ( .A1(n11716), .A2(n11715), .ZN(n15993) );
  OR2_X1 U10129 ( .A1(n15406), .A2(n15403), .ZN(n15404) );
  AND2_X1 U10130 ( .A1(n11472), .A2(n15409), .ZN(n15401) );
  XNOR2_X1 U10131 ( .A(n10920), .B(n10919), .ZN(n12628) );
  INV_X1 U10132 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11364) );
  XNOR2_X1 U10133 ( .A(n9054), .B(n9053), .ZN(n11845) );
  NAND2_X1 U10134 ( .A1(n11849), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16203) );
  INV_X1 U10135 ( .A(n15077), .ZN(n14952) );
  INV_X1 U10136 ( .A(n7185), .ZN(n14717) );
  INV_X1 U10137 ( .A(n14595), .ZN(n14745) );
  OR2_X1 U10138 ( .A1(n8805), .A2(n8804), .ZN(n14755) );
  INV_X1 U10139 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15875) );
  INV_X1 U10140 ( .A(n15526), .ZN(n15876) );
  OR2_X1 U10141 ( .A1(n15894), .A2(n16134), .ZN(n15003) );
  OR2_X1 U10142 ( .A1(n15894), .A2(n12153), .ZN(n15029) );
  OR3_X1 U10143 ( .A1(n15116), .A2(n15115), .A3(n15114), .ZN(n15146) );
  INV_X1 U10144 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11971) );
  INV_X1 U10145 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n11362) );
  XNOR2_X1 U10146 ( .A(n10345), .B(n10344), .ZN(n15608) );
  AND2_X2 U10147 ( .A1(n11845), .A2(n10969), .ZN(P1_U4016) );
  NAND2_X1 U10148 ( .A1(n8417), .A2(SI_1_), .ZN(n8420) );
  INV_X1 U10149 ( .A(n8551), .ZN(n8419) );
  INV_X1 U10150 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9095) );
  MUX2_X1 U10151 ( .A(n9095), .B(n10526), .S(n8424), .Z(n8418) );
  NOR2_X1 U10152 ( .A1(n8418), .A2(n15267), .ZN(n8549) );
  NAND2_X1 U10153 ( .A1(n8419), .A2(n8549), .ZN(n8553) );
  NAND2_X1 U10154 ( .A1(n8553), .A2(n8420), .ZN(n8571) );
  INV_X1 U10155 ( .A(n8572), .ZN(n8422) );
  NAND2_X1 U10156 ( .A1(n8571), .A2(n8422), .ZN(n8574) );
  NAND2_X1 U10157 ( .A1(n8574), .A2(n8423), .ZN(n8589) );
  INV_X1 U10158 ( .A(n8427), .ZN(n8616) );
  NAND2_X1 U10159 ( .A1(n8618), .A2(n8428), .ZN(n8632) );
  MUX2_X1 U10160 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8504), .Z(n8429) );
  NAND2_X1 U10161 ( .A1(n8429), .A2(SI_6_), .ZN(n8431) );
  OAI21_X1 U10162 ( .B1(SI_6_), .B2(n8429), .A(n8431), .ZN(n8430) );
  INV_X1 U10163 ( .A(n8430), .ZN(n8631) );
  MUX2_X1 U10164 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8504), .Z(n8432) );
  NAND2_X1 U10165 ( .A1(n8432), .A2(SI_7_), .ZN(n8434) );
  OAI21_X1 U10166 ( .B1(SI_7_), .B2(n8432), .A(n8434), .ZN(n8433) );
  INV_X1 U10167 ( .A(n8433), .ZN(n8648) );
  MUX2_X1 U10168 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n8504), .Z(n8435) );
  NAND2_X1 U10169 ( .A1(n8435), .A2(SI_8_), .ZN(n8437) );
  OAI21_X1 U10170 ( .B1(SI_8_), .B2(n8435), .A(n8437), .ZN(n8436) );
  INV_X1 U10171 ( .A(n8436), .ZN(n8665) );
  MUX2_X1 U10172 ( .A(n11040), .B(n11039), .S(n8504), .Z(n8683) );
  NOR2_X1 U10173 ( .A1(n8683), .A2(n8682), .ZN(n8441) );
  MUX2_X1 U10174 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8504), .Z(n8438) );
  NAND2_X1 U10175 ( .A1(n8438), .A2(SI_10_), .ZN(n8442) );
  OAI21_X1 U10176 ( .B1(SI_10_), .B2(n8438), .A(n8442), .ZN(n8701) );
  INV_X1 U10177 ( .A(n8683), .ZN(n8439) );
  NOR2_X1 U10178 ( .A1(n8439), .A2(SI_9_), .ZN(n8440) );
  MUX2_X1 U10179 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n8504), .Z(n8443) );
  XNOR2_X1 U10180 ( .A(n8443), .B(SI_11_), .ZN(n8719) );
  INV_X1 U10181 ( .A(n8443), .ZN(n8444) );
  NAND2_X1 U10182 ( .A1(n8444), .A2(n15313), .ZN(n8445) );
  MUX2_X1 U10183 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n8504), .Z(n8446) );
  XNOR2_X1 U10184 ( .A(n8446), .B(n15307), .ZN(n8737) );
  INV_X1 U10185 ( .A(n8446), .ZN(n8447) );
  MUX2_X1 U10186 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n8504), .Z(n8448) );
  OAI21_X1 U10187 ( .B1(SI_13_), .B2(n8448), .A(n8449), .ZN(n8752) );
  MUX2_X1 U10188 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n8504), .Z(n8450) );
  XNOR2_X1 U10189 ( .A(n8450), .B(SI_14_), .ZN(n8771) );
  INV_X1 U10190 ( .A(n8450), .ZN(n8451) );
  NAND2_X1 U10191 ( .A1(n8451), .A2(n11037), .ZN(n8452) );
  MUX2_X1 U10192 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n8504), .Z(n8453) );
  XNOR2_X1 U10193 ( .A(n8453), .B(n15305), .ZN(n8790) );
  INV_X1 U10194 ( .A(n8453), .ZN(n8454) );
  MUX2_X1 U10195 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n8504), .Z(n8455) );
  OAI21_X1 U10196 ( .B1(SI_16_), .B2(n8455), .A(n8456), .ZN(n8807) );
  MUX2_X1 U10197 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10986), .Z(n8458) );
  XNOR2_X1 U10198 ( .A(n8458), .B(SI_17_), .ZN(n8825) );
  INV_X1 U10199 ( .A(n8458), .ZN(n8459) );
  NAND2_X1 U10200 ( .A1(n8459), .A2(n15275), .ZN(n8460) );
  MUX2_X1 U10201 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10986), .Z(n8844) );
  NOR2_X1 U10202 ( .A1(n8844), .A2(SI_18_), .ZN(n8463) );
  MUX2_X1 U10203 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10986), .Z(n8464) );
  XNOR2_X1 U10204 ( .A(n8464), .B(SI_19_), .ZN(n8861) );
  INV_X1 U10205 ( .A(n8844), .ZN(n8842) );
  NOR2_X1 U10206 ( .A1(n8842), .A2(n11424), .ZN(n8461) );
  NOR2_X1 U10207 ( .A1(n8861), .A2(n8461), .ZN(n8462) );
  INV_X1 U10208 ( .A(n8464), .ZN(n8465) );
  MUX2_X1 U10209 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n10986), .Z(n8466) );
  XNOR2_X1 U10210 ( .A(n8466), .B(n11731), .ZN(n8880) );
  INV_X1 U10211 ( .A(n8466), .ZN(n8467) );
  MUX2_X1 U10212 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10986), .Z(n8468) );
  NAND2_X1 U10213 ( .A1(n8468), .A2(SI_21_), .ZN(n8469) );
  OAI21_X1 U10214 ( .B1(SI_21_), .B2(n8468), .A(n8469), .ZN(n8892) );
  MUX2_X1 U10215 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10986), .Z(n10789) );
  INV_X1 U10216 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8470) );
  MUX2_X1 U10217 ( .A(n8470), .B(n9501), .S(n10986), .Z(n8473) );
  NAND2_X1 U10218 ( .A1(n8473), .A2(n15172), .ZN(n8533) );
  OAI21_X1 U10219 ( .B1(SI_22_), .B2(n10789), .A(n8533), .ZN(n8471) );
  INV_X1 U10220 ( .A(n8471), .ZN(n8472) );
  NAND3_X1 U10221 ( .A1(n8533), .A2(n10789), .A3(SI_22_), .ZN(n8475) );
  INV_X1 U10222 ( .A(n8473), .ZN(n8474) );
  NAND2_X1 U10223 ( .A1(n8474), .A2(SI_23_), .ZN(n8532) );
  MUX2_X1 U10224 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8504), .Z(n8476) );
  NAND2_X1 U10225 ( .A1(n8476), .A2(SI_24_), .ZN(n8478) );
  OAI21_X1 U10226 ( .B1(SI_24_), .B2(n8476), .A(n8478), .ZN(n8477) );
  INV_X1 U10227 ( .A(n8477), .ZN(n8908) );
  MUX2_X1 U10228 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10986), .Z(n8479) );
  XNOR2_X1 U10229 ( .A(n8479), .B(SI_25_), .ZN(n8921) );
  INV_X1 U10230 ( .A(n8479), .ZN(n8480) );
  MUX2_X1 U10231 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10986), .Z(n8481) );
  NAND2_X1 U10232 ( .A1(n8481), .A2(SI_26_), .ZN(n8483) );
  OAI21_X1 U10233 ( .B1(SI_26_), .B2(n8481), .A(n8483), .ZN(n8933) );
  INV_X1 U10234 ( .A(n8933), .ZN(n8482) );
  INV_X1 U10235 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13008) );
  INV_X1 U10236 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13011) );
  MUX2_X1 U10237 ( .A(n13008), .B(n13011), .S(n10986), .Z(n8959) );
  INV_X1 U10238 ( .A(n8959), .ZN(n8484) );
  XNOR2_X1 U10239 ( .A(n8484), .B(SI_27_), .ZN(n8485) );
  NOR2_X1 U10240 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8489) );
  NOR2_X1 U10241 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8498) );
  NAND2_X1 U10242 ( .A1(n13007), .A2(n10171), .ZN(n8506) );
  NAND2_X1 U10243 ( .A1(n8972), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U10244 ( .A1(n10157), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8523) );
  INV_X1 U10245 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n13077) );
  OR2_X1 U10246 ( .A1(n8976), .A2(n13077), .ZN(n8522) );
  NAND2_X1 U10247 ( .A1(n8608), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8640) );
  NOR2_X1 U10248 ( .A1(n8640), .A2(n8639), .ZN(n8638) );
  NAND2_X1 U10249 ( .A1(n8638), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U10250 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n8513) );
  NAND2_X1 U10251 ( .A1(n8799), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8833) );
  INV_X1 U10252 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8832) );
  INV_X1 U10253 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14688) );
  NAND2_X1 U10254 ( .A1(n8538), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U10255 ( .A1(n8914), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U10256 ( .A1(n8926), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8925) );
  INV_X1 U10257 ( .A(n8947), .ZN(n8949) );
  INV_X1 U10258 ( .A(n8514), .ZN(n8940) );
  INV_X1 U10259 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10260 ( .A1(n8940), .A2(n8515), .ZN(n8516) );
  NAND2_X1 U10261 ( .A1(n8949), .A2(n8516), .ZN(n14536) );
  OR2_X1 U10262 ( .A1(n8609), .A2(n14536), .ZN(n8521) );
  INV_X1 U10263 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8519) );
  OR2_X1 U10264 ( .A1(n10161), .A2(n8519), .ZN(n8520) );
  OAI21_X1 U10265 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8538), .A(n8524), .ZN(
        n14935) );
  OR2_X1 U10266 ( .A1(n8977), .A2(n14935), .ZN(n8529) );
  NAND2_X1 U10267 ( .A1(n8951), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8528) );
  INV_X1 U10268 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8525) );
  OR2_X1 U10269 ( .A1(n8953), .A2(n8525), .ZN(n8527) );
  INV_X1 U10270 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14938) );
  OR2_X1 U10271 ( .A1(n8976), .A2(n14938), .ZN(n8526) );
  NAND4_X1 U10272 ( .A1(n8529), .A2(n8528), .A3(n8527), .A4(n8526), .ZN(n14912) );
  INV_X1 U10273 ( .A(n14912), .ZN(n14686) );
  NAND2_X1 U10274 ( .A1(n10788), .A2(n10789), .ZN(n10793) );
  NAND2_X1 U10275 ( .A1(n8530), .A2(SI_22_), .ZN(n8531) );
  NAND2_X1 U10276 ( .A1(n10793), .A2(n8531), .ZN(n8535) );
  NAND2_X1 U10277 ( .A1(n8533), .A2(n8532), .ZN(n8534) );
  NAND2_X1 U10278 ( .A1(n12731), .A2(n10171), .ZN(n8537) );
  NAND2_X1 U10279 ( .A1(n8972), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U10280 ( .A1(n8951), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8544) );
  AOI21_X1 U10281 ( .B1(n8899), .B2(n14688), .A(n8538), .ZN(n14948) );
  NAND2_X1 U10282 ( .A1(n8901), .A2(n14948), .ZN(n8543) );
  INV_X1 U10283 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8539) );
  OR2_X1 U10284 ( .A1(n8953), .A2(n8539), .ZN(n8542) );
  INV_X1 U10285 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8540) );
  OR2_X1 U10286 ( .A1(n8976), .A2(n8540), .ZN(n8541) );
  NAND4_X1 U10287 ( .A1(n8544), .A2(n8543), .A3(n8542), .A4(n8541), .ZN(n14748) );
  INV_X1 U10288 ( .A(n14748), .ZN(n14490) );
  NAND2_X1 U10289 ( .A1(n10788), .A2(n8421), .ZN(n8545) );
  XNOR2_X1 U10290 ( .A(n8545), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15163) );
  INV_X1 U10291 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8546) );
  INV_X1 U10292 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11148) );
  OR2_X1 U10293 ( .A1(n8976), .A2(n11148), .ZN(n8547) );
  INV_X1 U10294 ( .A(n8564), .ZN(n8555) );
  INV_X1 U10295 ( .A(n8549), .ZN(n8550) );
  NAND2_X1 U10296 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  NAND2_X1 U10297 ( .A1(n8553), .A2(n8552), .ZN(n11020) );
  INV_X1 U10298 ( .A(n8554), .ZN(n8576) );
  INV_X1 U10299 ( .A(n11147), .ZN(n14773) );
  NAND2_X1 U10300 ( .A1(n8951), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8561) );
  INV_X1 U10301 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8556) );
  INV_X1 U10302 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11748) );
  OR2_X1 U10303 ( .A1(n8977), .A2(n11748), .ZN(n8559) );
  INV_X1 U10304 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8557) );
  OR2_X1 U10305 ( .A1(n8976), .A2(n8557), .ZN(n8558) );
  NOR2_X1 U10306 ( .A1(n10986), .A2(n15267), .ZN(n8562) );
  XNOR2_X1 U10307 ( .A(n8562), .B(n9095), .ZN(n15399) );
  MUX2_X1 U10308 ( .A(n15398), .B(n15399), .S(n8563), .Z(n15914) );
  INV_X1 U10309 ( .A(n15914), .ZN(n15888) );
  NAND2_X1 U10310 ( .A1(n8555), .A2(n15934), .ZN(n8565) );
  NAND2_X1 U10311 ( .A1(n8951), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8570) );
  INV_X1 U10312 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8566) );
  INV_X1 U10313 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n12279) );
  OR2_X1 U10314 ( .A1(n8609), .A2(n12279), .ZN(n8568) );
  INV_X1 U10315 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U10316 ( .A1(n8573), .A2(n8572), .ZN(n8575) );
  NAND2_X1 U10317 ( .A1(n8575), .A2(n8574), .ZN(n11022) );
  NAND2_X1 U10318 ( .A1(n8576), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8577) );
  MUX2_X1 U10319 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8577), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n8579) );
  INV_X1 U10320 ( .A(n8578), .ZN(n8592) );
  NAND2_X1 U10321 ( .A1(n8579), .A2(n8592), .ZN(n11150) );
  INV_X1 U10322 ( .A(n11150), .ZN(n11436) );
  NAND2_X1 U10323 ( .A1(n11032), .A2(n11436), .ZN(n8580) );
  OR2_X1 U10324 ( .A1(n8609), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U10325 ( .A1(n8951), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8586) );
  INV_X1 U10326 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8583) );
  OR2_X1 U10327 ( .A1(n8953), .A2(n8583), .ZN(n8585) );
  INV_X1 U10328 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11152) );
  OR2_X1 U10329 ( .A1(n8976), .A2(n11152), .ZN(n8584) );
  OR2_X1 U10330 ( .A1(n8589), .A2(n8588), .ZN(n8590) );
  NAND2_X1 U10331 ( .A1(n15395), .A2(n10171), .ZN(n8595) );
  NAND2_X1 U10332 ( .A1(n8592), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8591) );
  MUX2_X1 U10333 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8591), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8593) );
  AND2_X1 U10334 ( .A1(n8593), .A2(n8602), .ZN(n15393) );
  AOI22_X1 U10335 ( .A1(n8972), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n11032), 
        .B2(n15393), .ZN(n8594) );
  XNOR2_X1 U10336 ( .A(n14767), .B(n14566), .ZN(n11584) );
  INV_X1 U10337 ( .A(n11584), .ZN(n11583) );
  INV_X1 U10338 ( .A(n14767), .ZN(n12276) );
  NAND2_X1 U10339 ( .A1(n12276), .A2(n11825), .ZN(n8596) );
  OR2_X1 U10340 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  AND2_X1 U10341 ( .A1(n8600), .A2(n8599), .ZN(n10981) );
  NAND2_X1 U10342 ( .A1(n10981), .A2(n10171), .ZN(n8607) );
  NAND2_X1 U10343 ( .A1(n8602), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8601) );
  MUX2_X1 U10344 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8601), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n8605) );
  INV_X1 U10345 ( .A(n8602), .ZN(n8604) );
  INV_X1 U10346 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U10347 ( .A1(n8604), .A2(n8603), .ZN(n8635) );
  NAND2_X1 U10348 ( .A1(n8605), .A2(n8635), .ZN(n15863) );
  INV_X1 U10349 ( .A(n15863), .ZN(n15861) );
  AOI22_X1 U10350 ( .A1(n8972), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11032), 
        .B2(n15861), .ZN(n8606) );
  INV_X1 U10351 ( .A(n8608), .ZN(n8623) );
  OAI21_X1 U10352 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n8623), .ZN(n11843) );
  OR2_X1 U10353 ( .A1(n8609), .A2(n11843), .ZN(n8614) );
  NAND2_X1 U10354 ( .A1(n8951), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8613) );
  INV_X1 U10355 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8610) );
  OR2_X1 U10356 ( .A1(n8953), .A2(n8610), .ZN(n8612) );
  INV_X1 U10357 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11155) );
  OR2_X1 U10358 ( .A1(n8976), .A2(n11155), .ZN(n8611) );
  NAND4_X1 U10359 ( .A1(n8614), .A2(n8613), .A3(n8612), .A4(n8611), .ZN(n14766) );
  NOR2_X1 U10360 ( .A1(n16008), .A2(n14766), .ZN(n8615) );
  INV_X1 U10361 ( .A(n16008), .ZN(n12299) );
  NAND2_X1 U10362 ( .A1(n8618), .A2(n8617), .ZN(n10984) );
  OR2_X1 U10363 ( .A1(n10984), .A2(n8937), .ZN(n8621) );
  NAND2_X1 U10364 ( .A1(n8635), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8619) );
  XNOR2_X1 U10365 ( .A(n8619), .B(P1_IR_REG_5__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U10366 ( .A1(n8972), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11032), 
        .B2(n11263), .ZN(n8620) );
  INV_X1 U10367 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U10368 ( .A1(n8623), .A2(n8622), .ZN(n8624) );
  NAND2_X1 U10369 ( .A1(n8640), .A2(n8624), .ZN(n12156) );
  OR2_X1 U10370 ( .A1(n8609), .A2(n12156), .ZN(n8629) );
  NAND2_X1 U10371 ( .A1(n8951), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8628) );
  INV_X1 U10372 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n8625) );
  OR2_X1 U10373 ( .A1(n8953), .A2(n8625), .ZN(n8627) );
  INV_X1 U10374 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n12160) );
  OR2_X1 U10375 ( .A1(n8976), .A2(n12160), .ZN(n8626) );
  XNOR2_X1 U10376 ( .A(n12159), .B(n14765), .ZN(n11628) );
  INV_X1 U10377 ( .A(n12159), .ZN(n9025) );
  INV_X1 U10378 ( .A(n14765), .ZN(n12292) );
  NAND2_X1 U10379 ( .A1(n9025), .A2(n12292), .ZN(n8630) );
  OR2_X1 U10380 ( .A1(n8632), .A2(n8631), .ZN(n8633) );
  NAND2_X1 U10381 ( .A1(n8652), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8636) );
  XNOR2_X1 U10382 ( .A(n8636), .B(P1_IR_REG_6__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U10383 ( .A1(n8972), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11032), 
        .B2(n11211), .ZN(n8637) );
  INV_X1 U10384 ( .A(n8638), .ZN(n8657) );
  NAND2_X1 U10385 ( .A1(n8640), .A2(n8639), .ZN(n8641) );
  NAND2_X1 U10386 ( .A1(n8657), .A2(n8641), .ZN(n12014) );
  OR2_X1 U10387 ( .A1(n8977), .A2(n12014), .ZN(n8646) );
  NAND2_X1 U10388 ( .A1(n8951), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8645) );
  INV_X1 U10389 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8642) );
  OR2_X1 U10390 ( .A1(n8953), .A2(n8642), .ZN(n8644) );
  INV_X1 U10391 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11160) );
  OR2_X1 U10392 ( .A1(n8976), .A2(n11160), .ZN(n8643) );
  NAND4_X1 U10393 ( .A1(n8646), .A2(n8645), .A3(n8644), .A4(n8643), .ZN(n14764) );
  XNOR2_X1 U10394 ( .A(n12437), .B(n14764), .ZN(n11803) );
  INV_X1 U10395 ( .A(n11803), .ZN(n11798) );
  OR2_X1 U10396 ( .A1(n12437), .A2(n14764), .ZN(n8647) );
  OR2_X1 U10397 ( .A1(n8649), .A2(n8648), .ZN(n8651) );
  NAND2_X1 U10398 ( .A1(n8651), .A2(n8650), .ZN(n11019) );
  OR2_X1 U10399 ( .A1(n11019), .A2(n8937), .ZN(n8655) );
  OAI21_X1 U10400 ( .B1(n8652), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8653) );
  XNOR2_X1 U10401 ( .A(n8653), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U10402 ( .A1(n8972), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11032), 
        .B2(n11295), .ZN(n8654) );
  NAND2_X1 U10403 ( .A1(n8655), .A2(n8654), .ZN(n12129) );
  INV_X1 U10404 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U10405 ( .A1(n8657), .A2(n8656), .ZN(n8658) );
  NAND2_X1 U10406 ( .A1(n8692), .A2(n8658), .ZN(n12241) );
  OR2_X1 U10407 ( .A1(n8609), .A2(n12241), .ZN(n8663) );
  NAND2_X1 U10408 ( .A1(n8951), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8662) );
  INV_X1 U10409 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8659) );
  OR2_X1 U10410 ( .A1(n8953), .A2(n8659), .ZN(n8661) );
  INV_X1 U10411 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n12242) );
  OR2_X1 U10412 ( .A1(n8976), .A2(n12242), .ZN(n8660) );
  NAND4_X1 U10413 ( .A1(n8663), .A2(n8662), .A3(n8661), .A4(n8660), .ZN(n14763) );
  XNOR2_X1 U10414 ( .A(n12129), .B(n14763), .ZN(n10211) );
  INV_X1 U10415 ( .A(n10211), .ZN(n12125) );
  OR2_X1 U10416 ( .A1(n12129), .A2(n14763), .ZN(n8664) );
  NAND2_X1 U10417 ( .A1(n8668), .A2(n8667), .ZN(n10483) );
  OR2_X1 U10418 ( .A1(n10483), .A2(n8937), .ZN(n8674) );
  INV_X1 U10419 ( .A(n8792), .ZN(n8669) );
  NAND2_X1 U10420 ( .A1(n8669), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8670) );
  MUX2_X1 U10421 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8670), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n8672) );
  INV_X1 U10422 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U10423 ( .A1(n8792), .A2(n8671), .ZN(n8687) );
  NAND2_X1 U10424 ( .A1(n8672), .A2(n8687), .ZN(n11321) );
  INV_X1 U10425 ( .A(n11321), .ZN(n11298) );
  AOI22_X1 U10426 ( .A1(n8972), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11032), 
        .B2(n11298), .ZN(n8673) );
  NAND2_X1 U10427 ( .A1(n8674), .A2(n8673), .ZN(n16076) );
  INV_X1 U10428 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8691) );
  XNOR2_X1 U10429 ( .A(n8692), .B(n8691), .ZN(n12350) );
  OR2_X1 U10430 ( .A1(n8977), .A2(n12350), .ZN(n8679) );
  NAND2_X1 U10431 ( .A1(n8951), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8678) );
  INV_X1 U10432 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8675) );
  OR2_X1 U10433 ( .A1(n8953), .A2(n8675), .ZN(n8677) );
  INV_X1 U10434 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n12260) );
  OR2_X1 U10435 ( .A1(n8976), .A2(n12260), .ZN(n8676) );
  NAND4_X1 U10436 ( .A1(n8679), .A2(n8678), .A3(n8677), .A4(n8676), .ZN(n14762) );
  INV_X1 U10437 ( .A(n14762), .ZN(n14656) );
  XNOR2_X1 U10438 ( .A(n16076), .B(n14656), .ZN(n12252) );
  NAND2_X1 U10439 ( .A1(n12253), .A2(n12252), .ZN(n12251) );
  OR2_X1 U10440 ( .A1(n16076), .A2(n14762), .ZN(n8680) );
  INV_X1 U10441 ( .A(SI_9_), .ZN(n8682) );
  NAND2_X1 U10442 ( .A1(n8684), .A2(n8683), .ZN(n8685) );
  NAND2_X1 U10443 ( .A1(n8687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8686) );
  MUX2_X1 U10444 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8686), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n8688) );
  AOI22_X1 U10445 ( .A1(n8972), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11032), 
        .B2(n11334), .ZN(n8689) );
  INV_X1 U10446 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8690) );
  OAI21_X1 U10447 ( .B1(n8692), .B2(n8691), .A(n8690), .ZN(n8693) );
  NAND2_X1 U10448 ( .A1(n8693), .A2(n8711), .ZN(n14659) );
  OR2_X1 U10449 ( .A1(n8609), .A2(n14659), .ZN(n8698) );
  NAND2_X1 U10450 ( .A1(n8951), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8697) );
  INV_X1 U10451 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8694) );
  OR2_X1 U10452 ( .A1(n8953), .A2(n8694), .ZN(n8696) );
  INV_X1 U10453 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n12326) );
  OR2_X1 U10454 ( .A1(n8976), .A2(n12326), .ZN(n8695) );
  NAND4_X1 U10455 ( .A1(n8698), .A2(n8697), .A3(n8696), .A4(n8695), .ZN(n14761) );
  INV_X1 U10456 ( .A(n14761), .ZN(n14397) );
  NAND2_X1 U10457 ( .A1(n14661), .A2(n14397), .ZN(n9004) );
  OR2_X1 U10458 ( .A1(n14661), .A2(n14397), .ZN(n8699) );
  OR2_X1 U10459 ( .A1(n14661), .A2(n14761), .ZN(n8700) );
  AND2_X1 U10460 ( .A1(n8702), .A2(n8701), .ZN(n8703) );
  NAND2_X1 U10461 ( .A1(n8721), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8707) );
  XNOR2_X1 U10462 ( .A(n8707), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U10463 ( .A1(n8972), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11032), 
        .B2(n11528), .ZN(n8708) );
  INV_X1 U10464 ( .A(n8710), .ZN(n8729) );
  NAND2_X1 U10465 ( .A1(n8711), .A2(n11332), .ZN(n8712) );
  NAND2_X1 U10466 ( .A1(n8729), .A2(n8712), .ZN(n14558) );
  OR2_X1 U10467 ( .A1(n8977), .A2(n14558), .ZN(n8717) );
  NAND2_X1 U10468 ( .A1(n8951), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8716) );
  INV_X1 U10469 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8713) );
  OR2_X1 U10470 ( .A1(n8953), .A2(n8713), .ZN(n8715) );
  INV_X1 U10471 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11335) );
  OR2_X1 U10472 ( .A1(n8976), .A2(n11335), .ZN(n8714) );
  NAND4_X1 U10473 ( .A1(n8717), .A2(n8716), .A3(n8715), .A4(n8714), .ZN(n14760) );
  OR2_X1 U10474 ( .A1(n14560), .A2(n14760), .ZN(n8718) );
  XNOR2_X1 U10475 ( .A(n8720), .B(n8719), .ZN(n11186) );
  NAND2_X1 U10476 ( .A1(n11186), .A2(n10171), .ZN(n8726) );
  INV_X1 U10477 ( .A(n8721), .ZN(n8723) );
  INV_X1 U10478 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U10479 ( .A1(n8723), .A2(n8722), .ZN(n8739) );
  NAND2_X1 U10480 ( .A1(n8739), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8724) );
  XNOR2_X1 U10481 ( .A(n8724), .B(P1_IR_REG_11__SCAN_IN), .ZN(n14805) );
  AOI22_X1 U10482 ( .A1(n8972), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11032), 
        .B2(n14805), .ZN(n8725) );
  NAND2_X1 U10483 ( .A1(n8726), .A2(n8725), .ZN(n14703) );
  INV_X1 U10484 ( .A(n8727), .ZN(n8744) );
  INV_X1 U10485 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U10486 ( .A1(n8729), .A2(n8728), .ZN(n8730) );
  NAND2_X1 U10487 ( .A1(n8744), .A2(n8730), .ZN(n14701) );
  OR2_X1 U10488 ( .A1(n8977), .A2(n14701), .ZN(n8735) );
  NAND2_X1 U10489 ( .A1(n8951), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8734) );
  INV_X1 U10490 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8731) );
  OR2_X1 U10491 ( .A1(n8953), .A2(n8731), .ZN(n8733) );
  INV_X1 U10492 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n12397) );
  OR2_X1 U10493 ( .A1(n8976), .A2(n12397), .ZN(n8732) );
  NAND4_X1 U10494 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n14759) );
  XNOR2_X1 U10495 ( .A(n14703), .B(n14759), .ZN(n10215) );
  INV_X1 U10496 ( .A(n10215), .ZN(n12401) );
  OR2_X1 U10497 ( .A1(n14703), .A2(n14759), .ZN(n8736) );
  XNOR2_X1 U10498 ( .A(n8738), .B(n8737), .ZN(n11361) );
  NAND2_X1 U10499 ( .A1(n11361), .A2(n10171), .ZN(n8742) );
  NAND2_X1 U10500 ( .A1(n8740), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8757) );
  XNOR2_X1 U10501 ( .A(n8757), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U10502 ( .A1(n8972), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11032), 
        .B2(n11815), .ZN(n8741) );
  INV_X1 U10503 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U10504 ( .A1(n8744), .A2(n8743), .ZN(n8745) );
  NAND2_X1 U10505 ( .A1(n8762), .A2(n8745), .ZN(n14613) );
  OR2_X1 U10506 ( .A1(n8609), .A2(n14613), .ZN(n8750) );
  NAND2_X1 U10507 ( .A1(n8951), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8749) );
  INV_X1 U10508 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8746) );
  OR2_X1 U10509 ( .A1(n8953), .A2(n8746), .ZN(n8748) );
  INV_X1 U10510 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12464) );
  OR2_X1 U10511 ( .A1(n8976), .A2(n12464), .ZN(n8747) );
  NAND4_X1 U10512 ( .A1(n8750), .A2(n8749), .A3(n8748), .A4(n8747), .ZN(n14758) );
  XNOR2_X1 U10513 ( .A(n14387), .B(n14758), .ZN(n12459) );
  INV_X1 U10514 ( .A(n12459), .ZN(n12455) );
  OR2_X1 U10515 ( .A1(n14387), .A2(n14758), .ZN(n8751) );
  NAND2_X1 U10516 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  NAND2_X1 U10517 ( .A1(n8755), .A2(n8754), .ZN(n11394) );
  OR2_X1 U10518 ( .A1(n11394), .A2(n8937), .ZN(n8760) );
  INV_X1 U10519 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U10520 ( .A1(n8757), .A2(n8756), .ZN(n8758) );
  NAND2_X1 U10521 ( .A1(n8758), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8774) );
  XNOR2_X1 U10522 ( .A(n8774), .B(P1_IR_REG_13__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U10523 ( .A1(n8972), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n12115), 
        .B2(n11032), .ZN(n8759) );
  NAND2_X1 U10524 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  NAND2_X1 U10525 ( .A1(n8780), .A2(n8763), .ZN(n14677) );
  OR2_X1 U10526 ( .A1(n8977), .A2(n14677), .ZN(n8769) );
  NAND2_X1 U10527 ( .A1(n8951), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8768) );
  INV_X1 U10528 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8764) );
  OR2_X1 U10529 ( .A1(n8953), .A2(n8764), .ZN(n8767) );
  INV_X1 U10530 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8765) );
  OR2_X1 U10531 ( .A1(n8976), .A2(n8765), .ZN(n8766) );
  NAND4_X1 U10532 ( .A1(n8769), .A2(n8768), .A3(n8767), .A4(n8766), .ZN(n14757) );
  INV_X1 U10533 ( .A(n14757), .ZN(n12457) );
  XNOR2_X1 U10534 ( .A(n14679), .B(n12457), .ZN(n12483) );
  OR2_X1 U10535 ( .A1(n14679), .A2(n14757), .ZN(n8770) );
  XNOR2_X1 U10536 ( .A(n8772), .B(n8771), .ZN(n11518) );
  NAND2_X1 U10537 ( .A1(n11518), .A2(n10171), .ZN(n8778) );
  INV_X1 U10538 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U10539 ( .A1(n8774), .A2(n8773), .ZN(n8775) );
  NAND2_X1 U10540 ( .A1(n8775), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8776) );
  XNOR2_X1 U10541 ( .A(n8776), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U10542 ( .A1(n12671), .A2(n11032), .B1(n8972), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U10543 ( .A1(n8951), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U10544 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  NAND2_X1 U10545 ( .A1(n8801), .A2(n8781), .ZN(n16180) );
  INV_X1 U10546 ( .A(n16180), .ZN(n12637) );
  NAND2_X1 U10547 ( .A1(n8901), .A2(n12637), .ZN(n8786) );
  INV_X1 U10548 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8782) );
  OR2_X1 U10549 ( .A1(n8953), .A2(n8782), .ZN(n8785) );
  INV_X1 U10550 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8783) );
  OR2_X1 U10551 ( .A1(n8976), .A2(n8783), .ZN(n8784) );
  NAND4_X1 U10552 ( .A1(n8787), .A2(n8786), .A3(n8785), .A4(n8784), .ZN(n14756) );
  XNOR2_X1 U10553 ( .A(n16177), .B(n14756), .ZN(n12633) );
  NAND2_X1 U10554 ( .A1(n16177), .A2(n14756), .ZN(n8789) );
  XNOR2_X1 U10555 ( .A(n8791), .B(n8790), .ZN(n11750) );
  NAND2_X1 U10556 ( .A1(n11750), .A2(n10171), .ZN(n8796) );
  NAND2_X1 U10557 ( .A1(n8811), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8793) );
  XNOR2_X1 U10558 ( .A(n8793), .B(n8810), .ZN(n15535) );
  INV_X1 U10559 ( .A(n15535), .ZN(n8794) );
  AOI22_X1 U10560 ( .A1(n8972), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11032), 
        .B2(n8794), .ZN(n8795) );
  INV_X1 U10561 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U10562 ( .A1(n10157), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8797) );
  OAI21_X1 U10563 ( .B1(n8798), .B2(n10161), .A(n8797), .ZN(n8805) );
  INV_X1 U10564 ( .A(n8799), .ZN(n8818) );
  NAND2_X1 U10565 ( .A1(n8801), .A2(n8800), .ZN(n8802) );
  NAND2_X1 U10566 ( .A1(n8818), .A2(n8802), .ZN(n14735) );
  NAND2_X1 U10567 ( .A1(n10156), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8803) );
  OAI21_X1 U10568 ( .B1(n14735), .B2(n8609), .A(n8803), .ZN(n8804) );
  XNOR2_X1 U10569 ( .A(n14738), .B(n14755), .ZN(n10218) );
  OR2_X1 U10570 ( .A1(n14738), .A2(n14755), .ZN(n8806) );
  INV_X1 U10571 ( .A(n8807), .ZN(n8808) );
  XNOR2_X1 U10572 ( .A(n8809), .B(n8808), .ZN(n11859) );
  NAND2_X1 U10573 ( .A1(n11859), .A2(n10171), .ZN(n8816) );
  NAND2_X1 U10574 ( .A1(n7323), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8812) );
  MUX2_X1 U10575 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8812), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8814) );
  NAND2_X1 U10576 ( .A1(n8814), .A2(n8828), .ZN(n12874) );
  INV_X1 U10577 ( .A(n12874), .ZN(n12871) );
  AOI22_X1 U10578 ( .A1(n8972), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11032), 
        .B2(n12871), .ZN(n8815) );
  INV_X1 U10579 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12866) );
  INV_X1 U10580 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U10581 ( .A1(n8818), .A2(n8817), .ZN(n8819) );
  NAND2_X1 U10582 ( .A1(n8833), .A2(n8819), .ZN(n16202) );
  OR2_X1 U10583 ( .A1(n16202), .A2(n8609), .ZN(n8823) );
  NAND2_X1 U10584 ( .A1(n8951), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U10585 ( .A1(n10157), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8820) );
  AND2_X1 U10586 ( .A1(n8821), .A2(n8820), .ZN(n8822) );
  OAI211_X1 U10587 ( .C1(n8976), .C2(n12866), .A(n8823), .B(n8822), .ZN(n14754) );
  INV_X1 U10588 ( .A(n14754), .ZN(n14438) );
  XNOR2_X1 U10589 ( .A(n16199), .B(n14438), .ZN(n12856) );
  OR2_X1 U10590 ( .A1(n16199), .A2(n14754), .ZN(n8824) );
  XNOR2_X1 U10591 ( .A(n8826), .B(n8825), .ZN(n11970) );
  NAND2_X1 U10592 ( .A1(n11970), .A2(n10171), .ZN(n8831) );
  NAND2_X1 U10593 ( .A1(n8828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8827) );
  MUX2_X1 U10594 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8827), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8829) );
  AND2_X1 U10595 ( .A1(n8829), .A2(n8863), .ZN(n14814) );
  AOI22_X1 U10596 ( .A1(n8972), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11032), 
        .B2(n14814), .ZN(n8830) );
  NAND2_X1 U10597 ( .A1(n8833), .A2(n8832), .ZN(n8834) );
  NAND2_X1 U10598 ( .A1(n8852), .A2(n8834), .ZN(n14636) );
  AOI22_X1 U10599 ( .A1(n8951), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n10157), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U10600 ( .A1(n10156), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8835) );
  OAI211_X1 U10601 ( .C1(n14636), .C2(n8977), .A(n8836), .B(n8835), .ZN(n14753) );
  XNOR2_X1 U10602 ( .A(n14449), .B(n14753), .ZN(n12934) );
  INV_X1 U10603 ( .A(n12934), .ZN(n8837) );
  NAND2_X1 U10604 ( .A1(n14449), .A2(n14753), .ZN(n8838) );
  NAND2_X1 U10605 ( .A1(n8839), .A2(n11424), .ZN(n8841) );
  NAND2_X1 U10606 ( .A1(n8840), .A2(SI_18_), .ZN(n8859) );
  INV_X1 U10607 ( .A(n8845), .ZN(n8843) );
  NAND2_X1 U10608 ( .A1(n8843), .A2(n8842), .ZN(n8846) );
  NAND2_X1 U10609 ( .A1(n8845), .A2(n8844), .ZN(n8860) );
  NAND2_X1 U10610 ( .A1(n12384), .A2(n10171), .ZN(n8849) );
  NAND2_X1 U10611 ( .A1(n8863), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8847) );
  XNOR2_X1 U10612 ( .A(n8847), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14826) );
  AOI22_X1 U10613 ( .A1(n8972), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11032), 
        .B2(n14826), .ZN(n8848) );
  INV_X1 U10614 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15020) );
  INV_X1 U10615 ( .A(n8850), .ZN(n8868) );
  NAND2_X1 U10616 ( .A1(n8852), .A2(n8851), .ZN(n8853) );
  NAND2_X1 U10617 ( .A1(n8868), .A2(n8853), .ZN(n15019) );
  OR2_X1 U10618 ( .A1(n15019), .A2(n8609), .ZN(n8855) );
  AOI22_X1 U10619 ( .A1(n8951), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n10157), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n8854) );
  OAI211_X1 U10620 ( .C1(n8976), .C2(n15020), .A(n8855), .B(n8854), .ZN(n14752) );
  XNOR2_X1 U10621 ( .A(n15025), .B(n14752), .ZN(n15004) );
  INV_X1 U10622 ( .A(n14752), .ZN(n8856) );
  NAND2_X1 U10623 ( .A1(n8860), .A2(n8859), .ZN(n8862) );
  XNOR2_X1 U10624 ( .A(n8862), .B(n8861), .ZN(n12469) );
  NAND2_X1 U10625 ( .A1(n12469), .A2(n10171), .ZN(n8866) );
  NAND2_X1 U10626 ( .A1(n7266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8864) );
  AOI22_X1 U10627 ( .A1(n8972), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14835), 
        .B2(n11032), .ZN(n8865) );
  INV_X1 U10628 ( .A(n8884), .ZN(n8870) );
  INV_X1 U10629 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U10630 ( .A1(n8868), .A2(n8867), .ZN(n8869) );
  NAND2_X1 U10631 ( .A1(n8870), .A2(n8869), .ZN(n14575) );
  OR2_X1 U10632 ( .A1(n14575), .A2(n8609), .ZN(n8876) );
  INV_X1 U10633 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U10634 ( .A1(n10156), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U10635 ( .A1(n10157), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8871) );
  OAI211_X1 U10636 ( .C1(n10161), .C2(n8873), .A(n8872), .B(n8871), .ZN(n8874)
         );
  INV_X1 U10637 ( .A(n8874), .ZN(n8875) );
  NAND2_X1 U10638 ( .A1(n8876), .A2(n8875), .ZN(n14751) );
  XNOR2_X1 U10639 ( .A(n15105), .B(n14751), .ZN(n10222) );
  NAND2_X1 U10640 ( .A1(n8878), .A2(n8877), .ZN(n8879) );
  XNOR2_X1 U10641 ( .A(n8881), .B(n8880), .ZN(n12388) );
  NAND2_X1 U10642 ( .A1(n12388), .A2(n10171), .ZN(n8883) );
  NAND2_X1 U10643 ( .A1(n8972), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8882) );
  NOR2_X1 U10644 ( .A1(n8884), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8885) );
  OR2_X1 U10645 ( .A1(n8898), .A2(n8885), .ZN(n14980) );
  INV_X1 U10646 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U10647 ( .A1(n10157), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U10648 ( .A1(n10156), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8886) );
  OAI211_X1 U10649 ( .C1(n8888), .C2(n10161), .A(n8887), .B(n8886), .ZN(n8889)
         );
  INV_X1 U10650 ( .A(n8889), .ZN(n8890) );
  OAI21_X1 U10651 ( .B1(n14980), .B2(n8977), .A(n8890), .ZN(n14750) );
  XNOR2_X1 U10652 ( .A(n15099), .B(n14750), .ZN(n14979) );
  NAND2_X1 U10653 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  NAND2_X1 U10654 ( .A1(n12478), .A2(n10171), .ZN(n8897) );
  NAND2_X1 U10655 ( .A1(n8972), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8896) );
  OR2_X1 U10656 ( .A1(n8898), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8900) );
  AND2_X1 U10657 ( .A1(n8900), .A2(n8899), .ZN(n14965) );
  NAND2_X1 U10658 ( .A1(n14965), .A2(n8901), .ZN(n8907) );
  INV_X1 U10659 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U10660 ( .A1(n10156), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U10661 ( .A1(n10157), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8902) );
  OAI211_X1 U10662 ( .C1(n10161), .C2(n8904), .A(n8903), .B(n8902), .ZN(n8905)
         );
  INV_X1 U10663 ( .A(n8905), .ZN(n8906) );
  NAND2_X1 U10664 ( .A1(n8907), .A2(n8906), .ZN(n14749) );
  INV_X1 U10665 ( .A(n14749), .ZN(n14666) );
  XNOR2_X1 U10666 ( .A(n15086), .B(n14666), .ZN(n14963) );
  XNOR2_X1 U10667 ( .A(n14952), .B(n14748), .ZN(n14945) );
  INV_X1 U10668 ( .A(n14945), .ZN(n14954) );
  XNOR2_X1 U10669 ( .A(n15073), .B(n14912), .ZN(n10225) );
  OR2_X1 U10670 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  NAND2_X1 U10671 ( .A1(n8972), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8912) );
  OAI21_X1 U10672 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8914), .A(n8913), .ZN(
        n14923) );
  OR2_X1 U10673 ( .A1(n8609), .A2(n14923), .ZN(n8919) );
  NAND2_X1 U10674 ( .A1(n8951), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8918) );
  INV_X1 U10675 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8915) );
  OR2_X1 U10676 ( .A1(n8953), .A2(n8915), .ZN(n8917) );
  INV_X1 U10677 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14924) );
  OR2_X1 U10678 ( .A1(n8976), .A2(n14924), .ZN(n8916) );
  NAND4_X1 U10679 ( .A1(n8919), .A2(n8918), .A3(n8917), .A4(n8916), .ZN(n14747) );
  INV_X1 U10680 ( .A(n15063), .ZN(n14922) );
  INV_X1 U10681 ( .A(n14747), .ZN(n14508) );
  XNOR2_X1 U10682 ( .A(n8922), .B(n8921), .ZN(n12648) );
  NAND2_X1 U10683 ( .A1(n12648), .A2(n10171), .ZN(n8924) );
  NAND2_X1 U10684 ( .A1(n8972), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8923) );
  OAI21_X1 U10685 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8926), .A(n8925), .ZN(
        n14904) );
  OR2_X1 U10686 ( .A1(n8609), .A2(n14904), .ZN(n8931) );
  NAND2_X1 U10687 ( .A1(n8951), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8930) );
  INV_X1 U10688 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8927) );
  OR2_X1 U10689 ( .A1(n8953), .A2(n8927), .ZN(n8929) );
  INV_X1 U10690 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14903) );
  OR2_X1 U10691 ( .A1(n8976), .A2(n14903), .ZN(n8928) );
  NAND4_X1 U10692 ( .A1(n8931), .A2(n8930), .A3(n8929), .A4(n8928), .ZN(n14913) );
  XNOR2_X1 U10693 ( .A(n15055), .B(n14516), .ZN(n14898) );
  INV_X1 U10694 ( .A(n15055), .ZN(n14517) );
  INV_X1 U10695 ( .A(n8932), .ZN(n8934) );
  NAND2_X1 U10696 ( .A1(n8934), .A2(n8933), .ZN(n8935) );
  NAND2_X1 U10697 ( .A1(n8936), .A2(n8935), .ZN(n12806) );
  OR2_X1 U10698 ( .A1(n12806), .A2(n8937), .ZN(n8939) );
  NAND2_X1 U10699 ( .A1(n8972), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8938) );
  OAI21_X1 U10700 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n8941), .A(n8940), .ZN(
        n14888) );
  OR2_X1 U10701 ( .A1(n8977), .A2(n14888), .ZN(n8946) );
  NAND2_X1 U10702 ( .A1(n8951), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8945) );
  INV_X1 U10703 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8942) );
  OR2_X1 U10704 ( .A1(n8953), .A2(n8942), .ZN(n8944) );
  INV_X1 U10705 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14887) );
  OR2_X1 U10706 ( .A1(n8976), .A2(n14887), .ZN(n8943) );
  NAND4_X1 U10707 ( .A1(n8946), .A2(n8945), .A3(n8944), .A4(n8943), .ZN(n14746) );
  XNOR2_X1 U10708 ( .A(n15047), .B(n14531), .ZN(n14884) );
  XNOR2_X1 U10709 ( .A(n15042), .B(n14745), .ZN(n13069) );
  NAND2_X1 U10710 ( .A1(n8947), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14851) );
  INV_X1 U10711 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U10712 ( .A1(n8949), .A2(n8948), .ZN(n8950) );
  NAND2_X1 U10713 ( .A1(n14851), .A2(n8950), .ZN(n14876) );
  OR2_X1 U10714 ( .A1(n8977), .A2(n14876), .ZN(n8958) );
  NAND2_X1 U10715 ( .A1(n8951), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8957) );
  INV_X1 U10716 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8952) );
  OR2_X1 U10717 ( .A1(n8953), .A2(n8952), .ZN(n8956) );
  INV_X1 U10718 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8954) );
  OR2_X1 U10719 ( .A1(n8976), .A2(n8954), .ZN(n8955) );
  NAND4_X1 U10720 ( .A1(n8958), .A2(n8957), .A3(n8956), .A4(n8955), .ZN(n14744) );
  NOR2_X1 U10721 ( .A1(n8959), .A2(n15283), .ZN(n8961) );
  NAND2_X1 U10722 ( .A1(n8959), .A2(n15283), .ZN(n8960) );
  MUX2_X1 U10723 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10986), .Z(n8968) );
  XNOR2_X1 U10724 ( .A(n8968), .B(n15177), .ZN(n8966) );
  NAND2_X1 U10725 ( .A1(n14374), .A2(n10171), .ZN(n8964) );
  NAND2_X1 U10726 ( .A1(n8972), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8963) );
  NOR2_X1 U10727 ( .A1(n14878), .A2(n14587), .ZN(n9018) );
  INV_X1 U10728 ( .A(n8968), .ZN(n8969) );
  NAND2_X1 U10729 ( .A1(n8969), .A2(n15177), .ZN(n8970) );
  INV_X1 U10730 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15154) );
  INV_X1 U10731 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14371) );
  MUX2_X1 U10732 ( .A(n15154), .B(n14371), .S(n10986), .Z(n10149) );
  XNOR2_X1 U10733 ( .A(n10149), .B(SI_29_), .ZN(n10147) );
  NAND2_X1 U10734 ( .A1(n14369), .A2(n10171), .ZN(n8974) );
  NAND2_X1 U10735 ( .A1(n8972), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U10736 ( .A1(n10157), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8982) );
  INV_X1 U10737 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8975) );
  OR2_X1 U10738 ( .A1(n8976), .A2(n8975), .ZN(n8981) );
  OR2_X1 U10739 ( .A1(n8977), .A2(n14851), .ZN(n8980) );
  INV_X1 U10740 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8978) );
  OR2_X1 U10741 ( .A1(n10161), .A2(n8978), .ZN(n8979) );
  XNOR2_X1 U10742 ( .A(n10181), .B(n14594), .ZN(n10227) );
  NAND2_X1 U10743 ( .A1(n8988), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U10744 ( .A1(n7260), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8987) );
  MUX2_X1 U10745 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8987), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8989) );
  NAND2_X1 U10746 ( .A1(n15162), .A2(n12471), .ZN(n8990) );
  NAND2_X1 U10747 ( .A1(n11438), .A2(n15162), .ZN(n8991) );
  NAND2_X1 U10748 ( .A1(n14589), .A2(n8991), .ZN(n12318) );
  NAND2_X1 U10749 ( .A1(n12389), .A2(n14835), .ZN(n8992) );
  NAND2_X1 U10750 ( .A1(n14862), .A2(n16139), .ZN(n9029) );
  NAND2_X1 U10751 ( .A1(n11441), .A2(n15914), .ZN(n10206) );
  NAND2_X1 U10752 ( .A1(n10037), .A2(n10035), .ZN(n12272) );
  INV_X1 U10753 ( .A(n12272), .ZN(n8994) );
  NAND2_X1 U10754 ( .A1(n8994), .A2(n12270), .ZN(n12274) );
  NAND2_X1 U10755 ( .A1(n7694), .A2(n12281), .ZN(n8995) );
  NAND2_X1 U10756 ( .A1(n11825), .A2(n14767), .ZN(n8996) );
  NAND2_X1 U10757 ( .A1(n12276), .A2(n14566), .ZN(n8997) );
  NAND2_X1 U10758 ( .A1(n16008), .A2(n11840), .ZN(n8998) );
  NAND2_X1 U10759 ( .A1(n8999), .A2(n8998), .ZN(n11629) );
  NAND2_X1 U10760 ( .A1(n9025), .A2(n14765), .ZN(n9000) );
  NAND2_X1 U10761 ( .A1(n7202), .A2(n9000), .ZN(n11804) );
  INV_X1 U10762 ( .A(n14764), .ZN(n12097) );
  OR2_X1 U10763 ( .A1(n12437), .A2(n12097), .ZN(n9001) );
  INV_X1 U10764 ( .A(n14763), .ZN(n12256) );
  NAND2_X1 U10765 ( .A1(n12129), .A2(n12256), .ZN(n9002) );
  INV_X1 U10766 ( .A(n12252), .ZN(n12254) );
  NOR2_X1 U10767 ( .A1(n16076), .A2(n14656), .ZN(n9003) );
  NAND2_X1 U10768 ( .A1(n12199), .A2(n12200), .ZN(n12198) );
  NAND2_X1 U10769 ( .A1(n12198), .A2(n9004), .ZN(n12312) );
  INV_X1 U10770 ( .A(n14760), .ZN(n14696) );
  OR2_X1 U10771 ( .A1(n14560), .A2(n14696), .ZN(n9005) );
  NAND2_X1 U10772 ( .A1(n12392), .A2(n10215), .ZN(n9007) );
  INV_X1 U10773 ( .A(n14759), .ZN(n14615) );
  OR2_X1 U10774 ( .A1(n14703), .A2(n14615), .ZN(n9006) );
  NAND2_X1 U10775 ( .A1(n9007), .A2(n9006), .ZN(n12458) );
  NAND2_X1 U10776 ( .A1(n12458), .A2(n12459), .ZN(n9009) );
  INV_X1 U10777 ( .A(n14758), .ZN(n14385) );
  OR2_X1 U10778 ( .A1(n14387), .A2(n14385), .ZN(n9008) );
  NAND2_X1 U10779 ( .A1(n9009), .A2(n9008), .ZN(n12480) );
  INV_X1 U10780 ( .A(n12483), .ZN(n12481) );
  OR2_X1 U10781 ( .A1(n14679), .A2(n12457), .ZN(n9010) );
  INV_X1 U10782 ( .A(n14756), .ZN(n14422) );
  NAND2_X1 U10783 ( .A1(n16177), .A2(n14422), .ZN(n9011) );
  INV_X1 U10784 ( .A(n10218), .ZN(n12688) );
  INV_X1 U10785 ( .A(n14755), .ZN(n14430) );
  OR2_X1 U10786 ( .A1(n14738), .A2(n14430), .ZN(n9012) );
  NAND2_X1 U10787 ( .A1(n16199), .A2(n14438), .ZN(n9013) );
  INV_X1 U10788 ( .A(n14753), .ZN(n15013) );
  NAND2_X1 U10789 ( .A1(n14449), .A2(n15013), .ZN(n9014) );
  NAND2_X1 U10790 ( .A1(n12933), .A2(n9014), .ZN(n15010) );
  INV_X1 U10791 ( .A(n14750), .ZN(n9015) );
  INV_X1 U10792 ( .A(n14963), .ZN(n14960) );
  OAI21_X1 U10793 ( .B1(n14508), .B2(n15063), .A(n14915), .ZN(n14896) );
  INV_X1 U10794 ( .A(n15047), .ZN(n14886) );
  INV_X1 U10795 ( .A(n14871), .ZN(n14868) );
  NOR2_X1 U10796 ( .A1(n14866), .A2(n9018), .ZN(n9019) );
  XNOR2_X1 U10797 ( .A(n9019), .B(n10227), .ZN(n14865) );
  NAND2_X1 U10798 ( .A1(n10042), .A2(n7860), .ZN(n10166) );
  NAND2_X1 U10799 ( .A1(n7861), .A2(n7860), .ZN(n10232) );
  OR2_X1 U10800 ( .A1(n10232), .A2(n15162), .ZN(n12154) );
  INV_X1 U10801 ( .A(n15161), .ZN(n11449) );
  INV_X1 U10802 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U10803 ( .A1(n10156), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U10804 ( .A1(n10157), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9020) );
  OAI211_X1 U10805 ( .C1(n10161), .C2(n9022), .A(n9021), .B(n9020), .ZN(n14742) );
  INV_X1 U10806 ( .A(P1_B_REG_SCAN_IN), .ZN(n9023) );
  OR2_X1 U10807 ( .A1(n13009), .A2(n9023), .ZN(n14839) );
  AND2_X1 U10808 ( .A1(n14742), .A2(n14839), .ZN(n9024) );
  NAND2_X1 U10809 ( .A1(n14914), .A2(n9024), .ZN(n14852) );
  AND2_X2 U10810 ( .A1(n11033), .A2(n11449), .ZN(n15925) );
  NAND2_X1 U10811 ( .A1(n15925), .A2(n14744), .ZN(n14854) );
  NAND2_X1 U10812 ( .A1(n14852), .A2(n14854), .ZN(n9027) );
  INV_X1 U10813 ( .A(n14738), .ZN(n14431) );
  INV_X1 U10814 ( .A(n12129), .ZN(n12240) );
  NAND2_X1 U10815 ( .A1(n12295), .A2(n9025), .ZN(n11632) );
  INV_X1 U10816 ( .A(n14703), .ZN(n14407) );
  INV_X1 U10817 ( .A(n15099), .ZN(n14984) );
  NAND2_X1 U10818 ( .A1(n15069), .A2(n14922), .ZN(n14919) );
  INV_X1 U10819 ( .A(n14874), .ZN(n9026) );
  AOI211_X1 U10820 ( .C1(n10181), .C2(n16009), .A(n9027), .B(n14861), .ZN(
        n9028) );
  INV_X1 U10821 ( .A(n8863), .ZN(n9030) );
  NAND2_X1 U10822 ( .A1(n9030), .A2(n8412), .ZN(n9033) );
  NOR2_X1 U10823 ( .A1(n12649), .A2(n9023), .ZN(n9037) );
  NAND2_X1 U10824 ( .A1(n9033), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9034) );
  MUX2_X1 U10825 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9034), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9036) );
  MUX2_X1 U10826 ( .A(n9037), .B(n9023), .S(n12608), .Z(n9038) );
  INV_X1 U10827 ( .A(n9038), .ZN(n9040) );
  NAND2_X1 U10828 ( .A1(n7267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U10829 ( .A1(n9040), .A2(n12804), .ZN(n11027) );
  OR2_X1 U10830 ( .A1(n12649), .A2(n12804), .ZN(n15150) );
  OAI21_X1 U10831 ( .B1(n11027), .B2(P1_D_REG_1__SCAN_IN), .A(n15150), .ZN(
        n11549) );
  INV_X1 U10832 ( .A(n11027), .ZN(n9052) );
  NOR4_X1 U10833 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9049) );
  NOR4_X1 U10834 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9048) );
  OR4_X1 U10835 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9046) );
  NOR4_X1 U10836 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9044) );
  NOR4_X1 U10837 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9043) );
  NOR4_X1 U10838 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9042) );
  NOR4_X1 U10839 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9041) );
  NAND4_X1 U10840 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(n9045)
         );
  NOR4_X1 U10841 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n9046), .A4(n9045), .ZN(n9047) );
  NAND3_X1 U10842 ( .A1(n9049), .A2(n9048), .A3(n9047), .ZN(n9050) );
  NAND2_X1 U10843 ( .A1(n9052), .A2(n9050), .ZN(n11548) );
  INV_X1 U10844 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9051) );
  NOR2_X1 U10845 ( .A1(n12608), .A2(n12804), .ZN(n11029) );
  NAND3_X2 U10846 ( .A1(n12649), .A2(n12804), .A3(n12608), .ZN(n11844) );
  NAND2_X1 U10847 ( .A1(n12389), .A2(n12471), .ZN(n9056) );
  NAND2_X1 U10848 ( .A1(n11033), .A2(n9056), .ZN(n11846) );
  AND2_X1 U10849 ( .A1(n11579), .A2(n11561), .ZN(n9057) );
  NAND2_X1 U10850 ( .A1(n15135), .A2(n16141), .ZN(n9059) );
  NAND2_X1 U10851 ( .A1(n16140), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U10852 ( .A1(n9059), .A2(n9058), .ZN(P1_U3557) );
  NOR2_X1 U10853 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n9062) );
  NOR2_X1 U10854 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9061) );
  NAND3_X1 U10855 ( .A1(n9067), .A2(n9066), .A3(n9065), .ZN(n9588) );
  NAND4_X1 U10856 ( .A1(n9596), .A2(n9068), .A3(n9592), .A4(n9645), .ZN(n9069)
         );
  NOR2_X1 U10857 ( .A1(n9588), .A2(n9069), .ZN(n9071) );
  INV_X1 U10858 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9070) );
  INV_X1 U10859 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U10860 ( .A1(n9088), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9075) );
  AND2_X2 U10861 ( .A1(n9078), .A2(n13881), .ZN(n9138) );
  NAND2_X1 U10862 ( .A1(n9138), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9082) );
  INV_X1 U10863 ( .A(n9078), .ZN(n9079) );
  AND2_X2 U10864 ( .A1(n9079), .A2(n13881), .ZN(n9140) );
  NAND2_X1 U10865 ( .A1(n9140), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U10866 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9083) );
  MUX2_X1 U10867 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9083), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n9085) );
  INV_X1 U10868 ( .A(n11410), .ZN(n13883) );
  XNOR2_X1 U10869 ( .A(n9109), .B(n9110), .ZN(n9086) );
  MUX2_X1 U10870 ( .A(n9086), .B(SI_1_), .S(n10986), .Z(n13884) );
  MUX2_X1 U10871 ( .A(n13883), .B(n13884), .S(n9928), .Z(n15908) );
  NAND2_X1 U10872 ( .A1(n9103), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U10873 ( .A1(n9138), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U10874 ( .A1(n9140), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U10875 ( .A1(n9139), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9091) );
  INV_X1 U10876 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11016) );
  INV_X1 U10877 ( .A(n9148), .ZN(n9099) );
  INV_X1 U10878 ( .A(n9109), .ZN(n9097) );
  NAND2_X1 U10879 ( .A1(n9095), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9096) );
  AND2_X1 U10880 ( .A1(n9097), .A2(n9096), .ZN(n11015) );
  INV_X1 U10881 ( .A(n11015), .ZN(n9098) );
  NAND2_X1 U10882 ( .A1(n9099), .A2(n9098), .ZN(n9100) );
  NAND2_X1 U10883 ( .A1(n11228), .A2(n11538), .ZN(n9101) );
  NAND2_X1 U10884 ( .A1(n9102), .A2(n9101), .ZN(n15956) );
  NAND2_X1 U10885 ( .A1(n9103), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U10886 ( .A1(n9138), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U10887 ( .A1(n9140), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U10888 ( .A1(n9139), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9104) );
  INV_X1 U10889 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U10890 ( .A1(n9111), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U10891 ( .A1(n10980), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9124) );
  INV_X1 U10892 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n11021) );
  NAND2_X1 U10893 ( .A1(n11021), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9113) );
  AND2_X1 U10894 ( .A1(n9124), .A2(n9113), .ZN(n9122) );
  XNOR2_X1 U10895 ( .A(n9123), .B(n9122), .ZN(n11007) );
  OR2_X1 U10896 ( .A1(n9148), .A2(n11007), .ZN(n9114) );
  INV_X1 U10897 ( .A(n15970), .ZN(n11351) );
  NAND2_X1 U10898 ( .A1(n11418), .A2(n11351), .ZN(n9760) );
  INV_X1 U10899 ( .A(n11418), .ZN(n13587) );
  NAND2_X1 U10900 ( .A1(n13587), .A2(n15970), .ZN(n9763) );
  NAND2_X1 U10901 ( .A1(n15956), .A2(n9713), .ZN(n9117) );
  NAND2_X1 U10902 ( .A1(n11418), .A2(n15970), .ZN(n9116) );
  INV_X1 U10903 ( .A(n11958), .ZN(n9136) );
  NAND2_X1 U10904 ( .A1(n9103), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U10905 ( .A1(n9138), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U10906 ( .A1(n9140), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9119) );
  INV_X1 U10907 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15343) );
  NAND2_X1 U10908 ( .A1(n9139), .A2(n15343), .ZN(n9118) );
  OR2_X1 U10909 ( .A1(n9262), .A2(SI_3_), .ZN(n9133) );
  NAND2_X1 U10910 ( .A1(n10989), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9151) );
  INV_X1 U10911 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9125) );
  NAND2_X1 U10912 ( .A1(n9125), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9126) );
  XNOR2_X1 U10913 ( .A(n9150), .B(n9149), .ZN(n10996) );
  OR2_X1 U10914 ( .A1(n9148), .A2(n10996), .ZN(n9132) );
  NOR2_X1 U10915 ( .A1(n9108), .A2(n9369), .ZN(n9127) );
  MUX2_X1 U10916 ( .A(n9369), .B(n9127), .S(P3_IR_REG_3__SCAN_IN), .Z(n9130)
         );
  NAND2_X1 U10917 ( .A1(n9108), .A2(n9128), .ZN(n9146) );
  INV_X1 U10918 ( .A(n9146), .ZN(n9129) );
  OR2_X1 U10919 ( .A1(n9928), .A2(n9980), .ZN(n9131) );
  AND3_X2 U10920 ( .A1(n9133), .A2(n9132), .A3(n9131), .ZN(n15986) );
  NAND2_X1 U10921 ( .A1(n15961), .A2(n15986), .ZN(n9768) );
  INV_X1 U10922 ( .A(n15961), .ZN(n13586) );
  INV_X1 U10923 ( .A(n15986), .ZN(n9134) );
  INV_X1 U10924 ( .A(n11957), .ZN(n9135) );
  NAND2_X1 U10925 ( .A1(n13586), .A2(n15986), .ZN(n9137) );
  NAND2_X1 U10926 ( .A1(n9177), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U10927 ( .A1(n9138), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9143) );
  NOR2_X1 U10928 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9157) );
  OR2_X1 U10929 ( .A1(n8414), .A2(n9157), .ZN(n11897) );
  NAND2_X1 U10930 ( .A1(n9139), .A2(n11897), .ZN(n9142) );
  NAND2_X1 U10931 ( .A1(n9477), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9141) );
  NAND4_X1 U10932 ( .A1(n9144), .A2(n9143), .A3(n9142), .A4(n9141), .ZN(n13585) );
  NAND2_X1 U10933 ( .A1(n9146), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9145) );
  MUX2_X1 U10934 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9145), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9147) );
  NAND2_X1 U10935 ( .A1(n9150), .A2(n9149), .ZN(n9152) );
  NAND2_X1 U10936 ( .A1(n10982), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9167) );
  INV_X1 U10937 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U10938 ( .A1(n11023), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9153) );
  XNOR2_X1 U10939 ( .A(n9166), .B(n9165), .ZN(n10998) );
  OR2_X1 U10940 ( .A1(n9148), .A2(n10998), .ZN(n9155) );
  OR2_X1 U10941 ( .A1(n9691), .A2(SI_4_), .ZN(n9154) );
  OAI211_X1 U10942 ( .C1(n15650), .C2(n9928), .A(n9155), .B(n9154), .ZN(n11569) );
  XNOR2_X1 U10943 ( .A(n13585), .B(n11569), .ZN(n11893) );
  INV_X1 U10944 ( .A(n11569), .ZN(n16001) );
  NAND2_X1 U10945 ( .A1(n13585), .A2(n16001), .ZN(n9156) );
  NAND2_X1 U10946 ( .A1(n9177), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U10947 ( .A1(n9138), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U10948 ( .A1(n9157), .A2(n9158), .ZN(n9178) );
  OR2_X1 U10949 ( .A1(n9158), .A2(n9157), .ZN(n9159) );
  NAND2_X1 U10950 ( .A1(n9178), .A2(n9159), .ZN(n11887) );
  NAND2_X1 U10951 ( .A1(n9139), .A2(n11887), .ZN(n9162) );
  NAND2_X1 U10952 ( .A1(n9477), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9161) );
  OR2_X1 U10953 ( .A1(n9691), .A2(SI_5_), .ZN(n9175) );
  NAND2_X1 U10954 ( .A1(n10983), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9187) );
  INV_X1 U10955 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U10956 ( .A1(n10985), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9168) );
  XNOR2_X1 U10957 ( .A(n9186), .B(n9185), .ZN(n11001) );
  OR2_X1 U10958 ( .A1(n9148), .A2(n11001), .ZN(n9174) );
  INV_X1 U10959 ( .A(n9200), .ZN(n9172) );
  NAND2_X1 U10960 ( .A1(n9169), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9170) );
  MUX2_X1 U10961 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9170), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n9171) );
  NAND2_X1 U10962 ( .A1(n9172), .A2(n9171), .ZN(n11002) );
  OR2_X1 U10963 ( .A1(n9928), .A2(n15664), .ZN(n9173) );
  NAND2_X1 U10964 ( .A1(n11994), .A2(n16022), .ZN(n9776) );
  INV_X1 U10965 ( .A(n16022), .ZN(n9191) );
  NAND2_X1 U10966 ( .A1(n13584), .A2(n9191), .ZN(n9775) );
  NAND2_X1 U10967 ( .A1(n9177), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U10968 ( .A1(n9138), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U10969 ( .A1(n9178), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U10970 ( .A1(n9194), .A2(n9179), .ZN(n11987) );
  NAND2_X1 U10971 ( .A1(n9139), .A2(n11987), .ZN(n9181) );
  NAND2_X1 U10972 ( .A1(n9477), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9180) );
  OR2_X1 U10973 ( .A1(n9200), .A2(n9369), .ZN(n9184) );
  XNOR2_X1 U10974 ( .A(n9184), .B(n7864), .ZN(n15683) );
  INV_X1 U10975 ( .A(SI_6_), .ZN(n10987) );
  OR2_X1 U10976 ( .A1(n9691), .A2(n10987), .ZN(n9190) );
  XNOR2_X1 U10977 ( .A(n10993), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n9188) );
  XNOR2_X1 U10978 ( .A(n9204), .B(n9188), .ZN(n10988) );
  OR2_X1 U10979 ( .A1(n9148), .A2(n10988), .ZN(n9189) );
  OAI211_X1 U10980 ( .C1(n9928), .C2(n15683), .A(n9190), .B(n9189), .ZN(n11996) );
  NAND2_X1 U10981 ( .A1(n12025), .A2(n11996), .ZN(n9780) );
  INV_X1 U10982 ( .A(n11996), .ZN(n16032) );
  NAND2_X1 U10983 ( .A1(n13583), .A2(n16032), .ZN(n9781) );
  NAND2_X1 U10984 ( .A1(n9780), .A2(n9781), .ZN(n11929) );
  NAND2_X1 U10985 ( .A1(n11994), .A2(n9191), .ZN(n11930) );
  AND2_X1 U10986 ( .A1(n11929), .A2(n11930), .ZN(n9192) );
  NAND2_X1 U10987 ( .A1(n13583), .A2(n11996), .ZN(n9193) );
  NAND2_X1 U10988 ( .A1(n11928), .A2(n9193), .ZN(n11904) );
  NAND2_X1 U10989 ( .A1(n9177), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U10990 ( .A1(n9601), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9198) );
  AND2_X1 U10991 ( .A1(n9194), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9195) );
  OR2_X1 U10992 ( .A1(n9195), .A2(n9214), .ZN(n12028) );
  NAND2_X1 U10993 ( .A1(n9139), .A2(n12028), .ZN(n9197) );
  NAND2_X1 U10994 ( .A1(n9477), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9196) );
  NAND4_X1 U10995 ( .A1(n9199), .A2(n9198), .A3(n9197), .A4(n9196), .ZN(n13582) );
  NAND2_X1 U10996 ( .A1(n9200), .A2(n7864), .ZN(n9220) );
  NAND2_X1 U10997 ( .A1(n9220), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9202) );
  INV_X1 U10998 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9201) );
  XNOR2_X1 U10999 ( .A(n9202), .B(n9201), .ZN(n11620) );
  INV_X1 U11000 ( .A(n11620), .ZN(n10001) );
  NAND2_X1 U11001 ( .A1(n10994), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U11002 ( .A1(n9204), .A2(n9203), .ZN(n9206) );
  NAND2_X1 U11003 ( .A1(n10993), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11004 ( .A1(n11018), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U11005 ( .A1(n11017), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U11006 ( .A1(n9222), .A2(n9207), .ZN(n9208) );
  NAND2_X1 U11007 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  AND2_X1 U11008 ( .A1(n9223), .A2(n9210), .ZN(n11012) );
  OR2_X1 U11009 ( .A1(n9148), .A2(n11012), .ZN(n9212) );
  OR2_X1 U11010 ( .A1(n9691), .A2(SI_7_), .ZN(n9211) );
  OAI211_X1 U11011 ( .C1(n10001), .C2(n9928), .A(n9212), .B(n9211), .ZN(n12024) );
  XNOR2_X1 U11012 ( .A(n13582), .B(n12024), .ZN(n11903) );
  INV_X1 U11013 ( .A(n12024), .ZN(n16052) );
  NAND2_X1 U11014 ( .A1(n13582), .A2(n16052), .ZN(n9213) );
  NAND2_X1 U11015 ( .A1(n9601), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U11016 ( .A1(n9177), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9218) );
  NOR2_X1 U11017 ( .A1(n9214), .A2(n15346), .ZN(n9215) );
  OR2_X1 U11018 ( .A1(n9232), .A2(n9215), .ZN(n12216) );
  NAND2_X1 U11019 ( .A1(n9139), .A2(n12216), .ZN(n9217) );
  NAND2_X1 U11020 ( .A1(n9477), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9216) );
  NAND4_X1 U11021 ( .A1(n9219), .A2(n9218), .A3(n9217), .A4(n9216), .ZN(n13581) );
  NAND2_X1 U11022 ( .A1(n9244), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11023 ( .A1(n11026), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U11024 ( .A1(n11025), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9224) );
  OR2_X1 U11025 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  NAND2_X1 U11026 ( .A1(n9239), .A2(n9227), .ZN(n11006) );
  OR2_X1 U11027 ( .A1(n9148), .A2(n11006), .ZN(n9229) );
  INV_X1 U11028 ( .A(SI_8_), .ZN(n15320) );
  OR2_X1 U11029 ( .A1(n9691), .A2(n15320), .ZN(n9228) );
  OAI211_X1 U11030 ( .C1(n9928), .C2(n11760), .A(n9229), .B(n9228), .ZN(n12106) );
  XNOR2_X1 U11031 ( .A(n13581), .B(n12106), .ZN(n12212) );
  INV_X1 U11032 ( .A(n13581), .ZN(n12376) );
  INV_X1 U11033 ( .A(n12106), .ZN(n16069) );
  NAND2_X1 U11034 ( .A1(n12376), .A2(n16069), .ZN(n9230) );
  NAND2_X1 U11035 ( .A1(n9177), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U11036 ( .A1(n9601), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9236) );
  OR2_X1 U11037 ( .A1(n9232), .A2(n9231), .ZN(n9233) );
  NAND2_X1 U11038 ( .A1(n9250), .A2(n9233), .ZN(n12236) );
  NAND2_X1 U11039 ( .A1(n9139), .A2(n12236), .ZN(n9235) );
  NAND2_X1 U11040 ( .A1(n9477), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9234) );
  NAND4_X1 U11041 ( .A1(n9237), .A2(n9236), .A3(n9235), .A4(n9234), .ZN(n13580) );
  NAND2_X1 U11042 ( .A1(n11040), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U11043 ( .A1(n11039), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9240) );
  NAND2_X1 U11044 ( .A1(n9242), .A2(n9241), .ZN(n9257) );
  OR2_X1 U11045 ( .A1(n9242), .A2(n9241), .ZN(n9243) );
  AND2_X1 U11046 ( .A1(n9257), .A2(n9243), .ZN(n11004) );
  OR2_X1 U11047 ( .A1(n9148), .A2(n11004), .ZN(n9248) );
  OR2_X1 U11048 ( .A1(n9691), .A2(SI_9_), .ZN(n9247) );
  OR2_X1 U11049 ( .A1(n9264), .A2(n9369), .ZN(n9245) );
  XNOR2_X1 U11050 ( .A(n9245), .B(n9263), .ZN(n12058) );
  INV_X1 U11051 ( .A(n12058), .ZN(n9904) );
  OR2_X1 U11052 ( .A1(n9928), .A2(n9904), .ZN(n9246) );
  NAND2_X1 U11053 ( .A1(n13580), .A2(n12379), .ZN(n9249) );
  NAND2_X1 U11054 ( .A1(n9601), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U11055 ( .A1(n9177), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U11056 ( .A1(n9250), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U11057 ( .A1(n9270), .A2(n9251), .ZN(n12513) );
  NAND2_X1 U11058 ( .A1(n9139), .A2(n12513), .ZN(n9253) );
  NAND2_X1 U11059 ( .A1(n9477), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11060 ( .A1(n11044), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11061 ( .A1(n11042), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9258) );
  OR2_X1 U11062 ( .A1(n9260), .A2(n9259), .ZN(n9261) );
  NAND2_X1 U11063 ( .A1(n9277), .A2(n9261), .ZN(n11011) );
  NAND2_X1 U11064 ( .A1(n9690), .A2(n11011), .ZN(n9268) );
  OR2_X1 U11065 ( .A1(n9691), .A2(SI_10_), .ZN(n9267) );
  NAND2_X1 U11066 ( .A1(n9264), .A2(n9263), .ZN(n9282) );
  NAND2_X1 U11067 ( .A1(n9282), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9265) );
  OR2_X1 U11068 ( .A1(n9928), .A2(n15705), .ZN(n9266) );
  NAND2_X1 U11069 ( .A1(n12497), .A2(n12516), .ZN(n9796) );
  INV_X1 U11070 ( .A(n12497), .ZN(n13579) );
  INV_X1 U11071 ( .A(n12516), .ZN(n16099) );
  NAND2_X1 U11072 ( .A1(n13579), .A2(n16099), .ZN(n9797) );
  NAND2_X1 U11073 ( .A1(n9796), .A2(n9797), .ZN(n12509) );
  NAND2_X1 U11074 ( .A1(n13579), .A2(n12516), .ZN(n9269) );
  NAND2_X1 U11075 ( .A1(n9177), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11076 ( .A1(n9601), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11077 ( .A1(n9270), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9271) );
  NAND2_X1 U11078 ( .A1(n9288), .A2(n9271), .ZN(n12500) );
  NAND2_X1 U11079 ( .A1(n9139), .A2(n12500), .ZN(n9273) );
  NAND2_X1 U11080 ( .A1(n9477), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9272) );
  NAND4_X1 U11081 ( .A1(n9275), .A2(n9274), .A3(n9273), .A4(n9272), .ZN(n13578) );
  NAND2_X1 U11082 ( .A1(n11188), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11083 ( .A1(n11187), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9278) );
  OR2_X1 U11084 ( .A1(n9280), .A2(n9279), .ZN(n9281) );
  NAND2_X1 U11085 ( .A1(n9295), .A2(n9281), .ZN(n10992) );
  NAND2_X1 U11086 ( .A1(n10992), .A2(n9690), .ZN(n9287) );
  OAI21_X1 U11087 ( .B1(n9282), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9284) );
  INV_X1 U11088 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9283) );
  XNOR2_X1 U11089 ( .A(n9284), .B(n9283), .ZN(n15721) );
  OAI22_X1 U11090 ( .A1(n9262), .A2(SI_11_), .B1(n10015), .B2(n9928), .ZN(
        n9285) );
  INV_X1 U11091 ( .A(n9285), .ZN(n9286) );
  NAND2_X1 U11092 ( .A1(n9287), .A2(n9286), .ZN(n12499) );
  INV_X1 U11093 ( .A(n13578), .ZN(n9615) );
  NAND2_X1 U11094 ( .A1(n9103), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11095 ( .A1(n9601), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9292) );
  AND2_X1 U11096 ( .A1(n9288), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9289) );
  OR2_X1 U11097 ( .A1(n9289), .A2(n9319), .ZN(n12658) );
  NAND2_X1 U11098 ( .A1(n9139), .A2(n12658), .ZN(n9291) );
  NAND2_X1 U11099 ( .A1(n9140), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11100 ( .A1(n11362), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9306) );
  NAND2_X1 U11101 ( .A1(n11364), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9296) );
  OR2_X1 U11102 ( .A1(n9298), .A2(n9297), .ZN(n9299) );
  NAND2_X1 U11103 ( .A1(n9307), .A2(n9299), .ZN(n11014) );
  NAND2_X1 U11104 ( .A1(n11014), .A2(n9690), .ZN(n9305) );
  NAND2_X1 U11105 ( .A1(n9300), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9301) );
  MUX2_X1 U11106 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9301), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9303) );
  AOI22_X1 U11107 ( .A1(n9426), .A2(n15307), .B1(n9425), .B2(n15737), .ZN(
        n9304) );
  NAND2_X1 U11108 ( .A1(n9311), .A2(n11393), .ZN(n9312) );
  NAND2_X1 U11109 ( .A1(n9328), .A2(n9312), .ZN(n11031) );
  NAND2_X1 U11110 ( .A1(n11031), .A2(n9690), .ZN(n9317) );
  INV_X1 U11111 ( .A(SI_13_), .ZN(n15304) );
  MUX2_X1 U11112 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9313), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n9315) );
  INV_X1 U11113 ( .A(n9590), .ZN(n9314) );
  NAND2_X1 U11114 ( .A1(n9315), .A2(n9314), .ZN(n11030) );
  AOI22_X1 U11115 ( .A1(n9426), .A2(n15304), .B1(n9425), .B2(n11030), .ZN(
        n9316) );
  NAND2_X1 U11116 ( .A1(n9317), .A2(n9316), .ZN(n16124) );
  NAND2_X1 U11117 ( .A1(n9177), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U11118 ( .A1(n9601), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U11119 ( .A1(n9319), .A2(n9318), .ZN(n9336) );
  OR2_X1 U11120 ( .A1(n9319), .A2(n9318), .ZN(n9320) );
  NAND2_X1 U11121 ( .A1(n9336), .A2(n9320), .ZN(n12786) );
  NAND2_X1 U11122 ( .A1(n9139), .A2(n12786), .ZN(n9322) );
  NAND2_X1 U11123 ( .A1(n9477), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9321) );
  NAND4_X1 U11124 ( .A1(n9324), .A2(n9323), .A3(n9322), .A4(n9321), .ZN(n13576) );
  XNOR2_X1 U11125 ( .A(n16124), .B(n13576), .ZN(n12748) );
  INV_X1 U11126 ( .A(n13576), .ZN(n12808) );
  OR2_X1 U11127 ( .A1(n16124), .A2(n12808), .ZN(n9325) );
  NAND2_X1 U11128 ( .A1(n11519), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U11129 ( .A1(n11521), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9329) );
  OR2_X1 U11130 ( .A1(n9331), .A2(n9330), .ZN(n9332) );
  NAND2_X1 U11131 ( .A1(n9343), .A2(n9332), .ZN(n11038) );
  NAND2_X1 U11132 ( .A1(n11038), .A2(n9690), .ZN(n9335) );
  OR2_X1 U11133 ( .A1(n9590), .A2(n9369), .ZN(n9333) );
  XNOR2_X1 U11134 ( .A(n9333), .B(n9348), .ZN(n11036) );
  AOI22_X1 U11135 ( .A1(n9426), .A2(n11037), .B1(n9425), .B2(n11036), .ZN(
        n9334) );
  NAND2_X1 U11136 ( .A1(n9335), .A2(n9334), .ZN(n16158) );
  NAND2_X1 U11137 ( .A1(n9601), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U11138 ( .A1(n9140), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U11139 ( .A1(n9336), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U11140 ( .A1(n9353), .A2(n9337), .ZN(n12819) );
  NAND2_X1 U11141 ( .A1(n9139), .A2(n12819), .ZN(n9339) );
  NAND2_X1 U11142 ( .A1(n9103), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9338) );
  NAND4_X1 U11143 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), .ZN(n13575) );
  OR2_X1 U11144 ( .A1(n16158), .A2(n13575), .ZN(n12973) );
  NAND2_X1 U11145 ( .A1(n16158), .A2(n13575), .ZN(n9753) );
  NAND2_X1 U11146 ( .A1(n12973), .A2(n9753), .ZN(n9707) );
  INV_X1 U11147 ( .A(n13575), .ZN(n12784) );
  NAND2_X1 U11148 ( .A1(n11752), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9361) );
  INV_X1 U11149 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11751) );
  NAND2_X1 U11150 ( .A1(n11751), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9344) );
  OR2_X1 U11151 ( .A1(n9346), .A2(n9345), .ZN(n9347) );
  NAND2_X1 U11152 ( .A1(n9362), .A2(n9347), .ZN(n11045) );
  OR2_X1 U11153 ( .A1(n11045), .A2(n9148), .ZN(n9351) );
  OR2_X1 U11154 ( .A1(n9368), .A2(n9369), .ZN(n9349) );
  XNOR2_X1 U11155 ( .A(n9349), .B(P3_IR_REG_15__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U11156 ( .A1(n9426), .A2(SI_15_), .B1(n9425), .B2(n10024), .ZN(
        n9350) );
  NAND2_X1 U11157 ( .A1(n9351), .A2(n9350), .ZN(n13815) );
  NAND2_X1 U11158 ( .A1(n9601), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U11159 ( .A1(n9103), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9358) );
  INV_X1 U11160 ( .A(n9373), .ZN(n9355) );
  NAND2_X1 U11161 ( .A1(n9353), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9354) );
  NAND2_X1 U11162 ( .A1(n9355), .A2(n9354), .ZN(n12977) );
  NAND2_X1 U11163 ( .A1(n9139), .A2(n12977), .ZN(n9357) );
  INV_X1 U11164 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15784) );
  OR2_X1 U11165 ( .A1(n9160), .A2(n15784), .ZN(n9356) );
  OR2_X1 U11166 ( .A1(n13815), .A2(n12983), .ZN(n9818) );
  NAND2_X1 U11167 ( .A1(n13815), .A2(n12983), .ZN(n9817) );
  INV_X1 U11168 ( .A(n12983), .ZN(n13574) );
  OR2_X1 U11169 ( .A1(n13815), .A2(n13574), .ZN(n13012) );
  NAND2_X1 U11170 ( .A1(n11861), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9381) );
  INV_X1 U11171 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U11172 ( .A1(n11860), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9363) );
  OR2_X1 U11173 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  NAND2_X1 U11174 ( .A1(n9382), .A2(n9366), .ZN(n11259) );
  OR2_X1 U11175 ( .A1(n11259), .A2(n9148), .ZN(n9372) );
  OR2_X1 U11176 ( .A1(n9388), .A2(n9369), .ZN(n9370) );
  XNOR2_X1 U11177 ( .A(n9370), .B(P3_IR_REG_16__SCAN_IN), .ZN(n15798) );
  AOI22_X1 U11178 ( .A1(n9426), .A2(SI_16_), .B1(n9425), .B2(n15798), .ZN(
        n9371) );
  NAND2_X1 U11179 ( .A1(n9372), .A2(n9371), .ZN(n13811) );
  NAND2_X1 U11180 ( .A1(n9601), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U11181 ( .A1(n9103), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9377) );
  NOR2_X1 U11182 ( .A1(n9373), .A2(n15357), .ZN(n9374) );
  OR2_X1 U11183 ( .A1(n9393), .A2(n9374), .ZN(n13019) );
  NAND2_X1 U11184 ( .A1(n9139), .A2(n13019), .ZN(n9376) );
  NAND2_X1 U11185 ( .A1(n9140), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9375) );
  OR2_X1 U11186 ( .A1(n13811), .A2(n13746), .ZN(n9822) );
  NAND2_X1 U11187 ( .A1(n13811), .A2(n13746), .ZN(n9821) );
  NAND2_X1 U11188 ( .A1(n9822), .A2(n9821), .ZN(n9719) );
  OR2_X1 U11189 ( .A1(n13811), .A2(n13573), .ZN(n9380) );
  NAND2_X1 U11190 ( .A1(n11971), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9399) );
  INV_X1 U11191 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11973) );
  NAND2_X1 U11192 ( .A1(n11973), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9383) );
  OR2_X1 U11193 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  NAND2_X1 U11194 ( .A1(n9400), .A2(n9386), .ZN(n11359) );
  OR2_X1 U11195 ( .A1(n11359), .A2(n9148), .ZN(n9391) );
  NAND2_X1 U11196 ( .A1(n9405), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9389) );
  XNOR2_X1 U11197 ( .A(n9389), .B(P3_IR_REG_17__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U11198 ( .A1(n9426), .A2(SI_17_), .B1(n9425), .B2(n9956), .ZN(n9390) );
  NAND2_X1 U11199 ( .A1(n9103), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9398) );
  NAND2_X1 U11200 ( .A1(n9601), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9397) );
  OR2_X1 U11201 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U11202 ( .A1(n9409), .A2(n9394), .ZN(n13752) );
  NAND2_X1 U11203 ( .A1(n9139), .A2(n13752), .ZN(n9396) );
  NAND2_X1 U11204 ( .A1(n9477), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9395) );
  OR2_X1 U11205 ( .A1(n13807), .A2(n13734), .ZN(n9826) );
  NAND2_X1 U11206 ( .A1(n13807), .A2(n13734), .ZN(n9833) );
  INV_X1 U11207 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n12385) );
  NAND2_X1 U11208 ( .A1(n12385), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9416) );
  INV_X1 U11209 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n12387) );
  NAND2_X1 U11210 ( .A1(n12387), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9401) );
  OR2_X1 U11211 ( .A1(n9403), .A2(n9402), .ZN(n9404) );
  NAND2_X1 U11212 ( .A1(n9417), .A2(n9404), .ZN(n11425) );
  OR2_X1 U11213 ( .A1(n11425), .A2(n9148), .ZN(n9408) );
  NAND2_X1 U11214 ( .A1(n9422), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9406) );
  XNOR2_X1 U11215 ( .A(n9406), .B(P3_IR_REG_18__SCAN_IN), .ZN(n15833) );
  AOI22_X1 U11216 ( .A1(n9426), .A2(SI_18_), .B1(n9425), .B2(n15833), .ZN(
        n9407) );
  NAND2_X1 U11217 ( .A1(n9408), .A2(n9407), .ZN(n13544) );
  NAND2_X1 U11218 ( .A1(n9103), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11219 ( .A1(n9601), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11220 ( .A1(n9409), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9410) );
  NAND2_X1 U11221 ( .A1(n9429), .A2(n9410), .ZN(n13739) );
  NAND2_X1 U11222 ( .A1(n9139), .A2(n13739), .ZN(n9412) );
  NAND2_X1 U11223 ( .A1(n9140), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9411) );
  OR2_X1 U11224 ( .A1(n13544), .A2(n13745), .ZN(n9834) );
  NAND2_X1 U11225 ( .A1(n13544), .A2(n13745), .ZN(n9830) );
  NAND2_X1 U11226 ( .A1(n9834), .A2(n9830), .ZN(n13730) );
  NAND2_X1 U11227 ( .A1(n13807), .A2(n13572), .ZN(n13731) );
  AND2_X1 U11228 ( .A1(n13730), .A2(n13731), .ZN(n9415) );
  INV_X1 U11229 ( .A(n13745), .ZN(n13571) );
  INV_X1 U11230 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12470) );
  NAND2_X1 U11231 ( .A1(n12470), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9439) );
  INV_X1 U11232 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13026) );
  NAND2_X1 U11233 ( .A1(n13026), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9418) );
  OR2_X1 U11234 ( .A1(n9420), .A2(n9419), .ZN(n9421) );
  NAND2_X1 U11235 ( .A1(n9440), .A2(n9421), .ZN(n11506) );
  NAND2_X1 U11236 ( .A1(n11506), .A2(n9690), .ZN(n9428) );
  AOI22_X1 U11237 ( .A1(n9426), .A2(n15192), .B1(n9425), .B2(n11505), .ZN(
        n9427) );
  AND2_X1 U11238 ( .A1(n9429), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9430) );
  OR2_X1 U11239 ( .A1(n9430), .A2(n9447), .ZN(n13724) );
  NAND2_X1 U11240 ( .A1(n13724), .A2(n9139), .ZN(n9435) );
  NAND2_X1 U11241 ( .A1(n9177), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11242 ( .A1(n9601), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9431) );
  AND2_X1 U11243 ( .A1(n9432), .A2(n9431), .ZN(n9434) );
  NAND2_X1 U11244 ( .A1(n9477), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9433) );
  OR2_X1 U11245 ( .A1(n13860), .A2(n13735), .ZN(n9436) );
  NAND2_X1 U11246 ( .A1(n13719), .A2(n9436), .ZN(n9438) );
  NAND2_X1 U11247 ( .A1(n13860), .A2(n13735), .ZN(n9437) );
  NAND2_X1 U11248 ( .A1(n9443), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U11249 ( .A1(n9454), .A2(n9444), .ZN(n11733) );
  OR2_X1 U11250 ( .A1(n9691), .A2(n11731), .ZN(n9445) );
  INV_X1 U11251 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n9451) );
  NOR2_X1 U11252 ( .A1(n9447), .A2(n15369), .ZN(n9448) );
  OR2_X1 U11253 ( .A1(n9461), .A2(n9448), .ZN(n13712) );
  NAND2_X1 U11254 ( .A1(n13712), .A2(n9139), .ZN(n9450) );
  AOI22_X1 U11255 ( .A1(n9601), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n9103), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n9449) );
  XNOR2_X1 U11256 ( .A(n13532), .B(n13687), .ZN(n13704) );
  NAND2_X1 U11257 ( .A1(n13532), .A2(n13687), .ZN(n9452) );
  INV_X1 U11258 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U11259 ( .A1(n12479), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9466) );
  INV_X1 U11260 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12520) );
  NAND2_X1 U11261 ( .A1(n12520), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9455) );
  AND2_X1 U11262 ( .A1(n9466), .A2(n9455), .ZN(n9456) );
  OR2_X1 U11263 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  NAND2_X1 U11264 ( .A1(n9467), .A2(n9458), .ZN(n11966) );
  OR2_X1 U11265 ( .A1(n11966), .A2(n9148), .ZN(n9460) );
  INV_X1 U11266 ( .A(SI_21_), .ZN(n15189) );
  OR2_X1 U11267 ( .A1(n9262), .A2(n15189), .ZN(n9459) );
  INV_X1 U11268 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n9465) );
  NOR2_X1 U11269 ( .A1(n9461), .A2(n15348), .ZN(n9462) );
  OR2_X1 U11270 ( .A1(n9475), .A2(n9462), .ZN(n13695) );
  NAND2_X1 U11271 ( .A1(n13695), .A2(n9139), .ZN(n9464) );
  AOI22_X1 U11272 ( .A1(n9601), .A2(P3_REG0_REG_21__SCAN_IN), .B1(n9177), .B2(
        P3_REG1_REG_21__SCAN_IN), .ZN(n9463) );
  OAI211_X1 U11273 ( .C1(n9160), .C2(n9465), .A(n9464), .B(n9463), .ZN(n13709)
         );
  AND2_X1 U11274 ( .A1(n13697), .A2(n13709), .ZN(n13096) );
  INV_X1 U11275 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U11276 ( .A1(n9468), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9487) );
  INV_X1 U11277 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12625) );
  NAND2_X1 U11278 ( .A1(n12625), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9469) );
  AND2_X1 U11279 ( .A1(n9487), .A2(n9469), .ZN(n9470) );
  OR2_X1 U11280 ( .A1(n9471), .A2(n9470), .ZN(n9472) );
  NAND2_X1 U11281 ( .A1(n9488), .A2(n9472), .ZN(n12002) );
  OR2_X1 U11282 ( .A1(n9691), .A2(n15295), .ZN(n9473) );
  INV_X1 U11283 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15374) );
  OR2_X1 U11284 ( .A1(n9475), .A2(n15374), .ZN(n9476) );
  NAND2_X1 U11285 ( .A1(n9476), .A2(n9492), .ZN(n13679) );
  NAND2_X1 U11286 ( .A1(n13679), .A2(n9139), .ZN(n9483) );
  INV_X1 U11287 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13846) );
  NAND2_X1 U11288 ( .A1(n9177), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U11289 ( .A1(n9477), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9478) );
  OAI211_X1 U11290 ( .C1(n9480), .C2(n13846), .A(n9479), .B(n9478), .ZN(n9481)
         );
  INV_X1 U11291 ( .A(n9481), .ZN(n9482) );
  NAND2_X1 U11292 ( .A1(n13539), .A2(n13688), .ZN(n9484) );
  NAND2_X1 U11293 ( .A1(n13673), .A2(n9484), .ZN(n9486) );
  OR2_X1 U11294 ( .A1(n13539), .A2(n13688), .ZN(n9485) );
  XNOR2_X1 U11295 ( .A(n9501), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n9499) );
  XNOR2_X1 U11296 ( .A(n9500), .B(n9499), .ZN(n12135) );
  NAND2_X1 U11297 ( .A1(n12135), .A2(n9690), .ZN(n9490) );
  OR2_X1 U11298 ( .A1(n9691), .A2(n15172), .ZN(n9489) );
  NAND2_X1 U11299 ( .A1(n9103), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11300 ( .A1(n9601), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9496) );
  INV_X1 U11301 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n13478) );
  INV_X1 U11302 ( .A(n9492), .ZN(n9491) );
  NAND2_X1 U11303 ( .A1(n13478), .A2(n9491), .ZN(n9507) );
  NAND2_X1 U11304 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(n9492), .ZN(n9493) );
  NAND2_X1 U11305 ( .A1(n9507), .A2(n9493), .ZN(n13668) );
  NAND2_X1 U11306 ( .A1(n9139), .A2(n13668), .ZN(n9495) );
  NAND2_X1 U11307 ( .A1(n9140), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9494) );
  NAND2_X1 U11308 ( .A1(n13474), .A2(n13676), .ZN(n9749) );
  INV_X1 U11309 ( .A(n13676), .ZN(n13570) );
  NAND2_X1 U11310 ( .A1(n13474), .A2(n13570), .ZN(n9498) );
  NAND2_X1 U11311 ( .A1(n9502), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9503) );
  XNOR2_X1 U11312 ( .A(n9514), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12560) );
  NAND2_X1 U11313 ( .A1(n12560), .A2(n9690), .ZN(n9505) );
  INV_X1 U11314 ( .A(SI_24_), .ZN(n15293) );
  OR2_X1 U11315 ( .A1(n9691), .A2(n15293), .ZN(n9504) );
  NAND2_X1 U11316 ( .A1(n9103), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U11317 ( .A1(n9601), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9511) );
  INV_X1 U11318 ( .A(n9507), .ZN(n9506) );
  INV_X1 U11319 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15246) );
  NAND2_X1 U11320 ( .A1(n9506), .A2(n15246), .ZN(n9523) );
  NAND2_X1 U11321 ( .A1(n9507), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9508) );
  NAND2_X1 U11322 ( .A1(n9523), .A2(n9508), .ZN(n13657) );
  NAND2_X1 U11323 ( .A1(n9139), .A2(n13657), .ZN(n9510) );
  NAND2_X1 U11324 ( .A1(n9140), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9509) );
  NAND2_X1 U11325 ( .A1(n13522), .A2(n13504), .ZN(n9739) );
  OR2_X1 U11326 ( .A1(n13522), .A2(n13665), .ZN(n9513) );
  INV_X1 U11327 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12626) );
  INV_X1 U11328 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9516) );
  NAND2_X1 U11329 ( .A1(n9516), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9529) );
  INV_X1 U11330 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U11331 ( .A1(n12685), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9517) );
  AND2_X1 U11332 ( .A1(n9529), .A2(n9517), .ZN(n9518) );
  NAND2_X1 U11333 ( .A1(n9530), .A2(n9520), .ZN(n12564) );
  OR2_X1 U11334 ( .A1(n9691), .A2(n15290), .ZN(n9521) );
  NAND2_X1 U11335 ( .A1(n9103), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U11336 ( .A1(n9601), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U11337 ( .A1(n9523), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9524) );
  NAND2_X1 U11338 ( .A1(n9539), .A2(n9524), .ZN(n13644) );
  NAND2_X1 U11339 ( .A1(n9139), .A2(n13644), .ZN(n9526) );
  NAND2_X1 U11340 ( .A1(n9140), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9525) );
  XNOR2_X1 U11341 ( .A(n13505), .B(n13656), .ZN(n13639) );
  INV_X1 U11342 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9531) );
  NAND2_X1 U11343 ( .A1(n9531), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9547) );
  INV_X1 U11344 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U11345 ( .A1(n9532), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9533) );
  AND2_X1 U11346 ( .A1(n9547), .A2(n9533), .ZN(n9534) );
  INV_X1 U11347 ( .A(SI_26_), .ZN(n15284) );
  OR2_X1 U11348 ( .A1(n9691), .A2(n15284), .ZN(n9535) );
  NAND2_X1 U11349 ( .A1(n9601), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9544) );
  NAND2_X1 U11350 ( .A1(n9140), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9543) );
  INV_X1 U11351 ( .A(n9539), .ZN(n9538) );
  INV_X1 U11352 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U11353 ( .A1(n9538), .A2(n9537), .ZN(n9552) );
  NAND2_X1 U11354 ( .A1(n9539), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U11355 ( .A1(n9552), .A2(n9540), .ZN(n13630) );
  NAND2_X1 U11356 ( .A1(n9139), .A2(n13630), .ZN(n9542) );
  NAND2_X1 U11357 ( .A1(n9177), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9541) );
  NAND4_X1 U11358 ( .A1(n9544), .A2(n9543), .A3(n9542), .A4(n9541), .ZN(n13637) );
  OR2_X1 U11359 ( .A1(n13560), .A2(n13637), .ZN(n9546) );
  AND2_X1 U11360 ( .A1(n13560), .A2(n13637), .ZN(n9545) );
  NAND2_X1 U11361 ( .A1(n13008), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U11362 ( .A1(n13011), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U11363 ( .A1(n9562), .A2(n9549), .ZN(n9559) );
  XNOR2_X1 U11364 ( .A(n9561), .B(n9559), .ZN(n13129) );
  NAND2_X1 U11365 ( .A1(n13129), .A2(n9690), .ZN(n9551) );
  OR2_X1 U11366 ( .A1(n9691), .A2(n15283), .ZN(n9550) );
  NAND2_X1 U11367 ( .A1(n9601), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U11368 ( .A1(n9103), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U11369 ( .A1(n9552), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9553) );
  NAND2_X1 U11370 ( .A1(n9572), .A2(n9553), .ZN(n13619) );
  NAND2_X1 U11371 ( .A1(n9139), .A2(n13619), .ZN(n9555) );
  NAND2_X1 U11372 ( .A1(n9140), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9554) );
  AND4_X2 U11373 ( .A1(n9557), .A2(n9556), .A3(n9555), .A4(n9554), .ZN(n13627)
         );
  XNOR2_X1 U11374 ( .A(n13117), .B(n13627), .ZN(n9877) );
  NAND2_X1 U11375 ( .A1(n9876), .A2(n9877), .ZN(n9875) );
  OR2_X1 U11376 ( .A1(n13117), .A2(n13568), .ZN(n9558) );
  INV_X1 U11377 ( .A(n9559), .ZN(n9560) );
  NAND2_X1 U11378 ( .A1(n9561), .A2(n9560), .ZN(n9563) );
  INV_X1 U11379 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15158) );
  NAND2_X1 U11380 ( .A1(n15158), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9579) );
  INV_X1 U11381 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U11382 ( .A1(n9564), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U11383 ( .A1(n9580), .A2(n9568), .ZN(n12801) );
  OR2_X1 U11384 ( .A1(n9691), .A2(n15177), .ZN(n9569) );
  NAND2_X1 U11385 ( .A1(n9601), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U11386 ( .A1(n9140), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9576) );
  INV_X1 U11387 ( .A(n9572), .ZN(n9571) );
  INV_X1 U11388 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U11389 ( .A1(n9571), .A2(n9570), .ZN(n13594) );
  NAND2_X1 U11390 ( .A1(n9572), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U11391 ( .A1(n13594), .A2(n9573), .ZN(n13613) );
  NAND2_X1 U11392 ( .A1(n9139), .A2(n13613), .ZN(n9575) );
  NAND2_X1 U11393 ( .A1(n9103), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9574) );
  XNOR2_X1 U11394 ( .A(n14371), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U11395 ( .A1(n13879), .A2(n9690), .ZN(n9582) );
  INV_X1 U11396 ( .A(SI_29_), .ZN(n15277) );
  OR2_X1 U11397 ( .A1(n9691), .A2(n15277), .ZN(n9581) );
  NAND2_X1 U11398 ( .A1(n9582), .A2(n9581), .ZN(n9669) );
  INV_X1 U11399 ( .A(n13594), .ZN(n9583) );
  NAND2_X1 U11400 ( .A1(n9139), .A2(n9583), .ZN(n9686) );
  NAND2_X1 U11401 ( .A1(n9601), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9586) );
  NAND2_X1 U11402 ( .A1(n9103), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U11403 ( .A1(n9140), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U11404 ( .A1(n9669), .A2(n13610), .ZN(n9695) );
  NAND2_X1 U11405 ( .A1(n9861), .A2(n9695), .ZN(n9706) );
  INV_X1 U11406 ( .A(n9595), .ZN(n9591) );
  NAND2_X1 U11407 ( .A1(n9644), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U11408 ( .A1(n9725), .A2(n12000), .ZN(n9887) );
  NAND2_X1 U11409 ( .A1(n9595), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9597) );
  INV_X1 U11410 ( .A(n11732), .ZN(n9702) );
  NAND2_X1 U11411 ( .A1(n11878), .A2(n9702), .ZN(n9728) );
  INV_X1 U11412 ( .A(n7187), .ZN(n9960) );
  NAND2_X1 U11413 ( .A1(n9960), .A2(n9966), .ZN(n9929) );
  NAND2_X1 U11414 ( .A1(n9929), .A2(n9928), .ZN(n11236) );
  INV_X1 U11415 ( .A(P3_B_REG_SCAN_IN), .ZN(n9599) );
  NOR2_X1 U11416 ( .A1(n7187), .A2(n9599), .ZN(n9600) );
  OR2_X1 U11417 ( .A1(n15962), .A2(n9600), .ZN(n13592) );
  NAND2_X1 U11418 ( .A1(n9177), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U11419 ( .A1(n9601), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U11420 ( .A1(n9140), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9602) );
  OAI22_X1 U11421 ( .A1(n13470), .A2(n15960), .B1(n13592), .B2(n12033), .ZN(
        n9605) );
  NAND2_X1 U11422 ( .A1(n13590), .A2(n11592), .ZN(n9709) );
  NAND2_X1 U11423 ( .A1(n9607), .A2(n9709), .ZN(n9756) );
  INV_X1 U11424 ( .A(n9713), .ZN(n15957) );
  NAND2_X1 U11425 ( .A1(n9609), .A2(n9768), .ZN(n11891) );
  INV_X1 U11426 ( .A(n11893), .ZN(n9767) );
  NAND2_X1 U11427 ( .A1(n11891), .A2(n9767), .ZN(n9610) );
  INV_X1 U11428 ( .A(n13585), .ZN(n11886) );
  NAND2_X1 U11429 ( .A1(n11886), .A2(n16001), .ZN(n9769) );
  INV_X1 U11430 ( .A(n11929), .ZN(n9778) );
  NAND2_X1 U11431 ( .A1(n9611), .A2(n9780), .ZN(n11901) );
  INV_X1 U11432 ( .A(n11903), .ZN(n9783) );
  NAND2_X1 U11433 ( .A1(n11901), .A2(n9783), .ZN(n9612) );
  NAND2_X1 U11434 ( .A1(n12214), .A2(n16052), .ZN(n9785) );
  NAND2_X1 U11435 ( .A1(n9612), .A2(n9785), .ZN(n12208) );
  NAND2_X1 U11436 ( .A1(n12208), .A2(n12212), .ZN(n9614) );
  NAND2_X1 U11437 ( .A1(n12376), .A2(n12106), .ZN(n9613) );
  NOR2_X1 U11438 ( .A1(n13580), .A2(n16084), .ZN(n9793) );
  NAND2_X1 U11439 ( .A1(n13580), .A2(n16084), .ZN(n9711) );
  INV_X1 U11440 ( .A(n12499), .ZN(n16108) );
  NAND2_X1 U11441 ( .A1(n9615), .A2(n16108), .ZN(n9802) );
  NAND2_X1 U11442 ( .A1(n13578), .A2(n12499), .ZN(n9803) );
  NAND2_X1 U11443 ( .A1(n12448), .A2(n9802), .ZN(n12654) );
  NAND2_X1 U11444 ( .A1(n12853), .A2(n13577), .ZN(n9806) );
  NAND2_X1 U11445 ( .A1(n12654), .A2(n12653), .ZN(n12652) );
  NAND2_X1 U11446 ( .A1(n12652), .A2(n9807), .ZN(n12747) );
  INV_X1 U11447 ( .A(n12748), .ZN(n12746) );
  OR2_X1 U11448 ( .A1(n16124), .A2(n13576), .ZN(n9752) );
  INV_X1 U11449 ( .A(n9707), .ZN(n12793) );
  NAND2_X1 U11450 ( .A1(n13749), .A2(n9833), .ZN(n13738) );
  INV_X1 U11451 ( .A(n13730), .ZN(n13737) );
  INV_X1 U11452 ( .A(n13860), .ZN(n9617) );
  NAND2_X1 U11453 ( .A1(n13860), .A2(n13707), .ZN(n9829) );
  INV_X1 U11454 ( .A(n13687), .ZN(n13721) );
  OR2_X1 U11455 ( .A1(n13532), .A2(n13721), .ZN(n9618) );
  NAND2_X1 U11456 ( .A1(n9619), .A2(n9618), .ZN(n13684) );
  INV_X1 U11457 ( .A(n13709), .ZN(n13675) );
  NAND2_X1 U11458 ( .A1(n13697), .A2(n13675), .ZN(n13099) );
  NAND2_X1 U11459 ( .A1(n13539), .A2(n13496), .ZN(n9751) );
  NAND2_X1 U11460 ( .A1(n13650), .A2(n13654), .ZN(n9620) );
  NAND2_X1 U11461 ( .A1(n9620), .A2(n9742), .ZN(n13636) );
  NAND2_X1 U11462 ( .A1(n13636), .A2(n13635), .ZN(n9622) );
  OR2_X1 U11463 ( .A1(n13505), .A2(n13656), .ZN(n9621) );
  NAND2_X1 U11464 ( .A1(n13560), .A2(n13115), .ZN(n9731) );
  AND2_X2 U11465 ( .A1(n9732), .A2(n9731), .ZN(n13628) );
  XNOR2_X1 U11466 ( .A(n9699), .B(n9706), .ZN(n13599) );
  NAND2_X1 U11467 ( .A1(n11505), .A2(n11732), .ZN(n9628) );
  NAND2_X1 U11468 ( .A1(n9628), .A2(n9887), .ZN(n9663) );
  OR2_X1 U11469 ( .A1(n9663), .A2(n9755), .ZN(n11658) );
  NAND2_X1 U11470 ( .A1(n11505), .A2(n11967), .ZN(n9625) );
  NAND2_X1 U11471 ( .A1(n11967), .A2(n11732), .ZN(n9664) );
  XNOR2_X1 U11472 ( .A(n12000), .B(n9664), .ZN(n9624) );
  NAND2_X1 U11473 ( .A1(n9625), .A2(n9624), .ZN(n11247) );
  INV_X1 U11474 ( .A(n9628), .ZN(n11245) );
  NAND3_X1 U11475 ( .A1(n11247), .A2(n11245), .A3(n16157), .ZN(n9626) );
  AND2_X1 U11476 ( .A1(n9725), .A2(n11732), .ZN(n11879) );
  OR2_X1 U11477 ( .A1(n11658), .A2(n9926), .ZN(n9629) );
  NAND2_X1 U11478 ( .A1(n9630), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U11479 ( .A1(n8172), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9632) );
  MUX2_X1 U11480 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9632), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9633) );
  XNOR2_X1 U11481 ( .A(n12562), .B(P3_B_REG_SCAN_IN), .ZN(n9636) );
  NAND2_X1 U11482 ( .A1(n7220), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9634) );
  MUX2_X1 U11483 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9634), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9635) );
  NAND2_X1 U11484 ( .A1(n9635), .A2(n9630), .ZN(n12563) );
  NAND2_X1 U11485 ( .A1(n9636), .A2(n12563), .ZN(n9637) );
  INV_X1 U11486 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U11487 ( .A1(n9649), .A2(n9638), .ZN(n9640) );
  INV_X1 U11488 ( .A(n9648), .ZN(n12647) );
  NAND2_X1 U11489 ( .A1(n12647), .A2(n12563), .ZN(n9639) );
  NAND2_X1 U11490 ( .A1(n11659), .A2(n13869), .ZN(n9668) );
  INV_X1 U11491 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9641) );
  NAND2_X1 U11492 ( .A1(n12647), .A2(n12562), .ZN(n9642) );
  NAND2_X1 U11493 ( .A1(n13871), .A2(n13869), .ZN(n9884) );
  NOR2_X1 U11494 ( .A1(n12563), .A2(n12562), .ZN(n9647) );
  NAND2_X1 U11495 ( .A1(n9648), .A2(n9647), .ZN(n11244) );
  NOR2_X1 U11496 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9653) );
  NOR4_X1 U11497 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9652) );
  NOR4_X1 U11498 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9651) );
  NOR4_X1 U11499 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9650) );
  NAND4_X1 U11500 ( .A1(n9653), .A2(n9652), .A3(n9651), .A4(n9650), .ZN(n9659)
         );
  NOR4_X1 U11501 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9657) );
  NOR4_X1 U11502 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9656) );
  NOR4_X1 U11503 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9655) );
  NOR4_X1 U11504 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9654) );
  NAND4_X1 U11505 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(n9658)
         );
  NOR2_X1 U11506 ( .A1(n9659), .A2(n9658), .ZN(n9660) );
  NOR2_X1 U11507 ( .A1(n11240), .A2(n9888), .ZN(n9662) );
  INV_X1 U11508 ( .A(n13871), .ZN(n9661) );
  NAND2_X1 U11509 ( .A1(n9661), .A2(n11662), .ZN(n9889) );
  NAND2_X1 U11510 ( .A1(n9663), .A2(n11967), .ZN(n9666) );
  NAND2_X1 U11511 ( .A1(n9755), .A2(n9664), .ZN(n9665) );
  NAND3_X1 U11512 ( .A1(n9666), .A2(n11662), .A3(n9665), .ZN(n9667) );
  INV_X1 U11513 ( .A(n9669), .ZN(n13601) );
  INV_X1 U11514 ( .A(n16157), .ZN(n16107) );
  INV_X1 U11515 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9671) );
  NOR2_X1 U11516 ( .A1(n16165), .A2(n9671), .ZN(n9672) );
  NOR2_X1 U11517 ( .A1(n9670), .A2(n9672), .ZN(n9673) );
  OAI21_X1 U11518 ( .B1(n10405), .B2(n9674), .A(n9673), .ZN(P3_U3488) );
  INV_X2 U11519 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U11520 ( .A(n9861), .ZN(n9698) );
  INV_X1 U11521 ( .A(n9675), .ZN(n9676) );
  NAND2_X1 U11522 ( .A1(n15154), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9678) );
  XNOR2_X1 U11523 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n9687) );
  INV_X1 U11524 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13128) );
  INV_X1 U11525 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9679) );
  XNOR2_X1 U11526 ( .A(n9679), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n9680) );
  XNOR2_X1 U11527 ( .A(n9681), .B(n9680), .ZN(n13877) );
  INV_X1 U11528 ( .A(SI_31_), .ZN(n13873) );
  OR2_X1 U11529 ( .A1(n9262), .A2(n13873), .ZN(n9682) );
  NAND2_X1 U11530 ( .A1(n9601), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U11531 ( .A1(n9140), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U11532 ( .A1(n9103), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n9683) );
  INV_X1 U11533 ( .A(n9687), .ZN(n9688) );
  XNOR2_X1 U11534 ( .A(n9689), .B(n9688), .ZN(n13460) );
  NAND2_X1 U11535 ( .A1(n13460), .A2(n9690), .ZN(n9693) );
  INV_X1 U11536 ( .A(SI_30_), .ZN(n15281) );
  OR2_X1 U11537 ( .A1(n9691), .A2(n15281), .ZN(n9692) );
  NAND2_X1 U11538 ( .A1(n13596), .A2(n12033), .ZN(n9694) );
  INV_X1 U11539 ( .A(n9695), .ZN(n9696) );
  NAND2_X1 U11540 ( .A1(n13596), .A2(n13593), .ZN(n9697) );
  NOR2_X1 U11541 ( .A1(n13596), .A2(n12033), .ZN(n9703) );
  OAI21_X1 U11542 ( .B1(n9703), .B2(n13593), .A(n13591), .ZN(n9700) );
  XNOR2_X1 U11543 ( .A(n9701), .B(n11505), .ZN(n9729) );
  NAND2_X1 U11544 ( .A1(n13591), .A2(n13593), .ZN(n9705) );
  INV_X1 U11545 ( .A(n9703), .ZN(n9704) );
  NAND2_X1 U11546 ( .A1(n9705), .A2(n9704), .ZN(n9863) );
  NOR2_X1 U11547 ( .A1(n9840), .A2(n7905), .ZN(n13722) );
  INV_X1 U11548 ( .A(n13750), .ZN(n9718) );
  NOR2_X1 U11549 ( .A1(n9707), .A2(n12748), .ZN(n9811) );
  INV_X1 U11550 ( .A(n9709), .ZN(n9710) );
  NOR2_X1 U11551 ( .A1(n9710), .A2(n11496), .ZN(n11502) );
  NAND4_X1 U11552 ( .A1(n11957), .A2(n11884), .A3(n9778), .A4(n11502), .ZN(
        n9712) );
  INV_X1 U11553 ( .A(n9711), .ZN(n9794) );
  OR2_X1 U11554 ( .A1(n9794), .A2(n9793), .ZN(n12232) );
  NOR4_X1 U11555 ( .A1(n9708), .A2(n9713), .A3(n9712), .A4(n12232), .ZN(n9715)
         );
  NOR3_X1 U11556 ( .A1(n11893), .A2(n12509), .A3(n11903), .ZN(n9714) );
  AND4_X1 U11557 ( .A1(n9715), .A2(n12449), .A3(n9714), .A4(n12212), .ZN(n9716) );
  NAND4_X1 U11558 ( .A1(n12969), .A2(n9811), .A3(n12653), .A4(n9716), .ZN(
        n9717) );
  NOR4_X1 U11559 ( .A1(n13730), .A2(n9719), .A3(n9718), .A4(n9717), .ZN(n9720)
         );
  AND4_X1 U11560 ( .A1(n13689), .A2(n13722), .A3(n9720), .A4(n13704), .ZN(
        n9721) );
  NAND4_X1 U11561 ( .A1(n9587), .A2(n13663), .A3(n13678), .A4(n9721), .ZN(
        n9723) );
  NAND2_X1 U11562 ( .A1(n13628), .A2(n13635), .ZN(n9722) );
  NAND3_X1 U11563 ( .A1(n9743), .A2(n13654), .A3(n13608), .ZN(n9747) );
  XNOR2_X1 U11564 ( .A(n9726), .B(n9725), .ZN(n9727) );
  NAND2_X1 U11565 ( .A1(n13505), .A2(n13656), .ZN(n9730) );
  NAND2_X1 U11566 ( .A1(n9731), .A2(n9730), .ZN(n9733) );
  NAND2_X1 U11567 ( .A1(n9733), .A2(n9732), .ZN(n9734) );
  NAND2_X1 U11568 ( .A1(n13117), .A2(n13627), .ZN(n9736) );
  NAND2_X1 U11569 ( .A1(n9737), .A2(n9736), .ZN(n9741) );
  INV_X1 U11570 ( .A(n9741), .ZN(n9738) );
  OAI21_X1 U11571 ( .B1(n9740), .B2(n9739), .A(n9738), .ZN(n9745) );
  NAND2_X1 U11572 ( .A1(n9746), .A2(n13608), .ZN(n9857) );
  INV_X1 U11573 ( .A(n9747), .ZN(n9855) );
  MUX2_X1 U11574 ( .A(n9749), .B(n9748), .S(n9926), .Z(n9854) );
  MUX2_X1 U11575 ( .A(n9751), .B(n9750), .S(n11657), .Z(n9852) );
  NAND2_X1 U11576 ( .A1(n9753), .A2(n7887), .ZN(n9754) );
  NAND2_X1 U11577 ( .A1(n9754), .A2(n12973), .ZN(n9814) );
  NOR2_X1 U11578 ( .A1(n9814), .A2(n9926), .ZN(n9813) );
  NAND2_X1 U11579 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  NAND3_X1 U11580 ( .A1(n15957), .A2(n11878), .A3(n9757), .ZN(n9759) );
  AOI22_X1 U11581 ( .A1(n15954), .A2(n9759), .B1(n9926), .B2(n9758), .ZN(n9762) );
  AOI21_X1 U11582 ( .B1(n9768), .B2(n9760), .A(n9926), .ZN(n9761) );
  OR2_X1 U11583 ( .A1(n9762), .A2(n9761), .ZN(n9766) );
  AOI21_X1 U11584 ( .B1(n9765), .B2(n9763), .A(n11657), .ZN(n9764) );
  AOI21_X1 U11585 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9773) );
  OAI21_X1 U11586 ( .B1(n11657), .B2(n9768), .A(n9767), .ZN(n9772) );
  NAND2_X1 U11587 ( .A1(n13585), .A2(n11569), .ZN(n9770) );
  MUX2_X1 U11588 ( .A(n9770), .B(n9769), .S(n11657), .Z(n9771) );
  OAI21_X1 U11589 ( .B1(n9773), .B2(n9772), .A(n9771), .ZN(n9774) );
  NAND2_X1 U11590 ( .A1(n9774), .A2(n11884), .ZN(n9779) );
  MUX2_X1 U11591 ( .A(n9776), .B(n9775), .S(n9926), .Z(n9777) );
  NAND3_X1 U11592 ( .A1(n9779), .A2(n9778), .A3(n9777), .ZN(n9784) );
  MUX2_X1 U11593 ( .A(n9781), .B(n9780), .S(n9926), .Z(n9782) );
  NAND3_X1 U11594 ( .A1(n9784), .A2(n9783), .A3(n9782), .ZN(n9788) );
  NAND2_X1 U11595 ( .A1(n13582), .A2(n12024), .ZN(n9786) );
  MUX2_X1 U11596 ( .A(n9786), .B(n9785), .S(n11657), .Z(n9787) );
  NAND3_X1 U11597 ( .A1(n9788), .A2(n12212), .A3(n9787), .ZN(n9792) );
  INV_X1 U11598 ( .A(n12232), .ZN(n9791) );
  MUX2_X1 U11599 ( .A(n13581), .B(n9926), .S(n12106), .Z(n9789) );
  OAI21_X1 U11600 ( .B1(n12376), .B2(n11657), .A(n9789), .ZN(n9790) );
  NAND3_X1 U11601 ( .A1(n9792), .A2(n9791), .A3(n9790), .ZN(n9801) );
  MUX2_X1 U11602 ( .A(n9794), .B(n9793), .S(n11657), .Z(n9795) );
  NOR2_X1 U11603 ( .A1(n9795), .A2(n12509), .ZN(n9800) );
  MUX2_X1 U11604 ( .A(n9797), .B(n9796), .S(n9926), .Z(n9798) );
  NAND2_X1 U11605 ( .A1(n9798), .A2(n12449), .ZN(n9799) );
  AOI21_X1 U11606 ( .B1(n9801), .B2(n9800), .A(n9799), .ZN(n9810) );
  NAND2_X1 U11607 ( .A1(n9807), .A2(n9802), .ZN(n9805) );
  NAND2_X1 U11608 ( .A1(n9806), .A2(n9803), .ZN(n9804) );
  MUX2_X1 U11609 ( .A(n9805), .B(n9804), .S(n9926), .Z(n9809) );
  MUX2_X1 U11610 ( .A(n9807), .B(n9806), .S(n11657), .Z(n9808) );
  OAI21_X1 U11611 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(n9812) );
  MUX2_X1 U11612 ( .A(n9813), .B(n9812), .S(n9811), .Z(n9816) );
  AND2_X1 U11613 ( .A1(n9814), .A2(n9926), .ZN(n9815) );
  OAI21_X1 U11614 ( .B1(n9816), .B2(n9815), .A(n12969), .ZN(n9820) );
  MUX2_X1 U11615 ( .A(n9818), .B(n9817), .S(n9926), .Z(n9819) );
  NAND3_X1 U11616 ( .A1(n9820), .A2(n13017), .A3(n9819), .ZN(n9824) );
  MUX2_X1 U11617 ( .A(n9822), .B(n9821), .S(n11657), .Z(n9823) );
  NAND2_X1 U11618 ( .A1(n9824), .A2(n9823), .ZN(n9825) );
  NAND4_X1 U11619 ( .A1(n9825), .A2(n13750), .A3(n9830), .A4(n9834), .ZN(n9839) );
  INV_X1 U11620 ( .A(n9834), .ZN(n9832) );
  INV_X1 U11621 ( .A(n9826), .ZN(n9827) );
  AOI21_X1 U11622 ( .B1(n9830), .B2(n9827), .A(n11657), .ZN(n9828) );
  NAND2_X1 U11623 ( .A1(n9829), .A2(n9828), .ZN(n9836) );
  OR3_X1 U11624 ( .A1(n9840), .A2(n9926), .A3(n7908), .ZN(n9831) );
  OAI21_X1 U11625 ( .B1(n9832), .B2(n9836), .A(n9831), .ZN(n9838) );
  INV_X1 U11626 ( .A(n9833), .ZN(n9835) );
  NAND3_X1 U11627 ( .A1(n9836), .A2(n9835), .A3(n9834), .ZN(n9837) );
  NAND3_X1 U11628 ( .A1(n9839), .A2(n9838), .A3(n9837), .ZN(n9843) );
  MUX2_X1 U11629 ( .A(n7905), .B(n9840), .S(n9926), .Z(n9841) );
  INV_X1 U11630 ( .A(n9841), .ZN(n9842) );
  NAND3_X1 U11631 ( .A1(n9843), .A2(n13704), .A3(n9842), .ZN(n9847) );
  NAND2_X1 U11632 ( .A1(n13687), .A2(n9926), .ZN(n9845) );
  NAND2_X1 U11633 ( .A1(n13721), .A2(n11657), .ZN(n9844) );
  MUX2_X1 U11634 ( .A(n9845), .B(n9844), .S(n13532), .Z(n9846) );
  NAND2_X1 U11635 ( .A1(n9847), .A2(n9846), .ZN(n9848) );
  NAND2_X1 U11636 ( .A1(n9848), .A2(n13689), .ZN(n9850) );
  MUX2_X1 U11637 ( .A(n13099), .B(n13097), .S(n9926), .Z(n9849) );
  NAND3_X1 U11638 ( .A1(n9850), .A2(n13678), .A3(n9849), .ZN(n9851) );
  NAND3_X1 U11639 ( .A1(n13663), .A2(n9852), .A3(n9851), .ZN(n9853) );
  NAND3_X1 U11640 ( .A1(n9855), .A2(n9854), .A3(n9853), .ZN(n9856) );
  INV_X1 U11641 ( .A(n9858), .ZN(n9859) );
  AND2_X1 U11642 ( .A1(n9862), .A2(n9863), .ZN(n9864) );
  INV_X1 U11643 ( .A(n11879), .ZN(n11664) );
  OR2_X1 U11644 ( .A1(n9925), .A2(P3_U3151), .ZN(n12136) );
  NOR2_X1 U11645 ( .A1(n11500), .A2(n11240), .ZN(n11253) );
  NAND3_X1 U11646 ( .A1(n11253), .A2(n9960), .A3(n13132), .ZN(n9871) );
  OAI211_X1 U11647 ( .C1(n12000), .C2(n12136), .A(n9871), .B(P3_B_REG_SCAN_IN), 
        .ZN(n9872) );
  NAND2_X1 U11648 ( .A1(n9873), .A2(n9872), .ZN(P3_U3296) );
  INV_X1 U11649 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n9893) );
  XNOR2_X1 U11650 ( .A(n9874), .B(n9877), .ZN(n13618) );
  OAI21_X1 U11651 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  INV_X1 U11652 ( .A(n9878), .ZN(n9883) );
  AOI21_X1 U11653 ( .B1(n13618), .B2(n16160), .A(n13622), .ZN(n13765) );
  INV_X1 U11654 ( .A(n9884), .ZN(n9886) );
  INV_X1 U11655 ( .A(n9888), .ZN(n9885) );
  NAND2_X1 U11656 ( .A1(n9886), .A2(n9885), .ZN(n11248) );
  OR2_X1 U11657 ( .A1(n9887), .A2(n11223), .ZN(n11250) );
  AND2_X1 U11658 ( .A1(n11500), .A2(n11250), .ZN(n9891) );
  NAND2_X1 U11659 ( .A1(n11251), .A2(n11247), .ZN(n9890) );
  OAI21_X1 U11660 ( .B1(n11248), .B2(n9891), .A(n9890), .ZN(n9892) );
  INV_X1 U11661 ( .A(n11240), .ZN(n11234) );
  MUX2_X1 U11662 ( .A(n9893), .B(n13765), .S(n16169), .Z(n9894) );
  NAND2_X1 U11663 ( .A1(n9894), .A2(n8407), .ZN(P3_U3454) );
  INV_X1 U11664 ( .A(n11244), .ZN(n9895) );
  INV_X1 U11665 ( .A(n15833), .ZN(n11423) );
  INV_X1 U11666 ( .A(n15798), .ZN(n11258) );
  INV_X1 U11667 ( .A(n11030), .ZN(n15745) );
  INV_X1 U11668 ( .A(n15705), .ZN(n11010) );
  INV_X1 U11669 ( .A(n15650), .ZN(n10999) );
  INV_X1 U11670 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9974) );
  XNOR2_X1 U11671 ( .A(n11391), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n11373) );
  INV_X1 U11672 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11672) );
  NOR2_X1 U11673 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11672), .ZN(n15609) );
  INV_X1 U11674 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U11675 ( .A1(n9930), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U11676 ( .A1(n11400), .A2(n9896), .ZN(n11372) );
  INV_X1 U11677 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n15622) );
  INV_X1 U11678 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9986) );
  XNOR2_X1 U11679 ( .A(n15650), .B(n9986), .ZN(n15639) );
  NOR2_X1 U11680 ( .A1(n9899), .A2(n15664), .ZN(n9900) );
  INV_X1 U11681 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15660) );
  NAND2_X1 U11682 ( .A1(n15683), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9999) );
  OR2_X1 U11683 ( .A1(n15683), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9901) );
  NAND2_X1 U11684 ( .A1(n9999), .A2(n9901), .ZN(n15676) );
  INV_X1 U11685 ( .A(n9999), .ZN(n9902) );
  NOR2_X1 U11686 ( .A1(n10001), .A2(n7241), .ZN(n9903) );
  INV_X1 U11687 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11908) );
  INV_X1 U11688 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U11689 ( .A1(n10005), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n12215), 
        .B2(n11760), .ZN(n11762) );
  INV_X1 U11690 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12053) );
  INV_X1 U11691 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n9907) );
  MUX2_X1 U11692 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n9907), .S(n15705), .Z(
        n15695) );
  NOR2_X1 U11693 ( .A1(n10015), .A2(n9908), .ZN(n9909) );
  INV_X1 U11694 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n15712) );
  INV_X1 U11695 ( .A(n15737), .ZN(n10018) );
  NAND2_X1 U11696 ( .A1(n10018), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9912) );
  INV_X1 U11697 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U11698 ( .A1(n15737), .A2(n9910), .ZN(n9911) );
  AND2_X1 U11699 ( .A1(n9912), .A2(n9911), .ZN(n15727) );
  NOR2_X1 U11700 ( .A1(n15745), .A2(n9913), .ZN(n9914) );
  INV_X1 U11701 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15755) );
  INV_X1 U11702 ( .A(n11036), .ZN(n15768) );
  NAND2_X1 U11703 ( .A1(n15768), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9916) );
  INV_X1 U11704 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12797) );
  NAND2_X1 U11705 ( .A1(n11036), .A2(n12797), .ZN(n9915) );
  AND2_X1 U11706 ( .A1(n9916), .A2(n9915), .ZN(n15763) );
  NAND2_X1 U11707 ( .A1(n11036), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U11708 ( .A1(n10024), .A2(n9918), .ZN(n9919) );
  INV_X1 U11709 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U11710 ( .A1(n15798), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n9920), 
        .B2(n11258), .ZN(n15808) );
  INV_X1 U11711 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n15816) );
  NOR2_X1 U11712 ( .A1(n15815), .A2(n15816), .ZN(n15814) );
  NOR2_X1 U11713 ( .A1(n9956), .A2(n9921), .ZN(n9922) );
  OR2_X1 U11714 ( .A1(n15833), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U11715 ( .A1(n15833), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9923) );
  AND2_X1 U11716 ( .A1(n9924), .A2(n9923), .ZN(n15846) );
  XNOR2_X1 U11717 ( .A(n11505), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n9967) );
  AND2_X1 U11718 ( .A1(n11240), .A2(n12136), .ZN(n9962) );
  NAND2_X1 U11719 ( .A1(n9926), .A2(n9925), .ZN(n9927) );
  NAND2_X1 U11720 ( .A1(n9928), .A2(n9927), .ZN(n9963) );
  INV_X1 U11721 ( .A(n9956), .ZN(n15821) );
  INV_X1 U11722 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U11723 ( .A1(n15798), .A2(n9955), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n11258), .ZN(n15804) );
  INV_X1 U11724 ( .A(n10024), .ZN(n15789) );
  INV_X1 U11725 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n16164) );
  INV_X1 U11726 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12851) );
  INV_X1 U11727 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n16104) );
  INV_X1 U11728 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n16073) );
  AOI22_X1 U11729 ( .A1(n10005), .A2(n16073), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n11760), .ZN(n11758) );
  NAND2_X1 U11730 ( .A1(n15683), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9998) );
  INV_X1 U11731 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9995) );
  MUX2_X1 U11732 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n9995), .S(n15683), .Z(
        n15688) );
  INV_X1 U11733 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9985) );
  INV_X1 U11734 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9973) );
  MUX2_X1 U11735 ( .A(n9973), .B(P3_REG1_REG_2__SCAN_IN), .S(n11391), .Z(
        n11375) );
  NAND2_X1 U11736 ( .A1(n9930), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U11737 ( .A1(n11410), .A2(n9934), .ZN(n9933) );
  NAND2_X1 U11738 ( .A1(n11016), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9931) );
  OR2_X1 U11739 ( .A1(n9931), .A2(n9930), .ZN(n9932) );
  NAND2_X1 U11740 ( .A1(n9933), .A2(n9932), .ZN(n11402) );
  NAND2_X1 U11741 ( .A1(n11402), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9935) );
  NAND2_X1 U11742 ( .A1(n9935), .A2(n9934), .ZN(n11376) );
  NAND2_X1 U11743 ( .A1(n11375), .A2(n11376), .ZN(n11380) );
  OR2_X1 U11744 ( .A1(n11391), .A2(n9973), .ZN(n9936) );
  NAND2_X1 U11745 ( .A1(n11380), .A2(n9936), .ZN(n9937) );
  XNOR2_X1 U11746 ( .A(n9937), .B(n9980), .ZN(n15633) );
  AND2_X1 U11747 ( .A1(n9937), .A2(n15630), .ZN(n9938) );
  AOI21_X1 U11748 ( .B1(n15633), .B2(P3_REG1_REG_3__SCAN_IN), .A(n9938), .ZN(
        n15652) );
  MUX2_X1 U11749 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n9985), .S(n15650), .Z(
        n15651) );
  NAND2_X1 U11750 ( .A1(n11002), .A2(n9939), .ZN(n9940) );
  NAND2_X1 U11751 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n15670), .ZN(n15669) );
  NAND2_X1 U11752 ( .A1(n9940), .A2(n15669), .ZN(n15689) );
  NAND2_X1 U11753 ( .A1(n15688), .A2(n15689), .ZN(n15687) );
  NAND2_X1 U11754 ( .A1(n9998), .A2(n15687), .ZN(n9941) );
  NAND2_X1 U11755 ( .A1(n11620), .A2(n9941), .ZN(n9942) );
  XNOR2_X1 U11756 ( .A(n9941), .B(n10001), .ZN(n11616) );
  NAND2_X1 U11757 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n11616), .ZN(n11615) );
  NAND2_X1 U11758 ( .A1(n12058), .A2(n9943), .ZN(n9944) );
  NAND2_X1 U11759 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n12056), .ZN(n12055) );
  MUX2_X1 U11760 ( .A(n16104), .B(P3_REG1_REG_10__SCAN_IN), .S(n15705), .Z(
        n15697) );
  NAND2_X1 U11761 ( .A1(n15721), .A2(n9945), .ZN(n9946) );
  NAND2_X1 U11762 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15716), .ZN(n15715) );
  NAND2_X1 U11763 ( .A1(n9946), .A2(n15715), .ZN(n15732) );
  NAND2_X1 U11764 ( .A1(n15737), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9947) );
  OAI21_X1 U11765 ( .B1(n15737), .B2(P3_REG1_REG_12__SCAN_IN), .A(n9947), .ZN(
        n9948) );
  INV_X1 U11766 ( .A(n9948), .ZN(n15733) );
  NAND2_X1 U11767 ( .A1(n15732), .A2(n15733), .ZN(n15731) );
  NAND2_X1 U11768 ( .A1(n11030), .A2(n9949), .ZN(n9950) );
  NAND2_X1 U11769 ( .A1(n11036), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9951) );
  OAI21_X1 U11770 ( .B1(n11036), .B2(P3_REG1_REG_14__SCAN_IN), .A(n9951), .ZN(
        n9952) );
  INV_X1 U11771 ( .A(n9952), .ZN(n15767) );
  NAND2_X1 U11772 ( .A1(n15766), .A2(n15767), .ZN(n15765) );
  NAND2_X1 U11773 ( .A1(n15789), .A2(n9953), .ZN(n9954) );
  NAND2_X1 U11774 ( .A1(n15804), .A2(n15803), .ZN(n15802) );
  NAND2_X1 U11775 ( .A1(n15821), .A2(n9957), .ZN(n9958) );
  XNOR2_X1 U11776 ( .A(n15833), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n15835) );
  AOI22_X1 U11777 ( .A1(n15836), .A2(n15835), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n11423), .ZN(n9959) );
  XNOR2_X1 U11778 ( .A(n11505), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n9968) );
  XNOR2_X1 U11779 ( .A(n9959), .B(n9968), .ZN(n10034) );
  INV_X1 U11780 ( .A(P3_U3897), .ZN(n13589) );
  MUX2_X1 U11781 ( .A(n9961), .B(n13589), .S(n9960), .Z(n15822) );
  NAND2_X1 U11782 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13485)
         );
  INV_X1 U11783 ( .A(n9962), .ZN(n9964) );
  NAND2_X1 U11784 ( .A1(n15832), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n9965) );
  OAI211_X1 U11785 ( .C1(n15822), .C2(n11505), .A(n13485), .B(n9965), .ZN(
        n10033) );
  MUX2_X1 U11786 ( .A(n9968), .B(n9967), .S(n9966), .Z(n10032) );
  MUX2_X1 U11787 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13132), .Z(n10029) );
  MUX2_X1 U11788 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13132), .Z(n10028) );
  MUX2_X1 U11789 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13132), .Z(n10020) );
  INV_X1 U11790 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U11791 ( .A1(n9971), .A2(n13883), .ZN(n11386) );
  INV_X1 U11792 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9972) );
  MUX2_X1 U11793 ( .A(n11672), .B(n9972), .S(n13132), .Z(n15610) );
  AND2_X1 U11794 ( .A1(n15610), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15613) );
  NAND2_X1 U11795 ( .A1(n11396), .A2(n15613), .ZN(n11395) );
  NAND2_X1 U11796 ( .A1(n11395), .A2(n11386), .ZN(n9978) );
  MUX2_X1 U11797 ( .A(n9974), .B(n9973), .S(n13132), .Z(n9975) );
  NAND2_X1 U11798 ( .A1(n9975), .A2(n11391), .ZN(n15625) );
  INV_X1 U11799 ( .A(n9975), .ZN(n9976) );
  INV_X1 U11800 ( .A(n11391), .ZN(n11008) );
  NAND2_X1 U11801 ( .A1(n9976), .A2(n11008), .ZN(n9977) );
  AND2_X1 U11802 ( .A1(n15625), .A2(n9977), .ZN(n11385) );
  NAND2_X1 U11803 ( .A1(n9978), .A2(n11385), .ZN(n15626) );
  NAND2_X1 U11804 ( .A1(n15626), .A2(n15625), .ZN(n9984) );
  INV_X1 U11805 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n9979) );
  MUX2_X1 U11806 ( .A(n15622), .B(n9979), .S(n13132), .Z(n9981) );
  NAND2_X1 U11807 ( .A1(n9981), .A2(n9980), .ZN(n15644) );
  INV_X1 U11808 ( .A(n9981), .ZN(n9982) );
  NAND2_X1 U11809 ( .A1(n9982), .A2(n15630), .ZN(n9983) );
  AND2_X1 U11810 ( .A1(n15644), .A2(n9983), .ZN(n15623) );
  NAND2_X1 U11811 ( .A1(n9984), .A2(n15623), .ZN(n15645) );
  NAND2_X1 U11812 ( .A1(n15645), .A2(n15644), .ZN(n9990) );
  MUX2_X1 U11813 ( .A(n9986), .B(n9985), .S(n13132), .Z(n9987) );
  NAND2_X1 U11814 ( .A1(n9987), .A2(n15650), .ZN(n9991) );
  INV_X1 U11815 ( .A(n9987), .ZN(n9988) );
  NAND2_X1 U11816 ( .A1(n9988), .A2(n10999), .ZN(n9989) );
  AND2_X1 U11817 ( .A1(n9991), .A2(n9989), .ZN(n15642) );
  NAND2_X1 U11818 ( .A1(n9990), .A2(n15642), .ZN(n15647) );
  NAND2_X1 U11819 ( .A1(n15647), .A2(n9991), .ZN(n15663) );
  MUX2_X1 U11820 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13132), .Z(n9992) );
  XNOR2_X1 U11821 ( .A(n9992), .B(n15664), .ZN(n15662) );
  INV_X1 U11822 ( .A(n9992), .ZN(n9993) );
  NAND2_X1 U11823 ( .A1(n9993), .A2(n15664), .ZN(n9994) );
  INV_X1 U11824 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11935) );
  MUX2_X1 U11825 ( .A(n11935), .B(n9995), .S(n13132), .Z(n9997) );
  INV_X1 U11826 ( .A(n15683), .ZN(n9996) );
  AND2_X1 U11827 ( .A1(n9997), .A2(n9996), .ZN(n15678) );
  MUX2_X1 U11828 ( .A(n9999), .B(n9998), .S(n13132), .Z(n15679) );
  MUX2_X1 U11829 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13132), .Z(n10000) );
  XNOR2_X1 U11830 ( .A(n10000), .B(n11620), .ZN(n11613) );
  OR2_X1 U11831 ( .A1(n11612), .A2(n11613), .ZN(n11610) );
  INV_X1 U11832 ( .A(n10000), .ZN(n10002) );
  NAND2_X1 U11833 ( .A1(n10002), .A2(n10001), .ZN(n10003) );
  NAND2_X1 U11834 ( .A1(n11610), .A2(n10003), .ZN(n11754) );
  MUX2_X1 U11835 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13132), .Z(n10004) );
  XNOR2_X1 U11836 ( .A(n10004), .B(n10005), .ZN(n11755) );
  NAND2_X1 U11837 ( .A1(n11754), .A2(n11755), .ZN(n10008) );
  INV_X1 U11838 ( .A(n10004), .ZN(n10006) );
  NAND2_X1 U11839 ( .A1(n10006), .A2(n10005), .ZN(n10007) );
  NAND2_X1 U11840 ( .A1(n10008), .A2(n10007), .ZN(n12061) );
  MUX2_X1 U11841 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13132), .Z(n10009) );
  XNOR2_X1 U11842 ( .A(n10009), .B(n12058), .ZN(n12062) );
  NAND2_X1 U11843 ( .A1(n10009), .A2(n12058), .ZN(n10010) );
  MUX2_X1 U11844 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13132), .Z(n10011) );
  XNOR2_X1 U11845 ( .A(n10011), .B(n15705), .ZN(n15703) );
  INV_X1 U11846 ( .A(n10011), .ZN(n10012) );
  NAND2_X1 U11847 ( .A1(n10012), .A2(n15705), .ZN(n10013) );
  MUX2_X1 U11848 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13132), .Z(n10014) );
  XNOR2_X1 U11849 ( .A(n10014), .B(n10015), .ZN(n15713) );
  INV_X1 U11850 ( .A(n10014), .ZN(n10016) );
  AND2_X1 U11851 ( .A1(n10016), .A2(n10015), .ZN(n10017) );
  AOI21_X1 U11852 ( .B1(n15714), .B2(n15713), .A(n10017), .ZN(n15730) );
  MUX2_X1 U11853 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13132), .Z(n10019) );
  XNOR2_X1 U11854 ( .A(n10019), .B(n10018), .ZN(n15729) );
  XNOR2_X1 U11855 ( .A(n10020), .B(n15745), .ZN(n15749) );
  MUX2_X1 U11856 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13132), .Z(n10021) );
  NAND2_X1 U11857 ( .A1(n10021), .A2(n11036), .ZN(n10022) );
  OAI21_X1 U11858 ( .B1(n10021), .B2(n11036), .A(n10022), .ZN(n15775) );
  INV_X1 U11859 ( .A(n10022), .ZN(n10023) );
  NOR2_X1 U11860 ( .A1(n15774), .A2(n10023), .ZN(n10025) );
  INV_X1 U11861 ( .A(n10025), .ZN(n10027) );
  INV_X1 U11862 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n10026) );
  MUX2_X1 U11863 ( .A(n15784), .B(n10026), .S(n13132), .Z(n15791) );
  XNOR2_X1 U11864 ( .A(n10028), .B(n15798), .ZN(n15800) );
  OAI21_X1 U11865 ( .B1(n10028), .B2(n11258), .A(n15799), .ZN(n15824) );
  XNOR2_X1 U11866 ( .A(n10029), .B(n15821), .ZN(n15825) );
  MUX2_X1 U11867 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13132), .Z(n15839) );
  AOI21_X1 U11868 ( .B1(n10030), .B2(n15833), .A(n15837), .ZN(n10031) );
  NAND2_X1 U11869 ( .A1(P3_U3897), .A2(n7187), .ZN(n15840) );
  INV_X1 U11870 ( .A(n10206), .ZN(n15922) );
  AOI22_X1 U11871 ( .A1(n15922), .A2(n10035), .B1(n10038), .B2(n7694), .ZN(
        n10044) );
  INV_X1 U11872 ( .A(n11441), .ZN(n15924) );
  NAND2_X1 U11873 ( .A1(n15924), .A2(n15888), .ZN(n10205) );
  NAND2_X1 U11874 ( .A1(n10205), .A2(n11438), .ZN(n10039) );
  AOI22_X1 U11875 ( .A1(n15921), .A2(n10039), .B1(n15978), .B2(n10038), .ZN(
        n10043) );
  MUX2_X1 U11876 ( .A(n15917), .B(n14769), .S(n10188), .Z(n10046) );
  NAND2_X1 U11877 ( .A1(n14769), .A2(n15917), .ZN(n10045) );
  NAND2_X1 U11878 ( .A1(n10046), .A2(n10045), .ZN(n10047) );
  NAND2_X1 U11879 ( .A1(n10109), .A2(n14768), .ZN(n10049) );
  NAND2_X1 U11880 ( .A1(n10188), .A2(n7694), .ZN(n10048) );
  MUX2_X1 U11881 ( .A(n14767), .B(n14566), .S(n10188), .Z(n10054) );
  INV_X4 U11882 ( .A(n10109), .ZN(n10191) );
  MUX2_X1 U11883 ( .A(n14566), .B(n14767), .S(n10191), .Z(n10051) );
  NAND2_X1 U11884 ( .A1(n10052), .A2(n10051), .ZN(n10058) );
  INV_X1 U11885 ( .A(n10053), .ZN(n10056) );
  INV_X1 U11886 ( .A(n10054), .ZN(n10055) );
  NAND2_X1 U11887 ( .A1(n10056), .A2(n10055), .ZN(n10057) );
  MUX2_X1 U11888 ( .A(n16008), .B(n14766), .S(n10191), .Z(n10060) );
  MUX2_X1 U11889 ( .A(n14766), .B(n16008), .S(n10191), .Z(n10059) );
  INV_X1 U11890 ( .A(n10060), .ZN(n10061) );
  MUX2_X1 U11891 ( .A(n14765), .B(n12159), .S(n10191), .Z(n10065) );
  NAND2_X1 U11892 ( .A1(n10064), .A2(n10065), .ZN(n10063) );
  MUX2_X1 U11893 ( .A(n12159), .B(n14765), .S(n10191), .Z(n10062) );
  INV_X1 U11894 ( .A(n10064), .ZN(n10067) );
  INV_X1 U11895 ( .A(n10065), .ZN(n10066) );
  MUX2_X1 U11896 ( .A(n12437), .B(n14764), .S(n10191), .Z(n10069) );
  MUX2_X1 U11897 ( .A(n14764), .B(n12437), .S(n10191), .Z(n10068) );
  INV_X1 U11898 ( .A(n10069), .ZN(n10070) );
  MUX2_X1 U11899 ( .A(n14763), .B(n12129), .S(n10191), .Z(n10074) );
  MUX2_X1 U11900 ( .A(n14763), .B(n12129), .S(n10182), .Z(n10071) );
  INV_X1 U11901 ( .A(n10073), .ZN(n10076) );
  INV_X1 U11902 ( .A(n10074), .ZN(n10075) );
  NAND2_X1 U11903 ( .A1(n10076), .A2(n10075), .ZN(n10077) );
  MUX2_X1 U11904 ( .A(n14762), .B(n16076), .S(n10182), .Z(n10079) );
  MUX2_X1 U11905 ( .A(n14762), .B(n16076), .S(n10191), .Z(n10078) );
  MUX2_X1 U11906 ( .A(n14761), .B(n14661), .S(n10191), .Z(n10082) );
  MUX2_X1 U11907 ( .A(n14761), .B(n14661), .S(n10182), .Z(n10080) );
  MUX2_X1 U11908 ( .A(n14760), .B(n14560), .S(n10182), .Z(n10084) );
  MUX2_X1 U11909 ( .A(n14760), .B(n14560), .S(n10191), .Z(n10083) );
  INV_X1 U11910 ( .A(n10084), .ZN(n10085) );
  MUX2_X1 U11911 ( .A(n14759), .B(n14703), .S(n10191), .Z(n10089) );
  NAND2_X1 U11912 ( .A1(n10088), .A2(n10089), .ZN(n10087) );
  MUX2_X1 U11913 ( .A(n14759), .B(n14703), .S(n10182), .Z(n10086) );
  INV_X1 U11914 ( .A(n10088), .ZN(n10091) );
  INV_X1 U11915 ( .A(n10089), .ZN(n10090) );
  NAND2_X1 U11916 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  MUX2_X1 U11917 ( .A(n14758), .B(n14387), .S(n10182), .Z(n10094) );
  MUX2_X1 U11918 ( .A(n14758), .B(n14387), .S(n10191), .Z(n10093) );
  MUX2_X1 U11919 ( .A(n14757), .B(n14679), .S(n10191), .Z(n10097) );
  MUX2_X1 U11920 ( .A(n14757), .B(n14679), .S(n10182), .Z(n10095) );
  MUX2_X1 U11921 ( .A(n14756), .B(n16177), .S(n10182), .Z(n10099) );
  MUX2_X1 U11922 ( .A(n14756), .B(n16177), .S(n10191), .Z(n10098) );
  INV_X1 U11923 ( .A(n10099), .ZN(n10100) );
  MUX2_X1 U11924 ( .A(n14755), .B(n14738), .S(n10191), .Z(n10104) );
  NAND2_X1 U11925 ( .A1(n10103), .A2(n10104), .ZN(n10102) );
  MUX2_X1 U11926 ( .A(n14755), .B(n14738), .S(n10182), .Z(n10101) );
  NAND2_X1 U11927 ( .A1(n10102), .A2(n10101), .ZN(n10108) );
  INV_X1 U11928 ( .A(n10103), .ZN(n10106) );
  INV_X1 U11929 ( .A(n10104), .ZN(n10105) );
  NAND2_X1 U11930 ( .A1(n10106), .A2(n10105), .ZN(n10107) );
  MUX2_X1 U11931 ( .A(n14754), .B(n16199), .S(n10182), .Z(n10111) );
  MUX2_X1 U11932 ( .A(n14754), .B(n16199), .S(n10191), .Z(n10110) );
  INV_X1 U11933 ( .A(n10111), .ZN(n10112) );
  MUX2_X1 U11934 ( .A(n14753), .B(n14449), .S(n10191), .Z(n10116) );
  NAND2_X1 U11935 ( .A1(n10115), .A2(n10116), .ZN(n10114) );
  MUX2_X1 U11936 ( .A(n14753), .B(n14449), .S(n10182), .Z(n10113) );
  MUX2_X1 U11937 ( .A(n15025), .B(n14752), .S(n10191), .Z(n10119) );
  MUX2_X1 U11938 ( .A(n15025), .B(n14752), .S(n10182), .Z(n10118) );
  MUX2_X1 U11939 ( .A(n14751), .B(n15105), .S(n10191), .Z(n10122) );
  MUX2_X1 U11940 ( .A(n15105), .B(n14751), .S(n10191), .Z(n10120) );
  MUX2_X1 U11941 ( .A(n14750), .B(n15099), .S(n10182), .Z(n10124) );
  MUX2_X1 U11942 ( .A(n14750), .B(n15099), .S(n10191), .Z(n10123) );
  INV_X1 U11943 ( .A(n10124), .ZN(n10125) );
  MUX2_X1 U11944 ( .A(n14749), .B(n15086), .S(n10191), .Z(n10129) );
  NAND2_X1 U11945 ( .A1(n10128), .A2(n10129), .ZN(n10127) );
  MUX2_X1 U11946 ( .A(n15086), .B(n14749), .S(n10191), .Z(n10126) );
  NAND2_X1 U11947 ( .A1(n10127), .A2(n10126), .ZN(n10133) );
  INV_X1 U11948 ( .A(n10128), .ZN(n10131) );
  INV_X1 U11949 ( .A(n10129), .ZN(n10130) );
  NAND2_X1 U11950 ( .A1(n10131), .A2(n10130), .ZN(n10132) );
  MUX2_X1 U11951 ( .A(n14748), .B(n15077), .S(n10182), .Z(n10135) );
  MUX2_X1 U11952 ( .A(n14748), .B(n15077), .S(n10191), .Z(n10134) );
  INV_X1 U11953 ( .A(n10135), .ZN(n10136) );
  MUX2_X1 U11954 ( .A(n14912), .B(n15073), .S(n10191), .Z(n10140) );
  NAND2_X1 U11955 ( .A1(n10139), .A2(n10140), .ZN(n10138) );
  MUX2_X1 U11956 ( .A(n14912), .B(n15073), .S(n10182), .Z(n10137) );
  MUX2_X1 U11957 ( .A(n15063), .B(n14747), .S(n10191), .Z(n10143) );
  MUX2_X1 U11958 ( .A(n14747), .B(n15063), .S(n10191), .Z(n10142) );
  MUX2_X1 U11959 ( .A(n14913), .B(n15055), .S(n10191), .Z(n10145) );
  MUX2_X1 U11960 ( .A(n14913), .B(n15055), .S(n10109), .Z(n10144) );
  INV_X1 U11961 ( .A(n10145), .ZN(n10146) );
  MUX2_X1 U11962 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10986), .Z(n10150) );
  XNOR2_X1 U11963 ( .A(n10150), .B(SI_30_), .ZN(n10169) );
  MUX2_X1 U11964 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10986), .Z(n10151) );
  XNOR2_X1 U11965 ( .A(n10151), .B(SI_31_), .ZN(n10152) );
  XNOR2_X1 U11966 ( .A(n10153), .B(n10152), .ZN(n14364) );
  NAND2_X1 U11967 ( .A1(n14364), .A2(n10171), .ZN(n10155) );
  NAND2_X1 U11968 ( .A1(n8972), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10154) );
  INV_X1 U11969 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U11970 ( .A1(n10156), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U11971 ( .A1(n10157), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n10158) );
  OAI211_X1 U11972 ( .C1(n10161), .C2(n10160), .A(n10159), .B(n10158), .ZN(
        n14840) );
  NAND2_X1 U11973 ( .A1(n10191), .A2(n14840), .ZN(n10237) );
  OR2_X1 U11974 ( .A1(n10245), .A2(n10237), .ZN(n10165) );
  NAND2_X1 U11975 ( .A1(n11438), .A2(n14835), .ZN(n12153) );
  OAI21_X1 U11976 ( .B1(n15162), .B2(n7860), .A(n11552), .ZN(n10162) );
  AND2_X1 U11977 ( .A1(n12153), .A2(n10162), .ZN(n10243) );
  INV_X1 U11978 ( .A(n10243), .ZN(n10163) );
  AND2_X1 U11979 ( .A1(n10163), .A2(n10232), .ZN(n10235) );
  INV_X1 U11980 ( .A(n14840), .ZN(n10236) );
  AND2_X1 U11981 ( .A1(n10182), .A2(n10236), .ZN(n10239) );
  NAND2_X1 U11982 ( .A1(n10245), .A2(n10239), .ZN(n10164) );
  OAI21_X1 U11983 ( .B1(n10166), .B2(n14840), .A(n14742), .ZN(n10167) );
  INV_X1 U11984 ( .A(n10167), .ZN(n10174) );
  INV_X1 U11985 ( .A(n10169), .ZN(n10170) );
  NAND2_X1 U11986 ( .A1(n13351), .A2(n10171), .ZN(n10173) );
  NAND2_X1 U11987 ( .A1(n8972), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n10172) );
  MUX2_X1 U11988 ( .A(n10174), .B(n14848), .S(n10182), .Z(n10196) );
  INV_X1 U11989 ( .A(n10196), .ZN(n10180) );
  AND2_X1 U11990 ( .A1(n14840), .A2(n7860), .ZN(n10176) );
  MUX2_X1 U11991 ( .A(n7861), .B(n10176), .S(n10175), .Z(n10177) );
  AND2_X1 U11992 ( .A1(n10177), .A2(n14742), .ZN(n10178) );
  AOI21_X1 U11993 ( .B1(n14848), .B2(n10191), .A(n10178), .ZN(n10195) );
  INV_X1 U11994 ( .A(n10195), .ZN(n10179) );
  NAND2_X1 U11995 ( .A1(n10180), .A2(n10179), .ZN(n10254) );
  AND2_X1 U11996 ( .A1(n10233), .A2(n10254), .ZN(n10252) );
  INV_X1 U11997 ( .A(n10252), .ZN(n10185) );
  INV_X1 U11998 ( .A(n14594), .ZN(n14743) );
  MUX2_X1 U11999 ( .A(n14743), .B(n10181), .S(n10182), .Z(n10197) );
  INV_X1 U12000 ( .A(n10197), .ZN(n10184) );
  MUX2_X1 U12001 ( .A(n14858), .B(n14594), .S(n10182), .Z(n10198) );
  INV_X1 U12002 ( .A(n10198), .ZN(n10183) );
  AND2_X1 U12003 ( .A1(n10184), .A2(n10183), .ZN(n10276) );
  OR2_X1 U12004 ( .A1(n10185), .A2(n10276), .ZN(n10259) );
  MUX2_X1 U12005 ( .A(n14878), .B(n14744), .S(n10191), .Z(n10200) );
  INV_X1 U12006 ( .A(n10200), .ZN(n10186) );
  MUX2_X1 U12007 ( .A(n14878), .B(n14744), .S(n10182), .Z(n10199) );
  NAND2_X1 U12008 ( .A1(n10186), .A2(n10199), .ZN(n10261) );
  INV_X1 U12009 ( .A(n10261), .ZN(n10187) );
  NOR2_X1 U12010 ( .A1(n10259), .A2(n10187), .ZN(n10275) );
  MUX2_X1 U12011 ( .A(n14745), .B(n15042), .S(n10182), .Z(n10202) );
  INV_X1 U12012 ( .A(n10202), .ZN(n10190) );
  MUX2_X1 U12013 ( .A(n14595), .B(n14383), .S(n10188), .Z(n10203) );
  INV_X1 U12014 ( .A(n10203), .ZN(n10189) );
  NAND2_X1 U12015 ( .A1(n10190), .A2(n10189), .ZN(n10273) );
  NAND2_X1 U12016 ( .A1(n10275), .A2(n10273), .ZN(n10271) );
  MUX2_X1 U12017 ( .A(n15047), .B(n14746), .S(n10191), .Z(n10269) );
  INV_X1 U12018 ( .A(n10269), .ZN(n10192) );
  MUX2_X1 U12019 ( .A(n14746), .B(n15047), .S(n10191), .Z(n10268) );
  NAND2_X1 U12020 ( .A1(n10192), .A2(n10268), .ZN(n10283) );
  INV_X1 U12021 ( .A(n10283), .ZN(n10193) );
  NOR2_X1 U12022 ( .A1(n10271), .A2(n10193), .ZN(n10194) );
  NAND2_X1 U12023 ( .A1(n10289), .A2(n10194), .ZN(n10285) );
  XNOR2_X1 U12024 ( .A(n10245), .B(n14840), .ZN(n10204) );
  NAND2_X1 U12025 ( .A1(n10204), .A2(n10243), .ZN(n10255) );
  AND2_X1 U12026 ( .A1(n10196), .A2(n10195), .ZN(n10234) );
  OR2_X1 U12027 ( .A1(n10255), .A2(n10234), .ZN(n10278) );
  AND2_X1 U12028 ( .A1(n10198), .A2(n10197), .ZN(n10253) );
  NOR2_X1 U12029 ( .A1(n10278), .A2(n10253), .ZN(n10260) );
  INV_X1 U12030 ( .A(n10199), .ZN(n10201) );
  NAND2_X1 U12031 ( .A1(n10201), .A2(n10200), .ZN(n10258) );
  AND2_X1 U12032 ( .A1(n10260), .A2(n10258), .ZN(n10272) );
  NAND2_X1 U12033 ( .A1(n10203), .A2(n10202), .ZN(n10279) );
  NAND2_X1 U12034 ( .A1(n10272), .A2(n10279), .ZN(n10287) );
  INV_X1 U12035 ( .A(n10204), .ZN(n10230) );
  XOR2_X1 U12036 ( .A(n14742), .B(n14848), .Z(n10229) );
  AND2_X1 U12037 ( .A1(n10206), .A2(n10205), .ZN(n15882) );
  NAND4_X1 U12038 ( .A1(n15882), .A2(n15920), .A3(n11584), .A4(n12270), .ZN(
        n10209) );
  NOR2_X1 U12039 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  NAND4_X1 U12040 ( .A1(n10211), .A2(n10210), .A3(n11803), .A4(n11628), .ZN(
        n10212) );
  NOR2_X1 U12041 ( .A1(n12252), .A2(n10212), .ZN(n10213) );
  NAND4_X1 U12042 ( .A1(n10214), .A2(n12200), .A3(n10215), .A4(n10213), .ZN(
        n10216) );
  NOR2_X1 U12043 ( .A1(n12483), .A2(n10216), .ZN(n10217) );
  NAND4_X1 U12044 ( .A1(n10218), .A2(n10217), .A3(n12633), .A4(n12459), .ZN(
        n10219) );
  NOR2_X1 U12045 ( .A1(n12856), .A2(n10219), .ZN(n10220) );
  NAND3_X1 U12046 ( .A1(n15004), .A2(n10220), .A3(n12934), .ZN(n10221) );
  NOR2_X1 U12047 ( .A1(n14963), .A2(n10221), .ZN(n10223) );
  NOR4_X1 U12048 ( .A1(n14884), .A2(n14898), .A3(n10224), .A4(n14945), .ZN(
        n10226) );
  NAND4_X1 U12049 ( .A1(n14871), .A2(n10226), .A3(n13069), .A4(n10225), .ZN(
        n10228) );
  NOR4_X1 U12050 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n10231) );
  XOR2_X1 U12051 ( .A(n14835), .B(n10231), .Z(n10266) );
  INV_X1 U12052 ( .A(n10232), .ZN(n10265) );
  INV_X1 U12053 ( .A(n10233), .ZN(n10250) );
  INV_X1 U12054 ( .A(n10234), .ZN(n10249) );
  INV_X1 U12055 ( .A(n10235), .ZN(n10240) );
  NOR2_X1 U12056 ( .A1(n10240), .A2(n10236), .ZN(n10238) );
  MUX2_X1 U12057 ( .A(n10243), .B(n10238), .S(n10237), .Z(n10247) );
  INV_X1 U12058 ( .A(n10239), .ZN(n10242) );
  OAI21_X1 U12059 ( .B1(n14840), .B2(n10240), .A(n10242), .ZN(n10241) );
  OAI21_X1 U12060 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(n10244) );
  NAND2_X1 U12061 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  OAI21_X1 U12062 ( .B1(n10245), .B2(n10247), .A(n10246), .ZN(n10248) );
  OAI21_X1 U12063 ( .B1(n10250), .B2(n10249), .A(n10248), .ZN(n10251) );
  OR2_X1 U12064 ( .A1(n10255), .A2(n10254), .ZN(n10256) );
  OAI211_X1 U12065 ( .C1(n10259), .C2(n10258), .A(n10257), .B(n10256), .ZN(
        n10264) );
  INV_X1 U12066 ( .A(n10260), .ZN(n10262) );
  NOR2_X1 U12067 ( .A1(n10262), .A2(n10261), .ZN(n10263) );
  AOI211_X1 U12068 ( .C1(n10266), .C2(n10265), .A(n10264), .B(n10263), .ZN(
        n10267) );
  INV_X1 U12069 ( .A(n10268), .ZN(n10270) );
  NAND2_X1 U12070 ( .A1(n10270), .A2(n10269), .ZN(n10286) );
  INV_X1 U12071 ( .A(n10272), .ZN(n10274) );
  NOR2_X1 U12072 ( .A1(n10274), .A2(n10273), .ZN(n10282) );
  INV_X1 U12073 ( .A(n10275), .ZN(n10280) );
  INV_X1 U12074 ( .A(n10276), .ZN(n10277) );
  OAI22_X1 U12075 ( .A1(n10280), .A2(n10279), .B1(n10278), .B2(n10277), .ZN(
        n10281) );
  NAND2_X1 U12076 ( .A1(n10285), .A2(n10284), .ZN(n10292) );
  INV_X1 U12077 ( .A(n10286), .ZN(n10288) );
  NOR3_X1 U12078 ( .A1(n10289), .A2(n10288), .A3(n10287), .ZN(n10291) );
  INV_X1 U12079 ( .A(n11845), .ZN(n10290) );
  NAND2_X1 U12080 ( .A1(n10290), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11034) );
  OAI21_X1 U12081 ( .B1(n10292), .B2(n10291), .A(n12732), .ZN(n10295) );
  INV_X1 U12082 ( .A(n13009), .ZN(n15518) );
  NAND3_X1 U12083 ( .A1(n11561), .A2(n15518), .A3(n15925), .ZN(n10293) );
  OAI211_X1 U12084 ( .C1(n15162), .C2(n11034), .A(n10293), .B(P1_B_REG_SCAN_IN), .ZN(n10294) );
  NAND2_X1 U12085 ( .A1(n10295), .A2(n10294), .ZN(P1_U3242) );
  INV_X1 U12086 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n10296) );
  NOR2_X1 U12087 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n10296), .ZN(n10328) );
  INV_X1 U12088 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15543) );
  AOI22_X1 U12089 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .B1(n15543), .B2(n10296), .ZN(n10334) );
  INV_X1 U12090 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10326) );
  XNOR2_X1 U12091 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10381) );
  INV_X1 U12092 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10324) );
  XNOR2_X1 U12093 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10380) );
  XNOR2_X1 U12094 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n10322), .ZN(n10375) );
  INV_X1 U12095 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n10297) );
  NOR2_X1 U12096 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n10297), .ZN(n10320) );
  INV_X1 U12097 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n10318) );
  INV_X1 U12098 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n10316) );
  INV_X1 U12099 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10314) );
  XNOR2_X1 U12100 ( .A(n10314), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n10364) );
  AND2_X1 U12101 ( .A1(n10306), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10305) );
  INV_X1 U12102 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U12103 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n10347), .ZN(n10346) );
  XNOR2_X1 U12104 ( .A(n10300), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n10340) );
  NOR2_X1 U12105 ( .A1(n10341), .A2(n10340), .ZN(n10299) );
  NOR2_X1 U12106 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n15875), .ZN(n10304) );
  NAND2_X1 U12107 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n10309), .ZN(n10312) );
  XOR2_X1 U12108 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n10309), .Z(n10361) );
  INV_X1 U12109 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U12110 ( .A1(n10361), .A2(n10310), .ZN(n10311) );
  NAND2_X1 U12111 ( .A1(n10312), .A2(n10311), .ZN(n10363) );
  NOR2_X1 U12112 ( .A1(n10364), .A2(n10363), .ZN(n10313) );
  XOR2_X1 U12113 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n10368) );
  XNOR2_X1 U12114 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10335) );
  NAND2_X1 U12115 ( .A1(n10336), .A2(n10335), .ZN(n10317) );
  INV_X1 U12116 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U12117 ( .A1(n10380), .A2(n10379), .ZN(n10323) );
  NAND2_X1 U12118 ( .A1(n10381), .A2(n10382), .ZN(n10325) );
  NOR2_X1 U12119 ( .A1(n10334), .A2(n10333), .ZN(n10327) );
  NOR2_X1 U12120 ( .A1(n10328), .A2(n10327), .ZN(n10329) );
  NAND2_X1 U12121 ( .A1(n10329), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n10331) );
  XNOR2_X1 U12122 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n10329), .ZN(n10332) );
  NAND2_X1 U12123 ( .A1(n10331), .A2(n10330), .ZN(n10390) );
  XOR2_X1 U12124 ( .A(n10390), .B(P1_ADDR_REG_17__SCAN_IN), .Z(n10392) );
  XOR2_X1 U12125 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n10392), .Z(n10388) );
  INV_X1 U12126 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10387) );
  NOR2_X1 U12127 ( .A1(n10388), .A2(n10387), .ZN(n10389) );
  XOR2_X1 U12128 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n10332), .Z(n10386) );
  XNOR2_X1 U12129 ( .A(n10334), .B(n10333), .ZN(n10384) );
  XOR2_X1 U12130 ( .A(n10336), .B(n10335), .Z(n15570) );
  AND2_X1 U12131 ( .A1(n10338), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10353) );
  XNOR2_X1 U12132 ( .A(n10338), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15554) );
  XOR2_X1 U12133 ( .A(n10341), .B(n10340), .Z(n15547) );
  INV_X1 U12134 ( .A(n10342), .ZN(n10343) );
  INV_X1 U12135 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10344) );
  NOR2_X1 U12136 ( .A1(n10345), .A2(n10344), .ZN(n10348) );
  OAI21_X1 U12137 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n10347), .A(n10346), .ZN(
        n15544) );
  NAND2_X1 U12138 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15544), .ZN(n15607) );
  NOR2_X1 U12139 ( .A1(n15608), .A2(n15607), .ZN(n15606) );
  NOR2_X1 U12140 ( .A1(n15547), .A2(n15546), .ZN(n10349) );
  NAND2_X1 U12141 ( .A1(n15547), .A2(n15546), .ZN(n15545) );
  OAI21_X1 U12142 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n10349), .A(n15545), .ZN(
        n10351) );
  NAND2_X1 U12143 ( .A1(n10350), .A2(n10351), .ZN(n10352) );
  INV_X1 U12144 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15550) );
  NAND2_X1 U12145 ( .A1(n15551), .A2(n15550), .ZN(n15549) );
  NAND2_X1 U12146 ( .A1(n10352), .A2(n15549), .ZN(n15553) );
  NOR2_X1 U12147 ( .A1(n15554), .A2(n15553), .ZN(n15552) );
  XNOR2_X1 U12148 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10355) );
  XOR2_X1 U12149 ( .A(n10355), .B(n10354), .Z(n10357) );
  INV_X1 U12150 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15556) );
  XNOR2_X1 U12151 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10359) );
  XNOR2_X1 U12152 ( .A(n10359), .B(n10358), .ZN(n15603) );
  INV_X1 U12153 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10360) );
  XNOR2_X1 U12154 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10361), .ZN(n15560) );
  XNOR2_X1 U12155 ( .A(n10364), .B(n10363), .ZN(n10366) );
  NOR2_X1 U12156 ( .A1(n10365), .A2(n10366), .ZN(n10367) );
  INV_X1 U12157 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15562) );
  XNOR2_X1 U12158 ( .A(n10369), .B(n10368), .ZN(n15565) );
  NAND2_X1 U12159 ( .A1(n15566), .A2(n15565), .ZN(n10370) );
  XNOR2_X1 U12160 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10372) );
  XOR2_X1 U12161 ( .A(n10372), .B(n10371), .Z(n15573) );
  XOR2_X1 U12162 ( .A(n10375), .B(n10374), .Z(n10376) );
  NAND2_X1 U12163 ( .A1(n10377), .A2(n10376), .ZN(n10378) );
  INV_X1 U12164 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15577) );
  XNOR2_X1 U12165 ( .A(n10380), .B(n10379), .ZN(n15580) );
  NAND2_X1 U12166 ( .A1(n15581), .A2(n15580), .ZN(n15579) );
  XNOR2_X1 U12167 ( .A(n10382), .B(n10381), .ZN(n15584) );
  INV_X1 U12168 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15591) );
  INV_X1 U12169 ( .A(n15593), .ZN(n15594) );
  INV_X1 U12170 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15596) );
  NAND2_X1 U12171 ( .A1(n15594), .A2(n15592), .ZN(n15599) );
  XNOR2_X1 U12172 ( .A(n10388), .B(n10387), .ZN(n15598) );
  NOR2_X1 U12173 ( .A1(n15599), .A2(n15598), .ZN(n15597) );
  XNOR2_X1 U12174 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n10396) );
  NAND2_X1 U12175 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n10390), .ZN(n10394) );
  INV_X1 U12176 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U12177 ( .A1(n10392), .A2(n10391), .ZN(n10393) );
  NAND2_X1 U12178 ( .A1(n10394), .A2(n10393), .ZN(n10395) );
  XNOR2_X1 U12179 ( .A(n10396), .B(n10395), .ZN(n15600) );
  INV_X1 U12180 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U12181 ( .A1(n10396), .A2(n10395), .ZN(n10397) );
  OAI21_X1 U12182 ( .B1(n10398), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n10397), 
        .ZN(n10399) );
  INV_X1 U12183 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10401) );
  OR2_X1 U12184 ( .A1(n16169), .A2(n10401), .ZN(n10402) );
  INV_X1 U12185 ( .A(n10403), .ZN(n10404) );
  OAI21_X1 U12186 ( .B1(n10405), .B2(n16166), .A(n10404), .ZN(P3_U3456) );
  NOR2_X1 U12187 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n10409) );
  INV_X2 U12188 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n10460) );
  NOR2_X1 U12189 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n10410) );
  INV_X1 U12190 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n10414) );
  INV_X1 U12191 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U12192 ( .A1(n13357), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10429) );
  NAND2_X2 U12193 ( .A1(n10417), .A2(n14372), .ZN(n10519) );
  INV_X1 U12194 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12406) );
  OR2_X1 U12195 ( .A1(n10519), .A2(n12406), .ZN(n10428) );
  NAND3_X1 U12196 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n10593) );
  INV_X1 U12197 ( .A(n10593), .ZN(n10418) );
  NAND2_X1 U12198 ( .A1(n10418), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10610) );
  INV_X1 U12199 ( .A(n10610), .ZN(n10419) );
  NAND2_X1 U12200 ( .A1(n10419), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10612) );
  INV_X1 U12201 ( .A(n10612), .ZN(n10420) );
  NAND2_X1 U12202 ( .A1(n10420), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10492) );
  INV_X1 U12203 ( .A(n10492), .ZN(n10422) );
  AND2_X1 U12204 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n10421) );
  NAND2_X1 U12205 ( .A1(n10422), .A2(n10421), .ZN(n10635) );
  NAND2_X1 U12206 ( .A1(n10637), .A2(n10423), .ZN(n10424) );
  NAND2_X1 U12207 ( .A1(n10655), .A2(n10424), .ZN(n12553) );
  OR2_X1 U12208 ( .A1(n10943), .A2(n12553), .ZN(n10427) );
  INV_X1 U12209 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n12420) );
  OR2_X1 U12210 ( .A1(n10553), .A2(n12420), .ZN(n10426) );
  NAND4_X1 U12211 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n14017) );
  NOR2_X1 U12212 ( .A1(n10431), .A2(n10415), .ZN(n10434) );
  NAND2_X1 U12213 ( .A1(n10431), .A2(n10430), .ZN(n10911) );
  NAND2_X1 U12214 ( .A1(n10911), .A2(n10432), .ZN(n10433) );
  NAND2_X1 U12215 ( .A1(n12624), .A2(n13452), .ZN(n15896) );
  NAND2_X1 U12216 ( .A1(n10442), .A2(n10441), .ZN(n10443) );
  XNOR2_X2 U12217 ( .A(n10446), .B(n10445), .ZN(n13024) );
  NAND2_X1 U12218 ( .A1(n14017), .A2(n10938), .ZN(n10644) );
  INV_X1 U12219 ( .A(n10644), .ZN(n10647) );
  NAND2_X1 U12220 ( .A1(n11361), .A2(n13350), .ZN(n10457) );
  INV_X2 U12221 ( .A(n10546), .ZN(n10741) );
  NAND2_X1 U12222 ( .A1(n7218), .A2(n10449), .ZN(n10571) );
  NOR2_X1 U12223 ( .A1(n10708), .A2(n10450), .ZN(n10453) );
  NOR2_X1 U12224 ( .A1(n10453), .A2(n10415), .ZN(n10451) );
  MUX2_X1 U12225 ( .A(n10415), .B(n10451), .S(P2_IR_REG_12__SCAN_IN), .Z(
        n10455) );
  INV_X1 U12226 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U12227 ( .A1(n10453), .A2(n10452), .ZN(n10649) );
  INV_X1 U12228 ( .A(n10649), .ZN(n10454) );
  OR2_X1 U12229 ( .A1(n10455), .A2(n10454), .ZN(n12421) );
  INV_X1 U12230 ( .A(n12421), .ZN(n15503) );
  AOI22_X1 U12231 ( .A1(n10741), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10740), 
        .B2(n15503), .ZN(n10456) );
  OR2_X1 U12232 ( .A1(n12624), .A2(n10458), .ZN(n10459) );
  NAND2_X4 U12233 ( .A1(n10459), .A2(n13136), .ZN(n10835) );
  XNOR2_X1 U12234 ( .A(n13237), .B(n10835), .ZN(n10646) );
  INV_X1 U12235 ( .A(n10708), .ZN(n10461) );
  NAND2_X1 U12236 ( .A1(n10461), .A2(n10460), .ZN(n10605) );
  INV_X1 U12237 ( .A(n10605), .ZN(n10463) );
  INV_X1 U12238 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U12239 ( .A1(n10463), .A2(n10462), .ZN(n10484) );
  NAND2_X1 U12240 ( .A1(n10631), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10464) );
  XNOR2_X1 U12241 ( .A(n10464), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U12242 ( .A1(n10740), .A2(n11193), .B1(n10741), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n10465) );
  XNOR2_X1 U12243 ( .A(n13216), .B(n10835), .ZN(n10627) );
  INV_X1 U12244 ( .A(n10627), .ZN(n10630) );
  NAND2_X1 U12245 ( .A1(n13357), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10472) );
  INV_X1 U12246 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10466) );
  OR2_X1 U12247 ( .A1(n10553), .A2(n10466), .ZN(n10471) );
  INV_X1 U12248 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10477) );
  INV_X1 U12249 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10467) );
  OAI21_X1 U12250 ( .B1(n10492), .B2(n10477), .A(n10467), .ZN(n10468) );
  NAND2_X1 U12251 ( .A1(n10468), .A2(n10635), .ZN(n12590) );
  OR2_X1 U12252 ( .A1(n10943), .A2(n12590), .ZN(n10470) );
  INV_X1 U12253 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11274) );
  OR2_X1 U12254 ( .A1(n10519), .A2(n11274), .ZN(n10469) );
  NAND4_X1 U12255 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .ZN(
        n14019) );
  NAND2_X1 U12256 ( .A1(n14019), .A2(n10938), .ZN(n10629) );
  NAND2_X1 U12257 ( .A1(n10486), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10473) );
  MUX2_X1 U12258 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10473), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n10474) );
  NAND2_X1 U12259 ( .A1(n10474), .A2(n10631), .ZN(n11201) );
  INV_X1 U12260 ( .A(n11201), .ZN(n11192) );
  AOI22_X1 U12261 ( .A1(n10740), .A2(n11192), .B1(n10741), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n10475) );
  INV_X1 U12262 ( .A(n10624), .ZN(n12143) );
  NAND2_X1 U12263 ( .A1(n13357), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10482) );
  INV_X1 U12264 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n12174) );
  OR2_X1 U12265 ( .A1(n10519), .A2(n12174), .ZN(n10481) );
  XNOR2_X1 U12266 ( .A(n10492), .B(n10477), .ZN(n12173) );
  OR2_X1 U12267 ( .A1(n10943), .A2(n12173), .ZN(n10480) );
  INV_X1 U12268 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10478) );
  OR2_X1 U12269 ( .A1(n10553), .A2(n10478), .ZN(n10479) );
  NAND4_X1 U12270 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n14020) );
  INV_X1 U12271 ( .A(n14020), .ZN(n13212) );
  NOR2_X1 U12272 ( .A1(n13212), .A2(n11781), .ZN(n10623) );
  INV_X1 U12273 ( .A(n10623), .ZN(n10626) );
  NAND2_X1 U12274 ( .A1(n10484), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10485) );
  MUX2_X1 U12275 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10485), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n10487) );
  AOI22_X1 U12276 ( .A1(n10741), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10740), 
        .B2(n11070), .ZN(n10488) );
  NAND2_X1 U12277 ( .A1(n13357), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n10497) );
  INV_X1 U12278 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n12084) );
  OR2_X1 U12279 ( .A1(n10519), .A2(n12084), .ZN(n10496) );
  INV_X1 U12280 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U12281 ( .A1(n10612), .A2(n10490), .ZN(n10491) );
  NAND2_X1 U12282 ( .A1(n10492), .A2(n10491), .ZN(n12083) );
  OR2_X1 U12283 ( .A1(n10943), .A2(n12083), .ZN(n10495) );
  INV_X1 U12284 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10493) );
  OR2_X1 U12285 ( .A1(n10553), .A2(n10493), .ZN(n10494) );
  NAND4_X1 U12286 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n14021) );
  NAND2_X1 U12287 ( .A1(n14021), .A2(n10938), .ZN(n10622) );
  NAND2_X1 U12288 ( .A1(n10981), .A2(n13350), .ZN(n10502) );
  NOR2_X1 U12289 ( .A1(n7218), .A2(n10415), .ZN(n10498) );
  MUX2_X1 U12290 ( .A(n10415), .B(n10498), .S(P2_IR_REG_4__SCAN_IN), .Z(n10500) );
  INV_X1 U12291 ( .A(n10571), .ZN(n10499) );
  NOR2_X1 U12292 ( .A1(n10500), .A2(n10499), .ZN(n15444) );
  AOI22_X1 U12293 ( .A1(n10741), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10740), 
        .B2(n15444), .ZN(n10501) );
  NAND2_X1 U12294 ( .A1(n10502), .A2(n10501), .ZN(n13176) );
  XNOR2_X1 U12295 ( .A(n13176), .B(n10835), .ZN(n10568) );
  INV_X1 U12296 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n11063) );
  OR2_X1 U12297 ( .A1(n10553), .A2(n11063), .ZN(n10507) );
  INV_X1 U12298 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10503) );
  OR2_X1 U12299 ( .A1(n10551), .A2(n10503), .ZN(n10506) );
  XNOR2_X1 U12300 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n12042) );
  OR2_X1 U12301 ( .A1(n10943), .A2(n12042), .ZN(n10505) );
  NAND2_X1 U12302 ( .A1(n10552), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10504) );
  NAND2_X1 U12303 ( .A1(n14025), .A2(n10938), .ZN(n10569) );
  XNOR2_X1 U12304 ( .A(n10568), .B(n10569), .ZN(n11600) );
  NAND2_X1 U12305 ( .A1(n15395), .A2(n13350), .ZN(n10511) );
  MUX2_X1 U12306 ( .A(n10415), .B(n10508), .S(P2_IR_REG_3__SCAN_IN), .Z(n10509) );
  NOR2_X1 U12307 ( .A1(n10509), .A2(n7218), .ZN(n11062) );
  AOI22_X1 U12308 ( .A1(n10741), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n10740), 
        .B2(n11062), .ZN(n10510) );
  XNOR2_X1 U12309 ( .A(n13168), .B(n10835), .ZN(n11597) );
  NAND2_X1 U12310 ( .A1(n10552), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10517) );
  INV_X1 U12311 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10512) );
  OR2_X1 U12312 ( .A1(n10551), .A2(n10512), .ZN(n10516) );
  INV_X1 U12313 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10513) );
  OR2_X1 U12314 ( .A1(n10553), .A2(n10513), .ZN(n10514) );
  NAND2_X1 U12315 ( .A1(n11597), .A2(n10518), .ZN(n10566) );
  AND2_X1 U12316 ( .A1(n11600), .A2(n10566), .ZN(n10567) );
  OR2_X1 U12317 ( .A1(n7192), .A2(n15901), .ZN(n10521) );
  INV_X1 U12318 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11130) );
  OR2_X1 U12319 ( .A1(n10519), .A2(n11130), .ZN(n10520) );
  AND2_X1 U12320 ( .A1(n10521), .A2(n10520), .ZN(n10525) );
  INV_X1 U12321 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10522) );
  OR2_X1 U12322 ( .A1(n10551), .A2(n10522), .ZN(n10524) );
  INV_X1 U12323 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11133) );
  INV_X1 U12324 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n15418) );
  NAND2_X1 U12325 ( .A1(n10986), .A2(SI_0_), .ZN(n10527) );
  XNOR2_X1 U12326 ( .A(n10526), .B(n10527), .ZN(n14379) );
  INV_X1 U12327 ( .A(n15895), .ZN(n13135) );
  NAND2_X1 U12328 ( .A1(n11452), .A2(n10938), .ZN(n11489) );
  NAND2_X1 U12329 ( .A1(n15895), .A2(n10857), .ZN(n10529) );
  AND2_X1 U12330 ( .A1(n11489), .A2(n10529), .ZN(n11366) );
  INV_X1 U12331 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11703) );
  OR2_X1 U12332 ( .A1(n10943), .A2(n11703), .ZN(n10534) );
  INV_X1 U12333 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10530) );
  OR2_X1 U12334 ( .A1(n10551), .A2(n10530), .ZN(n10532) );
  INV_X1 U12335 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n11058) );
  OR2_X1 U12336 ( .A1(n10553), .A2(n11058), .ZN(n10531) );
  INV_X1 U12337 ( .A(n10546), .ZN(n10535) );
  NAND2_X1 U12338 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10536) );
  MUX2_X1 U12339 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10536), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n10539) );
  INV_X1 U12340 ( .A(n10537), .ZN(n10538) );
  NAND2_X1 U12341 ( .A1(n10539), .A2(n10538), .ZN(n11059) );
  NAND2_X1 U12342 ( .A1(n11366), .A2(n11365), .ZN(n10970) );
  INV_X1 U12343 ( .A(n10540), .ZN(n10542) );
  NAND2_X1 U12344 ( .A1(n10542), .A2(n10541), .ZN(n10543) );
  NAND2_X1 U12345 ( .A1(n10970), .A2(n10543), .ZN(n10558) );
  OR2_X1 U12346 ( .A1(n10537), .A2(n10415), .ZN(n10544) );
  XNOR2_X1 U12347 ( .A(n10545), .B(n10544), .ZN(n15429) );
  OAI22_X1 U12348 ( .A1(n10546), .A2(n10980), .B1(n11054), .B2(n15429), .ZN(
        n10547) );
  XNOR2_X1 U12349 ( .A(n14248), .B(n10835), .ZN(n10559) );
  INV_X1 U12350 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n14245) );
  INV_X1 U12351 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10550) );
  OR2_X1 U12352 ( .A1(n10551), .A2(n10550), .ZN(n10556) );
  INV_X1 U12353 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n11060) );
  OR2_X1 U12354 ( .A1(n10553), .A2(n11060), .ZN(n10554) );
  XNOR2_X1 U12355 ( .A(n10559), .B(n10560), .ZN(n10971) );
  INV_X1 U12356 ( .A(n10559), .ZN(n10561) );
  NAND2_X1 U12357 ( .A1(n10561), .A2(n10560), .ZN(n10562) );
  INV_X1 U12358 ( .A(n11597), .ZN(n10564) );
  INV_X1 U12359 ( .A(n10568), .ZN(n11482) );
  NAND2_X1 U12360 ( .A1(n11482), .A2(n10569), .ZN(n10570) );
  OR2_X1 U12361 ( .A1(n10984), .A2(n7191), .ZN(n10575) );
  NAND2_X1 U12362 ( .A1(n10571), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10572) );
  MUX2_X1 U12363 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10572), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n10573) );
  AND2_X1 U12364 ( .A1(n10573), .A2(n10708), .ZN(n11066) );
  AOI22_X1 U12365 ( .A1(n10741), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10740), 
        .B2(n11066), .ZN(n10574) );
  NAND2_X1 U12366 ( .A1(n10575), .A2(n10574), .ZN(n13182) );
  XNOR2_X1 U12367 ( .A(n13182), .B(n10835), .ZN(n10584) );
  NAND2_X1 U12368 ( .A1(n10552), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10583) );
  INV_X1 U12369 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10576) );
  OR2_X1 U12370 ( .A1(n10551), .A2(n10576), .ZN(n10582) );
  INV_X1 U12371 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10578) );
  NAND2_X1 U12372 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10577) );
  NAND2_X1 U12373 ( .A1(n10578), .A2(n10577), .ZN(n10579) );
  NAND2_X1 U12374 ( .A1(n10593), .A2(n10579), .ZN(n11786) );
  OR2_X1 U12375 ( .A1(n10943), .A2(n11786), .ZN(n10581) );
  INV_X1 U12376 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11065) );
  OR2_X1 U12377 ( .A1(n10553), .A2(n11065), .ZN(n10580) );
  NAND4_X1 U12378 ( .A1(n10583), .A2(n10582), .A3(n10581), .A4(n10580), .ZN(
        n14024) );
  NAND2_X1 U12379 ( .A1(n14024), .A2(n10938), .ZN(n10585) );
  XNOR2_X1 U12380 ( .A(n10584), .B(n10585), .ZN(n11483) );
  INV_X1 U12381 ( .A(n10584), .ZN(n10586) );
  NAND2_X1 U12382 ( .A1(n10586), .A2(n10585), .ZN(n10587) );
  OR2_X1 U12383 ( .A1(n10995), .A2(n7191), .ZN(n10590) );
  NAND2_X1 U12384 ( .A1(n10708), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10588) );
  XNOR2_X1 U12385 ( .A(n10588), .B(P2_IR_REG_6__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U12386 ( .A1(n10741), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10740), 
        .B2(n11067), .ZN(n10589) );
  NAND2_X1 U12387 ( .A1(n10590), .A2(n10589), .ZN(n16043) );
  XNOR2_X1 U12388 ( .A(n16043), .B(n10835), .ZN(n11734) );
  NAND2_X1 U12389 ( .A1(n13357), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n10598) );
  INV_X1 U12390 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10591) );
  OR2_X1 U12391 ( .A1(n10553), .A2(n10591), .ZN(n10597) );
  INV_X1 U12392 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U12393 ( .A1(n10593), .A2(n10592), .ZN(n10594) );
  NAND2_X1 U12394 ( .A1(n10610), .A2(n10594), .ZN(n16039) );
  OR2_X1 U12395 ( .A1(n10943), .A2(n16039), .ZN(n10596) );
  INV_X1 U12396 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n16040) );
  OR2_X1 U12397 ( .A1(n10519), .A2(n16040), .ZN(n10595) );
  NAND4_X1 U12398 ( .A1(n10598), .A2(n10597), .A3(n10596), .A4(n10595), .ZN(
        n14023) );
  AND2_X1 U12399 ( .A1(n14023), .A2(n10938), .ZN(n10599) );
  NAND2_X1 U12400 ( .A1(n11734), .A2(n10599), .ZN(n10617) );
  INV_X1 U12401 ( .A(n11734), .ZN(n10601) );
  INV_X1 U12402 ( .A(n10599), .ZN(n10600) );
  NAND2_X1 U12403 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  NAND2_X1 U12404 ( .A1(n10617), .A2(n10602), .ZN(n11636) );
  OR2_X1 U12405 ( .A1(n11019), .A2(n7191), .ZN(n10608) );
  NAND2_X1 U12406 ( .A1(n10605), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10606) );
  XNOR2_X1 U12407 ( .A(n10606), .B(P2_IR_REG_7__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U12408 ( .A1(n10741), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10740), 
        .B2(n11069), .ZN(n10607) );
  NAND2_X1 U12409 ( .A1(n13357), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n10616) );
  INV_X1 U12410 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11051) );
  OR2_X1 U12411 ( .A1(n10519), .A2(n11051), .ZN(n10615) );
  INV_X1 U12412 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U12413 ( .A1(n10610), .A2(n10609), .ZN(n10611) );
  NAND2_X1 U12414 ( .A1(n10612), .A2(n10611), .ZN(n12185) );
  OR2_X1 U12415 ( .A1(n10943), .A2(n12185), .ZN(n10614) );
  INV_X1 U12416 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11068) );
  OR2_X1 U12417 ( .A1(n10553), .A2(n11068), .ZN(n10613) );
  NAND4_X1 U12418 ( .A1(n10616), .A2(n10615), .A3(n10614), .A4(n10613), .ZN(
        n14022) );
  NAND2_X1 U12419 ( .A1(n14022), .A2(n10938), .ZN(n10620) );
  XNOR2_X1 U12420 ( .A(n10619), .B(n10620), .ZN(n11736) );
  INV_X1 U12421 ( .A(n10619), .ZN(n11865) );
  NAND2_X1 U12422 ( .A1(n11865), .A2(n10620), .ZN(n10621) );
  XNOR2_X1 U12423 ( .A(n11981), .B(n10622), .ZN(n11867) );
  AOI21_X1 U12424 ( .B1(n11981), .B2(n10622), .A(n11980), .ZN(n10625) );
  XNOR2_X1 U12425 ( .A(n10624), .B(n10623), .ZN(n11983) );
  NOR2_X1 U12426 ( .A1(n10625), .A2(n11983), .ZN(n11974) );
  AOI21_X1 U12427 ( .B1(n12143), .B2(n10626), .A(n11974), .ZN(n10628) );
  XOR2_X1 U12428 ( .A(n10629), .B(n10627), .Z(n12145) );
  NAND2_X1 U12429 ( .A1(n11186), .A2(n13350), .ZN(n10634) );
  OAI21_X1 U12430 ( .B1(n10631), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10632) );
  XNOR2_X1 U12431 ( .A(n10632), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11278) );
  AOI22_X1 U12432 ( .A1(n11278), .A2(n10740), .B1(n10741), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n10633) );
  XNOR2_X1 U12433 ( .A(n13224), .B(n10857), .ZN(n12548) );
  NAND2_X1 U12434 ( .A1(n13357), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10641) );
  INV_X1 U12435 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11279) );
  OR2_X1 U12436 ( .A1(n10553), .A2(n11279), .ZN(n10640) );
  NAND2_X1 U12437 ( .A1(n10635), .A2(n12473), .ZN(n10636) );
  NAND2_X1 U12438 ( .A1(n10637), .A2(n10636), .ZN(n12541) );
  OR2_X1 U12439 ( .A1(n10943), .A2(n12541), .ZN(n10639) );
  INV_X1 U12440 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n12542) );
  OR2_X1 U12441 ( .A1(n10519), .A2(n12542), .ZN(n10638) );
  NAND4_X1 U12442 ( .A1(n10641), .A2(n10640), .A3(n10639), .A4(n10638), .ZN(
        n14018) );
  NAND2_X1 U12443 ( .A1(n14018), .A2(n10938), .ZN(n10642) );
  NOR2_X1 U12444 ( .A1(n12548), .A2(n10642), .ZN(n10643) );
  AOI21_X1 U12445 ( .B1(n12548), .B2(n10642), .A(n10643), .ZN(n12472) );
  INV_X1 U12446 ( .A(n10643), .ZN(n10645) );
  XNOR2_X1 U12447 ( .A(n10646), .B(n10644), .ZN(n12550) );
  OR2_X1 U12448 ( .A1(n11394), .A2(n7191), .ZN(n10652) );
  NAND2_X1 U12449 ( .A1(n10649), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10648) );
  MUX2_X1 U12450 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10648), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n10650) );
  AOI22_X1 U12451 ( .A1(n10741), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10740), 
        .B2(n15489), .ZN(n10651) );
  XNOR2_X1 U12452 ( .A(n16148), .B(n10835), .ZN(n10662) );
  NAND2_X1 U12453 ( .A1(n10552), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10660) );
  INV_X1 U12454 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10653) );
  OR2_X1 U12455 ( .A1(n10551), .A2(n10653), .ZN(n10659) );
  INV_X1 U12456 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n12601) );
  NAND2_X1 U12457 ( .A1(n10655), .A2(n12601), .ZN(n10656) );
  NAND2_X1 U12458 ( .A1(n10669), .A2(n10656), .ZN(n16144) );
  OR2_X1 U12459 ( .A1(n10943), .A2(n16144), .ZN(n10658) );
  INV_X1 U12460 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12422) );
  OR2_X1 U12461 ( .A1(n10553), .A2(n12422), .ZN(n10657) );
  NAND4_X1 U12462 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(
        n13244) );
  AND2_X1 U12463 ( .A1(n13244), .A2(n10938), .ZN(n10661) );
  NOR2_X1 U12464 ( .A1(n10662), .A2(n10661), .ZN(n12596) );
  NAND2_X1 U12465 ( .A1(n10662), .A2(n10661), .ZN(n12597) );
  NAND2_X1 U12466 ( .A1(n11518), .A2(n13350), .ZN(n10665) );
  NAND2_X1 U12467 ( .A1(n10678), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10663) );
  XNOR2_X1 U12468 ( .A(n10663), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U12469 ( .A1(n10741), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n12424), 
        .B2(n10740), .ZN(n10664) );
  XNOR2_X1 U12470 ( .A(n13249), .B(n10857), .ZN(n10676) );
  NAND2_X1 U12471 ( .A1(n10552), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10674) );
  INV_X1 U12472 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10666) );
  OR2_X1 U12473 ( .A1(n10551), .A2(n10666), .ZN(n10673) );
  INV_X1 U12474 ( .A(n10669), .ZN(n10667) );
  NAND2_X1 U12475 ( .A1(n10667), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n10683) );
  INV_X1 U12476 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U12477 ( .A1(n10669), .A2(n10668), .ZN(n10670) );
  NAND2_X1 U12478 ( .A1(n10683), .A2(n10670), .ZN(n12832) );
  OR2_X1 U12479 ( .A1(n10943), .A2(n12832), .ZN(n10672) );
  INV_X1 U12480 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12425) );
  OR2_X1 U12481 ( .A1(n10553), .A2(n12425), .ZN(n10671) );
  NAND4_X1 U12482 ( .A1(n10674), .A2(n10673), .A3(n10672), .A4(n10671), .ZN(
        n14016) );
  NAND2_X1 U12483 ( .A1(n14016), .A2(n10938), .ZN(n10675) );
  NAND2_X1 U12484 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  OAI21_X1 U12485 ( .B1(n10676), .B2(n10675), .A(n10677), .ZN(n12739) );
  NAND2_X1 U12486 ( .A1(n11750), .A2(n13350), .ZN(n10681) );
  OAI21_X1 U12487 ( .B1(n10678), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10679) );
  XNOR2_X1 U12488 ( .A(n10679), .B(P2_IR_REG_15__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U12489 ( .A1(n12426), .A2(n10740), .B1(n10741), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n10680) );
  XNOR2_X1 U12490 ( .A(n14342), .B(n10835), .ZN(n10693) );
  INV_X1 U12491 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10682) );
  NAND2_X1 U12492 ( .A1(n10683), .A2(n10682), .ZN(n10684) );
  AND2_X1 U12493 ( .A1(n10700), .A2(n10684), .ZN(n12911) );
  NAND2_X1 U12494 ( .A1(n10879), .A2(n12911), .ZN(n10691) );
  INV_X1 U12495 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10685) );
  OR2_X1 U12496 ( .A1(n10519), .A2(n10685), .ZN(n10690) );
  INV_X1 U12497 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10686) );
  OR2_X1 U12498 ( .A1(n10551), .A2(n10686), .ZN(n10689) );
  INV_X1 U12499 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10687) );
  OR2_X1 U12500 ( .A1(n10553), .A2(n10687), .ZN(n10688) );
  NAND4_X1 U12501 ( .A1(n10691), .A2(n10690), .A3(n10689), .A4(n10688), .ZN(
        n14015) );
  NAND2_X1 U12502 ( .A1(n14015), .A2(n10938), .ZN(n10692) );
  XNOR2_X1 U12503 ( .A(n10693), .B(n10692), .ZN(n12909) );
  INV_X1 U12504 ( .A(n10692), .ZN(n10694) );
  INV_X1 U12505 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12430) );
  INV_X1 U12506 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12995) );
  OR2_X1 U12507 ( .A1(n10519), .A2(n12995), .ZN(n10697) );
  INV_X1 U12508 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10695) );
  OR2_X1 U12509 ( .A1(n10551), .A2(n10695), .ZN(n10696) );
  AND2_X1 U12510 ( .A1(n10697), .A2(n10696), .ZN(n10703) );
  INV_X1 U12511 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10699) );
  NAND2_X1 U12512 ( .A1(n10700), .A2(n10699), .ZN(n10701) );
  NAND2_X1 U12513 ( .A1(n10717), .A2(n10701), .ZN(n13930) );
  OR2_X1 U12514 ( .A1(n13930), .A2(n10943), .ZN(n10702) );
  OAI211_X1 U12515 ( .C1(n10553), .C2(n12430), .A(n10703), .B(n10702), .ZN(
        n14014) );
  AND2_X1 U12516 ( .A1(n14014), .A2(n10938), .ZN(n10713) );
  NAND2_X1 U12517 ( .A1(n11859), .A2(n13350), .ZN(n10711) );
  NAND3_X1 U12518 ( .A1(n10704), .A2(n10706), .A3(n10705), .ZN(n10707) );
  OAI21_X1 U12519 ( .B1(n10708), .B2(n10707), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n10709) );
  XNOR2_X1 U12520 ( .A(n10709), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15481) );
  AOI22_X1 U12521 ( .A1(n10741), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10740), 
        .B2(n15481), .ZN(n10710) );
  XNOR2_X1 U12522 ( .A(n14337), .B(n10835), .ZN(n10712) );
  NOR2_X1 U12523 ( .A1(n10712), .A2(n10713), .ZN(n10714) );
  AOI21_X1 U12524 ( .B1(n10713), .B2(n10712), .A(n10714), .ZN(n13928) );
  INV_X1 U12525 ( .A(n10714), .ZN(n10715) );
  INV_X1 U12526 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10716) );
  NAND2_X1 U12527 ( .A1(n10717), .A2(n10716), .ZN(n10718) );
  NAND2_X1 U12528 ( .A1(n10733), .A2(n10718), .ZN(n14233) );
  AOI22_X1 U12529 ( .A1(n13357), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n10552), 
        .B2(P2_REG2_REG_17__SCAN_IN), .ZN(n10720) );
  INV_X1 U12530 ( .A(n10553), .ZN(n10747) );
  NAND2_X1 U12531 ( .A1(n10747), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n10719) );
  OAI211_X1 U12532 ( .C1(n14233), .C2(n10943), .A(n10720), .B(n10719), .ZN(
        n14013) );
  AND2_X1 U12533 ( .A1(n14013), .A2(n10938), .ZN(n10725) );
  NAND2_X1 U12534 ( .A1(n11970), .A2(n13350), .ZN(n10723) );
  XNOR2_X1 U12535 ( .A(n10721), .B(P2_IR_REG_17__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U12536 ( .A1(n10741), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n10740), 
        .B2(n12720), .ZN(n10722) );
  XNOR2_X1 U12537 ( .A(n14332), .B(n10835), .ZN(n10724) );
  NOR2_X1 U12538 ( .A1(n10724), .A2(n10725), .ZN(n10726) );
  AOI21_X1 U12539 ( .B1(n10725), .B2(n10724), .A(n10726), .ZN(n13939) );
  NAND2_X1 U12540 ( .A1(n12384), .A2(n13350), .ZN(n10730) );
  NAND2_X1 U12541 ( .A1(n10721), .A2(n7402), .ZN(n10727) );
  NAND2_X1 U12542 ( .A1(n10727), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10728) );
  XNOR2_X1 U12543 ( .A(n10728), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U12544 ( .A1(n10741), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n10740), 
        .B2(n12728), .ZN(n10729) );
  NAND2_X2 U12545 ( .A1(n10730), .A2(n10729), .ZN(n14327) );
  XNOR2_X1 U12546 ( .A(n14327), .B(n10835), .ZN(n10738) );
  INV_X1 U12547 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10737) );
  INV_X1 U12548 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10732) );
  NAND2_X1 U12549 ( .A1(n10733), .A2(n10732), .ZN(n10734) );
  NAND2_X1 U12550 ( .A1(n10745), .A2(n10734), .ZN(n13982) );
  OR2_X1 U12551 ( .A1(n13982), .A2(n10943), .ZN(n10736) );
  AOI22_X1 U12552 ( .A1(n10747), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n13357), 
        .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n10735) );
  OAI211_X1 U12553 ( .C1(n10519), .C2(n10737), .A(n10736), .B(n10735), .ZN(
        n14012) );
  INV_X1 U12554 ( .A(n14012), .ZN(n14190) );
  NOR2_X1 U12555 ( .A1(n14190), .A2(n11781), .ZN(n10739) );
  XNOR2_X1 U12556 ( .A(n10738), .B(n10739), .ZN(n13979) );
  NAND2_X1 U12557 ( .A1(n12469), .A2(n13350), .ZN(n10743) );
  AOI22_X1 U12558 ( .A1(n10741), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10740), 
        .B2(n10458), .ZN(n10742) );
  XNOR2_X1 U12559 ( .A(n14317), .B(n10835), .ZN(n10755) );
  INV_X1 U12560 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10744) );
  NAND2_X1 U12561 ( .A1(n10745), .A2(n10744), .ZN(n10746) );
  AND2_X1 U12562 ( .A1(n10759), .A2(n10746), .ZN(n14203) );
  NAND2_X1 U12563 ( .A1(n14203), .A2(n10879), .ZN(n10753) );
  INV_X1 U12564 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U12565 ( .A1(n10747), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n10749) );
  NAND2_X1 U12566 ( .A1(n13357), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n10748) );
  OAI211_X1 U12567 ( .C1(n10519), .C2(n10750), .A(n10749), .B(n10748), .ZN(
        n10751) );
  INV_X1 U12568 ( .A(n10751), .ZN(n10752) );
  NAND2_X1 U12569 ( .A1(n10753), .A2(n10752), .ZN(n14011) );
  NAND2_X1 U12570 ( .A1(n14011), .A2(n10938), .ZN(n10754) );
  XNOR2_X1 U12571 ( .A(n10755), .B(n10754), .ZN(n13903) );
  INV_X1 U12572 ( .A(n10754), .ZN(n10756) );
  INV_X1 U12573 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10758) );
  NAND2_X1 U12574 ( .A1(n10759), .A2(n10758), .ZN(n10760) );
  NAND2_X1 U12575 ( .A1(n10775), .A2(n10760), .ZN(n13963) );
  OR2_X1 U12576 ( .A1(n13963), .A2(n10943), .ZN(n10766) );
  INV_X1 U12577 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U12578 ( .A1(n13357), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n10762) );
  NAND2_X1 U12579 ( .A1(n10552), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n10761) );
  OAI211_X1 U12580 ( .C1(n10553), .C2(n10763), .A(n10762), .B(n10761), .ZN(
        n10764) );
  INV_X1 U12581 ( .A(n10764), .ZN(n10765) );
  NAND2_X1 U12582 ( .A1(n10766), .A2(n10765), .ZN(n14010) );
  AND2_X1 U12583 ( .A1(n14010), .A2(n10938), .ZN(n10770) );
  NAND2_X1 U12584 ( .A1(n12388), .A2(n13350), .ZN(n10768) );
  NAND2_X1 U12585 ( .A1(n10741), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n10767) );
  XNOR2_X1 U12586 ( .A(n14314), .B(n10835), .ZN(n10769) );
  NOR2_X1 U12587 ( .A1(n10769), .A2(n10770), .ZN(n10771) );
  AOI21_X1 U12588 ( .B1(n10770), .B2(n10769), .A(n10771), .ZN(n13959) );
  INV_X1 U12589 ( .A(n10771), .ZN(n10772) );
  INV_X1 U12590 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U12591 ( .A1(n10775), .A2(n10774), .ZN(n10776) );
  NAND2_X1 U12592 ( .A1(n10810), .A2(n10776), .ZN(n13914) );
  OR2_X1 U12593 ( .A1(n13914), .A2(n10943), .ZN(n10782) );
  INV_X1 U12594 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10779) );
  NAND2_X1 U12595 ( .A1(n10552), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n10778) );
  NAND2_X1 U12596 ( .A1(n13357), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n10777) );
  OAI211_X1 U12597 ( .C1(n10779), .C2(n10553), .A(n10778), .B(n10777), .ZN(
        n10780) );
  INV_X1 U12598 ( .A(n10780), .ZN(n10781) );
  NAND2_X1 U12599 ( .A1(n10782), .A2(n10781), .ZN(n14009) );
  NAND2_X1 U12600 ( .A1(n14009), .A2(n10938), .ZN(n10786) );
  NAND2_X1 U12601 ( .A1(n12478), .A2(n13350), .ZN(n10784) );
  NAND2_X1 U12602 ( .A1(n10741), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n10783) );
  XNOR2_X1 U12603 ( .A(n14309), .B(n10835), .ZN(n10785) );
  XOR2_X1 U12604 ( .A(n10786), .B(n10785), .Z(n13911) );
  INV_X1 U12605 ( .A(n10785), .ZN(n10787) );
  INV_X1 U12606 ( .A(n10788), .ZN(n10791) );
  INV_X1 U12607 ( .A(n10789), .ZN(n10790) );
  NAND2_X1 U12608 ( .A1(n10791), .A2(n10790), .ZN(n10792) );
  NAND2_X1 U12609 ( .A1(n10793), .A2(n10792), .ZN(n12623) );
  NAND2_X1 U12610 ( .A1(n10741), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n10794) );
  XNOR2_X1 U12611 ( .A(n14301), .B(n10835), .ZN(n10803) );
  XNOR2_X1 U12612 ( .A(n10810), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n14155) );
  NAND2_X1 U12613 ( .A1(n14155), .A2(n10879), .ZN(n10802) );
  INV_X1 U12614 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U12615 ( .A1(n13357), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n10798) );
  NAND2_X1 U12616 ( .A1(n10552), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n10797) );
  OAI211_X1 U12617 ( .C1(n10799), .C2(n10553), .A(n10798), .B(n10797), .ZN(
        n10800) );
  INV_X1 U12618 ( .A(n10800), .ZN(n10801) );
  NAND2_X1 U12619 ( .A1(n10802), .A2(n10801), .ZN(n14008) );
  AND2_X1 U12620 ( .A1(n14008), .A2(n10938), .ZN(n13969) );
  NAND2_X1 U12621 ( .A1(n12731), .A2(n13350), .ZN(n10807) );
  NAND2_X1 U12622 ( .A1(n10741), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n10806) );
  XNOR2_X1 U12623 ( .A(n14295), .B(n10835), .ZN(n10820) );
  XNOR2_X1 U12624 ( .A(n10819), .B(n10820), .ZN(n13898) );
  INV_X1 U12625 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10809) );
  INV_X1 U12626 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10808) );
  OAI21_X1 U12627 ( .B1(n10810), .B2(n10809), .A(n10808), .ZN(n10811) );
  AND2_X1 U12628 ( .A1(n10811), .A2(n10825), .ZN(n14136) );
  NAND2_X1 U12629 ( .A1(n14136), .A2(n10879), .ZN(n10817) );
  INV_X1 U12630 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U12631 ( .A1(n10552), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n10813) );
  NAND2_X1 U12632 ( .A1(n13357), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n10812) );
  OAI211_X1 U12633 ( .C1(n10814), .C2(n10553), .A(n10813), .B(n10812), .ZN(
        n10815) );
  INV_X1 U12634 ( .A(n10815), .ZN(n10816) );
  NAND2_X1 U12635 ( .A1(n10817), .A2(n10816), .ZN(n14007) );
  OR2_X1 U12636 ( .A1(n14145), .A2(n11781), .ZN(n10818) );
  NAND2_X1 U12637 ( .A1(n13898), .A2(n10818), .ZN(n13902) );
  INV_X1 U12638 ( .A(n10820), .ZN(n10821) );
  INV_X1 U12639 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10824) );
  NAND2_X1 U12640 ( .A1(n10825), .A2(n10824), .ZN(n10826) );
  NAND2_X1 U12641 ( .A1(n10860), .A2(n10826), .ZN(n13952) );
  OR2_X1 U12642 ( .A1(n13952), .A2(n10943), .ZN(n10832) );
  INV_X1 U12643 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10829) );
  NAND2_X1 U12644 ( .A1(n13357), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n10828) );
  NAND2_X1 U12645 ( .A1(n10552), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n10827) );
  OAI211_X1 U12646 ( .C1(n10553), .C2(n10829), .A(n10828), .B(n10827), .ZN(
        n10830) );
  INV_X1 U12647 ( .A(n10830), .ZN(n10831) );
  NAND2_X1 U12648 ( .A1(n10832), .A2(n10831), .ZN(n14006) );
  NAND2_X1 U12649 ( .A1(n14006), .A2(n10938), .ZN(n10838) );
  NAND2_X1 U12650 ( .A1(n12607), .A2(n13350), .ZN(n10834) );
  NAND2_X1 U12651 ( .A1(n10741), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n10833) );
  XNOR2_X1 U12652 ( .A(n14290), .B(n10835), .ZN(n10837) );
  XOR2_X1 U12653 ( .A(n10838), .B(n10837), .Z(n13948) );
  INV_X1 U12654 ( .A(n10838), .ZN(n10839) );
  NAND2_X1 U12655 ( .A1(n12648), .A2(n13350), .ZN(n10842) );
  NAND2_X1 U12656 ( .A1(n10741), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10841) );
  XNOR2_X1 U12657 ( .A(n14108), .B(n10835), .ZN(n10849) );
  XNOR2_X1 U12658 ( .A(n10860), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14105) );
  NAND2_X1 U12659 ( .A1(n14105), .A2(n10879), .ZN(n10848) );
  INV_X1 U12660 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10845) );
  NAND2_X1 U12661 ( .A1(n10552), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n10844) );
  NAND2_X1 U12662 ( .A1(n13357), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n10843) );
  OAI211_X1 U12663 ( .C1(n10845), .C2(n10553), .A(n10844), .B(n10843), .ZN(
        n10846) );
  INV_X1 U12664 ( .A(n10846), .ZN(n10847) );
  NOR2_X1 U12665 ( .A1(n14118), .A2(n11781), .ZN(n10850) );
  INV_X1 U12666 ( .A(n10849), .ZN(n10851) );
  NAND2_X1 U12667 ( .A1(n10851), .A2(n10850), .ZN(n10852) );
  OR2_X1 U12668 ( .A1(n12806), .A2(n7191), .ZN(n10856) );
  NAND2_X1 U12669 ( .A1(n10741), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n10855) );
  XNOR2_X1 U12670 ( .A(n14278), .B(n10857), .ZN(n10871) );
  INV_X1 U12671 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10859) );
  INV_X1 U12672 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10858) );
  OAI21_X1 U12673 ( .B1(n10860), .B2(n10859), .A(n10858), .ZN(n10863) );
  INV_X1 U12674 ( .A(n10860), .ZN(n10862) );
  AND2_X1 U12675 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n10861) );
  INV_X1 U12676 ( .A(n10875), .ZN(n10877) );
  NAND2_X1 U12677 ( .A1(n10863), .A2(n10877), .ZN(n13993) );
  OR2_X1 U12678 ( .A1(n13993), .A2(n10943), .ZN(n10869) );
  INV_X1 U12679 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10866) );
  NAND2_X1 U12680 ( .A1(n10552), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n10865) );
  NAND2_X1 U12681 ( .A1(n13357), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n10864) );
  OAI211_X1 U12682 ( .C1(n10866), .C2(n10553), .A(n10865), .B(n10864), .ZN(
        n10867) );
  INV_X1 U12683 ( .A(n10867), .ZN(n10868) );
  NAND2_X1 U12684 ( .A1(n14005), .A2(n10938), .ZN(n10870) );
  NAND2_X1 U12685 ( .A1(n10871), .A2(n10870), .ZN(n10872) );
  OAI21_X1 U12686 ( .B1(n10871), .B2(n10870), .A(n10872), .ZN(n13991) );
  NAND2_X1 U12687 ( .A1(n13007), .A2(n13350), .ZN(n10874) );
  NAND2_X1 U12688 ( .A1(n10741), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n10873) );
  XNOR2_X1 U12689 ( .A(n14271), .B(n10835), .ZN(n10886) );
  INV_X1 U12690 ( .A(n10892), .ZN(n10894) );
  INV_X1 U12691 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U12692 ( .A1(n10877), .A2(n10876), .ZN(n10878) );
  NAND2_X1 U12693 ( .A1(n13887), .A2(n10879), .ZN(n10885) );
  INV_X1 U12694 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U12695 ( .A1(n10552), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n10881) );
  NAND2_X1 U12696 ( .A1(n13357), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n10880) );
  OAI211_X1 U12697 ( .C1(n10882), .C2(n10553), .A(n10881), .B(n10880), .ZN(
        n10883) );
  INV_X1 U12698 ( .A(n10883), .ZN(n10884) );
  NOR2_X1 U12699 ( .A1(n14044), .A2(n11781), .ZN(n10887) );
  XNOR2_X1 U12700 ( .A(n10886), .B(n10887), .ZN(n13886) );
  INV_X1 U12701 ( .A(n10886), .ZN(n10889) );
  INV_X1 U12702 ( .A(n10887), .ZN(n10888) );
  NAND2_X1 U12703 ( .A1(n14374), .A2(n13350), .ZN(n10891) );
  NAND2_X1 U12704 ( .A1(n10741), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10890) );
  NAND2_X1 U12705 ( .A1(n10892), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n14059) );
  INV_X1 U12706 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U12707 ( .A1(n10894), .A2(n10893), .ZN(n10895) );
  NAND2_X1 U12708 ( .A1(n14059), .A2(n10895), .ZN(n10955) );
  INV_X1 U12709 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U12710 ( .A1(n13357), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n10897) );
  NAND2_X1 U12711 ( .A1(n10552), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n10896) );
  OAI211_X1 U12712 ( .C1(n10898), .C2(n10553), .A(n10897), .B(n10896), .ZN(
        n10899) );
  INV_X1 U12713 ( .A(n10899), .ZN(n10900) );
  NAND2_X1 U12714 ( .A1(n10901), .A2(n10900), .ZN(n14054) );
  NAND2_X1 U12715 ( .A1(n14267), .A2(n13889), .ZN(n10902) );
  XNOR2_X1 U12716 ( .A(n10937), .B(n14072), .ZN(n10966) );
  NOR4_X1 U12717 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n10906) );
  NOR4_X1 U12718 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n10905) );
  NOR4_X1 U12719 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n10904) );
  NOR4_X1 U12720 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10903) );
  NAND4_X1 U12721 ( .A1(n10906), .A2(n10905), .A3(n10904), .A4(n10903), .ZN(
        n10924) );
  NOR2_X1 U12722 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n10910) );
  NOR4_X1 U12723 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10909) );
  NOR4_X1 U12724 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n10908) );
  NOR4_X1 U12725 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n10907) );
  NAND4_X1 U12726 ( .A1(n10910), .A2(n10909), .A3(n10908), .A4(n10907), .ZN(
        n10923) );
  NAND2_X1 U12727 ( .A1(n10920), .A2(n10919), .ZN(n10913) );
  OR2_X1 U12728 ( .A1(n10916), .A2(n10915), .ZN(n10917) );
  NAND2_X1 U12729 ( .A1(n10918), .A2(n10917), .ZN(n12683) );
  XNOR2_X1 U12730 ( .A(P2_B_REG_SCAN_IN), .B(n12628), .ZN(n10921) );
  NAND2_X1 U12731 ( .A1(n12683), .A2(n10921), .ZN(n10922) );
  OAI21_X1 U12732 ( .B1(n10924), .B2(n10923), .A(n15403), .ZN(n11476) );
  NOR2_X1 U12733 ( .A1(n12683), .A2(n12628), .ZN(n10925) );
  NAND2_X1 U12734 ( .A1(n12802), .A2(n10925), .ZN(n10968) );
  NAND2_X1 U12735 ( .A1(n10911), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10927) );
  INV_X1 U12736 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15402) );
  NAND2_X1 U12737 ( .A1(n15403), .A2(n15402), .ZN(n10930) );
  INV_X1 U12738 ( .A(n12683), .ZN(n10928) );
  OR2_X1 U12739 ( .A1(n12802), .A2(n10928), .ZN(n10929) );
  AND2_X1 U12740 ( .A1(n15409), .A2(n11471), .ZN(n10931) );
  NAND2_X1 U12741 ( .A1(n11476), .A2(n10931), .ZN(n11695) );
  INV_X1 U12742 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15407) );
  NAND2_X1 U12743 ( .A1(n15403), .A2(n15407), .ZN(n10934) );
  INV_X1 U12744 ( .A(n12628), .ZN(n10932) );
  OR2_X1 U12745 ( .A1(n12802), .A2(n10932), .ZN(n10933) );
  INV_X1 U12746 ( .A(n11465), .ZN(n10935) );
  NAND2_X1 U12747 ( .A1(n13356), .A2(n13452), .ZN(n13443) );
  AND2_X1 U12748 ( .A1(n10935), .A2(n16182), .ZN(n10936) );
  INV_X2 U12749 ( .A(n13940), .ZN(n14001) );
  XNOR2_X1 U12750 ( .A(n10937), .B(n7758), .ZN(n10940) );
  NOR2_X1 U12751 ( .A1(n14001), .A2(n10938), .ZN(n10939) );
  NAND2_X1 U12752 ( .A1(n10940), .A2(n10939), .ZN(n10965) );
  NOR2_X1 U12753 ( .A1(n15896), .A2(n13399), .ZN(n11699) );
  NAND2_X1 U12754 ( .A1(n10954), .A2(n11699), .ZN(n10942) );
  OR2_X1 U12755 ( .A1(n14059), .A2(n10943), .ZN(n10949) );
  INV_X1 U12756 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10946) );
  NAND2_X1 U12757 ( .A1(n13357), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U12758 ( .A1(n10552), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n10944) );
  OAI211_X1 U12759 ( .C1(n7192), .C2(n10946), .A(n10945), .B(n10944), .ZN(
        n10947) );
  INV_X1 U12760 ( .A(n10947), .ZN(n10948) );
  NAND2_X1 U12761 ( .A1(n10949), .A2(n10948), .ZN(n14004) );
  NAND2_X1 U12762 ( .A1(n14004), .A2(n14091), .ZN(n10953) );
  INV_X1 U12763 ( .A(n10950), .ZN(n10951) );
  NAND2_X1 U12764 ( .A1(n14092), .A2(n14089), .ZN(n10952) );
  AND2_X1 U12765 ( .A1(n10953), .A2(n10952), .ZN(n14067) );
  INV_X1 U12766 ( .A(n13356), .ZN(n11464) );
  NAND2_X1 U12767 ( .A1(n10954), .A2(n11464), .ZN(n13984) );
  INV_X1 U12768 ( .A(n10955), .ZN(n14076) );
  NAND2_X1 U12769 ( .A1(n11471), .A2(n11476), .ZN(n10957) );
  INV_X1 U12770 ( .A(n11474), .ZN(n10956) );
  OAI21_X1 U12771 ( .B1(n15408), .B2(n10957), .A(n10956), .ZN(n10958) );
  NAND2_X1 U12772 ( .A1(n11465), .A2(n13356), .ZN(n11696) );
  NAND2_X1 U12773 ( .A1(n10958), .A2(n11696), .ZN(n10974) );
  INV_X1 U12774 ( .A(n10959), .ZN(n10960) );
  AOI22_X1 U12775 ( .A1(n14076), .A2(n13994), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10962) );
  OAI21_X1 U12776 ( .B1(n14067), .B2(n13984), .A(n10962), .ZN(n10963) );
  AOI21_X1 U12777 ( .B1(n14267), .B2(n13999), .A(n10963), .ZN(n10964) );
  OAI211_X1 U12778 ( .C1(n10966), .C2(n13897), .A(n10965), .B(n10964), .ZN(
        P2_U3192) );
  INV_X1 U12779 ( .A(n12734), .ZN(n10967) );
  NOR2_X1 U12780 ( .A1(n11844), .A2(P1_U3086), .ZN(n10969) );
  INV_X1 U12781 ( .A(n13897), .ZN(n13968) );
  AOI22_X1 U12782 ( .A1(n13968), .A2(n13144), .B1(n13940), .B2(n10540), .ZN(
        n10973) );
  INV_X1 U12783 ( .A(n10970), .ZN(n10972) );
  NOR3_X1 U12784 ( .A1(n10973), .A2(n10972), .A3(n10971), .ZN(n10978) );
  INV_X1 U12785 ( .A(n14026), .ZN(n11680) );
  OAI22_X1 U12786 ( .A1(n11680), .A2(n13996), .B1(n13992), .B2(n12036), .ZN(
        n10977) );
  INV_X1 U12787 ( .A(n14248), .ZN(n11673) );
  INV_X1 U12788 ( .A(n15409), .ZN(n15406) );
  NOR2_X1 U12789 ( .A1(n10974), .A2(n15406), .ZN(n11367) );
  OAI22_X1 U12790 ( .A1(n13978), .A2(n11673), .B1(n11367), .B2(n14245), .ZN(
        n10975) );
  OR4_X1 U12791 ( .A1(n10978), .A2(n10977), .A3(n10976), .A4(n10975), .ZN(
        P2_U3209) );
  NOR2_X1 U12792 ( .A1(n11059), .A2(P2_U3088), .ZN(n15417) );
  AOI21_X1 U12793 ( .B1(n14376), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n15417), 
        .ZN(n10979) );
  OAI21_X1 U12794 ( .B1(n11020), .B2(n14378), .A(n10979), .ZN(P2_U3326) );
  OAI222_X1 U12795 ( .A1(n14370), .A2(n10980), .B1(n14378), .B2(n11022), .C1(
        n15429), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U12796 ( .A(n15444), .ZN(n11064) );
  INV_X1 U12797 ( .A(n10981), .ZN(n11024) );
  OAI222_X1 U12798 ( .A1(P2_U3088), .A2(n11064), .B1(n14378), .B2(n11024), 
        .C1(n10982), .C2(n14370), .ZN(P2_U3323) );
  INV_X1 U12799 ( .A(n11066), .ZN(n11103) );
  OAI222_X1 U12800 ( .A1(n14370), .A2(n10983), .B1(n14378), .B2(n10984), .C1(
        n11103), .C2(P2_U3088), .ZN(P2_U3322) );
  AND2_X1 U12801 ( .A1(n8421), .A2(P1_U3086), .ZN(n15394) );
  INV_X2 U12802 ( .A(n15394), .ZN(n15160) );
  INV_X1 U12803 ( .A(n11263), .ZN(n11272) );
  OAI222_X1 U12804 ( .A1(n15157), .A2(n10985), .B1(n15160), .B2(n10984), .C1(
        P1_U3086), .C2(n11272), .ZN(P1_U3350) );
  NOR2_X1 U12805 ( .A1(n10986), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13876) );
  INV_X2 U12806 ( .A(n13876), .ZN(n13131) );
  OAI222_X1 U12807 ( .A1(n15683), .A2(P3_U3151), .B1(n13131), .B2(n10988), 
        .C1(n10987), .C2(n13880), .ZN(P3_U3289) );
  INV_X1 U12808 ( .A(n11062), .ZN(n11127) );
  OAI222_X1 U12809 ( .A1(n14370), .A2(n10989), .B1(n14378), .B2(n7378), .C1(
        n11127), .C2(P2_U3088), .ZN(P2_U3324) );
  AND2_X1 U12810 ( .A1(n10991), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12811 ( .A1(n10991), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12812 ( .A1(n10991), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12813 ( .A1(n10991), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12814 ( .A1(n10991), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12815 ( .A1(n10991), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12816 ( .A1(n10991), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12817 ( .A1(n10991), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12818 ( .A1(n10991), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12819 ( .A1(n10991), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12820 ( .A1(n10991), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12821 ( .A1(n10991), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12822 ( .A1(n10991), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12823 ( .A1(n10991), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12824 ( .A1(n10991), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12825 ( .A1(n10991), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12826 ( .A1(n10991), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12827 ( .A1(n10991), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12828 ( .A1(n10991), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12829 ( .A1(n10991), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12830 ( .A1(n10991), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12831 ( .A1(n10991), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12832 ( .A1(n10991), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12833 ( .A1(n10991), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12834 ( .A1(n10991), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12835 ( .A1(n10991), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12836 ( .A1(n10991), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12837 ( .A1(n10991), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12838 ( .A1(n10991), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12839 ( .A1(n10991), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  OAI222_X1 U12840 ( .A1(n13131), .A2(n10992), .B1(n15721), .B2(P3_U3151), 
        .C1(n13880), .C2(n15313), .ZN(P3_U3284) );
  INV_X1 U12841 ( .A(n11067), .ZN(n11115) );
  OAI222_X1 U12842 ( .A1(P2_U3088), .A2(n11115), .B1(n14378), .B2(n10995), 
        .C1(n10993), .C2(n14370), .ZN(P2_U3321) );
  INV_X1 U12843 ( .A(n11211), .ZN(n11171) );
  OAI222_X1 U12844 ( .A1(P1_U3086), .A2(n11171), .B1(n15160), .B2(n10995), 
        .C1(n10994), .C2(n15157), .ZN(P1_U3349) );
  INV_X1 U12845 ( .A(n10996), .ZN(n10997) );
  INV_X1 U12846 ( .A(SI_3_), .ZN(n15331) );
  OAI222_X1 U12847 ( .A1(n13131), .A2(n10997), .B1(n13880), .B2(n15331), .C1(
        n15630), .C2(P3_U3151), .ZN(P3_U3292) );
  INV_X1 U12848 ( .A(n10998), .ZN(n11000) );
  INV_X1 U12849 ( .A(SI_4_), .ZN(n15323) );
  OAI222_X1 U12850 ( .A1(n13131), .A2(n11000), .B1(n13880), .B2(n15323), .C1(
        n10999), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12851 ( .A(n11001), .ZN(n11003) );
  INV_X1 U12852 ( .A(SI_5_), .ZN(n15325) );
  OAI222_X1 U12853 ( .A1(n13131), .A2(n11003), .B1(n13880), .B2(n15325), .C1(
        n11002), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12854 ( .A(n11004), .ZN(n11005) );
  OAI222_X1 U12855 ( .A1(n13131), .A2(n11005), .B1(n13880), .B2(n8682), .C1(
        n12058), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12856 ( .A1(n13131), .A2(n11006), .B1(n13880), .B2(n15320), .C1(
        n11760), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U12857 ( .A(n11007), .ZN(n11009) );
  OAI222_X1 U12858 ( .A1(n13131), .A2(n11009), .B1(n13880), .B2(n7377), .C1(
        n11008), .C2(P3_U3151), .ZN(P3_U3293) );
  INV_X1 U12859 ( .A(SI_10_), .ZN(n15170) );
  OAI222_X1 U12860 ( .A1(n13131), .A2(n11011), .B1(n13880), .B2(n15170), .C1(
        n11010), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12861 ( .A(n11012), .ZN(n11013) );
  INV_X1 U12862 ( .A(SI_7_), .ZN(n15322) );
  OAI222_X1 U12863 ( .A1(n13131), .A2(n11013), .B1(n13880), .B2(n15322), .C1(
        n11620), .C2(P3_U3151), .ZN(P3_U3288) );
  OAI222_X1 U12864 ( .A1(n13131), .A2(n11014), .B1(n15737), .B2(P3_U3151), 
        .C1(n13880), .C2(n15307), .ZN(P3_U3283) );
  OAI222_X1 U12865 ( .A1(n11016), .A2(P3_U3151), .B1(n13131), .B2(n11015), 
        .C1(n15267), .C2(n13880), .ZN(P3_U3295) );
  INV_X1 U12866 ( .A(n11069), .ZN(n11185) );
  OAI222_X1 U12867 ( .A1(n14370), .A2(n11017), .B1(n14378), .B2(n11019), .C1(
        n11185), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U12868 ( .A(n11295), .ZN(n11220) );
  OAI222_X1 U12869 ( .A1(P1_U3086), .A2(n11220), .B1(n15160), .B2(n11019), 
        .C1(n11018), .C2(n15157), .ZN(P1_U3348) );
  OAI222_X1 U12870 ( .A1(n15157), .A2(n7665), .B1(n15160), .B2(n11020), .C1(
        P1_U3086), .C2(n11147), .ZN(P1_U3354) );
  OAI222_X1 U12871 ( .A1(P1_U3086), .A2(n11150), .B1(n15160), .B2(n11022), 
        .C1(n11021), .C2(n15157), .ZN(P1_U3353) );
  OAI222_X1 U12872 ( .A1(P1_U3086), .A2(n15863), .B1(n15160), .B2(n11024), 
        .C1(n11023), .C2(n15157), .ZN(P1_U3351) );
  INV_X1 U12873 ( .A(n11070), .ZN(n11083) );
  OAI222_X1 U12874 ( .A1(P2_U3088), .A2(n11083), .B1(n14378), .B2(n10483), 
        .C1(n11025), .C2(n14370), .ZN(P2_U3319) );
  OAI222_X1 U12875 ( .A1(n15157), .A2(n11026), .B1(n15160), .B2(n10483), .C1(
        P1_U3086), .C2(n11321), .ZN(P1_U3347) );
  NAND2_X2 U12876 ( .A1(n11557), .A2(n11027), .ZN(n15400) );
  NAND2_X1 U12877 ( .A1(n15400), .A2(P1_D_REG_0__SCAN_IN), .ZN(n11028) );
  OAI21_X1 U12878 ( .B1(n15400), .B2(n11029), .A(n11028), .ZN(P1_U3445) );
  OAI222_X1 U12879 ( .A1(n13131), .A2(n11031), .B1(n13880), .B2(n15304), .C1(
        n11030), .C2(P3_U3151), .ZN(P3_U3282) );
  AOI21_X1 U12880 ( .B1(n11033), .B2(n11845), .A(n11032), .ZN(n11138) );
  INV_X1 U12881 ( .A(n11138), .ZN(n11035) );
  INV_X1 U12882 ( .A(n11034), .ZN(n12732) );
  AND2_X1 U12883 ( .A1(n11035), .A2(n11137), .ZN(n15526) );
  NOR2_X1 U12884 ( .A1(n15526), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U12885 ( .A1(n13131), .A2(n11038), .B1(n13880), .B2(n11037), .C1(
        n11036), .C2(P3_U3151), .ZN(P3_U3281) );
  OAI222_X1 U12886 ( .A1(n14370), .A2(n11039), .B1(n14378), .B2(n11041), .C1(
        n11201), .C2(P2_U3088), .ZN(P2_U3318) );
  INV_X1 U12887 ( .A(n11334), .ZN(n11306) );
  OAI222_X1 U12888 ( .A1(P1_U3086), .A2(n11306), .B1(n15160), .B2(n11041), 
        .C1(n11040), .C2(n15157), .ZN(P1_U3346) );
  OAI222_X1 U12889 ( .A1(P2_U3088), .A2(n11277), .B1(n14378), .B2(n11043), 
        .C1(n11042), .C2(n14370), .ZN(P2_U3317) );
  INV_X1 U12890 ( .A(n11528), .ZN(n11344) );
  OAI222_X1 U12891 ( .A1(n15157), .A2(n11044), .B1(n15160), .B2(n11043), .C1(
        P1_U3086), .C2(n11344), .ZN(P1_U3345) );
  OAI222_X1 U12892 ( .A1(n13131), .A2(n11045), .B1(n15789), .B2(P3_U3151), 
        .C1(n15305), .C2(n13880), .ZN(P3_U3280) );
  MUX2_X1 U12893 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n12174), .S(n11201), .Z(
        n11053) );
  INV_X1 U12894 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11050) );
  INV_X1 U12895 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11049) );
  INV_X1 U12896 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11048) );
  INV_X1 U12897 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11047) );
  INV_X1 U12898 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11711) );
  MUX2_X1 U12899 ( .A(n11711), .B(P2_REG2_REG_1__SCAN_IN), .S(n11059), .Z(
        n15410) );
  AND2_X1 U12900 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n11046) );
  NAND2_X1 U12901 ( .A1(n15410), .A2(n11046), .ZN(n15411) );
  OAI21_X1 U12902 ( .B1(n11059), .B2(n11711), .A(n15411), .ZN(n15426) );
  XNOR2_X1 U12903 ( .A(n15429), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n15427) );
  NAND2_X1 U12904 ( .A1(n15426), .A2(n15427), .ZN(n15425) );
  OAI21_X1 U12905 ( .B1(n11047), .B2(n15429), .A(n15425), .ZN(n11123) );
  MUX2_X1 U12906 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11048), .S(n11062), .Z(
        n11124) );
  NAND2_X1 U12907 ( .A1(n11123), .A2(n11124), .ZN(n11122) );
  OAI21_X1 U12908 ( .B1(n11048), .B2(n11127), .A(n11122), .ZN(n15438) );
  XNOR2_X1 U12909 ( .A(n11064), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n15439) );
  NAND2_X1 U12910 ( .A1(n15438), .A2(n15439), .ZN(n15437) );
  OAI21_X1 U12911 ( .B1(n11064), .B2(n11049), .A(n15437), .ZN(n11099) );
  MUX2_X1 U12912 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11050), .S(n11066), .Z(
        n11100) );
  NAND2_X1 U12913 ( .A1(n11099), .A2(n11100), .ZN(n11098) );
  OAI21_X1 U12914 ( .B1(n11050), .B2(n11103), .A(n11098), .ZN(n11111) );
  XNOR2_X1 U12915 ( .A(n11115), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n11112) );
  NAND2_X1 U12916 ( .A1(n11111), .A2(n11112), .ZN(n11110) );
  OAI21_X1 U12917 ( .B1(n16040), .B2(n11115), .A(n11110), .ZN(n11181) );
  MUX2_X1 U12918 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11051), .S(n11069), .Z(
        n11182) );
  NAND2_X1 U12919 ( .A1(n11181), .A2(n11182), .ZN(n11180) );
  OAI21_X1 U12920 ( .B1(n11185), .B2(n11051), .A(n11180), .ZN(n11086) );
  XNOR2_X1 U12921 ( .A(n11070), .B(n12084), .ZN(n11087) );
  NAND2_X1 U12922 ( .A1(n11086), .A2(n11087), .ZN(n11085) );
  OAI21_X1 U12923 ( .B1(n11083), .B2(n12084), .A(n11085), .ZN(n11052) );
  NOR2_X1 U12924 ( .A1(n11052), .A2(n11053), .ZN(n11200) );
  AOI21_X1 U12925 ( .B1(n11053), .B2(n11052), .A(n11200), .ZN(n11079) );
  NAND2_X1 U12926 ( .A1(n11465), .A2(n12734), .ZN(n11055) );
  NAND2_X1 U12927 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  NAND2_X1 U12928 ( .A1(n11057), .A2(n11056), .ZN(n11074) );
  NOR2_X1 U12929 ( .A1(n10950), .A2(P2_U3088), .ZN(n14375) );
  INV_X1 U12930 ( .A(n13455), .ZN(n14029) );
  AND2_X1 U12931 ( .A1(n11073), .A2(n14029), .ZN(n15512) );
  MUX2_X1 U12932 ( .A(n11058), .B(P2_REG1_REG_1__SCAN_IN), .S(n11059), .Z(
        n15420) );
  NAND3_X1 U12933 ( .A1(n15420), .A2(P2_REG1_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n15419) );
  OAI21_X1 U12934 ( .B1(n11058), .B2(n11059), .A(n15419), .ZN(n15433) );
  MUX2_X1 U12935 ( .A(n11060), .B(P2_REG1_REG_2__SCAN_IN), .S(n15429), .Z(
        n15432) );
  NAND2_X1 U12936 ( .A1(n15433), .A2(n15432), .ZN(n15431) );
  INV_X1 U12937 ( .A(n15429), .ZN(n11061) );
  NAND2_X1 U12938 ( .A1(n11061), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n11117) );
  MUX2_X1 U12939 ( .A(n10513), .B(P2_REG1_REG_3__SCAN_IN), .S(n11062), .Z(
        n11118) );
  AOI21_X1 U12940 ( .B1(n15431), .B2(n11117), .A(n11118), .ZN(n11120) );
  AOI21_X1 U12941 ( .B1(n11062), .B2(P2_REG1_REG_3__SCAN_IN), .A(n11120), .ZN(
        n15447) );
  MUX2_X1 U12942 ( .A(n11063), .B(P2_REG1_REG_4__SCAN_IN), .S(n15444), .Z(
        n15446) );
  NOR2_X1 U12943 ( .A1(n15447), .A2(n15446), .ZN(n15445) );
  NOR2_X1 U12944 ( .A1(n11064), .A2(n11063), .ZN(n11093) );
  MUX2_X1 U12945 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n11065), .S(n11066), .Z(
        n11092) );
  OAI21_X1 U12946 ( .B1(n15445), .B2(n11093), .A(n11092), .ZN(n11106) );
  NAND2_X1 U12947 ( .A1(n11066), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11105) );
  MUX2_X1 U12948 ( .A(n10591), .B(P2_REG1_REG_6__SCAN_IN), .S(n11067), .Z(
        n11104) );
  AOI21_X1 U12949 ( .B1(n11106), .B2(n11105), .A(n11104), .ZN(n11175) );
  NOR2_X1 U12950 ( .A1(n11115), .A2(n10591), .ZN(n11174) );
  MUX2_X1 U12951 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n11068), .S(n11069), .Z(
        n11173) );
  OAI21_X1 U12952 ( .B1(n11175), .B2(n11174), .A(n11173), .ZN(n11172) );
  NAND2_X1 U12953 ( .A1(n11069), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11081) );
  MUX2_X1 U12954 ( .A(n10493), .B(P2_REG1_REG_8__SCAN_IN), .S(n11070), .Z(
        n11080) );
  AOI21_X1 U12955 ( .B1(n11172), .B2(n11081), .A(n11080), .ZN(n11091) );
  AOI21_X1 U12956 ( .B1(n11070), .B2(P2_REG1_REG_8__SCAN_IN), .A(n11091), .ZN(
        n11072) );
  MUX2_X1 U12957 ( .A(n10478), .B(P2_REG1_REG_9__SCAN_IN), .S(n11201), .Z(
        n11071) );
  NAND2_X1 U12958 ( .A1(n11072), .A2(n11071), .ZN(n11191) );
  OAI21_X1 U12959 ( .B1(n11072), .B2(n11071), .A(n11191), .ZN(n11077) );
  AND2_X1 U12960 ( .A1(n11074), .A2(n10950), .ZN(n15452) );
  OR2_X1 U12961 ( .A1(n11074), .A2(P2_U3088), .ZN(n15441) );
  INV_X1 U12962 ( .A(n15441), .ZN(n15502) );
  AND2_X1 U12963 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n11975) );
  AOI21_X1 U12964 ( .B1(n15502), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n11975), .ZN(
        n11075) );
  OAI21_X1 U12965 ( .B1(n15468), .B2(n11201), .A(n11075), .ZN(n11076) );
  AOI21_X1 U12966 ( .B1(n11077), .B2(n15494), .A(n11076), .ZN(n11078) );
  OAI21_X1 U12967 ( .B1(n11079), .B2(n15412), .A(n11078), .ZN(P2_U3223) );
  NAND3_X1 U12968 ( .A1(n11172), .A2(n11081), .A3(n11080), .ZN(n11082) );
  NAND2_X1 U12969 ( .A1(n11082), .A2(n15494), .ZN(n11090) );
  AND2_X1 U12970 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11869) );
  NOR2_X1 U12971 ( .A1(n15468), .A2(n11083), .ZN(n11084) );
  AOI211_X1 U12972 ( .C1(n15502), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n11869), .B(
        n11084), .ZN(n11089) );
  OAI211_X1 U12973 ( .C1(n11087), .C2(n11086), .A(n15512), .B(n11085), .ZN(
        n11088) );
  OAI211_X1 U12974 ( .C1(n11091), .C2(n11090), .A(n11089), .B(n11088), .ZN(
        P2_U3222) );
  NAND2_X1 U12975 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n11479) );
  INV_X1 U12976 ( .A(n11479), .ZN(n11097) );
  INV_X1 U12977 ( .A(n11106), .ZN(n11095) );
  NOR3_X1 U12978 ( .A1(n15445), .A2(n11093), .A3(n11092), .ZN(n11094) );
  NOR3_X1 U12979 ( .A1(n15508), .A2(n11095), .A3(n11094), .ZN(n11096) );
  AOI211_X1 U12980 ( .C1(n15502), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n11097), .B(
        n11096), .ZN(n11102) );
  OAI211_X1 U12981 ( .C1(n11100), .C2(n11099), .A(n15512), .B(n11098), .ZN(
        n11101) );
  OAI211_X1 U12982 ( .C1(n15468), .C2(n11103), .A(n11102), .B(n11101), .ZN(
        P2_U3219) );
  NAND2_X1 U12983 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n11642) );
  INV_X1 U12984 ( .A(n11642), .ZN(n11109) );
  AND3_X1 U12985 ( .A1(n11106), .A2(n11105), .A3(n11104), .ZN(n11107) );
  NOR3_X1 U12986 ( .A1(n15508), .A2(n11175), .A3(n11107), .ZN(n11108) );
  AOI211_X1 U12987 ( .C1(n15502), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n11109), .B(
        n11108), .ZN(n11114) );
  OAI211_X1 U12988 ( .C1(n11112), .C2(n11111), .A(n15512), .B(n11110), .ZN(
        n11113) );
  OAI211_X1 U12989 ( .C1(n15468), .C2(n11115), .A(n11114), .B(n11113), .ZN(
        P2_U3220) );
  INV_X1 U12990 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11116) );
  NOR2_X1 U12991 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11116), .ZN(n11510) );
  AND3_X1 U12992 ( .A1(n11118), .A2(n15431), .A3(n11117), .ZN(n11119) );
  NOR3_X1 U12993 ( .A1(n15508), .A2(n11120), .A3(n11119), .ZN(n11121) );
  AOI211_X1 U12994 ( .C1(n15502), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n11510), .B(
        n11121), .ZN(n11126) );
  OAI211_X1 U12995 ( .C1(n11124), .C2(n11123), .A(n15512), .B(n11122), .ZN(
        n11125) );
  OAI211_X1 U12996 ( .C1(n15468), .C2(n11127), .A(n11126), .B(n11125), .ZN(
        P2_U3217) );
  NAND2_X1 U12997 ( .A1(n15512), .A2(n11130), .ZN(n11129) );
  NAND2_X1 U12998 ( .A1(n15494), .A2(n15901), .ZN(n11128) );
  NAND3_X1 U12999 ( .A1(n15468), .A2(n11129), .A3(n11128), .ZN(n11132) );
  OAI22_X1 U13000 ( .A1(n11130), .A2(n15412), .B1(n15508), .B2(n15901), .ZN(
        n11131) );
  MUX2_X1 U13001 ( .A(n11132), .B(n11131), .S(n15418), .Z(n11136) );
  INV_X1 U13002 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n11134) );
  OAI22_X1 U13003 ( .A1(n15441), .A2(n11134), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11133), .ZN(n11135) );
  OR2_X1 U13004 ( .A1(n11136), .A2(n11135), .ZN(P2_U3214) );
  NAND2_X1 U13005 ( .A1(n11138), .A2(n11137), .ZN(n15529) );
  INV_X1 U13006 ( .A(n15862), .ZN(n15534) );
  INV_X1 U13007 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11139) );
  MUX2_X1 U13008 ( .A(n11139), .B(P1_REG1_REG_6__SCAN_IN), .S(n11211), .Z(
        n11145) );
  INV_X1 U13009 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n11141) );
  INV_X1 U13010 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n11140) );
  INV_X1 U13011 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15885) );
  NAND3_X1 U13012 ( .A1(n14772), .A2(n15398), .A3(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14770) );
  OAI21_X1 U13013 ( .B1(n11147), .B2(n11140), .A(n14770), .ZN(n11428) );
  MUX2_X1 U13014 ( .A(n11141), .B(P1_REG1_REG_2__SCAN_IN), .S(n11150), .Z(
        n11429) );
  NAND2_X1 U13015 ( .A1(n11428), .A2(n11429), .ZN(n11427) );
  OAI21_X1 U13016 ( .B1(n11150), .B2(n11141), .A(n11427), .ZN(n14781) );
  INV_X1 U13017 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11793) );
  MUX2_X1 U13018 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n11793), .S(n15393), .Z(
        n14782) );
  NAND2_X1 U13019 ( .A1(n14781), .A2(n14782), .ZN(n15856) );
  NAND2_X1 U13020 ( .A1(n15393), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n15854) );
  INV_X1 U13021 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11142) );
  MUX2_X1 U13022 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n11142), .S(n15863), .Z(
        n15855) );
  AOI21_X1 U13023 ( .B1(n15856), .B2(n15854), .A(n15855), .ZN(n15858) );
  AOI21_X1 U13024 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n15861), .A(n15858), .ZN(
        n11261) );
  XOR2_X1 U13025 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n11263), .Z(n11262) );
  NAND2_X1 U13026 ( .A1(n11261), .A2(n11262), .ZN(n11260) );
  OAI21_X1 U13027 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n11263), .A(n11260), .ZN(
        n11144) );
  NOR2_X1 U13028 ( .A1(n11144), .A2(n11145), .ZN(n11206) );
  INV_X1 U13029 ( .A(n15529), .ZN(n11143) );
  NAND2_X1 U13030 ( .A1(n11143), .A2(n13009), .ZN(n15859) );
  AOI211_X1 U13031 ( .C1(n11145), .C2(n11144), .A(n11206), .B(n15859), .ZN(
        n11167) );
  NAND2_X1 U13032 ( .A1(n11449), .A2(n15518), .ZN(n11146) );
  NOR2_X2 U13033 ( .A1(n15529), .A2(n11146), .ZN(n15869) );
  MUX2_X1 U13034 ( .A(n11148), .B(P1_REG2_REG_1__SCAN_IN), .S(n11147), .Z(
        n14775) );
  AND2_X1 U13035 ( .A1(n15398), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U13036 ( .A1(n14775), .A2(n14776), .ZN(n14774) );
  NAND2_X1 U13037 ( .A1(n14773), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n11149) );
  NAND2_X1 U13038 ( .A1(n14774), .A2(n11149), .ZN(n11430) );
  MUX2_X1 U13039 ( .A(n11151), .B(P1_REG2_REG_2__SCAN_IN), .S(n11150), .Z(
        n11431) );
  NAND2_X1 U13040 ( .A1(n11430), .A2(n11431), .ZN(n14786) );
  NAND2_X1 U13041 ( .A1(n11436), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14785) );
  NAND2_X1 U13042 ( .A1(n14786), .A2(n14785), .ZN(n11154) );
  MUX2_X1 U13043 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11152), .S(n15393), .Z(
        n11153) );
  NAND2_X1 U13044 ( .A1(n11154), .A2(n11153), .ZN(n15865) );
  NAND2_X1 U13045 ( .A1(n15393), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n15864) );
  NAND2_X1 U13046 ( .A1(n15865), .A2(n15864), .ZN(n11157) );
  MUX2_X1 U13047 ( .A(n11155), .B(P1_REG2_REG_4__SCAN_IN), .S(n15863), .Z(
        n11156) );
  NAND2_X1 U13048 ( .A1(n11157), .A2(n11156), .ZN(n15868) );
  NAND2_X1 U13049 ( .A1(n15861), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n11265) );
  NAND2_X1 U13050 ( .A1(n15868), .A2(n11265), .ZN(n11159) );
  MUX2_X1 U13051 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n12160), .S(n11263), .Z(
        n11158) );
  NAND2_X1 U13052 ( .A1(n11159), .A2(n11158), .ZN(n11267) );
  NAND2_X1 U13053 ( .A1(n11263), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n11164) );
  NAND2_X1 U13054 ( .A1(n11267), .A2(n11164), .ZN(n11162) );
  MUX2_X1 U13055 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11160), .S(n11211), .Z(
        n11161) );
  NAND2_X1 U13056 ( .A1(n11162), .A2(n11161), .ZN(n11216) );
  MUX2_X1 U13057 ( .A(n11160), .B(P1_REG2_REG_6__SCAN_IN), .S(n11211), .Z(
        n11163) );
  NAND3_X1 U13058 ( .A1(n11267), .A2(n11164), .A3(n11163), .ZN(n11165) );
  AND3_X1 U13059 ( .A1(n15869), .A2(n11216), .A3(n11165), .ZN(n11166) );
  NOR2_X1 U13060 ( .A1(n11167), .A2(n11166), .ZN(n11170) );
  NAND2_X1 U13061 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n12015) );
  INV_X1 U13062 ( .A(n12015), .ZN(n11168) );
  AOI21_X1 U13063 ( .B1(n15526), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n11168), .ZN(
        n11169) );
  OAI211_X1 U13064 ( .C1(n11171), .C2(n15534), .A(n11170), .B(n11169), .ZN(
        P1_U3249) );
  NAND2_X1 U13065 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11737) );
  INV_X1 U13066 ( .A(n11737), .ZN(n11179) );
  INV_X1 U13067 ( .A(n11172), .ZN(n11177) );
  NOR3_X1 U13068 ( .A1(n11175), .A2(n11174), .A3(n11173), .ZN(n11176) );
  NOR3_X1 U13069 ( .A1(n11177), .A2(n11176), .A3(n15508), .ZN(n11178) );
  AOI211_X1 U13070 ( .C1(n15502), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n11179), .B(
        n11178), .ZN(n11184) );
  OAI211_X1 U13071 ( .C1(n11182), .C2(n11181), .A(n15512), .B(n11180), .ZN(
        n11183) );
  OAI211_X1 U13072 ( .C1(n15468), .C2(n11185), .A(n11184), .B(n11183), .ZN(
        P2_U3221) );
  INV_X1 U13073 ( .A(n11186), .ZN(n11189) );
  INV_X1 U13074 ( .A(n11278), .ZN(n12419) );
  OAI222_X1 U13075 ( .A1(n14370), .A2(n11187), .B1(n14378), .B2(n11189), .C1(
        P2_U3088), .C2(n12419), .ZN(P2_U3316) );
  INV_X1 U13076 ( .A(n14805), .ZN(n11190) );
  OAI222_X1 U13077 ( .A1(n11190), .A2(P1_U3086), .B1(n15160), .B2(n11189), 
        .C1(n11188), .C2(n15157), .ZN(P1_U3344) );
  OAI21_X1 U13078 ( .B1(n11192), .B2(P2_REG1_REG_9__SCAN_IN), .A(n11191), .ZN(
        n11195) );
  MUX2_X1 U13079 ( .A(n10466), .B(P2_REG1_REG_10__SCAN_IN), .S(n11193), .Z(
        n11194) );
  NOR2_X1 U13080 ( .A1(n11195), .A2(n11194), .ZN(n11282) );
  AOI211_X1 U13081 ( .C1(n11195), .C2(n11194), .A(n15508), .B(n11282), .ZN(
        n11199) );
  NAND2_X1 U13082 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n12139)
         );
  INV_X1 U13083 ( .A(n12139), .ZN(n11196) );
  AOI21_X1 U13084 ( .B1(n15502), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n11196), 
        .ZN(n11197) );
  OAI21_X1 U13085 ( .B1(n15468), .B2(n11277), .A(n11197), .ZN(n11198) );
  NOR2_X1 U13086 ( .A1(n11199), .A2(n11198), .ZN(n11205) );
  AOI21_X1 U13087 ( .B1(n12174), .B2(n11201), .A(n11200), .ZN(n11203) );
  XNOR2_X1 U13088 ( .A(n11277), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U13089 ( .A1(n11203), .A2(n11202), .ZN(n11273) );
  OAI211_X1 U13090 ( .C1(n11203), .C2(n11202), .A(n11273), .B(n15512), .ZN(
        n11204) );
  NAND2_X1 U13091 ( .A1(n11205), .A2(n11204), .ZN(P2_U3224) );
  AOI21_X1 U13092 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n11211), .A(n11206), .ZN(
        n11209) );
  INV_X1 U13093 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n11207) );
  MUX2_X1 U13094 ( .A(n11207), .B(P1_REG1_REG_7__SCAN_IN), .S(n11295), .Z(
        n11208) );
  NOR2_X1 U13095 ( .A1(n11209), .A2(n11208), .ZN(n11290) );
  AOI211_X1 U13096 ( .C1(n11209), .C2(n11208), .A(n15859), .B(n11290), .ZN(
        n11222) );
  NAND2_X1 U13097 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n12096) );
  INV_X1 U13098 ( .A(n12096), .ZN(n11210) );
  AOI21_X1 U13099 ( .B1(n15526), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n11210), .ZN(
        n11219) );
  NAND2_X1 U13100 ( .A1(n11211), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U13101 ( .A1(n11216), .A2(n11215), .ZN(n11213) );
  MUX2_X1 U13102 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n12242), .S(n11295), .Z(
        n11212) );
  NAND2_X1 U13103 ( .A1(n11213), .A2(n11212), .ZN(n11316) );
  MUX2_X1 U13104 ( .A(n12242), .B(P1_REG2_REG_7__SCAN_IN), .S(n11295), .Z(
        n11214) );
  NAND3_X1 U13105 ( .A1(n11216), .A2(n11215), .A3(n11214), .ZN(n11217) );
  NAND3_X1 U13106 ( .A1(n15869), .A2(n11316), .A3(n11217), .ZN(n11218) );
  OAI211_X1 U13107 ( .C1(n15534), .C2(n11220), .A(n11219), .B(n11218), .ZN(
        n11221) );
  OR2_X1 U13108 ( .A1(n11222), .A2(n11221), .ZN(P1_U3250) );
  INV_X1 U13109 ( .A(n11223), .ZN(n11224) );
  NAND2_X1 U13110 ( .A1(n13871), .A2(n11224), .ZN(n11225) );
  XNOR2_X1 U13111 ( .A(n15908), .B(n11350), .ZN(n11227) );
  OAI21_X1 U13112 ( .B1(n12498), .B2(n11669), .A(n11494), .ZN(n11229) );
  AOI21_X1 U13113 ( .B1(n11230), .B2(n11229), .A(n11349), .ZN(n11257) );
  NAND2_X1 U13114 ( .A1(n11247), .A2(n16157), .ZN(n11233) );
  INV_X1 U13115 ( .A(n11250), .ZN(n11231) );
  NAND2_X1 U13116 ( .A1(n11251), .A2(n11231), .ZN(n11232) );
  OAI21_X1 U13117 ( .B1(n11248), .B2(n11233), .A(n11232), .ZN(n11235) );
  AND2_X1 U13118 ( .A1(n11251), .A2(n11253), .ZN(n11237) );
  INV_X1 U13119 ( .A(n11236), .ZN(n11238) );
  INV_X1 U13120 ( .A(n11237), .ZN(n11239) );
  NAND2_X1 U13121 ( .A1(n11248), .A2(n11664), .ZN(n11242) );
  INV_X1 U13122 ( .A(n11665), .ZN(n11241) );
  OAI22_X1 U13123 ( .A1(n11418), .A2(n13551), .B1(n11538), .B2(n13561), .ZN(
        n11243) );
  AOI21_X1 U13124 ( .B1(n13549), .B2(n13590), .A(n11243), .ZN(n11256) );
  OAI21_X1 U13125 ( .B1(n11245), .B2(n11657), .A(n11244), .ZN(n11246) );
  AOI21_X1 U13126 ( .B1(n11248), .B2(n11247), .A(n11246), .ZN(n11249) );
  OAI21_X1 U13127 ( .B1(n11251), .B2(n11250), .A(n11249), .ZN(n11254) );
  INV_X1 U13128 ( .A(n11251), .ZN(n11252) );
  AOI22_X1 U13129 ( .A1(n11254), .A2(P3_STATE_REG_SCAN_IN), .B1(n11253), .B2(
        n11252), .ZN(n11411) );
  NAND2_X1 U13130 ( .A1(n11411), .A2(n13870), .ZN(n11356) );
  NAND2_X1 U13131 ( .A1(n11356), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n11255) );
  OAI211_X1 U13132 ( .C1(n11257), .C2(n13566), .A(n11256), .B(n11255), .ZN(
        P3_U3162) );
  INV_X1 U13133 ( .A(SI_16_), .ZN(n15196) );
  OAI222_X1 U13134 ( .A1(n13131), .A2(n11259), .B1(n13880), .B2(n15196), .C1(
        n11258), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U13135 ( .A(n15859), .ZN(n15539) );
  OAI21_X1 U13136 ( .B1(n11262), .B2(n11261), .A(n11260), .ZN(n11269) );
  MUX2_X1 U13137 ( .A(n12160), .B(P1_REG2_REG_5__SCAN_IN), .S(n11263), .Z(
        n11264) );
  NAND3_X1 U13138 ( .A1(n15868), .A2(n11265), .A3(n11264), .ZN(n11266) );
  AND3_X1 U13139 ( .A1(n15869), .A2(n11267), .A3(n11266), .ZN(n11268) );
  AOI21_X1 U13140 ( .B1(n15539), .B2(n11269), .A(n11268), .ZN(n11271) );
  AND2_X1 U13141 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11920) );
  AOI21_X1 U13142 ( .B1(n15526), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n11920), .ZN(
        n11270) );
  OAI211_X1 U13143 ( .C1(n11272), .C2(n15534), .A(n11271), .B(n11270), .ZN(
        P1_U3248) );
  MUX2_X1 U13144 ( .A(n12542), .B(P2_REG2_REG_11__SCAN_IN), .S(n11278), .Z(
        n11276) );
  OAI21_X1 U13145 ( .B1(n11274), .B2(n11277), .A(n11273), .ZN(n11275) );
  NOR2_X1 U13146 ( .A1(n11275), .A2(n11276), .ZN(n12405) );
  AOI21_X1 U13147 ( .B1(n11276), .B2(n11275), .A(n12405), .ZN(n11288) );
  NOR2_X1 U13148 ( .A1(n11277), .A2(n10466), .ZN(n11281) );
  MUX2_X1 U13149 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11279), .S(n11278), .Z(
        n11280) );
  OAI21_X1 U13150 ( .B1(n11282), .B2(n11281), .A(n11280), .ZN(n12418) );
  OR3_X1 U13151 ( .A1(n11282), .A2(n11281), .A3(n11280), .ZN(n11283) );
  NAND3_X1 U13152 ( .A1(n12418), .A2(n15494), .A3(n11283), .ZN(n11287) );
  NOR2_X1 U13153 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12473), .ZN(n11285) );
  NOR2_X1 U13154 ( .A1(n15468), .A2(n12419), .ZN(n11284) );
  AOI211_X1 U13155 ( .C1(n15502), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11285), 
        .B(n11284), .ZN(n11286) );
  OAI211_X1 U13156 ( .C1(n11288), .C2(n15412), .A(n11287), .B(n11286), .ZN(
        P2_U3225) );
  INV_X1 U13157 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11289) );
  MUX2_X1 U13158 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n11289), .S(n11334), .Z(
        n11293) );
  INV_X1 U13159 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n11291) );
  MUX2_X1 U13160 ( .A(n11291), .B(P1_REG1_REG_8__SCAN_IN), .S(n11321), .Z(
        n11311) );
  OAI21_X1 U13161 ( .B1(n11293), .B2(n11292), .A(n11329), .ZN(n11308) );
  NAND2_X1 U13162 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n14655) );
  INV_X1 U13163 ( .A(n14655), .ZN(n11294) );
  AOI21_X1 U13164 ( .B1(n15526), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n11294), .ZN(
        n11305) );
  NAND2_X1 U13165 ( .A1(n11295), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n11315) );
  NAND2_X1 U13166 ( .A1(n11316), .A2(n11315), .ZN(n11297) );
  MUX2_X1 U13167 ( .A(n12260), .B(P1_REG2_REG_8__SCAN_IN), .S(n11321), .Z(
        n11296) );
  NAND2_X1 U13168 ( .A1(n11297), .A2(n11296), .ZN(n11318) );
  NAND2_X1 U13169 ( .A1(n11298), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11302) );
  NAND2_X1 U13170 ( .A1(n11318), .A2(n11302), .ZN(n11300) );
  MUX2_X1 U13171 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n12326), .S(n11334), .Z(
        n11299) );
  NAND2_X1 U13172 ( .A1(n11300), .A2(n11299), .ZN(n11340) );
  MUX2_X1 U13173 ( .A(n12326), .B(P1_REG2_REG_9__SCAN_IN), .S(n11334), .Z(
        n11301) );
  NAND3_X1 U13174 ( .A1(n11318), .A2(n11302), .A3(n11301), .ZN(n11303) );
  NAND3_X1 U13175 ( .A1(n15869), .A2(n11340), .A3(n11303), .ZN(n11304) );
  OAI211_X1 U13176 ( .C1(n15534), .C2(n11306), .A(n11305), .B(n11304), .ZN(
        n11307) );
  AOI21_X1 U13177 ( .B1(n11308), .B2(n15539), .A(n11307), .ZN(n11309) );
  INV_X1 U13178 ( .A(n11309), .ZN(P1_U3252) );
  OAI21_X1 U13179 ( .B1(n11312), .B2(n11311), .A(n11310), .ZN(n11323) );
  NAND2_X1 U13180 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n12351) );
  INV_X1 U13181 ( .A(n12351), .ZN(n11313) );
  AOI21_X1 U13182 ( .B1(n15526), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n11313), .ZN(
        n11320) );
  MUX2_X1 U13183 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n12260), .S(n11321), .Z(
        n11314) );
  NAND3_X1 U13184 ( .A1(n11316), .A2(n11315), .A3(n11314), .ZN(n11317) );
  NAND3_X1 U13185 ( .A1(n15869), .A2(n11318), .A3(n11317), .ZN(n11319) );
  OAI211_X1 U13186 ( .C1(n15534), .C2(n11321), .A(n11320), .B(n11319), .ZN(
        n11322) );
  AOI21_X1 U13187 ( .B1(n11323), .B2(n15539), .A(n11322), .ZN(n11324) );
  INV_X1 U13188 ( .A(n11324), .ZN(P1_U3251) );
  OAI22_X1 U13189 ( .A1(n11228), .A2(n13551), .B1(n11592), .B2(n13561), .ZN(
        n11326) );
  NOR2_X1 U13190 ( .A1(n11502), .A2(n13566), .ZN(n11325) );
  AOI211_X1 U13191 ( .C1(P3_REG3_REG_0__SCAN_IN), .C2(n11356), .A(n11326), .B(
        n11325), .ZN(n11327) );
  INV_X1 U13192 ( .A(n11327), .ZN(P3_U3172) );
  INV_X1 U13193 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11328) );
  MUX2_X1 U13194 ( .A(n11328), .B(P1_REG1_REG_10__SCAN_IN), .S(n11528), .Z(
        n11331) );
  OAI21_X1 U13195 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n11334), .A(n11329), .ZN(
        n11330) );
  AOI211_X1 U13196 ( .C1(n11331), .C2(n11330), .A(n15859), .B(n11523), .ZN(
        n11346) );
  NOR2_X1 U13197 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11332), .ZN(n11333) );
  AOI21_X1 U13198 ( .B1(n15526), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11333), 
        .ZN(n11343) );
  NAND2_X1 U13199 ( .A1(n11334), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11339) );
  NAND2_X1 U13200 ( .A1(n11340), .A2(n11339), .ZN(n11337) );
  MUX2_X1 U13201 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11335), .S(n11528), .Z(
        n11336) );
  NAND2_X1 U13202 ( .A1(n11337), .A2(n11336), .ZN(n14802) );
  MUX2_X1 U13203 ( .A(n11335), .B(P1_REG2_REG_10__SCAN_IN), .S(n11528), .Z(
        n11338) );
  NAND3_X1 U13204 ( .A1(n11340), .A2(n11339), .A3(n11338), .ZN(n11341) );
  NAND3_X1 U13205 ( .A1(n15869), .A2(n14802), .A3(n11341), .ZN(n11342) );
  OAI211_X1 U13206 ( .C1(n15534), .C2(n11344), .A(n11343), .B(n11342), .ZN(
        n11345) );
  OR2_X1 U13207 ( .A1(n11346), .A2(n11345), .ZN(P1_U3253) );
  INV_X1 U13208 ( .A(n11347), .ZN(n11348) );
  XNOR2_X1 U13209 ( .A(n11412), .B(n11418), .ZN(n11352) );
  AOI21_X1 U13210 ( .B1(n11353), .B2(n11352), .A(n11416), .ZN(n11358) );
  NOR2_X1 U13211 ( .A1(n11228), .A2(n13559), .ZN(n11355) );
  OAI22_X1 U13212 ( .A1(n15961), .A2(n13551), .B1(n15970), .B2(n13561), .ZN(
        n11354) );
  AOI211_X1 U13213 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n11356), .A(n11355), .B(
        n11354), .ZN(n11357) );
  OAI21_X1 U13214 ( .B1(n11358), .B2(n13566), .A(n11357), .ZN(P3_U3177) );
  OAI222_X1 U13215 ( .A1(n13131), .A2(n11359), .B1(n15821), .B2(P3_U3151), 
        .C1(n15275), .C2(n13880), .ZN(P3_U3278) );
  NAND2_X1 U13216 ( .A1(n13138), .A2(P2_U3947), .ZN(n11360) );
  OAI21_X1 U13217 ( .B1(n15405), .B2(n9095), .A(n11360), .ZN(P2_U3531) );
  INV_X1 U13218 ( .A(n11815), .ZN(n11532) );
  INV_X1 U13219 ( .A(n11361), .ZN(n11363) );
  OAI222_X1 U13220 ( .A1(P1_U3086), .A2(n11532), .B1(n15160), .B2(n11363), 
        .C1(n11362), .C2(n15157), .ZN(P1_U3343) );
  OAI222_X1 U13221 ( .A1(n14370), .A2(n11364), .B1(n14378), .B2(n11363), .C1(
        n12421), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U13222 ( .A(n13996), .ZN(n13975) );
  AOI22_X1 U13223 ( .A1(n13975), .A2(n14027), .B1(n13143), .B2(n13999), .ZN(
        n11370) );
  OAI21_X1 U13224 ( .B1(n11366), .B2(n11365), .A(n10970), .ZN(n11368) );
  INV_X1 U13225 ( .A(n11367), .ZN(n11491) );
  AOI22_X1 U13226 ( .A1(n13940), .A2(n11368), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n11491), .ZN(n11369) );
  OAI211_X1 U13227 ( .C1(n13133), .C2(n13992), .A(n11370), .B(n11369), .ZN(
        P2_U3194) );
  OAI21_X1 U13228 ( .B1(n11373), .B2(n11372), .A(n11371), .ZN(n11374) );
  NAND2_X1 U13229 ( .A1(n15845), .A2(n11374), .ZN(n11384) );
  AOI22_X1 U13230 ( .A1(n15832), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11383) );
  INV_X1 U13231 ( .A(n11375), .ZN(n11378) );
  INV_X1 U13232 ( .A(n11376), .ZN(n11377) );
  NAND2_X1 U13233 ( .A1(n11378), .A2(n11377), .ZN(n11379) );
  NAND2_X1 U13234 ( .A1(n11380), .A2(n11379), .ZN(n11381) );
  NAND2_X1 U13235 ( .A1(n15844), .A2(n11381), .ZN(n11382) );
  NAND3_X1 U13236 ( .A1(n11384), .A2(n11383), .A3(n11382), .ZN(n11390) );
  INV_X1 U13237 ( .A(n11385), .ZN(n11387) );
  NAND3_X1 U13238 ( .A1(n11395), .A2(n11387), .A3(n11386), .ZN(n11388) );
  AOI21_X1 U13239 ( .B1(n15626), .B2(n11388), .A(n15840), .ZN(n11389) );
  AOI211_X1 U13240 ( .C1(n15834), .C2(n11391), .A(n11390), .B(n11389), .ZN(
        n11392) );
  INV_X1 U13241 ( .A(n11392), .ZN(P3_U3184) );
  INV_X1 U13242 ( .A(n15489), .ZN(n12423) );
  OAI222_X1 U13243 ( .A1(n14370), .A2(n11393), .B1(n14378), .B2(n11394), .C1(
        n12423), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U13244 ( .A(n12115), .ZN(n11821) );
  OAI222_X1 U13245 ( .A1(n11821), .A2(P1_U3086), .B1(n15157), .B2(n9308), .C1(
        n11394), .C2(n15160), .ZN(P1_U3342) );
  INV_X1 U13246 ( .A(n15840), .ZN(n15806) );
  OAI21_X1 U13247 ( .B1(n11396), .B2(n15613), .A(n11395), .ZN(n11408) );
  NAND2_X1 U13248 ( .A1(n11398), .A2(n11397), .ZN(n11399) );
  NAND2_X1 U13249 ( .A1(n11400), .A2(n11399), .ZN(n11401) );
  NAND2_X1 U13250 ( .A1(n15845), .A2(n11401), .ZN(n11406) );
  AOI22_X1 U13251 ( .A1(n15832), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11405) );
  XNOR2_X1 U13252 ( .A(n11402), .B(P3_REG1_REG_1__SCAN_IN), .ZN(n11403) );
  NAND2_X1 U13253 ( .A1(n15844), .A2(n11403), .ZN(n11404) );
  NAND3_X1 U13254 ( .A1(n11406), .A2(n11405), .A3(n11404), .ZN(n11407) );
  AOI21_X1 U13255 ( .B1(n15806), .B2(n11408), .A(n11407), .ZN(n11409) );
  OAI21_X1 U13256 ( .B1(n11410), .B2(n15822), .A(n11409), .ZN(P3_U3183) );
  INV_X1 U13257 ( .A(n11412), .ZN(n11413) );
  NOR2_X1 U13258 ( .A1(n13587), .A2(n11413), .ZN(n11415) );
  XNOR2_X1 U13259 ( .A(n15986), .B(n11350), .ZN(n11566) );
  XNOR2_X1 U13260 ( .A(n15961), .B(n11566), .ZN(n11414) );
  OAI21_X1 U13261 ( .B1(n11416), .B2(n11415), .A(n11414), .ZN(n11417) );
  NAND3_X1 U13262 ( .A1(n7527), .A2(n13476), .A3(n11417), .ZN(n11421) );
  NOR2_X1 U13263 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15343), .ZN(n15628) );
  OAI22_X1 U13264 ( .A1(n11418), .A2(n13559), .B1(n11886), .B2(n13551), .ZN(
        n11419) );
  AOI211_X1 U13265 ( .C1(n12504), .C2(n15986), .A(n15628), .B(n11419), .ZN(
        n11420) );
  OAI211_X1 U13266 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12382), .A(n11421), .B(
        n11420), .ZN(P3_U3158) );
  NAND2_X1 U13267 ( .A1(n13244), .A2(n15405), .ZN(n11422) );
  OAI21_X1 U13268 ( .B1(n9308), .B2(n15405), .A(n11422), .ZN(P2_U3544) );
  OAI222_X1 U13269 ( .A1(n13131), .A2(n11425), .B1(n13880), .B2(n11424), .C1(
        n11423), .C2(P3_U3151), .ZN(P3_U3277) );
  NAND2_X1 U13270 ( .A1(n15526), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n11426) );
  OAI21_X1 U13271 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n12279), .A(n11426), .ZN(
        n11435) );
  OAI211_X1 U13272 ( .C1(n11429), .C2(n11428), .A(n15539), .B(n11427), .ZN(
        n11433) );
  OAI211_X1 U13273 ( .C1(n11431), .C2(n11430), .A(n15869), .B(n14786), .ZN(
        n11432) );
  NAND2_X1 U13274 ( .A1(n11433), .A2(n11432), .ZN(n11434) );
  AOI211_X1 U13275 ( .C1(n11436), .C2(n15862), .A(n11435), .B(n11434), .ZN(
        n11451) );
  NAND2_X2 U13276 ( .A1(n11437), .A2(n11844), .ZN(n14585) );
  OR2_X4 U13277 ( .A1(n16012), .A2(n14585), .ZN(n14586) );
  NAND2_X4 U13278 ( .A1(n11438), .A2(n11844), .ZN(n14588) );
  INV_X2 U13279 ( .A(n14588), .ZN(n11917) );
  INV_X1 U13280 ( .A(n11844), .ZN(n11439) );
  AOI22_X1 U13281 ( .A1(n11917), .A2(n15914), .B1(n11439), .B2(n15398), .ZN(
        n11440) );
  OAI21_X1 U13282 ( .B1(n14586), .B2(n11441), .A(n11440), .ZN(n11445) );
  NOR2_X1 U13283 ( .A1(n11844), .A2(n15885), .ZN(n11442) );
  AOI21_X1 U13284 ( .B1(n11917), .B2(n15924), .A(n11442), .ZN(n11444) );
  NAND2_X1 U13285 ( .A1(n14526), .A2(n15914), .ZN(n11443) );
  NAND2_X1 U13286 ( .A1(n11444), .A2(n11443), .ZN(n11545) );
  NAND2_X1 U13287 ( .A1(n11445), .A2(n11545), .ZN(n11544) );
  OR2_X1 U13288 ( .A1(n11445), .A2(n11545), .ZN(n11446) );
  NAND2_X1 U13289 ( .A1(n11544), .A2(n11446), .ZN(n11745) );
  MUX2_X1 U13290 ( .A(n11745), .B(n14776), .S(n15518), .Z(n11447) );
  INV_X1 U13291 ( .A(n11447), .ZN(n11450) );
  OR2_X1 U13292 ( .A1(n13009), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U13293 ( .A1(n11449), .A2(n11448), .ZN(n15519) );
  INV_X1 U13294 ( .A(n15398), .ZN(n15521) );
  NAND2_X1 U13295 ( .A1(n15519), .A2(n15521), .ZN(n15524) );
  OAI211_X1 U13296 ( .C1(n11450), .C2(n15161), .A(P1_U4016), .B(n15524), .ZN(
        n15872) );
  NAND2_X1 U13297 ( .A1(n11451), .A2(n15872), .ZN(P1_U3245) );
  NAND3_X1 U13298 ( .A1(n12624), .A2(n10458), .A3(n13399), .ZN(n15897) );
  INV_X1 U13299 ( .A(n15897), .ZN(n16121) );
  XNOR2_X1 U13300 ( .A(n13144), .B(n13143), .ZN(n13404) );
  INV_X1 U13301 ( .A(n13404), .ZN(n11454) );
  INV_X1 U13302 ( .A(n11452), .ZN(n11453) );
  NAND2_X1 U13303 ( .A1(n11454), .A2(n11453), .ZN(n11694) );
  NAND2_X1 U13304 ( .A1(n12036), .A2(n15948), .ZN(n11455) );
  NAND2_X1 U13305 ( .A1(n11694), .A2(n11455), .ZN(n11456) );
  XNOR2_X1 U13306 ( .A(n14027), .B(n14248), .ZN(n13403) );
  INV_X1 U13307 ( .A(n13403), .ZN(n11462) );
  NAND2_X1 U13308 ( .A1(n11456), .A2(n11462), .ZN(n11675) );
  OR2_X1 U13309 ( .A1(n11456), .A2(n11462), .ZN(n11457) );
  NAND2_X1 U13310 ( .A1(n11675), .A2(n11457), .ZN(n14249) );
  INV_X1 U13311 ( .A(n11701), .ZN(n11458) );
  OR2_X1 U13312 ( .A1(n11701), .A2(n14248), .ZN(n11717) );
  OAI211_X1 U13313 ( .C1(n11458), .C2(n11673), .A(n14302), .B(n11717), .ZN(
        n14246) );
  OAI21_X1 U13314 ( .B1(n11673), .B2(n16182), .A(n14246), .ZN(n11470) );
  OR2_X1 U13315 ( .A1(n13399), .A2(n13452), .ZN(n11459) );
  NOR2_X1 U13316 ( .A1(n13138), .A2(n15895), .ZN(n11706) );
  NAND2_X1 U13317 ( .A1(n13404), .A2(n11706), .ZN(n11705) );
  NAND2_X1 U13318 ( .A1(n12036), .A2(n13143), .ZN(n11461) );
  NAND2_X1 U13319 ( .A1(n11705), .A2(n11461), .ZN(n11460) );
  NAND2_X1 U13320 ( .A1(n11460), .A2(n13403), .ZN(n11724) );
  NAND3_X1 U13321 ( .A1(n11705), .A2(n11462), .A3(n11461), .ZN(n11463) );
  AND2_X1 U13322 ( .A1(n11724), .A2(n11463), .ZN(n11469) );
  NAND2_X1 U13323 ( .A1(n11465), .A2(n11464), .ZN(n13454) );
  AND2_X1 U13324 ( .A1(n13454), .A2(n13024), .ZN(n11466) );
  NAND2_X1 U13325 ( .A1(n14249), .A2(n14121), .ZN(n11468) );
  AOI22_X1 U13326 ( .A1(n14091), .A2(n14026), .B1(n13144), .B2(n14089), .ZN(
        n11467) );
  OAI211_X1 U13327 ( .C1(n14214), .C2(n11469), .A(n11468), .B(n11467), .ZN(
        n14250) );
  AOI211_X1 U13328 ( .C1(n16121), .C2(n14249), .A(n11470), .B(n14250), .ZN(
        n11508) );
  INV_X1 U13329 ( .A(n11471), .ZN(n11472) );
  INV_X1 U13330 ( .A(n11696), .ZN(n11473) );
  NOR2_X1 U13331 ( .A1(n11474), .A2(n11473), .ZN(n11475) );
  NAND2_X1 U13332 ( .A1(n16188), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n11478) );
  OAI21_X1 U13333 ( .B1(n11508), .B2(n16188), .A(n11478), .ZN(P2_U3501) );
  INV_X1 U13334 ( .A(n13994), .ZN(n13931) );
  OAI21_X1 U13335 ( .B1(n13931), .B2(n11786), .A(n11479), .ZN(n11481) );
  INV_X1 U13336 ( .A(n14025), .ZN(n13178) );
  INV_X1 U13337 ( .A(n14023), .ZN(n12069) );
  OAI22_X1 U13338 ( .A1(n13178), .A2(n13992), .B1(n13996), .B2(n12069), .ZN(
        n11480) );
  AOI211_X1 U13339 ( .C1(n13182), .C2(n13999), .A(n11481), .B(n11480), .ZN(
        n11487) );
  OAI22_X1 U13340 ( .A1(n13897), .A2(n13178), .B1(n11482), .B2(n14001), .ZN(
        n11485) );
  NAND3_X1 U13341 ( .A1(n11485), .A2(n7411), .A3(n11484), .ZN(n11486) );
  OAI211_X1 U13342 ( .C1(n14001), .C2(n11488), .A(n11487), .B(n11486), .ZN(
        P2_U3199) );
  OAI22_X1 U13343 ( .A1(n13897), .A2(n13133), .B1(n15895), .B2(n14001), .ZN(
        n11490) );
  NAND2_X1 U13344 ( .A1(n11490), .A2(n11489), .ZN(n11493) );
  AOI22_X1 U13345 ( .A1(n13999), .A2(n13135), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n11491), .ZN(n11492) );
  OAI211_X1 U13346 ( .C1(n12036), .C2(n13996), .A(n11493), .B(n11492), .ZN(
        P2_U3204) );
  XNOR2_X1 U13347 ( .A(n11494), .B(n9708), .ZN(n11495) );
  INV_X1 U13348 ( .A(n15960), .ZN(n13708) );
  AOI222_X1 U13349 ( .A1(n13705), .A2(n11495), .B1(n13587), .B2(n9880), .C1(
        n13590), .C2(n13708), .ZN(n15905) );
  NAND2_X1 U13350 ( .A1(n9708), .A2(n11496), .ZN(n15903) );
  NAND3_X1 U13351 ( .A1(n15904), .A2(n15903), .A3(n16160), .ZN(n11497) );
  NAND2_X1 U13352 ( .A1(n15905), .A2(n11497), .ZN(n11540) );
  OAI22_X1 U13353 ( .A1(n13806), .A2(n11538), .B1(n16165), .B2(n9970), .ZN(
        n11498) );
  AOI21_X1 U13354 ( .B1(n11540), .B2(n16165), .A(n11498), .ZN(n11499) );
  INV_X1 U13355 ( .A(n11499), .ZN(P3_U3460) );
  NAND2_X1 U13356 ( .A1(n11500), .A2(n16157), .ZN(n11501) );
  OAI22_X1 U13357 ( .A1(n11502), .A2(n11501), .B1(n11228), .B2(n15962), .ZN(
        n11666) );
  OAI22_X1 U13358 ( .A1(n13806), .A2(n11592), .B1(n16165), .B2(n9972), .ZN(
        n11503) );
  AOI21_X1 U13359 ( .B1(n11666), .B2(n16165), .A(n11503), .ZN(n11504) );
  INV_X1 U13360 ( .A(n11504), .ZN(P3_U3459) );
  OAI222_X1 U13361 ( .A1(n13131), .A2(n11506), .B1(P3_U3151), .B2(n11505), 
        .C1(n13880), .C2(n15192), .ZN(P3_U3276) );
  INV_X2 U13362 ( .A(n16190), .ZN(n16192) );
  OR2_X1 U13363 ( .A1(n11508), .A2(n16190), .ZN(n11509) );
  OAI21_X1 U13364 ( .B1(n16192), .B2(n10550), .A(n11509), .ZN(P2_U3436) );
  INV_X1 U13365 ( .A(n13168), .ZN(n15995) );
  INV_X1 U13366 ( .A(n13992), .ZN(n13955) );
  AOI22_X1 U13367 ( .A1(n13975), .A2(n14025), .B1(n13955), .B2(n14027), .ZN(
        n11512) );
  AOI21_X1 U13368 ( .B1(n13994), .B2(n11116), .A(n11510), .ZN(n11511) );
  OAI211_X1 U13369 ( .C1(n15995), .C2(n13978), .A(n11512), .B(n11511), .ZN(
        n11517) );
  INV_X1 U13370 ( .A(n11599), .ZN(n11513) );
  AOI211_X1 U13371 ( .C1(n11515), .C2(n11514), .A(n11513), .B(n14001), .ZN(
        n11516) );
  OR2_X1 U13372 ( .A1(n11517), .A2(n11516), .ZN(P2_U3190) );
  INV_X1 U13373 ( .A(n11518), .ZN(n11520) );
  OAI222_X1 U13374 ( .A1(n7793), .A2(P1_U3086), .B1(n15160), .B2(n11520), .C1(
        n11519), .C2(n15157), .ZN(P1_U3341) );
  INV_X1 U13375 ( .A(n12424), .ZN(n15453) );
  OAI222_X1 U13376 ( .A1(n14370), .A2(n11521), .B1(n14378), .B2(n11520), .C1(
        P2_U3088), .C2(n15453), .ZN(P2_U3313) );
  INV_X1 U13377 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11522) );
  MUX2_X1 U13378 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n11522), .S(n11815), .Z(
        n11526) );
  INV_X1 U13379 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11524) );
  MUX2_X1 U13380 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11524), .S(n14805), .Z(
        n14794) );
  NAND2_X1 U13381 ( .A1(n11525), .A2(n11526), .ZN(n11811) );
  OAI21_X1 U13382 ( .B1(n11526), .B2(n11525), .A(n11811), .ZN(n11527) );
  NAND2_X1 U13383 ( .A1(n11527), .A2(n15539), .ZN(n11536) );
  MUX2_X1 U13384 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n12464), .S(n11815), .Z(
        n11530) );
  NAND2_X1 U13385 ( .A1(n11528), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n14801) );
  MUX2_X1 U13386 ( .A(n12397), .B(P1_REG2_REG_11__SCAN_IN), .S(n14805), .Z(
        n14800) );
  AOI21_X1 U13387 ( .B1(n14802), .B2(n14801), .A(n14800), .ZN(n14799) );
  AOI21_X1 U13388 ( .B1(n14805), .B2(P1_REG2_REG_11__SCAN_IN), .A(n14799), 
        .ZN(n11529) );
  NAND2_X1 U13389 ( .A1(n11529), .A2(n11530), .ZN(n11814) );
  OAI21_X1 U13390 ( .B1(n11530), .B2(n11529), .A(n11814), .ZN(n11534) );
  NAND2_X1 U13391 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14614)
         );
  NAND2_X1 U13392 ( .A1(n15526), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11531) );
  OAI211_X1 U13393 ( .C1(n15534), .C2(n11532), .A(n14614), .B(n11531), .ZN(
        n11533) );
  AOI21_X1 U13394 ( .B1(n11534), .B2(n15869), .A(n11533), .ZN(n11535) );
  NAND2_X1 U13395 ( .A1(n11536), .A2(n11535), .ZN(P1_U3255) );
  INV_X1 U13396 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n11537) );
  OAI22_X1 U13397 ( .A1(n13864), .A2(n11538), .B1(n16169), .B2(n11537), .ZN(
        n11539) );
  AOI21_X1 U13398 ( .B1(n11540), .B2(n16169), .A(n11539), .ZN(n11541) );
  INV_X1 U13399 ( .A(n11541), .ZN(P3_U3393) );
  OAI22_X1 U13400 ( .A1(n14586), .A2(n7694), .B1(n15978), .B2(n14588), .ZN(
        n11828) );
  OAI22_X1 U13401 ( .A1(n14585), .A2(n15978), .B1(n7694), .B2(n14588), .ZN(
        n11542) );
  XNOR2_X1 U13402 ( .A(n11542), .B(n14589), .ZN(n11827) );
  XOR2_X1 U13403 ( .A(n11828), .B(n11827), .Z(n11831) );
  OAI22_X1 U13404 ( .A1(n14586), .A2(n8555), .B1(n15934), .B2(n14588), .ZN(
        n11547) );
  OAI22_X1 U13405 ( .A1(n14585), .A2(n15934), .B1(n8555), .B2(n14588), .ZN(
        n11543) );
  XNOR2_X1 U13406 ( .A(n11543), .B(n14589), .ZN(n11546) );
  XNOR2_X1 U13407 ( .A(n11547), .B(n11546), .ZN(n11605) );
  OAI21_X1 U13408 ( .B1(n11545), .B2(n14589), .A(n11544), .ZN(n11606) );
  XOR2_X1 U13409 ( .A(n11831), .B(n11832), .Z(n11565) );
  INV_X1 U13410 ( .A(n11548), .ZN(n11550) );
  OR2_X1 U13411 ( .A1(n11550), .A2(n11549), .ZN(n12150) );
  INV_X1 U13412 ( .A(n11579), .ZN(n11551) );
  INV_X1 U13413 ( .A(n11562), .ZN(n11555) );
  NAND2_X1 U13414 ( .A1(n11557), .A2(n11552), .ZN(n11553) );
  NOR2_X1 U13415 ( .A1(n16009), .A2(n11553), .ZN(n11554) );
  INV_X1 U13416 ( .A(n12154), .ZN(n11556) );
  NAND2_X1 U13417 ( .A1(n11557), .A2(n11556), .ZN(n11559) );
  INV_X1 U13418 ( .A(n11557), .ZN(n11558) );
  NAND2_X1 U13419 ( .A1(n11562), .A2(n11560), .ZN(n11848) );
  NAND2_X1 U13420 ( .A1(n11848), .A2(n11561), .ZN(n11744) );
  AOI22_X1 U13421 ( .A1(n7185), .A2(n12281), .B1(n11744), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n11564) );
  INV_X1 U13422 ( .A(n11561), .ZN(n11580) );
  NOR2_X2 U13423 ( .A1(n11562), .A2(n11580), .ZN(n16197) );
  NAND2_X1 U13424 ( .A1(n16197), .A2(n14914), .ZN(n14538) );
  INV_X1 U13425 ( .A(n14538), .ZN(n14699) );
  AND2_X1 U13426 ( .A1(n16197), .A2(n15925), .ZN(n14714) );
  AOI22_X1 U13427 ( .A1(n14699), .A2(n14767), .B1(n14714), .B2(n14769), .ZN(
        n11563) );
  OAI211_X1 U13428 ( .C1(n11565), .C2(n14740), .A(n11564), .B(n11563), .ZN(
        P1_U3237) );
  INV_X1 U13429 ( .A(n11897), .ZN(n11578) );
  INV_X1 U13430 ( .A(n11566), .ZN(n11568) );
  CLKBUF_X3 U13431 ( .A(n11350), .Z(n13119) );
  XNOR2_X1 U13432 ( .A(n11569), .B(n13119), .ZN(n11570) );
  NOR2_X1 U13433 ( .A1(n11570), .A2(n13585), .ZN(n11647) );
  AOI21_X1 U13434 ( .B1(n13585), .B2(n11570), .A(n11647), .ZN(n11571) );
  OAI21_X1 U13435 ( .B1(n11572), .B2(n11571), .A(n11649), .ZN(n11573) );
  NAND2_X1 U13436 ( .A1(n11573), .A2(n13476), .ZN(n11577) );
  INV_X1 U13437 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11574) );
  NOR2_X1 U13438 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11574), .ZN(n15640) );
  OAI22_X1 U13439 ( .A1(n15961), .A2(n13559), .B1(n11994), .B2(n13551), .ZN(
        n11575) );
  AOI211_X1 U13440 ( .C1(n12504), .C2(n16001), .A(n15640), .B(n11575), .ZN(
        n11576) );
  OAI211_X1 U13441 ( .C1(n11578), .C2(n12382), .A(n11577), .B(n11576), .ZN(
        P3_U3170) );
  INV_X2 U13442 ( .A(n16142), .ZN(n15984) );
  XNOR2_X1 U13443 ( .A(n11583), .B(n11582), .ZN(n12225) );
  INV_X1 U13444 ( .A(n12225), .ZN(n11589) );
  XNOR2_X1 U13445 ( .A(n11585), .B(n11584), .ZN(n11586) );
  AOI222_X1 U13446 ( .A1(n16019), .A2(n11586), .B1(n14766), .B2(n14914), .C1(
        n14768), .C2(n15925), .ZN(n12228) );
  OAI21_X1 U13447 ( .B1(n12280), .B2(n11825), .A(n12293), .ZN(n12222) );
  INV_X1 U13448 ( .A(n12222), .ZN(n11587) );
  AOI22_X1 U13449 ( .A1(n11587), .A2(n16012), .B1(n14566), .B2(n16009), .ZN(
        n11588) );
  OAI211_X1 U13450 ( .C1(n16015), .C2(n11589), .A(n12228), .B(n11588), .ZN(
        n11791) );
  NAND2_X1 U13451 ( .A1(n11791), .A2(n15984), .ZN(n11590) );
  OAI21_X1 U13452 ( .B1(n15984), .B2(n8583), .A(n11590), .ZN(P1_U3468) );
  INV_X1 U13453 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11591) );
  OAI22_X1 U13454 ( .A1(n13864), .A2(n11592), .B1(n16169), .B2(n11591), .ZN(
        n11593) );
  AOI21_X1 U13455 ( .B1(n11666), .B2(n16169), .A(n11593), .ZN(n11594) );
  INV_X1 U13456 ( .A(n11594), .ZN(P3_U3390) );
  NAND2_X1 U13457 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n15450) );
  OAI21_X1 U13458 ( .B1(n13931), .B2(n12042), .A(n15450), .ZN(n11596) );
  INV_X1 U13459 ( .A(n14024), .ZN(n11944) );
  OAI22_X1 U13460 ( .A1(n11680), .A2(n13992), .B1(n13996), .B2(n11944), .ZN(
        n11595) );
  AOI211_X1 U13461 ( .C1(n13176), .C2(n13999), .A(n11596), .B(n11595), .ZN(
        n11604) );
  NAND3_X1 U13462 ( .A1(n13968), .A2(n11597), .A3(n14026), .ZN(n11598) );
  OAI21_X1 U13463 ( .B1(n14001), .B2(n11599), .A(n11598), .ZN(n11602) );
  INV_X1 U13464 ( .A(n11600), .ZN(n11601) );
  NAND2_X1 U13465 ( .A1(n11602), .A2(n11601), .ZN(n11603) );
  OAI211_X1 U13466 ( .C1(n14001), .C2(n11484), .A(n11604), .B(n11603), .ZN(
        P2_U3202) );
  XOR2_X1 U13467 ( .A(n11606), .B(n11605), .Z(n11609) );
  AOI22_X1 U13468 ( .A1(n7185), .A2(n15917), .B1(n11744), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U13469 ( .A1(n14699), .A2(n14768), .B1(n14714), .B2(n15924), .ZN(
        n11607) );
  OAI211_X1 U13470 ( .C1(n11609), .C2(n14740), .A(n11608), .B(n11607), .ZN(
        P1_U3222) );
  INV_X1 U13471 ( .A(n11610), .ZN(n11611) );
  AOI21_X1 U13472 ( .B1(n11613), .B2(n11612), .A(n11611), .ZN(n11624) );
  XNOR2_X1 U13473 ( .A(n11614), .B(n11908), .ZN(n11622) );
  OAI21_X1 U13474 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11616), .A(n11615), .ZN(
        n11617) );
  NAND2_X1 U13475 ( .A1(n11617), .A2(n15844), .ZN(n11619) );
  INV_X1 U13476 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15263) );
  NOR2_X1 U13477 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15263), .ZN(n12027) );
  AOI21_X1 U13478 ( .B1(n15832), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12027), .ZN(
        n11618) );
  OAI211_X1 U13479 ( .C1(n15822), .C2(n11620), .A(n11619), .B(n11618), .ZN(
        n11621) );
  AOI21_X1 U13480 ( .B1(n15845), .B2(n11622), .A(n11621), .ZN(n11623) );
  OAI21_X1 U13481 ( .B1(n11624), .B2(n15840), .A(n11623), .ZN(P3_U3189) );
  INV_X1 U13482 ( .A(n11625), .ZN(n11626) );
  AOI21_X1 U13483 ( .B1(n11628), .B2(n11627), .A(n11626), .ZN(n12164) );
  AOI21_X1 U13484 ( .B1(n11629), .B2(n7677), .A(n16134), .ZN(n11631) );
  NAND2_X1 U13485 ( .A1(n15925), .A2(n14766), .ZN(n11630) );
  OAI21_X1 U13486 ( .B1(n12097), .B2(n15916), .A(n11630), .ZN(n11921) );
  AOI21_X1 U13487 ( .B1(n11631), .B2(n7202), .A(n11921), .ZN(n12161) );
  INV_X1 U13488 ( .A(n12295), .ZN(n11633) );
  INV_X1 U13489 ( .A(n11632), .ZN(n11801) );
  AOI211_X1 U13490 ( .C1(n12159), .C2(n11633), .A(n16077), .B(n11801), .ZN(
        n12155) );
  AOI21_X1 U13491 ( .B1(n12159), .B2(n16009), .A(n12155), .ZN(n11634) );
  OAI211_X1 U13492 ( .C1(n12164), .C2(n16015), .A(n12161), .B(n11634), .ZN(
        n11794) );
  NAND2_X1 U13493 ( .A1(n11794), .A2(n15984), .ZN(n11635) );
  OAI21_X1 U13494 ( .B1(n15984), .B2(n8625), .A(n11635), .ZN(P1_U3474) );
  INV_X1 U13495 ( .A(n16043), .ZN(n11646) );
  AOI21_X1 U13496 ( .B1(n11637), .B2(n11636), .A(n14001), .ZN(n11639) );
  NAND2_X1 U13497 ( .A1(n11639), .A2(n11638), .ZN(n11645) );
  INV_X1 U13498 ( .A(n13984), .ZN(n12603) );
  NAND2_X1 U13499 ( .A1(n14022), .A2(n14091), .ZN(n11641) );
  NAND2_X1 U13500 ( .A1(n14024), .A2(n14089), .ZN(n11640) );
  NAND2_X1 U13501 ( .A1(n11641), .A2(n11640), .ZN(n11948) );
  OAI21_X1 U13502 ( .B1(n13931), .B2(n16039), .A(n11642), .ZN(n11643) );
  AOI21_X1 U13503 ( .B1(n12603), .B2(n11948), .A(n11643), .ZN(n11644) );
  OAI211_X1 U13504 ( .C1(n11646), .C2(n13978), .A(n11645), .B(n11644), .ZN(
        P2_U3211) );
  INV_X1 U13505 ( .A(n11887), .ZN(n11656) );
  XNOR2_X1 U13506 ( .A(n16022), .B(n13119), .ZN(n11988) );
  XNOR2_X1 U13507 ( .A(n13584), .B(n11988), .ZN(n11651) );
  INV_X1 U13508 ( .A(n11647), .ZN(n11648) );
  NAND2_X1 U13509 ( .A1(n11650), .A2(n11651), .ZN(n11990) );
  OAI21_X1 U13510 ( .B1(n11651), .B2(n11650), .A(n11990), .ZN(n11652) );
  NAND2_X1 U13511 ( .A1(n11652), .A2(n13476), .ZN(n11655) );
  NOR2_X1 U13512 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9158), .ZN(n15668) );
  OAI22_X1 U13513 ( .A1(n11886), .A2(n13559), .B1(n12025), .B2(n13551), .ZN(
        n11653) );
  AOI211_X1 U13514 ( .C1(n12504), .C2(n16022), .A(n15668), .B(n11653), .ZN(
        n11654) );
  OAI211_X1 U13515 ( .C1(n11656), .C2(n12382), .A(n11655), .B(n11654), .ZN(
        P3_U3167) );
  NAND2_X1 U13516 ( .A1(n11659), .A2(n11662), .ZN(n11661) );
  NAND2_X1 U13517 ( .A1(n11666), .A2(n13715), .ZN(n11671) );
  INV_X1 U13518 ( .A(n11667), .ZN(n11668) );
  NOR2_X1 U13519 ( .A1(n11879), .A2(n16157), .ZN(n15966) );
  INV_X1 U13520 ( .A(n13754), .ZN(n13696) );
  AOI22_X1 U13521 ( .A1(n13696), .A2(n11669), .B1(n15909), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11670) );
  OAI211_X1 U13522 ( .C1(n11672), .C2(n13715), .A(n11671), .B(n11670), .ZN(
        P3_U3233) );
  INV_X1 U13523 ( .A(n14027), .ZN(n11707) );
  NAND2_X1 U13524 ( .A1(n11707), .A2(n11673), .ZN(n11674) );
  NAND2_X1 U13525 ( .A1(n11675), .A2(n11674), .ZN(n11714) );
  NAND2_X1 U13526 ( .A1(n11714), .A2(n13405), .ZN(n11716) );
  NAND2_X1 U13527 ( .A1(n11680), .A2(n15995), .ZN(n11676) );
  XNOR2_X1 U13528 ( .A(n13176), .B(n14025), .ZN(n13407) );
  INV_X1 U13529 ( .A(n13407), .ZN(n11683) );
  OAI21_X1 U13530 ( .B1(n11677), .B2(n11683), .A(n11771), .ZN(n12049) );
  INV_X1 U13531 ( .A(n12049), .ZN(n11689) );
  OAI22_X1 U13532 ( .A1(n11680), .A2(n14189), .B1(n11944), .B2(n14191), .ZN(
        n11686) );
  NAND2_X1 U13533 ( .A1(n11707), .A2(n14248), .ZN(n11723) );
  NAND2_X1 U13534 ( .A1(n11724), .A2(n11723), .ZN(n11679) );
  INV_X1 U13535 ( .A(n13405), .ZN(n11678) );
  NAND2_X1 U13536 ( .A1(n11679), .A2(n11678), .ZN(n11722) );
  NAND2_X1 U13537 ( .A1(n11680), .A2(n13168), .ZN(n11682) );
  NAND2_X1 U13538 ( .A1(n11722), .A2(n11682), .ZN(n11681) );
  NAND2_X1 U13539 ( .A1(n11681), .A2(n13407), .ZN(n11775) );
  NAND3_X1 U13540 ( .A1(n11722), .A2(n11683), .A3(n11682), .ZN(n11684) );
  AOI21_X1 U13541 ( .B1(n11775), .B2(n11684), .A(n14214), .ZN(n11685) );
  AOI211_X1 U13542 ( .C1(n12049), .C2(n14121), .A(n11686), .B(n11685), .ZN(
        n12051) );
  INV_X1 U13543 ( .A(n11687), .ZN(n11719) );
  INV_X1 U13544 ( .A(n13176), .ZN(n12047) );
  NAND2_X1 U13545 ( .A1(n11687), .A2(n12047), .ZN(n11784) );
  INV_X1 U13546 ( .A(n11784), .ZN(n11785) );
  AOI211_X1 U13547 ( .C1(n13176), .C2(n11719), .A(n14319), .B(n11785), .ZN(
        n12044) );
  AOI21_X1 U13548 ( .B1(n14343), .B2(n13176), .A(n12044), .ZN(n11688) );
  OAI211_X1 U13549 ( .C1(n11689), .C2(n15897), .A(n12051), .B(n11688), .ZN(
        n11691) );
  NAND2_X1 U13550 ( .A1(n11691), .A2(n16192), .ZN(n11690) );
  OAI21_X1 U13551 ( .B1(n16192), .B2(n10503), .A(n11690), .ZN(P2_U3442) );
  NAND2_X1 U13552 ( .A1(n11691), .A2(n16189), .ZN(n11692) );
  OAI21_X1 U13553 ( .B1(n16189), .B2(n11063), .A(n11692), .ZN(P2_U3503) );
  NAND2_X1 U13554 ( .A1(n13404), .A2(n11452), .ZN(n11693) );
  AND2_X1 U13555 ( .A1(n11694), .A2(n11693), .ZN(n15946) );
  INV_X1 U13556 ( .A(n11695), .ZN(n11783) );
  AND2_X1 U13557 ( .A1(n15408), .A2(n11696), .ZN(n11697) );
  NAND2_X1 U13558 ( .A1(n11783), .A2(n11697), .ZN(n11700) );
  AOI21_X1 U13559 ( .B1(n13135), .B2(n13143), .A(n14319), .ZN(n11702) );
  NAND2_X1 U13560 ( .A1(n11702), .A2(n11701), .ZN(n15947) );
  OAI22_X1 U13561 ( .A1(n16045), .A2(n15947), .B1(n11703), .B2(n16038), .ZN(
        n11704) );
  AOI21_X1 U13562 ( .B1(n16147), .B2(n13143), .A(n11704), .ZN(n11713) );
  OAI21_X1 U13563 ( .B1(n11706), .B2(n13404), .A(n11705), .ZN(n11710) );
  OAI22_X1 U13564 ( .A1(n13133), .A2(n14189), .B1(n11707), .B2(n14191), .ZN(
        n11709) );
  NOR2_X1 U13565 ( .A1(n15946), .A2(n14197), .ZN(n11708) );
  AOI211_X1 U13566 ( .C1(n14236), .C2(n11710), .A(n11709), .B(n11708), .ZN(
        n15949) );
  MUX2_X1 U13567 ( .A(n11711), .B(n15949), .S(n16041), .Z(n11712) );
  OAI211_X1 U13568 ( .C1(n15946), .C2(n12713), .A(n11713), .B(n11712), .ZN(
        P2_U3264) );
  OR2_X1 U13569 ( .A1(n11714), .A2(n13405), .ZN(n11715) );
  OAI22_X1 U13570 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n16038), .B1(n16041), 
        .B2(n11048), .ZN(n11721) );
  AOI21_X1 U13571 ( .B1(n11717), .B2(n13168), .A(n14319), .ZN(n11718) );
  NAND2_X1 U13572 ( .A1(n11719), .A2(n11718), .ZN(n15994) );
  NOR2_X1 U13573 ( .A1(n16045), .A2(n15994), .ZN(n11720) );
  AOI211_X1 U13574 ( .C1(n16147), .C2(n13168), .A(n11721), .B(n11720), .ZN(
        n11730) );
  AOI22_X1 U13575 ( .A1(n14091), .A2(n14025), .B1(n14027), .B2(n14089), .ZN(
        n11728) );
  INV_X1 U13576 ( .A(n11722), .ZN(n11726) );
  AND3_X1 U13577 ( .A1(n11724), .A2(n13405), .A3(n11723), .ZN(n11725) );
  OAI21_X1 U13578 ( .B1(n11726), .B2(n11725), .A(n14236), .ZN(n11727) );
  OAI211_X1 U13579 ( .C1(n15993), .C2(n14197), .A(n11728), .B(n11727), .ZN(
        n15996) );
  NAND2_X1 U13580 ( .A1(n15996), .A2(n16041), .ZN(n11729) );
  OAI211_X1 U13581 ( .C1(n15993), .C2(n12713), .A(n11730), .B(n11729), .ZN(
        P2_U3262) );
  OAI222_X1 U13582 ( .A1(n13131), .A2(n11733), .B1(P3_U3151), .B2(n11732), 
        .C1(n11731), .C2(n13880), .ZN(P3_U3275) );
  NAND3_X1 U13583 ( .A1(n13968), .A2(n11734), .A3(n14023), .ZN(n11735) );
  OAI21_X1 U13584 ( .B1(n11638), .B2(n14001), .A(n11735), .ZN(n11742) );
  INV_X1 U13585 ( .A(n11736), .ZN(n11741) );
  NAND2_X1 U13586 ( .A1(n13999), .A2(n13195), .ZN(n11738) );
  OAI211_X1 U13587 ( .C1(n13931), .C2(n12185), .A(n11738), .B(n11737), .ZN(
        n11740) );
  OAI22_X1 U13588 ( .A1(n12169), .A2(n13996), .B1(n13992), .B2(n12069), .ZN(
        n11739) );
  AOI211_X1 U13589 ( .C1(n11742), .C2(n11741), .A(n11740), .B(n11739), .ZN(
        n11743) );
  OAI21_X1 U13590 ( .B1(n11868), .B2(n14001), .A(n11743), .ZN(P2_U3185) );
  INV_X1 U13591 ( .A(n11744), .ZN(n11749) );
  INV_X1 U13592 ( .A(n16197), .ZN(n14711) );
  NAND2_X1 U13593 ( .A1(n14914), .A2(n14769), .ZN(n15878) );
  OAI22_X1 U13594 ( .A1(n14711), .A2(n15878), .B1(n14740), .B2(n11745), .ZN(
        n11746) );
  AOI21_X1 U13595 ( .B1(n15914), .B2(n7185), .A(n11746), .ZN(n11747) );
  OAI21_X1 U13596 ( .B1(n11749), .B2(n11748), .A(n11747), .ZN(P1_U3232) );
  INV_X1 U13597 ( .A(n11750), .ZN(n11753) );
  INV_X1 U13598 ( .A(n12426), .ZN(n15467) );
  OAI222_X1 U13599 ( .A1(n14370), .A2(n11751), .B1(n14378), .B2(n11753), .C1(
        n15467), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI222_X1 U13600 ( .A1(P1_U3086), .A2(n15535), .B1(n15160), .B2(n11753), 
        .C1(n11752), .C2(n15157), .ZN(P1_U3340) );
  XOR2_X1 U13601 ( .A(n11755), .B(n11754), .Z(n11769) );
  OAI21_X1 U13602 ( .B1(n11758), .B2(n11757), .A(n11756), .ZN(n11767) );
  NOR2_X1 U13603 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15346), .ZN(n12105) );
  AOI21_X1 U13604 ( .B1(n15832), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12105), .ZN(
        n11759) );
  OAI21_X1 U13605 ( .B1(n15822), .B2(n11760), .A(n11759), .ZN(n11766) );
  AOI21_X1 U13606 ( .B1(n11763), .B2(n11762), .A(n11761), .ZN(n11764) );
  NOR2_X1 U13607 ( .A1(n11764), .A2(n15830), .ZN(n11765) );
  AOI211_X1 U13608 ( .C1(n15844), .C2(n11767), .A(n11766), .B(n11765), .ZN(
        n11768) );
  OAI21_X1 U13609 ( .B1(n11769), .B2(n15840), .A(n11768), .ZN(P3_U3190) );
  OR2_X1 U13610 ( .A1(n13176), .A2(n14025), .ZN(n11770) );
  XNOR2_X1 U13611 ( .A(n13182), .B(n14024), .ZN(n13408) );
  INV_X1 U13612 ( .A(n13408), .ZN(n11776) );
  OR2_X1 U13613 ( .A1(n11772), .A2(n11776), .ZN(n11773) );
  NAND2_X1 U13614 ( .A1(n11939), .A2(n11773), .ZN(n11857) );
  INV_X1 U13615 ( .A(n11857), .ZN(n11790) );
  NAND2_X1 U13616 ( .A1(n13176), .A2(n13178), .ZN(n11774) );
  XNOR2_X1 U13617 ( .A(n11943), .B(n11776), .ZN(n11779) );
  NAND2_X1 U13618 ( .A1(n11857), .A2(n14121), .ZN(n11778) );
  AOI22_X1 U13619 ( .A1(n14089), .A2(n14025), .B1(n14023), .B2(n14091), .ZN(
        n11777) );
  OAI211_X1 U13620 ( .C1(n14214), .C2(n11779), .A(n11778), .B(n11777), .ZN(
        n11855) );
  MUX2_X1 U13621 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11855), .S(n16041), .Z(
        n11780) );
  INV_X1 U13622 ( .A(n11780), .ZN(n11789) );
  AND2_X1 U13623 ( .A1(n15408), .A2(n11781), .ZN(n11782) );
  NAND2_X1 U13624 ( .A1(n11783), .A2(n11782), .ZN(n14206) );
  INV_X1 U13625 ( .A(n13182), .ZN(n11941) );
  OR2_X1 U13626 ( .A1(n11784), .A2(n13182), .ZN(n11949) );
  OAI21_X1 U13627 ( .B1(n11941), .B2(n11785), .A(n11949), .ZN(n11854) );
  OAI22_X1 U13628 ( .A1(n14206), .A2(n11854), .B1(n11786), .B2(n16038), .ZN(
        n11787) );
  AOI21_X1 U13629 ( .B1(n16147), .B2(n13182), .A(n11787), .ZN(n11788) );
  OAI211_X1 U13630 ( .C1(n11790), .C2(n12713), .A(n11789), .B(n11788), .ZN(
        P2_U3260) );
  NAND2_X1 U13631 ( .A1(n11791), .A2(n16141), .ZN(n11792) );
  OAI21_X1 U13632 ( .B1(n16141), .B2(n11793), .A(n11792), .ZN(P1_U3531) );
  INV_X1 U13633 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U13634 ( .A1(n11794), .A2(n16141), .ZN(n11795) );
  OAI21_X1 U13635 ( .B1(n16141), .B2(n11796), .A(n11795), .ZN(P1_U3533) );
  OAI21_X1 U13636 ( .B1(n11799), .B2(n11798), .A(n11797), .ZN(n12443) );
  INV_X1 U13637 ( .A(n12437), .ZN(n12017) );
  INV_X1 U13638 ( .A(n11800), .ZN(n12128) );
  OAI21_X1 U13639 ( .B1(n12017), .B2(n11801), .A(n12128), .ZN(n12439) );
  OAI22_X1 U13640 ( .A1(n12439), .A2(n16077), .B1(n12017), .B2(n16133), .ZN(
        n11808) );
  INV_X1 U13641 ( .A(n12443), .ZN(n11807) );
  AOI22_X1 U13642 ( .A1(n14914), .A2(n14763), .B1(n15925), .B2(n14765), .ZN(
        n11806) );
  OAI211_X1 U13643 ( .C1(n11804), .C2(n11803), .A(n11802), .B(n16019), .ZN(
        n11805) );
  OAI211_X1 U13644 ( .C1(n11807), .C2(n15927), .A(n11806), .B(n11805), .ZN(
        n12440) );
  AOI211_X1 U13645 ( .C1(n7680), .C2(n12443), .A(n11808), .B(n12440), .ZN(
        n11968) );
  NAND2_X1 U13646 ( .A1(n16140), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n11809) );
  OAI21_X1 U13647 ( .B1(n11968), .B2(n16140), .A(n11809), .ZN(P1_U3534) );
  INV_X1 U13648 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11810) );
  MUX2_X1 U13649 ( .A(n11810), .B(P1_REG1_REG_13__SCAN_IN), .S(n12115), .Z(
        n11813) );
  AOI211_X1 U13650 ( .C1(n11813), .C2(n11812), .A(n15859), .B(n12114), .ZN(
        n11824) );
  OAI21_X1 U13651 ( .B1(n11815), .B2(P1_REG2_REG_12__SCAN_IN), .A(n11814), 
        .ZN(n11818) );
  MUX2_X1 U13652 ( .A(n8765), .B(P1_REG2_REG_13__SCAN_IN), .S(n12115), .Z(
        n11817) );
  INV_X1 U13653 ( .A(n15869), .ZN(n15536) );
  INV_X1 U13654 ( .A(n12112), .ZN(n11816) );
  AOI211_X1 U13655 ( .C1(n11818), .C2(n11817), .A(n15536), .B(n11816), .ZN(
        n11823) );
  NAND2_X1 U13656 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14676)
         );
  INV_X1 U13657 ( .A(n14676), .ZN(n11819) );
  AOI21_X1 U13658 ( .B1(n15526), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11819), 
        .ZN(n11820) );
  OAI21_X1 U13659 ( .B1(n15534), .B2(n11821), .A(n11820), .ZN(n11822) );
  OR3_X1 U13660 ( .A1(n11824), .A2(n11823), .A3(n11822), .ZN(P1_U3256) );
  OAI22_X1 U13661 ( .A1(n14586), .A2(n12276), .B1(n11825), .B2(n14588), .ZN(
        n11834) );
  INV_X1 U13662 ( .A(n11834), .ZN(n11836) );
  OAI22_X1 U13663 ( .A1(n14585), .A2(n11825), .B1(n12276), .B2(n14588), .ZN(
        n11826) );
  XNOR2_X1 U13664 ( .A(n11826), .B(n14589), .ZN(n11833) );
  INV_X1 U13665 ( .A(n11833), .ZN(n11835) );
  INV_X1 U13666 ( .A(n11827), .ZN(n11830) );
  INV_X1 U13667 ( .A(n11828), .ZN(n11829) );
  AOI22_X1 U13668 ( .A1(n11832), .A2(n11831), .B1(n11830), .B2(n11829), .ZN(
        n14565) );
  XOR2_X1 U13669 ( .A(n11834), .B(n11833), .Z(n14564) );
  NAND2_X1 U13670 ( .A1(n14565), .A2(n14564), .ZN(n14563) );
  OAI22_X1 U13671 ( .A1(n14586), .A2(n11840), .B1(n12299), .B2(n14588), .ZN(
        n11837) );
  INV_X1 U13672 ( .A(n11913), .ZN(n11839) );
  NAND2_X1 U13673 ( .A1(n11839), .A2(n11911), .ZN(n11842) );
  OAI22_X1 U13674 ( .A1(n14585), .A2(n12299), .B1(n11840), .B2(n14588), .ZN(
        n11841) );
  XOR2_X1 U13675 ( .A(n14589), .B(n11841), .Z(n11912) );
  XNOR2_X1 U13676 ( .A(n11842), .B(n11912), .ZN(n11853) );
  INV_X1 U13677 ( .A(n11843), .ZN(n12296) );
  AND3_X1 U13678 ( .A1(n11846), .A2(n11845), .A3(n11844), .ZN(n11847) );
  NAND2_X1 U13679 ( .A1(n11848), .A2(n11847), .ZN(n11849) );
  INV_X1 U13680 ( .A(n16203), .ZN(n14690) );
  AOI22_X1 U13681 ( .A1(n14699), .A2(n14765), .B1(n14714), .B2(n14767), .ZN(
        n11850) );
  NAND2_X1 U13682 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15873) );
  OAI211_X1 U13683 ( .C1(n12299), .C2(n14717), .A(n11850), .B(n15873), .ZN(
        n11851) );
  AOI21_X1 U13684 ( .B1(n12296), .B2(n14690), .A(n11851), .ZN(n11852) );
  OAI21_X1 U13685 ( .B1(n11853), .B2(n14740), .A(n11852), .ZN(P1_U3230) );
  OAI22_X1 U13686 ( .A1(n11854), .A2(n14319), .B1(n11941), .B2(n16182), .ZN(
        n11856) );
  AOI211_X1 U13687 ( .C1(n16121), .C2(n11857), .A(n11856), .B(n11855), .ZN(
        n11863) );
  OR2_X1 U13688 ( .A1(n11863), .A2(n16190), .ZN(n11858) );
  OAI21_X1 U13689 ( .B1(n16192), .B2(n10576), .A(n11858), .ZN(P2_U3445) );
  INV_X1 U13690 ( .A(n15481), .ZN(n12429) );
  INV_X1 U13691 ( .A(n11859), .ZN(n11862) );
  OAI222_X1 U13692 ( .A1(P2_U3088), .A2(n12429), .B1(n14378), .B2(n11862), 
        .C1(n11860), .C2(n14370), .ZN(P2_U3311) );
  OAI222_X1 U13693 ( .A1(P1_U3086), .A2(n12874), .B1(n15160), .B2(n11862), 
        .C1(n11861), .C2(n15157), .ZN(P1_U3339) );
  OR2_X1 U13694 ( .A1(n11863), .A2(n16188), .ZN(n11864) );
  OAI21_X1 U13695 ( .B1(n16189), .B2(n11065), .A(n11864), .ZN(P2_U3504) );
  INV_X1 U13696 ( .A(n13202), .ZN(n12305) );
  INV_X1 U13697 ( .A(n14022), .ZN(n13197) );
  OAI22_X1 U13698 ( .A1(n13897), .A2(n13197), .B1(n11865), .B2(n14001), .ZN(
        n11866) );
  NAND3_X1 U13699 ( .A1(n11868), .A2(n11867), .A3(n11866), .ZN(n11875) );
  OR2_X1 U13700 ( .A1(n13996), .A2(n13212), .ZN(n11872) );
  INV_X1 U13701 ( .A(n12083), .ZN(n11870) );
  AOI21_X1 U13702 ( .B1(n13994), .B2(n11870), .A(n11869), .ZN(n11871) );
  OAI211_X1 U13703 ( .C1(n13197), .C2(n13992), .A(n11872), .B(n11871), .ZN(
        n11873) );
  INV_X1 U13704 ( .A(n11873), .ZN(n11874) );
  OAI211_X1 U13705 ( .C1(n12305), .C2(n13978), .A(n11875), .B(n11874), .ZN(
        n11876) );
  AOI21_X1 U13706 ( .B1(n11980), .B2(n13940), .A(n11876), .ZN(n11877) );
  INV_X1 U13707 ( .A(n11877), .ZN(P2_U3193) );
  AND2_X1 U13708 ( .A1(n11879), .A2(n11878), .ZN(n12230) );
  OR2_X1 U13709 ( .A1(n16057), .A2(n12230), .ZN(n15974) );
  XOR2_X1 U13710 ( .A(n11880), .B(n11884), .Z(n16024) );
  INV_X1 U13711 ( .A(n11881), .ZN(n11882) );
  AOI21_X1 U13712 ( .B1(n11884), .B2(n11883), .A(n11882), .ZN(n11885) );
  OAI222_X1 U13713 ( .A1(n15960), .A2(n11886), .B1(n15962), .B2(n12025), .C1(
        n15959), .C2(n11885), .ZN(n16021) );
  AOI22_X1 U13714 ( .A1(n13696), .A2(n16022), .B1(n15909), .B2(n11887), .ZN(
        n11888) );
  OAI21_X1 U13715 ( .B1(n15660), .B2(n13715), .A(n11888), .ZN(n11889) );
  AOI21_X1 U13716 ( .B1(n16021), .B2(n13715), .A(n11889), .ZN(n11890) );
  OAI21_X1 U13717 ( .B1(n13717), .B2(n16024), .A(n11890), .ZN(P3_U3228) );
  XNOR2_X1 U13718 ( .A(n11891), .B(n11893), .ZN(n16003) );
  OAI211_X1 U13719 ( .C1(n11894), .C2(n11893), .A(n11892), .B(n13705), .ZN(
        n11896) );
  OR2_X1 U13720 ( .A1(n15961), .A2(n15960), .ZN(n11895) );
  OAI211_X1 U13721 ( .C1(n11994), .C2(n15962), .A(n11896), .B(n11895), .ZN(
        n16000) );
  AOI22_X1 U13722 ( .A1(n13696), .A2(n16001), .B1(n15909), .B2(n11897), .ZN(
        n11898) );
  OAI21_X1 U13723 ( .B1(n9986), .B2(n13715), .A(n11898), .ZN(n11899) );
  AOI21_X1 U13724 ( .B1(n16000), .B2(n13715), .A(n11899), .ZN(n11900) );
  OAI21_X1 U13725 ( .B1(n13717), .B2(n16003), .A(n11900), .ZN(P3_U3229) );
  XNOR2_X1 U13726 ( .A(n11901), .B(n11903), .ZN(n16054) );
  OAI211_X1 U13727 ( .C1(n11904), .C2(n11903), .A(n11902), .B(n13705), .ZN(
        n11906) );
  AOI22_X1 U13728 ( .A1(n13583), .A2(n13708), .B1(n9880), .B2(n13581), .ZN(
        n11905) );
  NAND2_X1 U13729 ( .A1(n11906), .A2(n11905), .ZN(n16051) );
  AOI22_X1 U13730 ( .A1(n13696), .A2(n16052), .B1(n15909), .B2(n12028), .ZN(
        n11907) );
  OAI21_X1 U13731 ( .B1(n11908), .B2(n13715), .A(n11907), .ZN(n11909) );
  AOI21_X1 U13732 ( .B1(n16051), .B2(n13715), .A(n11909), .ZN(n11910) );
  OAI21_X1 U13733 ( .B1(n13717), .B2(n16054), .A(n11910), .ZN(P3_U3226) );
  NAND2_X1 U13734 ( .A1(n12159), .A2(n14526), .ZN(n11915) );
  NAND2_X1 U13735 ( .A1(n11917), .A2(n14765), .ZN(n11914) );
  NAND2_X1 U13736 ( .A1(n11915), .A2(n11914), .ZN(n11916) );
  XNOR2_X1 U13737 ( .A(n11916), .B(n14589), .ZN(n12004) );
  NAND2_X1 U13738 ( .A1(n12159), .A2(n11917), .ZN(n11918) );
  OAI21_X1 U13739 ( .B1(n14586), .B2(n12292), .A(n11918), .ZN(n12003) );
  XNOR2_X1 U13740 ( .A(n12004), .B(n12003), .ZN(n11919) );
  XNOR2_X1 U13741 ( .A(n12005), .B(n11919), .ZN(n11925) );
  AOI21_X1 U13742 ( .B1(n16197), .B2(n11921), .A(n11920), .ZN(n11923) );
  NAND2_X1 U13743 ( .A1(n7185), .A2(n12159), .ZN(n11922) );
  OAI211_X1 U13744 ( .C1(n16203), .C2(n12156), .A(n11923), .B(n11922), .ZN(
        n11924) );
  AOI21_X1 U13745 ( .B1(n11925), .B2(n16195), .A(n11924), .ZN(n11926) );
  INV_X1 U13746 ( .A(n11926), .ZN(P1_U3227) );
  XNOR2_X1 U13747 ( .A(n11927), .B(n11929), .ZN(n16030) );
  INV_X1 U13748 ( .A(n11928), .ZN(n11932) );
  AOI21_X1 U13749 ( .B1(n11881), .B2(n11930), .A(n11929), .ZN(n11931) );
  NOR3_X1 U13750 ( .A1(n11932), .A2(n11931), .A3(n15959), .ZN(n11934) );
  OAI22_X1 U13751 ( .A1(n12214), .A2(n15962), .B1(n11994), .B2(n15960), .ZN(
        n11933) );
  NOR2_X1 U13752 ( .A1(n11934), .A2(n11933), .ZN(n16031) );
  MUX2_X1 U13753 ( .A(n11935), .B(n16031), .S(n13715), .Z(n11937) );
  AOI22_X1 U13754 ( .A1(n13696), .A2(n11996), .B1(n15909), .B2(n11987), .ZN(
        n11936) );
  OAI211_X1 U13755 ( .C1(n13717), .C2(n16030), .A(n11937), .B(n11936), .ZN(
        P3_U3227) );
  INV_X1 U13756 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11953) );
  NAND2_X1 U13757 ( .A1(n11941), .A2(n11944), .ZN(n11938) );
  NAND2_X1 U13758 ( .A1(n11939), .A2(n11938), .ZN(n11940) );
  XNOR2_X1 U13759 ( .A(n16043), .B(n14023), .ZN(n13410) );
  NAND2_X1 U13760 ( .A1(n11940), .A2(n11945), .ZN(n12077) );
  OAI21_X1 U13761 ( .B1(n11940), .B2(n11945), .A(n12077), .ZN(n16048) );
  INV_X1 U13762 ( .A(n16048), .ZN(n11951) );
  NAND2_X1 U13763 ( .A1(n11941), .A2(n14024), .ZN(n11942) );
  XNOR2_X1 U13764 ( .A(n12068), .B(n11945), .ZN(n11946) );
  NOR2_X1 U13765 ( .A1(n11946), .A2(n14214), .ZN(n11947) );
  AOI211_X1 U13766 ( .C1(n14121), .C2(n16048), .A(n11948), .B(n11947), .ZN(
        n16050) );
  AOI211_X1 U13767 ( .C1(n16043), .C2(n11949), .A(n14319), .B(n12184), .ZN(
        n16037) );
  AOI21_X1 U13768 ( .B1(n14343), .B2(n16043), .A(n16037), .ZN(n11950) );
  OAI211_X1 U13769 ( .C1(n11951), .C2(n15897), .A(n16050), .B(n11950), .ZN(
        n11954) );
  NAND2_X1 U13770 ( .A1(n11954), .A2(n16192), .ZN(n11952) );
  OAI21_X1 U13771 ( .B1(n16192), .B2(n11953), .A(n11952), .ZN(P2_U3448) );
  NAND2_X1 U13772 ( .A1(n11954), .A2(n16189), .ZN(n11955) );
  OAI21_X1 U13773 ( .B1(n16189), .B2(n10591), .A(n11955), .ZN(P2_U3505) );
  XOR2_X1 U13774 ( .A(n11956), .B(n11957), .Z(n15988) );
  AOI22_X1 U13775 ( .A1(n13696), .A2(n15986), .B1(n15909), .B2(n15343), .ZN(
        n11965) );
  NAND2_X1 U13776 ( .A1(n11958), .A2(n11957), .ZN(n11959) );
  NAND3_X1 U13777 ( .A1(n11960), .A2(n13705), .A3(n11959), .ZN(n11962) );
  AOI22_X1 U13778 ( .A1(n13587), .A2(n13708), .B1(n9880), .B2(n13585), .ZN(
        n11961) );
  NAND2_X1 U13779 ( .A1(n11962), .A2(n11961), .ZN(n15985) );
  MUX2_X1 U13780 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n15985), .S(n13715), .Z(
        n11963) );
  INV_X1 U13781 ( .A(n11963), .ZN(n11964) );
  OAI211_X1 U13782 ( .C1(n15988), .C2(n13717), .A(n11965), .B(n11964), .ZN(
        P3_U3230) );
  OAI222_X1 U13783 ( .A1(n11967), .A2(P3_U3151), .B1(n13880), .B2(n15189), 
        .C1(n13131), .C2(n11966), .ZN(P3_U3274) );
  OR2_X1 U13784 ( .A1(n11968), .A2(n16142), .ZN(n11969) );
  OAI21_X1 U13785 ( .B1(n15984), .B2(n8642), .A(n11969), .ZN(P1_U3477) );
  INV_X1 U13786 ( .A(n14814), .ZN(n14811) );
  INV_X1 U13787 ( .A(n11970), .ZN(n11972) );
  OAI222_X1 U13788 ( .A1(n14811), .A2(P1_U3086), .B1(n15160), .B2(n11972), 
        .C1(n11971), .C2(n15157), .ZN(P1_U3338) );
  INV_X1 U13789 ( .A(n12720), .ZN(n12435) );
  OAI222_X1 U13790 ( .A1(n14370), .A2(n11973), .B1(n14378), .B2(n11972), .C1(
        P2_U3088), .C2(n12435), .ZN(P2_U3310) );
  INV_X1 U13791 ( .A(n11974), .ZN(n12146) );
  INV_X1 U13792 ( .A(n14019), .ZN(n12537) );
  OR2_X1 U13793 ( .A1(n13992), .A2(n12169), .ZN(n11978) );
  INV_X1 U13794 ( .A(n12173), .ZN(n11976) );
  AOI21_X1 U13795 ( .B1(n13994), .B2(n11976), .A(n11975), .ZN(n11977) );
  OAI211_X1 U13796 ( .C1(n12537), .C2(n13996), .A(n11978), .B(n11977), .ZN(
        n11979) );
  AOI21_X1 U13797 ( .B1(n13210), .B2(n13999), .A(n11979), .ZN(n11986) );
  INV_X1 U13798 ( .A(n11980), .ZN(n11984) );
  OAI22_X1 U13799 ( .A1(n13897), .A2(n12169), .B1(n11981), .B2(n14001), .ZN(
        n11982) );
  NAND3_X1 U13800 ( .A1(n11984), .A2(n11983), .A3(n11982), .ZN(n11985) );
  OAI211_X1 U13801 ( .C1(n12146), .C2(n14001), .A(n11986), .B(n11985), .ZN(
        P2_U3203) );
  INV_X1 U13802 ( .A(n11987), .ZN(n11999) );
  XNOR2_X1 U13803 ( .A(n11996), .B(n13119), .ZN(n12021) );
  XNOR2_X1 U13804 ( .A(n12025), .B(n12021), .ZN(n11992) );
  AOI211_X1 U13805 ( .C1(n11992), .C2(n11991), .A(n13566), .B(n12022), .ZN(
        n11993) );
  INV_X1 U13806 ( .A(n11993), .ZN(n11998) );
  INV_X1 U13807 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15165) );
  NOR2_X1 U13808 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15165), .ZN(n15686) );
  OAI22_X1 U13809 ( .A1(n11994), .A2(n13559), .B1(n12214), .B2(n13551), .ZN(
        n11995) );
  AOI211_X1 U13810 ( .C1(n12504), .C2(n11996), .A(n15686), .B(n11995), .ZN(
        n11997) );
  OAI211_X1 U13811 ( .C1(n11999), .C2(n12382), .A(n11998), .B(n11997), .ZN(
        P3_U3179) );
  OAI22_X1 U13812 ( .A1(n12000), .A2(P3_U3151), .B1(SI_22_), .B2(n13880), .ZN(
        n12001) );
  AOI21_X1 U13813 ( .B1(n12002), .B2(n13876), .A(n12001), .ZN(P3_U3273) );
  NAND2_X1 U13814 ( .A1(n12437), .A2(n14526), .ZN(n12007) );
  NAND2_X1 U13815 ( .A1(n11917), .A2(n14764), .ZN(n12006) );
  NAND2_X1 U13816 ( .A1(n12007), .A2(n12006), .ZN(n12008) );
  XNOR2_X1 U13817 ( .A(n12008), .B(n14589), .ZN(n12012) );
  NAND2_X1 U13818 ( .A1(n12437), .A2(n14533), .ZN(n12010) );
  NAND2_X1 U13819 ( .A1(n14480), .A2(n14764), .ZN(n12009) );
  NAND2_X1 U13820 ( .A1(n12010), .A2(n12009), .ZN(n12011) );
  NAND2_X1 U13821 ( .A1(n12012), .A2(n12011), .ZN(n12090) );
  NAND2_X1 U13822 ( .A1(n7400), .A2(n12090), .ZN(n12013) );
  XNOR2_X1 U13823 ( .A(n12091), .B(n12013), .ZN(n12020) );
  INV_X1 U13824 ( .A(n12014), .ZN(n12436) );
  AOI22_X1 U13825 ( .A1(n14699), .A2(n14763), .B1(n14714), .B2(n14765), .ZN(
        n12016) );
  OAI211_X1 U13826 ( .C1(n12017), .C2(n14717), .A(n12016), .B(n12015), .ZN(
        n12018) );
  AOI21_X1 U13827 ( .B1(n12436), .B2(n14690), .A(n12018), .ZN(n12019) );
  OAI21_X1 U13828 ( .B1(n12020), .B2(n14740), .A(n12019), .ZN(P1_U3239) );
  INV_X1 U13829 ( .A(n12021), .ZN(n12023) );
  XNOR2_X1 U13830 ( .A(n12024), .B(n13119), .ZN(n12102) );
  XNOR2_X1 U13831 ( .A(n12102), .B(n13582), .ZN(n12103) );
  XNOR2_X1 U13832 ( .A(n7337), .B(n12103), .ZN(n12031) );
  OAI22_X1 U13833 ( .A1(n12025), .A2(n13559), .B1(n12376), .B2(n13551), .ZN(
        n12026) );
  AOI211_X1 U13834 ( .C1(n12504), .C2(n16052), .A(n12027), .B(n12026), .ZN(
        n12030) );
  NAND2_X1 U13835 ( .A1(n13564), .A2(n12028), .ZN(n12029) );
  OAI211_X1 U13836 ( .C1(n12031), .C2(n13566), .A(n12030), .B(n12029), .ZN(
        P3_U3153) );
  NAND2_X1 U13837 ( .A1(n13589), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n12032) );
  OAI21_X1 U13838 ( .B1(n12033), .B2(n13589), .A(n12032), .ZN(P3_U3521) );
  NAND2_X1 U13839 ( .A1(n13589), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n12034) );
  OAI21_X1 U13840 ( .B1(n13610), .B2(n13589), .A(n12034), .ZN(P3_U3520) );
  NAND2_X1 U13841 ( .A1(n13589), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(n12035) );
  OAI21_X1 U13842 ( .B1(n13593), .B2(n13589), .A(n12035), .ZN(P3_U3522) );
  XNOR2_X1 U13843 ( .A(n13138), .B(n13135), .ZN(n15898) );
  INV_X1 U13844 ( .A(n16038), .ZN(n16146) );
  NOR2_X1 U13845 ( .A1(n14121), .A2(n14236), .ZN(n12037) );
  OAI22_X1 U13846 ( .A1(n12037), .A2(n15898), .B1(n12036), .B2(n14191), .ZN(
        n15900) );
  AOI21_X1 U13847 ( .B1(n16146), .B2(P2_REG3_REG_0__SCAN_IN), .A(n15900), .ZN(
        n12038) );
  NOR2_X1 U13848 ( .A1(n16156), .A2(n12038), .ZN(n12039) );
  AOI21_X1 U13849 ( .B1(n16156), .B2(P2_REG2_REG_0__SCAN_IN), .A(n12039), .ZN(
        n12041) );
  INV_X1 U13850 ( .A(n14206), .ZN(n14159) );
  OAI21_X1 U13851 ( .B1(n16147), .B2(n14159), .A(n13135), .ZN(n12040) );
  OAI211_X1 U13852 ( .C1(n15898), .C2(n12713), .A(n12041), .B(n12040), .ZN(
        P2_U3265) );
  INV_X1 U13853 ( .A(n12713), .ZN(n16151) );
  INV_X1 U13854 ( .A(n12042), .ZN(n12043) );
  AOI22_X1 U13855 ( .A1(n16150), .A2(n12044), .B1(n12043), .B2(n16146), .ZN(
        n12046) );
  NAND2_X1 U13856 ( .A1(n16156), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n12045) );
  OAI211_X1 U13857 ( .C1(n14231), .C2(n12047), .A(n12046), .B(n12045), .ZN(
        n12048) );
  AOI21_X1 U13858 ( .B1(n16151), .B2(n12049), .A(n12048), .ZN(n12050) );
  OAI21_X1 U13859 ( .B1(n16156), .B2(n12051), .A(n12050), .ZN(P2_U3261) );
  AOI21_X1 U13860 ( .B1(n12054), .B2(n12053), .A(n12052), .ZN(n12067) );
  OAI21_X1 U13861 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n12056), .A(n12055), .ZN(
        n12065) );
  NOR2_X1 U13862 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9231), .ZN(n12378) );
  AOI21_X1 U13863 ( .B1(n15832), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12378), .ZN(
        n12057) );
  OAI21_X1 U13864 ( .B1(n15822), .B2(n12058), .A(n12057), .ZN(n12064) );
  INV_X1 U13865 ( .A(n12059), .ZN(n12060) );
  AOI211_X1 U13866 ( .C1(n12062), .C2(n12061), .A(n15840), .B(n12060), .ZN(
        n12063) );
  AOI211_X1 U13867 ( .C1(n15844), .C2(n12065), .A(n12064), .B(n12063), .ZN(
        n12066) );
  OAI21_X1 U13868 ( .B1(n12067), .B2(n15830), .A(n12066), .ZN(P3_U3191) );
  NAND2_X1 U13869 ( .A1(n16043), .A2(n12069), .ZN(n12070) );
  NAND2_X1 U13870 ( .A1(n12071), .A2(n12070), .ZN(n12188) );
  AND2_X1 U13871 ( .A1(n13195), .A2(n13197), .ZN(n12073) );
  OR2_X1 U13872 ( .A1(n13195), .A2(n13197), .ZN(n12072) );
  NAND2_X1 U13873 ( .A1(n13202), .A2(n12169), .ZN(n12167) );
  OR2_X1 U13874 ( .A1(n13202), .A2(n12169), .ZN(n12074) );
  NAND2_X1 U13875 ( .A1(n12167), .A2(n12074), .ZN(n13413) );
  INV_X1 U13876 ( .A(n13413), .ZN(n12081) );
  OAI21_X1 U13877 ( .B1(n7339), .B2(n12081), .A(n12168), .ZN(n12075) );
  AOI222_X1 U13878 ( .A1(n14236), .A2(n12075), .B1(n14022), .B2(n14089), .C1(
        n14020), .C2(n14091), .ZN(n12304) );
  INV_X1 U13879 ( .A(n13195), .ZN(n16063) );
  OAI211_X1 U13880 ( .C1(n12305), .C2(n12182), .A(n14302), .B(n12175), .ZN(
        n12303) );
  OR2_X1 U13881 ( .A1(n16043), .A2(n14023), .ZN(n12076) );
  XNOR2_X1 U13882 ( .A(n13195), .B(n13197), .ZN(n13412) );
  OR2_X1 U13883 ( .A1(n13195), .A2(n14022), .ZN(n12078) );
  INV_X1 U13884 ( .A(n12166), .ZN(n12079) );
  AOI21_X1 U13885 ( .B1(n12081), .B2(n12080), .A(n12079), .ZN(n12307) );
  AND2_X1 U13886 ( .A1(n10835), .A2(n13454), .ZN(n12082) );
  NAND2_X1 U13887 ( .A1(n12307), .A2(n14151), .ZN(n12087) );
  OAI22_X1 U13888 ( .A1(n16041), .A2(n12084), .B1(n12083), .B2(n16038), .ZN(
        n12085) );
  AOI21_X1 U13889 ( .B1(n16147), .B2(n13202), .A(n12085), .ZN(n12086) );
  OAI211_X1 U13890 ( .C1(n12303), .C2(n16045), .A(n12087), .B(n12086), .ZN(
        n12088) );
  INV_X1 U13891 ( .A(n12088), .ZN(n12089) );
  OAI21_X1 U13892 ( .B1(n16156), .B2(n12304), .A(n12089), .ZN(P2_U3257) );
  OAI22_X1 U13893 ( .A1(n12240), .A2(n14585), .B1(n12256), .B2(n14588), .ZN(
        n12092) );
  XNOR2_X1 U13894 ( .A(n12092), .B(n14589), .ZN(n12345) );
  NOR2_X1 U13895 ( .A1(n14586), .A2(n12256), .ZN(n12093) );
  AOI21_X1 U13896 ( .B1(n12129), .B2(n14533), .A(n12093), .ZN(n12347) );
  XNOR2_X1 U13897 ( .A(n12345), .B(n12347), .ZN(n12094) );
  OAI211_X1 U13898 ( .C1(n12095), .C2(n12094), .A(n12346), .B(n16195), .ZN(
        n12101) );
  OAI22_X1 U13899 ( .A1(n14717), .A2(n12240), .B1(n16203), .B2(n12241), .ZN(
        n12099) );
  INV_X1 U13900 ( .A(n14714), .ZN(n14697) );
  OAI21_X1 U13901 ( .B1(n14697), .B2(n12097), .A(n12096), .ZN(n12098) );
  AOI211_X1 U13902 ( .C1(n14699), .C2(n14762), .A(n12099), .B(n12098), .ZN(
        n12100) );
  NAND2_X1 U13903 ( .A1(n12101), .A2(n12100), .ZN(P1_U3213) );
  XNOR2_X1 U13904 ( .A(n12106), .B(n13119), .ZN(n12357) );
  XNOR2_X1 U13905 ( .A(n12357), .B(n13581), .ZN(n12359) );
  XNOR2_X1 U13906 ( .A(n12360), .B(n12359), .ZN(n12109) );
  INV_X1 U13907 ( .A(n13580), .ZN(n12362) );
  OAI22_X1 U13908 ( .A1(n12214), .A2(n13559), .B1(n12362), .B2(n13551), .ZN(
        n12104) );
  AOI211_X1 U13909 ( .C1(n12504), .C2(n12106), .A(n12105), .B(n12104), .ZN(
        n12108) );
  NAND2_X1 U13910 ( .A1(n13564), .A2(n12216), .ZN(n12107) );
  OAI211_X1 U13911 ( .C1(n12109), .C2(n13566), .A(n12108), .B(n12107), .ZN(
        P3_U3161) );
  NAND2_X1 U13912 ( .A1(n12115), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n12111) );
  MUX2_X1 U13913 ( .A(n8783), .B(P1_REG2_REG_14__SCAN_IN), .S(n12671), .Z(
        n12110) );
  AOI21_X1 U13914 ( .B1(n12112), .B2(n12111), .A(n12110), .ZN(n12670) );
  NAND3_X1 U13915 ( .A1(n12112), .A2(n12111), .A3(n12110), .ZN(n12113) );
  NAND2_X1 U13916 ( .A1(n12113), .A2(n15869), .ZN(n12122) );
  INV_X1 U13917 ( .A(n12116), .ZN(n12117) );
  INV_X1 U13918 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n12773) );
  OAI211_X1 U13919 ( .C1(P1_REG1_REG_14__SCAN_IN), .C2(n12117), .A(n12663), 
        .B(n15539), .ZN(n12121) );
  NAND2_X1 U13920 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n16178)
         );
  INV_X1 U13921 ( .A(n16178), .ZN(n12119) );
  NOR2_X1 U13922 ( .A1(n15534), .A2(n7793), .ZN(n12118) );
  AOI211_X1 U13923 ( .C1(n15526), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n12119), 
        .B(n12118), .ZN(n12120) );
  OAI211_X1 U13924 ( .C1(n12670), .C2(n12122), .A(n12121), .B(n12120), .ZN(
        P1_U3257) );
  OAI21_X1 U13925 ( .B1(n12124), .B2(n12125), .A(n12123), .ZN(n12247) );
  INV_X1 U13926 ( .A(n12247), .ZN(n12131) );
  XNOR2_X1 U13927 ( .A(n12126), .B(n12125), .ZN(n12127) );
  AOI222_X1 U13928 ( .A1(n14764), .A2(n15925), .B1(n14762), .B2(n14914), .C1(
        n16019), .C2(n12127), .ZN(n12250) );
  AOI21_X1 U13929 ( .B1(n12129), .B2(n12128), .A(n8319), .ZN(n12245) );
  AOI22_X1 U13930 ( .A1(n12245), .A2(n16012), .B1(n12129), .B2(n16009), .ZN(
        n12130) );
  OAI211_X1 U13931 ( .C1(n16015), .C2(n12131), .A(n12250), .B(n12130), .ZN(
        n12133) );
  NAND2_X1 U13932 ( .A1(n12133), .A2(n15984), .ZN(n12132) );
  OAI21_X1 U13933 ( .B1(n15984), .B2(n8659), .A(n12132), .ZN(P1_U3480) );
  NAND2_X1 U13934 ( .A1(n12133), .A2(n16141), .ZN(n12134) );
  OAI21_X1 U13935 ( .B1(n16141), .B2(n11207), .A(n12134), .ZN(P1_U3535) );
  NAND2_X1 U13936 ( .A1(n12135), .A2(n13876), .ZN(n12137) );
  OAI211_X1 U13937 ( .C1(n15172), .C2(n13880), .A(n12137), .B(n12136), .ZN(
        P3_U3272) );
  INV_X1 U13938 ( .A(n12138), .ZN(n12149) );
  OAI21_X1 U13939 ( .B1(n13931), .B2(n12590), .A(n12139), .ZN(n12140) );
  AOI21_X1 U13940 ( .B1(n13955), .B2(n14020), .A(n12140), .ZN(n12141) );
  OAI21_X1 U13941 ( .B1(n13226), .B2(n13996), .A(n12141), .ZN(n12142) );
  AOI21_X1 U13942 ( .B1(n13216), .B2(n13999), .A(n12142), .ZN(n12148) );
  OAI22_X1 U13943 ( .A1(n12143), .A2(n14001), .B1(n13212), .B2(n13897), .ZN(
        n12144) );
  NAND3_X1 U13944 ( .A1(n12146), .A2(n12145), .A3(n12144), .ZN(n12147) );
  OAI211_X1 U13945 ( .C1(n12149), .C2(n14001), .A(n12148), .B(n12147), .ZN(
        P2_U3189) );
  INV_X1 U13946 ( .A(n12150), .ZN(n12151) );
  NAND2_X1 U13947 ( .A1(n12152), .A2(n12151), .ZN(n14853) );
  OAI21_X1 U13948 ( .B1(n15894), .B2(n15927), .A(n15029), .ZN(n12246) );
  INV_X1 U13949 ( .A(n12246), .ZN(n12287) );
  INV_X1 U13950 ( .A(n12155), .ZN(n12157) );
  NOR2_X1 U13951 ( .A1(n14853), .A2(n14835), .ZN(n14860) );
  INV_X1 U13952 ( .A(n14860), .ZN(n14880) );
  OAI22_X1 U13953 ( .A1(n12157), .A2(n14880), .B1(n12156), .B2(n15931), .ZN(
        n12158) );
  AOI21_X1 U13954 ( .B1(n15026), .B2(n12159), .A(n12158), .ZN(n12163) );
  MUX2_X1 U13955 ( .A(n12161), .B(n12160), .S(n15894), .Z(n12162) );
  OAI211_X1 U13956 ( .C1(n12164), .C2(n12287), .A(n12163), .B(n12162), .ZN(
        P1_U3288) );
  NAND2_X1 U13957 ( .A1(n13202), .A2(n14021), .ZN(n12165) );
  XNOR2_X1 U13958 ( .A(n13210), .B(n14020), .ZN(n13415) );
  INV_X1 U13959 ( .A(n13415), .ZN(n12521) );
  XNOR2_X1 U13960 ( .A(n12522), .B(n12521), .ZN(n16091) );
  XNOR2_X1 U13961 ( .A(n12533), .B(n13415), .ZN(n12171) );
  OAI22_X1 U13962 ( .A1(n12169), .A2(n14189), .B1(n12537), .B2(n14191), .ZN(
        n12170) );
  AOI21_X1 U13963 ( .B1(n12171), .B2(n14236), .A(n12170), .ZN(n12172) );
  OAI21_X1 U13964 ( .B1(n16091), .B2(n14197), .A(n12172), .ZN(n16093) );
  NAND2_X1 U13965 ( .A1(n16093), .A2(n16041), .ZN(n12179) );
  OAI22_X1 U13966 ( .A1(n16041), .A2(n12174), .B1(n12173), .B2(n16038), .ZN(
        n12177) );
  OAI211_X1 U13967 ( .C1(n7756), .C2(n7755), .A(n14302), .B(n12589), .ZN(
        n16092) );
  NOR2_X1 U13968 ( .A1(n16092), .A2(n16045), .ZN(n12176) );
  AOI211_X1 U13969 ( .C1(n16147), .C2(n13210), .A(n12177), .B(n12176), .ZN(
        n12178) );
  OAI211_X1 U13970 ( .C1(n16091), .C2(n12713), .A(n12179), .B(n12178), .ZN(
        P2_U3256) );
  OAI21_X1 U13971 ( .B1(n12181), .B2(n13412), .A(n12180), .ZN(n16066) );
  INV_X1 U13972 ( .A(n12182), .ZN(n12183) );
  OAI211_X1 U13973 ( .C1(n16063), .C2(n12184), .A(n12183), .B(n14302), .ZN(
        n16062) );
  INV_X1 U13974 ( .A(n12185), .ZN(n12186) );
  AOI22_X1 U13975 ( .A1(n16147), .A2(n13195), .B1(n12186), .B2(n16146), .ZN(
        n12187) );
  OAI21_X1 U13976 ( .B1(n16045), .B2(n16062), .A(n12187), .ZN(n12193) );
  XNOR2_X1 U13977 ( .A(n12188), .B(n13412), .ZN(n12191) );
  NAND2_X1 U13978 ( .A1(n16066), .A2(n14121), .ZN(n12190) );
  AOI22_X1 U13979 ( .A1(n14091), .A2(n14021), .B1(n14023), .B2(n14089), .ZN(
        n12189) );
  OAI211_X1 U13980 ( .C1(n14214), .C2(n12191), .A(n12190), .B(n12189), .ZN(
        n16064) );
  MUX2_X1 U13981 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n16064), .S(n16041), .Z(
        n12192) );
  AOI211_X1 U13982 ( .C1(n16151), .C2(n16066), .A(n12193), .B(n12192), .ZN(
        n12194) );
  INV_X1 U13983 ( .A(n12194), .ZN(P2_U3258) );
  OAI21_X1 U13984 ( .B1(n12197), .B2(n12196), .A(n12195), .ZN(n12330) );
  INV_X1 U13985 ( .A(n12330), .ZN(n12204) );
  OAI21_X1 U13986 ( .B1(n12200), .B2(n12199), .A(n12198), .ZN(n12201) );
  AOI222_X1 U13987 ( .A1(n16019), .A2(n12201), .B1(n14760), .B2(n14914), .C1(
        n14762), .C2(n15925), .ZN(n12333) );
  INV_X1 U13988 ( .A(n12316), .ZN(n12202) );
  AOI21_X1 U13989 ( .B1(n14661), .B2(n12263), .A(n12202), .ZN(n12329) );
  AOI22_X1 U13990 ( .A1(n12329), .A2(n16012), .B1(n14661), .B2(n16009), .ZN(
        n12203) );
  OAI211_X1 U13991 ( .C1(n16015), .C2(n12204), .A(n12333), .B(n12203), .ZN(
        n12206) );
  NAND2_X1 U13992 ( .A1(n12206), .A2(n15984), .ZN(n12205) );
  OAI21_X1 U13993 ( .B1(n15984), .B2(n8694), .A(n12205), .ZN(P1_U3486) );
  NAND2_X1 U13994 ( .A1(n12206), .A2(n16141), .ZN(n12207) );
  OAI21_X1 U13995 ( .B1(n16141), .B2(n11289), .A(n12207), .ZN(P1_U3537) );
  XNOR2_X1 U13996 ( .A(n12208), .B(n12212), .ZN(n16072) );
  INV_X1 U13997 ( .A(n16072), .ZN(n12221) );
  INV_X1 U13998 ( .A(n12209), .ZN(n12210) );
  AOI21_X1 U13999 ( .B1(n12212), .B2(n12211), .A(n12210), .ZN(n12213) );
  OAI222_X1 U14000 ( .A1(n15960), .A2(n12214), .B1(n15962), .B2(n12362), .C1(
        n15959), .C2(n12213), .ZN(n16070) );
  NOR2_X1 U14001 ( .A1(n13715), .A2(n12215), .ZN(n12219) );
  INV_X1 U14002 ( .A(n12216), .ZN(n12217) );
  OAI22_X1 U14003 ( .A1(n13754), .A2(n16069), .B1(n12217), .B2(n15967), .ZN(
        n12218) );
  AOI211_X1 U14004 ( .C1(n16070), .C2(n13715), .A(n12219), .B(n12218), .ZN(
        n12220) );
  OAI21_X1 U14005 ( .B1(n12221), .B2(n13717), .A(n12220), .ZN(P3_U3225) );
  OAI22_X1 U14006 ( .A1(n15942), .A2(n11152), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15931), .ZN(n12224) );
  NOR2_X1 U14007 ( .A1(n15936), .A2(n12222), .ZN(n12223) );
  AOI211_X1 U14008 ( .C1(n15026), .C2(n14566), .A(n12224), .B(n12223), .ZN(
        n12227) );
  NAND2_X1 U14009 ( .A1(n12246), .A2(n12225), .ZN(n12226) );
  OAI211_X1 U14010 ( .C1(n15894), .C2(n12228), .A(n12227), .B(n12226), .ZN(
        P1_U3290) );
  XNOR2_X1 U14011 ( .A(n12229), .B(n12232), .ZN(n16083) );
  NAND2_X1 U14012 ( .A1(n13715), .A2(n12230), .ZN(n13700) );
  INV_X1 U14013 ( .A(n16057), .ZN(n13694) );
  XNOR2_X1 U14014 ( .A(n12231), .B(n12232), .ZN(n12234) );
  OAI22_X1 U14015 ( .A1(n12376), .A2(n15960), .B1(n12497), .B2(n15962), .ZN(
        n12233) );
  AOI21_X1 U14016 ( .B1(n12234), .B2(n13705), .A(n12233), .ZN(n12235) );
  OAI21_X1 U14017 ( .B1(n16083), .B2(n13694), .A(n12235), .ZN(n16085) );
  NAND2_X1 U14018 ( .A1(n16085), .A2(n13715), .ZN(n12239) );
  INV_X1 U14019 ( .A(n12236), .ZN(n12383) );
  OAI22_X1 U14020 ( .A1(n13754), .A2(n16084), .B1(n12383), .B2(n15967), .ZN(
        n12237) );
  AOI21_X1 U14021 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n7188), .A(n12237), .ZN(
        n12238) );
  OAI211_X1 U14022 ( .C1(n16083), .C2(n13700), .A(n12239), .B(n12238), .ZN(
        P3_U3224) );
  NOR2_X1 U14023 ( .A1(n15933), .A2(n12240), .ZN(n12244) );
  OAI22_X1 U14024 ( .A1(n15942), .A2(n12242), .B1(n12241), .B2(n15931), .ZN(
        n12243) );
  AOI211_X1 U14025 ( .C1(n12245), .C2(n14958), .A(n12244), .B(n12243), .ZN(
        n12249) );
  NAND2_X1 U14026 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  OAI211_X1 U14027 ( .C1(n12250), .C2(n14997), .A(n12249), .B(n12248), .ZN(
        P1_U3286) );
  OAI21_X1 U14028 ( .B1(n12253), .B2(n12252), .A(n12251), .ZN(n16081) );
  INV_X1 U14029 ( .A(n16081), .ZN(n12268) );
  XNOR2_X1 U14030 ( .A(n12255), .B(n12254), .ZN(n12259) );
  INV_X1 U14031 ( .A(n15927), .ZN(n15877) );
  OAI22_X1 U14032 ( .A1(n15012), .A2(n12256), .B1(n14397), .B2(n15916), .ZN(
        n12257) );
  AOI21_X1 U14033 ( .B1(n16081), .B2(n15877), .A(n12257), .ZN(n12258) );
  OAI21_X1 U14034 ( .B1(n16134), .B2(n12259), .A(n12258), .ZN(n16079) );
  NAND2_X1 U14035 ( .A1(n16079), .A2(n15942), .ZN(n12267) );
  OAI22_X1 U14036 ( .A1(n15942), .A2(n12260), .B1(n12350), .B2(n15931), .ZN(
        n12265) );
  NAND2_X1 U14037 ( .A1(n12261), .A2(n16076), .ZN(n12262) );
  NAND2_X1 U14038 ( .A1(n12263), .A2(n12262), .ZN(n16078) );
  NOR2_X1 U14039 ( .A1(n15936), .A2(n16078), .ZN(n12264) );
  AOI211_X1 U14040 ( .C1(n15026), .C2(n16076), .A(n12265), .B(n12264), .ZN(
        n12266) );
  OAI211_X1 U14041 ( .C1(n12268), .C2(n15029), .A(n12267), .B(n12266), .ZN(
        P1_U3285) );
  XNOR2_X1 U14042 ( .A(n12269), .B(n12270), .ZN(n15976) );
  NAND2_X1 U14043 ( .A1(n12272), .A2(n12271), .ZN(n12273) );
  NAND2_X1 U14044 ( .A1(n12274), .A2(n12273), .ZN(n12278) );
  NAND2_X1 U14045 ( .A1(n15925), .A2(n14769), .ZN(n12275) );
  OAI21_X1 U14046 ( .B1(n12276), .B2(n15916), .A(n12275), .ZN(n12277) );
  AOI21_X1 U14047 ( .B1(n12278), .B2(n16019), .A(n12277), .ZN(n15979) );
  OAI22_X1 U14048 ( .A1(n14997), .A2(n15979), .B1(n12279), .B2(n15931), .ZN(
        n12285) );
  INV_X1 U14049 ( .A(n12280), .ZN(n12283) );
  OAI21_X1 U14050 ( .B1(n15917), .B2(n15914), .A(n12281), .ZN(n12282) );
  NAND2_X1 U14051 ( .A1(n12283), .A2(n12282), .ZN(n15977) );
  OAI22_X1 U14052 ( .A1(n15936), .A2(n15977), .B1(n15978), .B2(n15933), .ZN(
        n12284) );
  AOI211_X1 U14053 ( .C1(n15894), .C2(P1_REG2_REG_2__SCAN_IN), .A(n12285), .B(
        n12284), .ZN(n12286) );
  OAI21_X1 U14054 ( .B1(n12287), .B2(n15976), .A(n12286), .ZN(P1_U3291) );
  OR2_X1 U14055 ( .A1(n15894), .A2(n12318), .ZN(n14974) );
  XNOR2_X1 U14056 ( .A(n12288), .B(n12290), .ZN(n16016) );
  INV_X1 U14057 ( .A(n15003), .ZN(n14972) );
  XNOR2_X1 U14058 ( .A(n12289), .B(n12290), .ZN(n16018) );
  NAND2_X1 U14059 ( .A1(n15925), .A2(n14767), .ZN(n12291) );
  OAI21_X1 U14060 ( .B1(n12292), .B2(n15916), .A(n12291), .ZN(n16010) );
  MUX2_X1 U14061 ( .A(n16010), .B(P1_REG2_REG_4__SCAN_IN), .S(n15894), .Z(
        n12301) );
  AND2_X1 U14062 ( .A1(n12293), .A2(n16008), .ZN(n12294) );
  NOR2_X1 U14063 ( .A1(n12295), .A2(n12294), .ZN(n16013) );
  NAND2_X1 U14064 ( .A1(n14958), .A2(n16013), .ZN(n12298) );
  INV_X1 U14065 ( .A(n15931), .ZN(n15887) );
  NAND2_X1 U14066 ( .A1(n15887), .A2(n12296), .ZN(n12297) );
  OAI211_X1 U14067 ( .C1(n12299), .C2(n15933), .A(n12298), .B(n12297), .ZN(
        n12300) );
  AOI211_X1 U14068 ( .C1(n14972), .C2(n16018), .A(n12301), .B(n12300), .ZN(
        n12302) );
  OAI21_X1 U14069 ( .B1(n14974), .B2(n16016), .A(n12302), .ZN(P1_U3289) );
  NAND2_X1 U14070 ( .A1(n14197), .A2(n15897), .ZN(n16186) );
  OAI211_X1 U14071 ( .C1(n12305), .C2(n16182), .A(n12304), .B(n12303), .ZN(
        n12306) );
  AOI21_X1 U14072 ( .B1(n12307), .B2(n16186), .A(n12306), .ZN(n12311) );
  INV_X1 U14073 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n12308) );
  OR2_X1 U14074 ( .A1(n16192), .A2(n12308), .ZN(n12309) );
  OAI21_X1 U14075 ( .B1(n12311), .B2(n16190), .A(n12309), .ZN(P2_U3454) );
  OR2_X1 U14076 ( .A1(n16189), .A2(n10493), .ZN(n12310) );
  OAI21_X1 U14077 ( .B1(n12311), .B2(n16188), .A(n12310), .ZN(P2_U3507) );
  XNOR2_X1 U14078 ( .A(n12312), .B(n12314), .ZN(n12340) );
  OAI21_X1 U14079 ( .B1(n12315), .B2(n12314), .A(n12313), .ZN(n12337) );
  INV_X1 U14080 ( .A(n12337), .ZN(n12319) );
  NAND2_X1 U14081 ( .A1(n14914), .A2(n14759), .ZN(n12335) );
  AOI211_X1 U14082 ( .C1(n14560), .C2(n12316), .A(n16077), .B(n12394), .ZN(
        n12336) );
  INV_X1 U14083 ( .A(n12336), .ZN(n12317) );
  OAI211_X1 U14084 ( .C1(n12319), .C2(n12318), .A(n12335), .B(n12317), .ZN(
        n12324) );
  INV_X1 U14085 ( .A(n15029), .ZN(n15941) );
  NAND2_X1 U14086 ( .A1(n12337), .A2(n15941), .ZN(n12322) );
  NAND2_X1 U14087 ( .A1(n15925), .A2(n14761), .ZN(n12334) );
  OAI22_X1 U14088 ( .A1(n15894), .A2(n12334), .B1(n14558), .B2(n15931), .ZN(
        n12320) );
  AOI21_X1 U14089 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n14997), .A(n12320), 
        .ZN(n12321) );
  OAI211_X1 U14090 ( .C1(n7777), .C2(n15933), .A(n12322), .B(n12321), .ZN(
        n12323) );
  AOI21_X1 U14091 ( .B1(n12324), .B2(n14860), .A(n12323), .ZN(n12325) );
  OAI21_X1 U14092 ( .B1(n12340), .B2(n15003), .A(n12325), .ZN(P1_U3283) );
  NOR2_X1 U14093 ( .A1(n7778), .A2(n15933), .ZN(n12328) );
  OAI22_X1 U14094 ( .A1(n15942), .A2(n12326), .B1(n14659), .B2(n15931), .ZN(
        n12327) );
  AOI211_X1 U14095 ( .C1(n12329), .C2(n14958), .A(n12328), .B(n12327), .ZN(
        n12332) );
  NAND2_X1 U14096 ( .A1(n12330), .A2(n15001), .ZN(n12331) );
  OAI211_X1 U14097 ( .C1(n12333), .C2(n14997), .A(n12332), .B(n12331), .ZN(
        P1_U3284) );
  NAND2_X1 U14098 ( .A1(n12335), .A2(n12334), .ZN(n14556) );
  AOI211_X1 U14099 ( .C1(n14560), .C2(n16009), .A(n14556), .B(n12336), .ZN(
        n12339) );
  NAND2_X1 U14100 ( .A1(n12337), .A2(n16139), .ZN(n12338) );
  OAI211_X1 U14101 ( .C1(n16134), .C2(n12340), .A(n12339), .B(n12338), .ZN(
        n12342) );
  NAND2_X1 U14102 ( .A1(n12342), .A2(n15984), .ZN(n12341) );
  OAI21_X1 U14103 ( .B1(n15984), .B2(n8713), .A(n12341), .ZN(P1_U3489) );
  NAND2_X1 U14104 ( .A1(n12342), .A2(n16141), .ZN(n12343) );
  OAI21_X1 U14105 ( .B1(n16141), .B2(n11328), .A(n12343), .ZN(P1_U3538) );
  AOI22_X1 U14106 ( .A1(n16076), .A2(n14526), .B1(n14533), .B2(n14762), .ZN(
        n12344) );
  XNOR2_X1 U14107 ( .A(n12344), .B(n14589), .ZN(n14392) );
  AOI22_X1 U14108 ( .A1(n16076), .A2(n14533), .B1(n14480), .B2(n14762), .ZN(
        n14393) );
  XNOR2_X1 U14109 ( .A(n14392), .B(n14393), .ZN(n12349) );
  AOI21_X1 U14110 ( .B1(n12349), .B2(n12348), .A(n14391), .ZN(n12356) );
  NOR2_X1 U14111 ( .A1(n16203), .A2(n12350), .ZN(n12354) );
  NAND2_X1 U14112 ( .A1(n14714), .A2(n14763), .ZN(n12352) );
  OAI211_X1 U14113 ( .C1(n14397), .C2(n14538), .A(n12352), .B(n12351), .ZN(
        n12353) );
  AOI211_X1 U14114 ( .C1(n16076), .C2(n7185), .A(n12354), .B(n12353), .ZN(
        n12355) );
  OAI21_X1 U14115 ( .B1(n12356), .B2(n14740), .A(n12355), .ZN(P1_U3221) );
  INV_X1 U14116 ( .A(n12357), .ZN(n12358) );
  XNOR2_X1 U14117 ( .A(n12379), .B(n13119), .ZN(n12361) );
  XNOR2_X1 U14118 ( .A(n12361), .B(n13580), .ZN(n12374) );
  XNOR2_X1 U14119 ( .A(n12516), .B(n12498), .ZN(n12494) );
  XNOR2_X1 U14120 ( .A(n12494), .B(n12497), .ZN(n12363) );
  NAND2_X1 U14121 ( .A1(n12362), .A2(n12361), .ZN(n12364) );
  NAND2_X1 U14122 ( .A1(n12495), .A2(n13476), .ZN(n12371) );
  AOI21_X1 U14123 ( .B1(n12372), .B2(n12364), .A(n12363), .ZN(n12370) );
  NAND2_X1 U14124 ( .A1(n13564), .A2(n12513), .ZN(n12368) );
  INV_X1 U14125 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15339) );
  NOR2_X1 U14126 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15339), .ZN(n15701) );
  AOI21_X1 U14127 ( .B1(n13580), .B2(n13549), .A(n15701), .ZN(n12367) );
  NAND2_X1 U14128 ( .A1(n12504), .A2(n12516), .ZN(n12366) );
  INV_X1 U14129 ( .A(n13551), .ZN(n13557) );
  NAND2_X1 U14130 ( .A1(n13557), .A2(n13578), .ZN(n12365) );
  AND4_X1 U14131 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12369) );
  OAI21_X1 U14132 ( .B1(n12371), .B2(n12370), .A(n12369), .ZN(P3_U3157) );
  OAI21_X1 U14133 ( .B1(n12374), .B2(n12373), .A(n12372), .ZN(n12375) );
  NAND2_X1 U14134 ( .A1(n12375), .A2(n13476), .ZN(n12381) );
  OAI22_X1 U14135 ( .A1(n12376), .A2(n13559), .B1(n12497), .B2(n13551), .ZN(
        n12377) );
  AOI211_X1 U14136 ( .C1(n12504), .C2(n12379), .A(n12378), .B(n12377), .ZN(
        n12380) );
  OAI211_X1 U14137 ( .C1(n12383), .C2(n12382), .A(n12381), .B(n12380), .ZN(
        P3_U3171) );
  INV_X1 U14138 ( .A(n14826), .ZN(n14815) );
  INV_X1 U14139 ( .A(n12384), .ZN(n12386) );
  OAI222_X1 U14140 ( .A1(P1_U3086), .A2(n14815), .B1(n15160), .B2(n12386), 
        .C1(n12385), .C2(n15157), .ZN(P1_U3337) );
  INV_X1 U14141 ( .A(n12728), .ZN(n12923) );
  OAI222_X1 U14142 ( .A1(n14370), .A2(n12387), .B1(n14378), .B2(n12386), .C1(
        n12923), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U14143 ( .A(n12388), .ZN(n12390) );
  OAI222_X1 U14144 ( .A1(n12389), .A2(P1_U3086), .B1(n15160), .B2(n12390), 
        .C1(n8015), .C2(n15157), .ZN(P1_U3335) );
  INV_X1 U14145 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12391) );
  OAI222_X1 U14146 ( .A1(n14370), .A2(n12391), .B1(P2_U3088), .B2(n13399), 
        .C1(n14378), .C2(n12390), .ZN(P2_U3307) );
  XNOR2_X1 U14147 ( .A(n12392), .B(n12401), .ZN(n12393) );
  AOI222_X1 U14148 ( .A1(n14760), .A2(n15925), .B1(n14758), .B2(n14914), .C1(
        n16019), .C2(n12393), .ZN(n12568) );
  INV_X1 U14149 ( .A(n12394), .ZN(n12396) );
  INV_X1 U14150 ( .A(n12463), .ZN(n12395) );
  AOI21_X1 U14151 ( .B1(n14703), .B2(n12396), .A(n12395), .ZN(n12566) );
  NOR2_X1 U14152 ( .A1(n14407), .A2(n15933), .ZN(n12399) );
  OAI22_X1 U14153 ( .A1(n15942), .A2(n12397), .B1(n14701), .B2(n15931), .ZN(
        n12398) );
  AOI211_X1 U14154 ( .C1(n12566), .C2(n14958), .A(n12399), .B(n12398), .ZN(
        n12404) );
  OAI21_X1 U14155 ( .B1(n12402), .B2(n12401), .A(n12400), .ZN(n12565) );
  NAND2_X1 U14156 ( .A1(n12565), .A2(n15001), .ZN(n12403) );
  OAI211_X1 U14157 ( .C1(n12568), .C2(n14997), .A(n12404), .B(n12403), .ZN(
        P1_U3282) );
  INV_X1 U14158 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12414) );
  NOR2_X1 U14159 ( .A1(n12435), .A2(n12414), .ZN(n12413) );
  NAND2_X1 U14160 ( .A1(n15481), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U14161 ( .A1(n15481), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12995), 
        .B2(n12429), .ZN(n15480) );
  AOI21_X1 U14162 ( .B1(n12419), .B2(n12542), .A(n12405), .ZN(n15511) );
  XNOR2_X1 U14163 ( .A(n12421), .B(n12406), .ZN(n15510) );
  OAI22_X1 U14164 ( .A1(n15511), .A2(n15510), .B1(n15503), .B2(
        P2_REG2_REG_12__SCAN_IN), .ZN(n15492) );
  INV_X1 U14165 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U14166 ( .A1(n15489), .A2(n12407), .B1(P2_REG2_REG_13__SCAN_IN), 
        .B2(n12423), .ZN(n15491) );
  NOR2_X1 U14167 ( .A1(n15492), .A2(n15491), .ZN(n15490) );
  AOI21_X1 U14168 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n15489), .A(n15490), 
        .ZN(n15459) );
  AND2_X1 U14169 ( .A1(n12424), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n15456) );
  INV_X1 U14170 ( .A(n15456), .ZN(n12408) );
  NOR2_X1 U14171 ( .A1(n12424), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n15457) );
  AOI21_X1 U14172 ( .B1(n15459), .B2(n12408), .A(n15457), .ZN(n12409) );
  NAND2_X1 U14173 ( .A1(n12426), .A2(n12409), .ZN(n12410) );
  XNOR2_X1 U14174 ( .A(n12409), .B(n15467), .ZN(n15472) );
  NAND2_X1 U14175 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15472), .ZN(n15471) );
  NAND2_X1 U14176 ( .A1(n12410), .A2(n15471), .ZN(n15479) );
  NAND2_X1 U14177 ( .A1(n15480), .A2(n15479), .ZN(n15478) );
  NAND2_X1 U14178 ( .A1(n12411), .A2(n15478), .ZN(n12415) );
  INV_X1 U14179 ( .A(n12415), .ZN(n12412) );
  AOI211_X1 U14180 ( .C1(n12414), .C2(n12435), .A(n12413), .B(n12412), .ZN(
        n12717) );
  NOR2_X1 U14181 ( .A1(n12435), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12416) );
  AOI211_X1 U14182 ( .C1(n12435), .C2(P2_REG2_REG_17__SCAN_IN), .A(n12416), 
        .B(n12415), .ZN(n12417) );
  OR3_X1 U14183 ( .A1(n12717), .A2(n12417), .A3(n15412), .ZN(n12434) );
  AND2_X1 U14184 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13944) );
  XNOR2_X1 U14185 ( .A(n12435), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n12722) );
  XNOR2_X1 U14186 ( .A(n12429), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15483) );
  OAI21_X1 U14187 ( .B1(n11279), .B2(n12419), .A(n12418), .ZN(n15506) );
  MUX2_X1 U14188 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n12420), .S(n12421), .Z(
        n15507) );
  NOR2_X1 U14189 ( .A1(n15506), .A2(n15507), .ZN(n15505) );
  AOI21_X1 U14190 ( .B1(n12420), .B2(n12421), .A(n15505), .ZN(n15497) );
  MUX2_X1 U14191 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n12422), .S(n15489), .Z(
        n15496) );
  NAND2_X1 U14192 ( .A1(n15497), .A2(n15496), .ZN(n15495) );
  OAI21_X1 U14193 ( .B1(n12422), .B2(n12423), .A(n15495), .ZN(n15463) );
  MUX2_X1 U14194 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n12425), .S(n12424), .Z(
        n15462) );
  NAND2_X1 U14195 ( .A1(n15463), .A2(n15462), .ZN(n15461) );
  OAI21_X1 U14196 ( .B1(n12425), .B2(n15453), .A(n15461), .ZN(n12427) );
  NAND2_X1 U14197 ( .A1(n12426), .A2(n12427), .ZN(n12428) );
  XNOR2_X1 U14198 ( .A(n12427), .B(n15467), .ZN(n15474) );
  NAND2_X1 U14199 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15474), .ZN(n15473) );
  NAND2_X1 U14200 ( .A1(n12428), .A2(n15473), .ZN(n15484) );
  NAND2_X1 U14201 ( .A1(n15483), .A2(n15484), .ZN(n15482) );
  OAI21_X1 U14202 ( .B1(n12430), .B2(n12429), .A(n15482), .ZN(n12721) );
  XNOR2_X1 U14203 ( .A(n12722), .B(n12721), .ZN(n12431) );
  NOR2_X1 U14204 ( .A1(n15508), .A2(n12431), .ZN(n12432) );
  AOI211_X1 U14205 ( .C1(n15502), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n13944), 
        .B(n12432), .ZN(n12433) );
  OAI211_X1 U14206 ( .C1(n15468), .C2(n12435), .A(n12434), .B(n12433), .ZN(
        P2_U3231) );
  AOI22_X1 U14207 ( .A1(n15026), .A2(n12437), .B1(n15887), .B2(n12436), .ZN(
        n12438) );
  OAI21_X1 U14208 ( .B1(n15936), .B2(n12439), .A(n12438), .ZN(n12442) );
  MUX2_X1 U14209 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n12440), .S(n15942), .Z(
        n12441) );
  AOI211_X1 U14210 ( .C1(n15941), .C2(n12443), .A(n12442), .B(n12441), .ZN(
        n12444) );
  INV_X1 U14211 ( .A(n12444), .ZN(P1_U3287) );
  XNOR2_X1 U14212 ( .A(n12445), .B(n12449), .ZN(n12447) );
  OAI22_X1 U14213 ( .A1(n12497), .A2(n15960), .B1(n12776), .B2(n15962), .ZN(
        n12446) );
  AOI21_X1 U14214 ( .B1(n12447), .B2(n13705), .A(n12446), .ZN(n16110) );
  OAI21_X1 U14215 ( .B1(n12450), .B2(n12449), .A(n12448), .ZN(n16109) );
  AOI22_X1 U14216 ( .A1(n7188), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15909), 
        .B2(n12500), .ZN(n12451) );
  OAI21_X1 U14217 ( .B1(n12499), .B2(n13754), .A(n12451), .ZN(n12452) );
  AOI21_X1 U14218 ( .B1(n16109), .B2(n13757), .A(n12452), .ZN(n12453) );
  OAI21_X1 U14219 ( .B1(n16110), .B2(n7188), .A(n12453), .ZN(P3_U3222) );
  OAI21_X1 U14220 ( .B1(n12456), .B2(n12455), .A(n12454), .ZN(n12573) );
  OAI22_X1 U14221 ( .A1(n15012), .A2(n14615), .B1(n12457), .B2(n15916), .ZN(
        n12462) );
  XNOR2_X1 U14222 ( .A(n12458), .B(n12459), .ZN(n12460) );
  NOR2_X1 U14223 ( .A1(n12460), .A2(n16134), .ZN(n12461) );
  AOI211_X1 U14224 ( .C1(n15877), .C2(n12573), .A(n12462), .B(n12461), .ZN(
        n12576) );
  AOI21_X1 U14225 ( .B1(n14387), .B2(n12463), .A(n8323), .ZN(n12574) );
  INV_X1 U14226 ( .A(n14387), .ZN(n14620) );
  NOR2_X1 U14227 ( .A1(n14620), .A2(n15933), .ZN(n12466) );
  OAI22_X1 U14228 ( .A1(n15942), .A2(n12464), .B1(n14613), .B2(n15931), .ZN(
        n12465) );
  AOI211_X1 U14229 ( .C1(n12574), .C2(n14958), .A(n12466), .B(n12465), .ZN(
        n12468) );
  NAND2_X1 U14230 ( .A1(n12573), .A2(n15941), .ZN(n12467) );
  OAI211_X1 U14231 ( .C1(n12576), .C2(n14997), .A(n12468), .B(n12467), .ZN(
        P1_U3281) );
  INV_X1 U14232 ( .A(n12469), .ZN(n13025) );
  OAI222_X1 U14233 ( .A1(P1_U3086), .A2(n12471), .B1(n15160), .B2(n13025), 
        .C1(n12470), .C2(n15157), .ZN(P1_U3336) );
  INV_X1 U14234 ( .A(n13224), .ZN(n16117) );
  OAI211_X1 U14235 ( .C1(n7343), .C2(n12472), .A(n12549), .B(n13940), .ZN(
        n12477) );
  OAI22_X1 U14236 ( .A1(n13931), .A2(n12541), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12473), .ZN(n12475) );
  NOR2_X1 U14237 ( .A1(n13992), .A2(n12537), .ZN(n12474) );
  AOI211_X1 U14238 ( .C1(n13975), .C2(n14017), .A(n12475), .B(n12474), .ZN(
        n12476) );
  OAI211_X1 U14239 ( .C1(n16117), .C2(n13978), .A(n12477), .B(n12476), .ZN(
        P2_U3208) );
  INV_X1 U14240 ( .A(n12478), .ZN(n12519) );
  OAI222_X1 U14241 ( .A1(n7861), .A2(P1_U3086), .B1(n15160), .B2(n12519), .C1(
        n12479), .C2(n15157), .ZN(P1_U3334) );
  XNOR2_X1 U14242 ( .A(n12480), .B(n12481), .ZN(n16135) );
  OAI21_X1 U14243 ( .B1(n12484), .B2(n12483), .A(n12482), .ZN(n16138) );
  AOI21_X1 U14244 ( .B1(n12485), .B2(n14679), .A(n16077), .ZN(n12486) );
  NAND2_X1 U14245 ( .A1(n12486), .A2(n12634), .ZN(n16132) );
  NAND2_X1 U14246 ( .A1(n14914), .A2(n14756), .ZN(n12488) );
  NAND2_X1 U14247 ( .A1(n15925), .A2(n14758), .ZN(n12487) );
  NAND2_X1 U14248 ( .A1(n12488), .A2(n12487), .ZN(n14674) );
  INV_X1 U14249 ( .A(n14674), .ZN(n16131) );
  OAI22_X1 U14250 ( .A1(n15894), .A2(n16131), .B1(n14677), .B2(n15931), .ZN(
        n12490) );
  NOR2_X1 U14251 ( .A1(n8322), .A2(n15933), .ZN(n12489) );
  AOI211_X1 U14252 ( .C1(n15894), .C2(P1_REG2_REG_13__SCAN_IN), .A(n12490), 
        .B(n12489), .ZN(n12491) );
  OAI21_X1 U14253 ( .B1(n14880), .B2(n16132), .A(n12491), .ZN(n12492) );
  AOI21_X1 U14254 ( .B1(n16138), .B2(n15001), .A(n12492), .ZN(n12493) );
  OAI21_X1 U14255 ( .B1(n15003), .B2(n16135), .A(n12493), .ZN(P1_U3280) );
  INV_X1 U14256 ( .A(n12494), .ZN(n12496) );
  XNOR2_X1 U14257 ( .A(n12499), .B(n12498), .ZN(n12611) );
  XNOR2_X1 U14258 ( .A(n12611), .B(n13578), .ZN(n12613) );
  XNOR2_X1 U14259 ( .A(n12614), .B(n12613), .ZN(n12506) );
  NAND2_X1 U14260 ( .A1(n13564), .A2(n12500), .ZN(n12502) );
  INV_X1 U14261 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15377) );
  NOR2_X1 U14262 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15377), .ZN(n15718) );
  AOI21_X1 U14263 ( .B1(n13579), .B2(n13549), .A(n15718), .ZN(n12501) );
  OAI211_X1 U14264 ( .C1(n12776), .C2(n13551), .A(n12502), .B(n12501), .ZN(
        n12503) );
  AOI21_X1 U14265 ( .B1(n16108), .B2(n12504), .A(n12503), .ZN(n12505) );
  OAI21_X1 U14266 ( .B1(n12506), .B2(n13566), .A(n12505), .ZN(P3_U3176) );
  AOI21_X1 U14267 ( .B1(n12509), .B2(n12507), .A(n7317), .ZN(n16098) );
  AOI22_X1 U14268 ( .A1(n13708), .A2(n13580), .B1(n13578), .B2(n9880), .ZN(
        n12512) );
  XOR2_X1 U14269 ( .A(n12509), .B(n12508), .Z(n12510) );
  NAND2_X1 U14270 ( .A1(n12510), .A2(n13705), .ZN(n12511) );
  OAI211_X1 U14271 ( .C1(n16098), .C2(n13694), .A(n12512), .B(n12511), .ZN(
        n16100) );
  NAND2_X1 U14272 ( .A1(n16100), .A2(n13715), .ZN(n12518) );
  INV_X1 U14273 ( .A(n12513), .ZN(n12514) );
  OAI22_X1 U14274 ( .A1(n13715), .A2(n9907), .B1(n12514), .B2(n15967), .ZN(
        n12515) );
  AOI21_X1 U14275 ( .B1(n12516), .B2(n13696), .A(n12515), .ZN(n12517) );
  OAI211_X1 U14276 ( .C1(n16098), .C2(n13700), .A(n12518), .B(n12517), .ZN(
        P3_U3223) );
  OAI222_X1 U14277 ( .A1(n14370), .A2(n12520), .B1(P2_U3088), .B2(n13452), 
        .C1(n14378), .C2(n12519), .ZN(P2_U3306) );
  NAND2_X1 U14278 ( .A1(n12522), .A2(n12521), .ZN(n12524) );
  NAND2_X1 U14279 ( .A1(n13210), .A2(n14020), .ZN(n12523) );
  NAND2_X1 U14280 ( .A1(n12524), .A2(n12523), .ZN(n12584) );
  INV_X1 U14281 ( .A(n12584), .ZN(n12526) );
  XNOR2_X1 U14282 ( .A(n13216), .B(n14019), .ZN(n13414) );
  OR2_X1 U14283 ( .A1(n13216), .A2(n14019), .ZN(n12527) );
  NAND2_X1 U14284 ( .A1(n13224), .A2(n13226), .ZN(n12699) );
  OR2_X1 U14285 ( .A1(n13224), .A2(n13226), .ZN(n12528) );
  NAND2_X1 U14286 ( .A1(n12530), .A2(n13417), .ZN(n12531) );
  NAND2_X1 U14287 ( .A1(n12704), .A2(n12531), .ZN(n16115) );
  OR2_X1 U14288 ( .A1(n13210), .A2(n13212), .ZN(n12532) );
  NAND2_X1 U14289 ( .A1(n13210), .A2(n13212), .ZN(n12534) );
  NAND2_X1 U14290 ( .A1(n12535), .A2(n12534), .ZN(n12581) );
  AND2_X1 U14291 ( .A1(n13216), .A2(n12537), .ZN(n12536) );
  OAI21_X1 U14292 ( .B1(n7313), .B2(n13417), .A(n12700), .ZN(n12539) );
  INV_X1 U14293 ( .A(n14017), .ZN(n12697) );
  OAI22_X1 U14294 ( .A1(n12537), .A2(n14189), .B1(n12697), .B2(n14191), .ZN(
        n12538) );
  AOI21_X1 U14295 ( .B1(n12539), .B2(n14236), .A(n12538), .ZN(n12540) );
  OAI21_X1 U14296 ( .B1(n16115), .B2(n14197), .A(n12540), .ZN(n16118) );
  NAND2_X1 U14297 ( .A1(n16118), .A2(n16041), .ZN(n12546) );
  OAI22_X1 U14298 ( .A1(n16041), .A2(n12542), .B1(n12541), .B2(n16038), .ZN(
        n12544) );
  NAND2_X1 U14299 ( .A1(n12588), .A2(n16117), .ZN(n12709) );
  OAI211_X1 U14300 ( .C1(n12588), .C2(n16117), .A(n12709), .B(n14302), .ZN(
        n16116) );
  NOR2_X1 U14301 ( .A1(n16116), .A2(n16045), .ZN(n12543) );
  AOI211_X1 U14302 ( .C1(n16147), .C2(n13224), .A(n12544), .B(n12543), .ZN(
        n12545) );
  OAI211_X1 U14303 ( .C1(n16115), .C2(n12713), .A(n12546), .B(n12545), .ZN(
        P2_U3254) );
  NAND2_X1 U14304 ( .A1(n13968), .A2(n14018), .ZN(n12547) );
  OAI22_X1 U14305 ( .A1(n12549), .A2(n14001), .B1(n12548), .B2(n12547), .ZN(
        n12552) );
  INV_X1 U14306 ( .A(n12550), .ZN(n12551) );
  NAND2_X1 U14307 ( .A1(n12552), .A2(n12551), .ZN(n12558) );
  INV_X1 U14308 ( .A(n13244), .ZN(n12822) );
  NOR2_X1 U14309 ( .A1(n13996), .A2(n12822), .ZN(n12556) );
  NAND2_X1 U14310 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15516)
         );
  INV_X1 U14311 ( .A(n12553), .ZN(n12710) );
  NAND2_X1 U14312 ( .A1(n13994), .A2(n12710), .ZN(n12554) );
  OAI211_X1 U14313 ( .C1(n13992), .C2(n13226), .A(n15516), .B(n12554), .ZN(
        n12555) );
  AOI211_X1 U14314 ( .C1(n13237), .C2(n13999), .A(n12556), .B(n12555), .ZN(
        n12557) );
  OAI211_X1 U14315 ( .C1(n12559), .C2(n14001), .A(n12558), .B(n12557), .ZN(
        P2_U3196) );
  INV_X1 U14316 ( .A(n12560), .ZN(n12561) );
  OAI222_X1 U14317 ( .A1(n12562), .A2(P3_U3151), .B1(n13880), .B2(n15293), 
        .C1(n13131), .C2(n12561), .ZN(P3_U3271) );
  OAI222_X1 U14318 ( .A1(n13131), .A2(n12564), .B1(P3_U3151), .B2(n12563), 
        .C1(n15290), .C2(n13880), .ZN(P3_U3270) );
  INV_X1 U14319 ( .A(n12565), .ZN(n12569) );
  AOI22_X1 U14320 ( .A1(n12566), .A2(n16012), .B1(n14703), .B2(n16009), .ZN(
        n12567) );
  OAI211_X1 U14321 ( .C1(n16015), .C2(n12569), .A(n12568), .B(n12567), .ZN(
        n12571) );
  NAND2_X1 U14322 ( .A1(n12571), .A2(n16141), .ZN(n12570) );
  OAI21_X1 U14323 ( .B1(n16141), .B2(n11524), .A(n12570), .ZN(P1_U3539) );
  NAND2_X1 U14324 ( .A1(n12571), .A2(n15984), .ZN(n12572) );
  OAI21_X1 U14325 ( .B1(n15984), .B2(n8731), .A(n12572), .ZN(P1_U3492) );
  INV_X1 U14326 ( .A(n12573), .ZN(n12577) );
  AOI22_X1 U14327 ( .A1(n12574), .A2(n16012), .B1(n14387), .B2(n16009), .ZN(
        n12575) );
  OAI211_X1 U14328 ( .C1(n12577), .C2(n15881), .A(n12576), .B(n12575), .ZN(
        n12579) );
  NAND2_X1 U14329 ( .A1(n12579), .A2(n15984), .ZN(n12578) );
  OAI21_X1 U14330 ( .B1(n15984), .B2(n8746), .A(n12578), .ZN(P1_U3495) );
  NAND2_X1 U14331 ( .A1(n12579), .A2(n16141), .ZN(n12580) );
  OAI21_X1 U14332 ( .B1(n16141), .B2(n11522), .A(n12580), .ZN(P1_U3540) );
  XNOR2_X1 U14333 ( .A(n12581), .B(n13414), .ZN(n12587) );
  OAI22_X1 U14334 ( .A1(n13226), .A2(n14191), .B1(n13212), .B2(n14189), .ZN(
        n12586) );
  INV_X1 U14335 ( .A(n12582), .ZN(n12583) );
  AOI21_X1 U14336 ( .B1(n13414), .B2(n12584), .A(n12583), .ZN(n12760) );
  NOR2_X1 U14337 ( .A1(n12760), .A2(n14197), .ZN(n12585) );
  AOI211_X1 U14338 ( .C1(n14236), .C2(n12587), .A(n12586), .B(n12585), .ZN(
        n12759) );
  AOI21_X1 U14339 ( .B1(n13216), .B2(n12589), .A(n12588), .ZN(n12757) );
  INV_X1 U14340 ( .A(n12590), .ZN(n12591) );
  AOI22_X1 U14341 ( .A1(n16156), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12591), 
        .B2(n16146), .ZN(n12592) );
  OAI21_X1 U14342 ( .B1(n7492), .B2(n14231), .A(n12592), .ZN(n12594) );
  NOR2_X1 U14343 ( .A1(n12760), .A2(n12713), .ZN(n12593) );
  AOI211_X1 U14344 ( .C1(n12757), .C2(n14159), .A(n12594), .B(n12593), .ZN(
        n12595) );
  OAI21_X1 U14345 ( .B1(n12759), .B2(n16156), .A(n12595), .ZN(P2_U3255) );
  INV_X1 U14346 ( .A(n12596), .ZN(n12598) );
  NAND2_X1 U14347 ( .A1(n12598), .A2(n12597), .ZN(n12599) );
  XNOR2_X1 U14348 ( .A(n12600), .B(n12599), .ZN(n12606) );
  INV_X1 U14349 ( .A(n14016), .ZN(n13251) );
  OAI22_X1 U14350 ( .A1(n12697), .A2(n14189), .B1(n13251), .B2(n14191), .ZN(
        n12960) );
  OAI22_X1 U14351 ( .A1(n13931), .A2(n16144), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12601), .ZN(n12602) );
  AOI21_X1 U14352 ( .B1(n12603), .B2(n12960), .A(n12602), .ZN(n12605) );
  NAND2_X1 U14353 ( .A1(n16148), .A2(n13999), .ZN(n12604) );
  OAI211_X1 U14354 ( .C1(n12606), .C2(n14001), .A(n12605), .B(n12604), .ZN(
        P2_U3206) );
  INV_X1 U14355 ( .A(n12607), .ZN(n12627) );
  INV_X1 U14356 ( .A(n15157), .ZN(n15392) );
  AOI22_X1 U14357 ( .A1(n12608), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n15392), .ZN(n12609) );
  OAI21_X1 U14358 ( .B1(n12627), .B2(n15160), .A(n12609), .ZN(P1_U3331) );
  XNOR2_X1 U14359 ( .A(n12610), .B(n13119), .ZN(n12777) );
  XNOR2_X1 U14360 ( .A(n12777), .B(n13577), .ZN(n12616) );
  INV_X1 U14361 ( .A(n12611), .ZN(n12612) );
  NAND2_X1 U14362 ( .A1(n12615), .A2(n12616), .ZN(n12779) );
  OAI21_X1 U14363 ( .B1(n12616), .B2(n12615), .A(n12779), .ZN(n12621) );
  NOR2_X1 U14364 ( .A1(n12853), .A2(n13561), .ZN(n12620) );
  NAND2_X1 U14365 ( .A1(n13564), .A2(n12658), .ZN(n12618) );
  INV_X1 U14366 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n15230) );
  NOR2_X1 U14367 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15230), .ZN(n15735) );
  AOI21_X1 U14368 ( .B1(n13578), .B2(n13549), .A(n15735), .ZN(n12617) );
  OAI211_X1 U14369 ( .C1(n12808), .C2(n13551), .A(n12618), .B(n12617), .ZN(
        n12619) );
  AOI211_X1 U14370 ( .C1(n12621), .C2(n13476), .A(n12620), .B(n12619), .ZN(
        n12622) );
  INV_X1 U14371 ( .A(n12622), .ZN(P3_U3164) );
  OAI222_X1 U14372 ( .A1(n14370), .A2(n12625), .B1(P2_U3088), .B2(n12624), 
        .C1(n14378), .C2(n12623), .ZN(P2_U3305) );
  OAI222_X1 U14373 ( .A1(P2_U3088), .A2(n12628), .B1(n14378), .B2(n12627), 
        .C1(n12626), .C2(n14370), .ZN(P2_U3303) );
  XNOR2_X1 U14374 ( .A(n12629), .B(n12633), .ZN(n12771) );
  INV_X1 U14375 ( .A(n12630), .ZN(n12631) );
  AOI21_X1 U14376 ( .B1(n12633), .B2(n12632), .A(n12631), .ZN(n12769) );
  NAND2_X1 U14377 ( .A1(n12634), .A2(n16177), .ZN(n12765) );
  NAND2_X1 U14378 ( .A1(n12765), .A2(n14958), .ZN(n12643) );
  NAND2_X1 U14379 ( .A1(n14914), .A2(n14755), .ZN(n12636) );
  NAND2_X1 U14380 ( .A1(n15925), .A2(n14757), .ZN(n12635) );
  NAND2_X1 U14381 ( .A1(n12636), .A2(n12635), .ZN(n16176) );
  INV_X1 U14382 ( .A(n16176), .ZN(n12640) );
  NAND2_X1 U14383 ( .A1(n14997), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12639) );
  NAND2_X1 U14384 ( .A1(n15887), .A2(n12637), .ZN(n12638) );
  OAI211_X1 U14385 ( .C1(n15894), .C2(n12640), .A(n12639), .B(n12638), .ZN(
        n12641) );
  AOI21_X1 U14386 ( .B1(n16177), .B2(n15026), .A(n12641), .ZN(n12642) );
  OAI21_X1 U14387 ( .B1(n7298), .B2(n12643), .A(n12642), .ZN(n12644) );
  AOI21_X1 U14388 ( .B1(n12769), .B2(n15001), .A(n12644), .ZN(n12645) );
  OAI21_X1 U14389 ( .B1(n15003), .B2(n12771), .A(n12645), .ZN(P1_U3279) );
  OAI222_X1 U14390 ( .A1(n12647), .A2(P3_U3151), .B1(n13880), .B2(n15284), 
        .C1(n13131), .C2(n12646), .ZN(P3_U3269) );
  INV_X1 U14391 ( .A(n12648), .ZN(n12684) );
  AOI22_X1 U14392 ( .A1(n12649), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n15392), .ZN(n12650) );
  OAI21_X1 U14393 ( .B1(n12684), .B2(n15160), .A(n12650), .ZN(P1_U3330) );
  XNOR2_X1 U14394 ( .A(n12651), .B(n12653), .ZN(n12657) );
  OAI21_X1 U14395 ( .B1(n12654), .B2(n12653), .A(n12652), .ZN(n12847) );
  NAND2_X1 U14396 ( .A1(n12847), .A2(n16057), .ZN(n12656) );
  AOI22_X1 U14397 ( .A1(n13708), .A2(n13578), .B1(n13576), .B2(n9880), .ZN(
        n12655) );
  OAI211_X1 U14398 ( .C1(n12657), .C2(n15959), .A(n12656), .B(n12655), .ZN(
        n12846) );
  INV_X1 U14399 ( .A(n12846), .ZN(n12662) );
  INV_X1 U14400 ( .A(n13700), .ZN(n13647) );
  AOI22_X1 U14401 ( .A1(n7188), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15909), 
        .B2(n12658), .ZN(n12659) );
  OAI21_X1 U14402 ( .B1(n12853), .B2(n13754), .A(n12659), .ZN(n12660) );
  AOI21_X1 U14403 ( .B1(n12847), .B2(n13647), .A(n12660), .ZN(n12661) );
  OAI21_X1 U14404 ( .B1(n12662), .B2(n7188), .A(n12661), .ZN(P3_U3221) );
  OAI21_X1 U14405 ( .B1(n12664), .B2(n7793), .A(n12663), .ZN(n12665) );
  NAND2_X1 U14406 ( .A1(n12666), .A2(n15535), .ZN(n12667) );
  XNOR2_X1 U14407 ( .A(n12871), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12668) );
  NOR2_X1 U14408 ( .A1(n12669), .A2(n12668), .ZN(n12870) );
  AOI211_X1 U14409 ( .C1(n12669), .C2(n12668), .A(n15859), .B(n12870), .ZN(
        n12682) );
  MUX2_X1 U14410 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n12866), .S(n12874), .Z(
        n12677) );
  AOI21_X1 U14411 ( .B1(n12671), .B2(P1_REG2_REG_14__SCAN_IN), .A(n12670), 
        .ZN(n12672) );
  NAND2_X1 U14412 ( .A1(n12672), .A2(n15535), .ZN(n12675) );
  XNOR2_X1 U14413 ( .A(n12672), .B(n15535), .ZN(n15533) );
  NOR2_X1 U14414 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15533), .ZN(n15532) );
  INV_X1 U14415 ( .A(n15532), .ZN(n12673) );
  NAND2_X1 U14416 ( .A1(n12675), .A2(n12673), .ZN(n12676) );
  AOI21_X1 U14417 ( .B1(n12874), .B2(n12866), .A(n15532), .ZN(n12674) );
  OAI211_X1 U14418 ( .C1(n12866), .C2(n12874), .A(n12675), .B(n12674), .ZN(
        n12880) );
  INV_X1 U14419 ( .A(n12880), .ZN(n12877) );
  AOI211_X1 U14420 ( .C1(n12677), .C2(n12676), .A(n15536), .B(n12877), .ZN(
        n12681) );
  NAND2_X1 U14421 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n16200)
         );
  INV_X1 U14422 ( .A(n16200), .ZN(n12678) );
  AOI21_X1 U14423 ( .B1(n15526), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n12678), 
        .ZN(n12679) );
  OAI21_X1 U14424 ( .B1(n15534), .B2(n12874), .A(n12679), .ZN(n12680) );
  OR3_X1 U14425 ( .A1(n12682), .A2(n12681), .A3(n12680), .ZN(P1_U3259) );
  OAI222_X1 U14426 ( .A1(n14370), .A2(n12685), .B1(n14378), .B2(n12684), .C1(
        P2_U3088), .C2(n12683), .ZN(P2_U3302) );
  XNOR2_X1 U14427 ( .A(n12686), .B(n12688), .ZN(n12844) );
  AOI21_X1 U14428 ( .B1(n12688), .B2(n12687), .A(n7316), .ZN(n12842) );
  OAI21_X1 U14429 ( .B1(n14431), .B2(n7298), .A(n12858), .ZN(n12840) );
  NAND2_X1 U14430 ( .A1(n14914), .A2(n14754), .ZN(n12690) );
  NAND2_X1 U14431 ( .A1(n15925), .A2(n14756), .ZN(n12689) );
  NAND2_X1 U14432 ( .A1(n12690), .A2(n12689), .ZN(n14733) );
  INV_X1 U14433 ( .A(n14733), .ZN(n12691) );
  OAI22_X1 U14434 ( .A1(n15894), .A2(n12691), .B1(n14735), .B2(n15931), .ZN(
        n12693) );
  NOR2_X1 U14435 ( .A1(n14431), .A2(n15933), .ZN(n12692) );
  AOI211_X1 U14436 ( .C1(n15894), .C2(P1_REG2_REG_15__SCAN_IN), .A(n12693), 
        .B(n12692), .ZN(n12694) );
  OAI21_X1 U14437 ( .B1(n15936), .B2(n12840), .A(n12694), .ZN(n12695) );
  AOI21_X1 U14438 ( .B1(n12842), .B2(n14972), .A(n12695), .ZN(n12696) );
  OAI21_X1 U14439 ( .B1(n12844), .B2(n14974), .A(n12696), .ZN(P1_U3278) );
  NAND2_X1 U14440 ( .A1(n13237), .A2(n12697), .ZN(n12955) );
  OR2_X1 U14441 ( .A1(n13237), .A2(n12697), .ZN(n12698) );
  NAND2_X1 U14442 ( .A1(n12955), .A2(n12698), .ZN(n13419) );
  INV_X1 U14443 ( .A(n13419), .ZN(n12702) );
  OAI21_X1 U14444 ( .B1(n12702), .B2(n12701), .A(n12957), .ZN(n12707) );
  OAI22_X1 U14445 ( .A1(n13226), .A2(n14189), .B1(n12822), .B2(n14191), .ZN(
        n12706) );
  NAND2_X1 U14446 ( .A1(n13224), .A2(n14018), .ZN(n12703) );
  XNOR2_X1 U14447 ( .A(n12826), .B(n13419), .ZN(n12947) );
  NOR2_X1 U14448 ( .A1(n12947), .A2(n14197), .ZN(n12705) );
  AOI211_X1 U14449 ( .C1(n14236), .C2(n12707), .A(n12706), .B(n12705), .ZN(
        n12946) );
  OR2_X1 U14450 ( .A1(n12709), .A2(n13237), .ZN(n12963) );
  INV_X1 U14451 ( .A(n12963), .ZN(n12708) );
  AOI211_X1 U14452 ( .C1(n13237), .C2(n12709), .A(n14319), .B(n12708), .ZN(
        n12944) );
  INV_X1 U14453 ( .A(n13237), .ZN(n12712) );
  AOI22_X1 U14454 ( .A1(n16156), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12710), 
        .B2(n16146), .ZN(n12711) );
  OAI21_X1 U14455 ( .B1(n12712), .B2(n14231), .A(n12711), .ZN(n12715) );
  NOR2_X1 U14456 ( .A1(n12947), .A2(n12713), .ZN(n12714) );
  AOI211_X1 U14457 ( .C1(n12944), .C2(n16150), .A(n12715), .B(n12714), .ZN(
        n12716) );
  OAI21_X1 U14458 ( .B1(n12946), .B2(n16156), .A(n12716), .ZN(P2_U3253) );
  AOI21_X1 U14459 ( .B1(n12720), .B2(P2_REG2_REG_17__SCAN_IN), .A(n12717), 
        .ZN(n12718) );
  NAND2_X1 U14460 ( .A1(n12718), .A2(n12923), .ZN(n12919) );
  OAI21_X1 U14461 ( .B1(n12718), .B2(n12923), .A(n12919), .ZN(n12719) );
  NOR2_X1 U14462 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n12719), .ZN(n12917) );
  AOI21_X1 U14463 ( .B1(n12719), .B2(P2_REG2_REG_18__SCAN_IN), .A(n12917), 
        .ZN(n12730) );
  INV_X1 U14464 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U14465 ( .A1(n12722), .A2(n12721), .B1(n12720), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n12924) );
  XNOR2_X1 U14466 ( .A(n12924), .B(n12728), .ZN(n12723) );
  NAND2_X1 U14467 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n12723), .ZN(n12922) );
  OAI211_X1 U14468 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n12723), .A(n15494), 
        .B(n12922), .ZN(n12725) );
  NAND2_X1 U14469 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n12724)
         );
  OAI211_X1 U14470 ( .C1(n15441), .C2(n12726), .A(n12725), .B(n12724), .ZN(
        n12727) );
  AOI21_X1 U14471 ( .B1(n12728), .B2(n15504), .A(n12727), .ZN(n12729) );
  OAI21_X1 U14472 ( .B1(n12730), .B2(n15412), .A(n12729), .ZN(P2_U3232) );
  INV_X1 U14473 ( .A(n12731), .ZN(n12736) );
  AOI21_X1 U14474 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15392), .A(n12732), 
        .ZN(n12733) );
  OAI21_X1 U14475 ( .B1(n12736), .B2(n15160), .A(n12733), .ZN(P1_U3332) );
  NAND2_X1 U14476 ( .A1(n14376), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12735) );
  OR2_X1 U14477 ( .A1(n12734), .A2(P2_U3088), .ZN(n13458) );
  OAI211_X1 U14478 ( .C1(n12736), .C2(n14378), .A(n12735), .B(n13458), .ZN(
        P2_U3304) );
  AOI21_X1 U14479 ( .B1(n12739), .B2(n12738), .A(n12737), .ZN(n12744) );
  AOI22_X1 U14480 ( .A1(n14089), .A2(n13244), .B1(n14015), .B2(n14091), .ZN(
        n12824) );
  INV_X1 U14481 ( .A(n12832), .ZN(n12740) );
  AOI22_X1 U14482 ( .A1(n13994), .A2(n12740), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12741) );
  OAI21_X1 U14483 ( .B1(n13984), .B2(n12824), .A(n12741), .ZN(n12742) );
  AOI21_X1 U14484 ( .B1(n13249), .B2(n13999), .A(n12742), .ZN(n12743) );
  OAI21_X1 U14485 ( .B1(n12744), .B2(n14001), .A(n12743), .ZN(P2_U3187) );
  OAI21_X1 U14486 ( .B1(n12747), .B2(n12746), .A(n12745), .ZN(n16127) );
  INV_X1 U14487 ( .A(n16127), .ZN(n12756) );
  XNOR2_X1 U14488 ( .A(n12749), .B(n12748), .ZN(n12750) );
  OAI222_X1 U14489 ( .A1(n15962), .A2(n12784), .B1(n15960), .B2(n12776), .C1(
        n12750), .C2(n15959), .ZN(n16125) );
  NAND2_X1 U14490 ( .A1(n16125), .A2(n13715), .ZN(n12755) );
  INV_X1 U14491 ( .A(n16124), .ZN(n12753) );
  INV_X1 U14492 ( .A(n12786), .ZN(n12751) );
  OAI22_X1 U14493 ( .A1(n13715), .A2(n15755), .B1(n12751), .B2(n15967), .ZN(
        n12752) );
  AOI21_X1 U14494 ( .B1(n12753), .B2(n13696), .A(n12752), .ZN(n12754) );
  OAI211_X1 U14495 ( .C1(n13717), .C2(n12756), .A(n12755), .B(n12754), .ZN(
        P3_U3220) );
  INV_X1 U14496 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U14497 ( .A1(n12757), .A2(n14302), .B1(n14343), .B2(n13216), .ZN(
        n12758) );
  OAI211_X1 U14498 ( .C1(n12760), .C2(n15897), .A(n12759), .B(n12758), .ZN(
        n12763) );
  NAND2_X1 U14499 ( .A1(n12763), .A2(n16192), .ZN(n12761) );
  OAI21_X1 U14500 ( .B1(n16192), .B2(n12762), .A(n12761), .ZN(P2_U3460) );
  NAND2_X1 U14501 ( .A1(n12763), .A2(n16189), .ZN(n12764) );
  OAI21_X1 U14502 ( .B1(n16189), .B2(n10466), .A(n12764), .ZN(P2_U3509) );
  NAND2_X1 U14503 ( .A1(n12765), .A2(n16012), .ZN(n12767) );
  AOI21_X1 U14504 ( .B1(n16177), .B2(n15126), .A(n16176), .ZN(n12766) );
  OAI21_X1 U14505 ( .B1(n7298), .B2(n12767), .A(n12766), .ZN(n12768) );
  AOI21_X1 U14506 ( .B1(n12769), .B2(n16139), .A(n12768), .ZN(n12770) );
  OAI21_X1 U14507 ( .B1(n16134), .B2(n12771), .A(n12770), .ZN(n12774) );
  NAND2_X1 U14508 ( .A1(n12774), .A2(n16141), .ZN(n12772) );
  OAI21_X1 U14509 ( .B1(n16141), .B2(n12773), .A(n12772), .ZN(P1_U3542) );
  NAND2_X1 U14510 ( .A1(n12774), .A2(n15984), .ZN(n12775) );
  OAI21_X1 U14511 ( .B1(n15984), .B2(n8782), .A(n12775), .ZN(P1_U3501) );
  XNOR2_X1 U14512 ( .A(n16124), .B(n13119), .ZN(n12807) );
  XNOR2_X1 U14513 ( .A(n12807), .B(n12808), .ZN(n12780) );
  NAND2_X1 U14514 ( .A1(n12777), .A2(n12776), .ZN(n12781) );
  NAND2_X1 U14515 ( .A1(n12779), .A2(n12778), .ZN(n12814) );
  INV_X1 U14516 ( .A(n12814), .ZN(n12810) );
  AOI21_X1 U14517 ( .B1(n12779), .B2(n12781), .A(n12780), .ZN(n12782) );
  OR3_X1 U14518 ( .A1(n12810), .A2(n12782), .A3(n13566), .ZN(n12788) );
  NOR2_X1 U14519 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9318), .ZN(n15753) );
  AOI21_X1 U14520 ( .B1(n13577), .B2(n13549), .A(n15753), .ZN(n12783) );
  OAI21_X1 U14521 ( .B1(n12784), .B2(n13551), .A(n12783), .ZN(n12785) );
  AOI21_X1 U14522 ( .B1(n12786), .B2(n13564), .A(n12785), .ZN(n12787) );
  OAI211_X1 U14523 ( .C1(n13561), .C2(n16124), .A(n12788), .B(n12787), .ZN(
        P3_U3174) );
  XNOR2_X1 U14524 ( .A(n12789), .B(n12793), .ZN(n12792) );
  NAND2_X1 U14525 ( .A1(n13576), .A2(n13708), .ZN(n12790) );
  OAI21_X1 U14526 ( .B1(n12983), .B2(n15962), .A(n12790), .ZN(n12791) );
  AOI21_X1 U14527 ( .B1(n12792), .B2(n13705), .A(n12791), .ZN(n16163) );
  OR2_X1 U14528 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  NAND2_X1 U14529 ( .A1(n12974), .A2(n12795), .ZN(n16161) );
  NOR2_X1 U14530 ( .A1(n16158), .A2(n13754), .ZN(n12799) );
  INV_X1 U14531 ( .A(n12819), .ZN(n12796) );
  OAI22_X1 U14532 ( .A1(n13715), .A2(n12797), .B1(n12796), .B2(n15967), .ZN(
        n12798) );
  AOI211_X1 U14533 ( .C1(n16161), .C2(n13757), .A(n12799), .B(n12798), .ZN(
        n12800) );
  OAI21_X1 U14534 ( .B1(n16163), .B2(n7188), .A(n12800), .ZN(P3_U3219) );
  OAI222_X1 U14535 ( .A1(n13131), .A2(n12801), .B1(n7187), .B2(P3_U3151), .C1(
        n15177), .C2(n13880), .ZN(P3_U3267) );
  AOI22_X1 U14536 ( .A1(n12802), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14376), .ZN(n12803) );
  OAI21_X1 U14537 ( .B1(n12806), .B2(n14378), .A(n12803), .ZN(P2_U3301) );
  AOI22_X1 U14538 ( .A1(n12804), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n15392), .ZN(n12805) );
  OAI21_X1 U14539 ( .B1(n12806), .B2(n15160), .A(n12805), .ZN(P1_U3329) );
  INV_X1 U14540 ( .A(n12807), .ZN(n12809) );
  NOR2_X1 U14541 ( .A1(n12809), .A2(n12808), .ZN(n12811) );
  XNOR2_X1 U14542 ( .A(n16158), .B(n13119), .ZN(n12886) );
  XNOR2_X1 U14543 ( .A(n12886), .B(n13575), .ZN(n12812) );
  OAI21_X1 U14544 ( .B1(n12810), .B2(n12811), .A(n12812), .ZN(n12815) );
  NOR2_X1 U14545 ( .A1(n12812), .A2(n12811), .ZN(n12813) );
  AOI21_X1 U14546 ( .B1(n12815), .B2(n12888), .A(n13566), .ZN(n12816) );
  INV_X1 U14547 ( .A(n12816), .ZN(n12821) );
  INV_X1 U14548 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U14549 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15335), .ZN(n15769) );
  AOI21_X1 U14550 ( .B1(n13576), .B2(n13549), .A(n15769), .ZN(n12817) );
  OAI21_X1 U14551 ( .B1(n12983), .B2(n13551), .A(n12817), .ZN(n12818) );
  AOI21_X1 U14552 ( .B1(n13564), .B2(n12819), .A(n12818), .ZN(n12820) );
  OAI211_X1 U14553 ( .C1(n13561), .C2(n16158), .A(n12821), .B(n12820), .ZN(
        P3_U3155) );
  XNOR2_X1 U14554 ( .A(n16148), .B(n13244), .ZN(n13420) );
  NAND2_X1 U14555 ( .A1(n16148), .A2(n12822), .ZN(n12823) );
  XNOR2_X1 U14556 ( .A(n13249), .B(n14016), .ZN(n13421) );
  XNOR2_X1 U14557 ( .A(n12900), .B(n12830), .ZN(n12825) );
  OAI21_X1 U14558 ( .B1(n12825), .B2(n14214), .A(n12824), .ZN(n16184) );
  INV_X1 U14559 ( .A(n16184), .ZN(n12838) );
  AND2_X1 U14560 ( .A1(n13237), .A2(n14017), .ZN(n12827) );
  OR2_X1 U14561 ( .A1(n13237), .A2(n14017), .ZN(n12828) );
  NAND2_X1 U14562 ( .A1(n16148), .A2(n13244), .ZN(n12829) );
  OAI21_X1 U14563 ( .B1(n12831), .B2(n12830), .A(n12898), .ZN(n16187) );
  INV_X1 U14564 ( .A(n13249), .ZN(n16183) );
  OAI211_X1 U14565 ( .C1(n16183), .C2(n12962), .A(n14302), .B(n12903), .ZN(
        n16181) );
  INV_X1 U14566 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12833) );
  OAI22_X1 U14567 ( .A1(n16041), .A2(n12833), .B1(n12832), .B2(n16038), .ZN(
        n12834) );
  AOI21_X1 U14568 ( .B1(n13249), .B2(n16147), .A(n12834), .ZN(n12835) );
  OAI21_X1 U14569 ( .B1(n16181), .B2(n16045), .A(n12835), .ZN(n12836) );
  AOI21_X1 U14570 ( .B1(n16187), .B2(n14151), .A(n12836), .ZN(n12837) );
  OAI21_X1 U14571 ( .B1(n16156), .B2(n12838), .A(n12837), .ZN(P2_U3251) );
  AOI21_X1 U14572 ( .B1(n14738), .B2(n15126), .A(n14733), .ZN(n12839) );
  OAI21_X1 U14573 ( .B1(n12840), .B2(n16077), .A(n12839), .ZN(n12841) );
  AOI21_X1 U14574 ( .B1(n12842), .B2(n16019), .A(n12841), .ZN(n12843) );
  OAI21_X1 U14575 ( .B1(n16015), .B2(n12844), .A(n12843), .ZN(n15149) );
  NAND2_X1 U14576 ( .A1(n15149), .A2(n16141), .ZN(n12845) );
  OAI21_X1 U14577 ( .B1(n16141), .B2(n8798), .A(n12845), .ZN(P1_U3543) );
  INV_X1 U14578 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n12848) );
  AOI21_X1 U14579 ( .B1(n16103), .B2(n12847), .A(n12846), .ZN(n12850) );
  MUX2_X1 U14580 ( .A(n12848), .B(n12850), .S(n16169), .Z(n12849) );
  OAI21_X1 U14581 ( .B1(n13864), .B2(n12853), .A(n12849), .ZN(P3_U3426) );
  MUX2_X1 U14582 ( .A(n12851), .B(n12850), .S(n16165), .Z(n12852) );
  OAI21_X1 U14583 ( .B1(n13806), .B2(n12853), .A(n12852), .ZN(P3_U3471) );
  XOR2_X1 U14584 ( .A(n12856), .B(n12854), .Z(n15132) );
  OAI21_X1 U14585 ( .B1(n12857), .B2(n12856), .A(n12855), .ZN(n15130) );
  NAND2_X1 U14586 ( .A1(n12858), .A2(n16199), .ZN(n12859) );
  NAND2_X1 U14587 ( .A1(n12936), .A2(n12859), .ZN(n15128) );
  NOR2_X1 U14588 ( .A1(n15128), .A2(n15936), .ZN(n12868) );
  NAND2_X1 U14589 ( .A1(n16199), .A2(n15026), .ZN(n12865) );
  NAND2_X1 U14590 ( .A1(n14914), .A2(n14753), .ZN(n12861) );
  NAND2_X1 U14591 ( .A1(n15925), .A2(n14755), .ZN(n12860) );
  NAND2_X1 U14592 ( .A1(n12861), .A2(n12860), .ZN(n16198) );
  INV_X1 U14593 ( .A(n16198), .ZN(n12862) );
  OAI22_X1 U14594 ( .A1(n15894), .A2(n12862), .B1(n16202), .B2(n15931), .ZN(
        n12863) );
  INV_X1 U14595 ( .A(n12863), .ZN(n12864) );
  OAI211_X1 U14596 ( .C1(n15942), .C2(n12866), .A(n12865), .B(n12864), .ZN(
        n12867) );
  AOI211_X1 U14597 ( .C1(n15130), .C2(n15001), .A(n12868), .B(n12867), .ZN(
        n12869) );
  OAI21_X1 U14598 ( .B1(n15003), .B2(n15132), .A(n12869), .ZN(P1_U3277) );
  AOI21_X1 U14599 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n12871), .A(n12870), 
        .ZN(n12873) );
  XNOR2_X1 U14600 ( .A(n14814), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n12872) );
  AOI211_X1 U14601 ( .C1(n12873), .C2(n12872), .A(n15859), .B(n14813), .ZN(
        n12885) );
  NOR2_X1 U14602 ( .A1(n12874), .A2(n12866), .ZN(n12878) );
  NAND2_X1 U14603 ( .A1(n14814), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n12876) );
  INV_X1 U14604 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14812) );
  NAND2_X1 U14605 ( .A1(n14811), .A2(n14812), .ZN(n12875) );
  OAI211_X1 U14606 ( .C1(n12877), .C2(n12878), .A(n12876), .B(n12875), .ZN(
        n14810) );
  AOI21_X1 U14607 ( .B1(n14811), .B2(P1_REG2_REG_17__SCAN_IN), .A(n12878), 
        .ZN(n12879) );
  OAI211_X1 U14608 ( .C1(P1_REG2_REG_17__SCAN_IN), .C2(n14811), .A(n12880), 
        .B(n12879), .ZN(n12881) );
  NAND3_X1 U14609 ( .A1(n14810), .A2(n15869), .A3(n12881), .ZN(n12883) );
  AND2_X1 U14610 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14638) );
  AOI21_X1 U14611 ( .B1(n15526), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14638), 
        .ZN(n12882) );
  OAI211_X1 U14612 ( .C1(n15534), .C2(n14811), .A(n12883), .B(n12882), .ZN(
        n12884) );
  OR2_X1 U14613 ( .A1(n12885), .A2(n12884), .ZN(P1_U3260) );
  INV_X1 U14614 ( .A(n13815), .ZN(n12979) );
  XNOR2_X1 U14615 ( .A(n13815), .B(n13119), .ZN(n12982) );
  XNOR2_X1 U14616 ( .A(n12982), .B(n12983), .ZN(n12890) );
  AOI21_X1 U14617 ( .B1(n12889), .B2(n12890), .A(n13566), .ZN(n12892) );
  INV_X1 U14618 ( .A(n12890), .ZN(n12891) );
  NAND2_X1 U14619 ( .A1(n12892), .A2(n12985), .ZN(n12896) );
  INV_X1 U14620 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15384) );
  NOR2_X1 U14621 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15384), .ZN(n15787) );
  AOI21_X1 U14622 ( .B1(n13575), .B2(n13549), .A(n15787), .ZN(n12893) );
  OAI21_X1 U14623 ( .B1(n13746), .B2(n13551), .A(n12893), .ZN(n12894) );
  AOI21_X1 U14624 ( .B1(n13564), .B2(n12977), .A(n12894), .ZN(n12895) );
  OAI211_X1 U14625 ( .C1(n12979), .C2(n13561), .A(n12896), .B(n12895), .ZN(
        P3_U3181) );
  OR2_X1 U14626 ( .A1(n13249), .A2(n14016), .ZN(n12897) );
  XNOR2_X1 U14627 ( .A(n14342), .B(n14015), .ZN(n13423) );
  XNOR2_X1 U14628 ( .A(n12992), .B(n13423), .ZN(n14345) );
  OR2_X1 U14629 ( .A1(n13249), .A2(n13251), .ZN(n12899) );
  INV_X1 U14630 ( .A(n13423), .ZN(n12991) );
  OAI211_X1 U14631 ( .C1(n7318), .C2(n13423), .A(n14236), .B(n13000), .ZN(
        n12901) );
  AOI22_X1 U14632 ( .A1(n14014), .A2(n14091), .B1(n14016), .B2(n14089), .ZN(
        n12913) );
  NAND2_X1 U14633 ( .A1(n12901), .A2(n12913), .ZN(n14340) );
  INV_X1 U14634 ( .A(n14342), .ZN(n12906) );
  INV_X1 U14635 ( .A(n12994), .ZN(n12902) );
  AOI211_X1 U14636 ( .C1(n14342), .C2(n12903), .A(n14319), .B(n12902), .ZN(
        n14341) );
  NAND2_X1 U14637 ( .A1(n14341), .A2(n16150), .ZN(n12905) );
  AOI22_X1 U14638 ( .A1(n16156), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12911), 
        .B2(n16146), .ZN(n12904) );
  OAI211_X1 U14639 ( .C1(n12906), .C2(n14231), .A(n12905), .B(n12904), .ZN(
        n12907) );
  AOI21_X1 U14640 ( .B1(n14340), .B2(n16041), .A(n12907), .ZN(n12908) );
  OAI21_X1 U14641 ( .B1(n14345), .B2(n14244), .A(n12908), .ZN(P2_U3250) );
  XNOR2_X1 U14642 ( .A(n12910), .B(n12909), .ZN(n12916) );
  AND2_X1 U14643 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n15470) );
  AOI21_X1 U14644 ( .B1(n13994), .B2(n12911), .A(n15470), .ZN(n12912) );
  OAI21_X1 U14645 ( .B1(n13984), .B2(n12913), .A(n12912), .ZN(n12914) );
  AOI21_X1 U14646 ( .B1(n14342), .B2(n13999), .A(n12914), .ZN(n12915) );
  OAI21_X1 U14647 ( .B1(n12916), .B2(n14001), .A(n12915), .ZN(P2_U3213) );
  MUX2_X1 U14648 ( .A(n10750), .B(P2_REG2_REG_19__SCAN_IN), .S(n13024), .Z(
        n12921) );
  INV_X1 U14649 ( .A(n12917), .ZN(n12918) );
  NAND2_X1 U14650 ( .A1(n12919), .A2(n12918), .ZN(n12920) );
  XOR2_X1 U14651 ( .A(n12921), .B(n12920), .Z(n12931) );
  OAI21_X1 U14652 ( .B1(n12924), .B2(n12923), .A(n12922), .ZN(n12926) );
  XNOR2_X1 U14653 ( .A(n13024), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n12925) );
  XNOR2_X1 U14654 ( .A(n12926), .B(n12925), .ZN(n12928) );
  NAND2_X1 U14655 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13905)
         );
  NAND2_X1 U14656 ( .A1(n15502), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n12927) );
  OAI211_X1 U14657 ( .C1(n15508), .C2(n12928), .A(n13905), .B(n12927), .ZN(
        n12929) );
  AOI21_X1 U14658 ( .B1(n10458), .B2(n15504), .A(n12929), .ZN(n12930) );
  OAI21_X1 U14659 ( .B1(n12931), .B2(n15412), .A(n12930), .ZN(P2_U3233) );
  OAI21_X1 U14660 ( .B1(n7333), .B2(n8837), .A(n12932), .ZN(n15125) );
  OAI21_X1 U14661 ( .B1(n12935), .B2(n12934), .A(n12933), .ZN(n15123) );
  INV_X1 U14662 ( .A(n14449), .ZN(n15121) );
  NAND2_X1 U14663 ( .A1(n14449), .A2(n12936), .ZN(n15117) );
  NAND3_X1 U14664 ( .A1(n15118), .A2(n14958), .A3(n15117), .ZN(n12941) );
  NAND2_X1 U14665 ( .A1(n14752), .A2(n14914), .ZN(n12938) );
  NAND2_X1 U14666 ( .A1(n15925), .A2(n14754), .ZN(n12937) );
  NAND2_X1 U14667 ( .A1(n12938), .A2(n12937), .ZN(n14639) );
  INV_X1 U14668 ( .A(n14639), .ZN(n15119) );
  OAI22_X1 U14669 ( .A1(n15894), .A2(n15119), .B1(n14636), .B2(n15931), .ZN(
        n12939) );
  AOI21_X1 U14670 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14997), .A(n12939), 
        .ZN(n12940) );
  OAI211_X1 U14671 ( .C1(n15121), .C2(n15933), .A(n12941), .B(n12940), .ZN(
        n12942) );
  AOI21_X1 U14672 ( .B1(n15123), .B2(n14972), .A(n12942), .ZN(n12943) );
  OAI21_X1 U14673 ( .B1(n15125), .B2(n14974), .A(n12943), .ZN(P1_U3276) );
  INV_X1 U14674 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n12949) );
  AOI21_X1 U14675 ( .B1(n14343), .B2(n13237), .A(n12944), .ZN(n12945) );
  OAI211_X1 U14676 ( .C1(n15897), .C2(n12947), .A(n12946), .B(n12945), .ZN(
        n12950) );
  NAND2_X1 U14677 ( .A1(n12950), .A2(n16192), .ZN(n12948) );
  OAI21_X1 U14678 ( .B1(n16192), .B2(n12949), .A(n12948), .ZN(P2_U3466) );
  NAND2_X1 U14679 ( .A1(n12950), .A2(n16189), .ZN(n12951) );
  OAI21_X1 U14680 ( .B1(n16189), .B2(n12420), .A(n12951), .ZN(P2_U3511) );
  INV_X1 U14681 ( .A(n12952), .ZN(n12953) );
  AOI21_X1 U14682 ( .B1(n13420), .B2(n12954), .A(n12953), .ZN(n16152) );
  INV_X1 U14683 ( .A(n16152), .ZN(n12965) );
  INV_X1 U14684 ( .A(n13420), .ZN(n12956) );
  NAND3_X1 U14685 ( .A1(n12957), .A2(n12956), .A3(n12955), .ZN(n12958) );
  AOI21_X1 U14686 ( .B1(n12959), .B2(n12958), .A(n14214), .ZN(n12961) );
  AOI211_X1 U14687 ( .C1(n16152), .C2(n14121), .A(n12961), .B(n12960), .ZN(
        n16155) );
  AOI211_X1 U14688 ( .C1(n16148), .C2(n12963), .A(n14319), .B(n12962), .ZN(
        n16149) );
  AOI21_X1 U14689 ( .B1(n14343), .B2(n16148), .A(n16149), .ZN(n12964) );
  OAI211_X1 U14690 ( .C1(n15897), .C2(n12965), .A(n16155), .B(n12964), .ZN(
        n12967) );
  NAND2_X1 U14691 ( .A1(n12967), .A2(n16192), .ZN(n12966) );
  OAI21_X1 U14692 ( .B1(n16192), .B2(n10653), .A(n12966), .ZN(P2_U3469) );
  NAND2_X1 U14693 ( .A1(n12967), .A2(n16189), .ZN(n12968) );
  OAI21_X1 U14694 ( .B1(n16189), .B2(n12422), .A(n12968), .ZN(P2_U3512) );
  OAI21_X1 U14695 ( .B1(n12971), .B2(n9360), .A(n12970), .ZN(n12972) );
  AOI222_X1 U14696 ( .A1(n13705), .A2(n12972), .B1(n13575), .B2(n13708), .C1(
        n13573), .C2(n9880), .ZN(n13818) );
  NAND3_X1 U14697 ( .A1(n12974), .A2(n9360), .A3(n12973), .ZN(n12975) );
  NAND2_X1 U14698 ( .A1(n12976), .A2(n12975), .ZN(n13816) );
  AOI22_X1 U14699 ( .A1(n7188), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15909), 
        .B2(n12977), .ZN(n12978) );
  OAI21_X1 U14700 ( .B1(n12979), .B2(n13754), .A(n12978), .ZN(n12980) );
  AOI21_X1 U14701 ( .B1(n13816), .B2(n13757), .A(n12980), .ZN(n12981) );
  OAI21_X1 U14702 ( .B1(n13818), .B2(n7188), .A(n12981), .ZN(P3_U3218) );
  INV_X1 U14703 ( .A(n12982), .ZN(n12984) );
  XNOR2_X1 U14704 ( .A(n13811), .B(n13119), .ZN(n13084) );
  XNOR2_X1 U14705 ( .A(n13084), .B(n13573), .ZN(n13082) );
  XNOR2_X1 U14706 ( .A(n13083), .B(n13082), .ZN(n12990) );
  NAND2_X1 U14707 ( .A1(n13574), .A2(n13549), .ZN(n12986) );
  NAND2_X1 U14708 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n15811)
         );
  OAI211_X1 U14709 ( .C1(n13734), .C2(n13551), .A(n12986), .B(n15811), .ZN(
        n12988) );
  INV_X1 U14710 ( .A(n13811), .ZN(n13021) );
  NOR2_X1 U14711 ( .A1(n13021), .A2(n13561), .ZN(n12987) );
  AOI211_X1 U14712 ( .C1(n13019), .C2(n13564), .A(n12988), .B(n12987), .ZN(
        n12989) );
  OAI21_X1 U14713 ( .B1(n12990), .B2(n13566), .A(n12989), .ZN(P3_U3166) );
  OR2_X1 U14714 ( .A1(n14342), .A2(n14015), .ZN(n12993) );
  INV_X1 U14715 ( .A(n14014), .ZN(n13040) );
  XNOR2_X1 U14716 ( .A(n14337), .B(n13040), .ZN(n13425) );
  INV_X1 U14717 ( .A(n13425), .ZN(n13001) );
  OAI21_X1 U14718 ( .B1(n7213), .B2(n13425), .A(n7315), .ZN(n14339) );
  AOI211_X1 U14719 ( .C1(n14337), .C2(n12994), .A(n14319), .B(n14228), .ZN(
        n14336) );
  NOR2_X1 U14720 ( .A1(n7762), .A2(n14231), .ZN(n12997) );
  OAI22_X1 U14721 ( .A1(n16041), .A2(n12995), .B1(n13930), .B2(n16038), .ZN(
        n12996) );
  AOI211_X1 U14722 ( .C1(n14336), .C2(n16150), .A(n12997), .B(n12996), .ZN(
        n13006) );
  INV_X1 U14723 ( .A(n14015), .ZN(n12998) );
  OR2_X1 U14724 ( .A1(n14342), .A2(n12998), .ZN(n12999) );
  NAND2_X1 U14725 ( .A1(n13000), .A2(n12999), .ZN(n13002) );
  NAND2_X1 U14726 ( .A1(n13002), .A2(n13001), .ZN(n13042) );
  OAI211_X1 U14727 ( .C1(n13002), .C2(n13001), .A(n13042), .B(n14236), .ZN(
        n13004) );
  AND2_X1 U14728 ( .A1(n14015), .A2(n14089), .ZN(n13003) );
  AOI21_X1 U14729 ( .B1(n14013), .B2(n14091), .A(n13003), .ZN(n13932) );
  NAND2_X1 U14730 ( .A1(n13004), .A2(n13932), .ZN(n14335) );
  NAND2_X1 U14731 ( .A1(n14335), .A2(n16041), .ZN(n13005) );
  OAI211_X1 U14732 ( .C1(n14339), .C2(n14244), .A(n13006), .B(n13005), .ZN(
        P2_U3249) );
  INV_X1 U14733 ( .A(n13007), .ZN(n13010) );
  OAI222_X1 U14734 ( .A1(n13009), .A2(P1_U3086), .B1(n15160), .B2(n13010), 
        .C1(n13008), .C2(n15157), .ZN(P1_U3328) );
  OAI222_X1 U14735 ( .A1(n14370), .A2(n13011), .B1(n14378), .B2(n13010), .C1(
        n13455), .C2(P2_U3088), .ZN(P2_U3300) );
  NAND3_X1 U14736 ( .A1(n12970), .A2(n13017), .A3(n13012), .ZN(n13013) );
  NAND2_X1 U14737 ( .A1(n13014), .A2(n13013), .ZN(n13015) );
  AOI222_X1 U14738 ( .A1(n13705), .A2(n13015), .B1(n13572), .B2(n9880), .C1(
        n13574), .C2(n13708), .ZN(n13814) );
  OAI21_X1 U14739 ( .B1(n13018), .B2(n13017), .A(n13016), .ZN(n13812) );
  AOI22_X1 U14740 ( .A1(n7188), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15909), 
        .B2(n13019), .ZN(n13020) );
  OAI21_X1 U14741 ( .B1(n13021), .B2(n13754), .A(n13020), .ZN(n13022) );
  AOI21_X1 U14742 ( .B1(n13812), .B2(n13757), .A(n13022), .ZN(n13023) );
  OAI21_X1 U14743 ( .B1(n13814), .B2(n7188), .A(n13023), .ZN(P3_U3217) );
  OAI222_X1 U14744 ( .A1(n14370), .A2(n13026), .B1(n14378), .B2(n13025), .C1(
        n13024), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U14745 ( .A(n14332), .B(n14013), .ZN(n14238) );
  INV_X1 U14746 ( .A(n14238), .ZN(n14225) );
  OR2_X1 U14747 ( .A1(n14332), .A2(n14013), .ZN(n13027) );
  NAND2_X1 U14748 ( .A1(n14224), .A2(n13027), .ZN(n14210) );
  XNOR2_X1 U14749 ( .A(n14327), .B(n14012), .ZN(n14211) );
  INV_X1 U14750 ( .A(n14211), .ZN(n13028) );
  OR2_X1 U14751 ( .A1(n14327), .A2(n14012), .ZN(n13029) );
  NAND2_X1 U14752 ( .A1(n14317), .A2(n14011), .ZN(n13031) );
  OR2_X1 U14753 ( .A1(n14317), .A2(n14011), .ZN(n13030) );
  NAND2_X1 U14754 ( .A1(n13031), .A2(n13030), .ZN(n14194) );
  NAND2_X1 U14755 ( .A1(n14196), .A2(n13031), .ZN(n14175) );
  OR2_X1 U14756 ( .A1(n14314), .A2(n14010), .ZN(n13032) );
  NAND2_X1 U14757 ( .A1(n14314), .A2(n14010), .ZN(n13033) );
  AND2_X1 U14758 ( .A1(n14309), .A2(n14009), .ZN(n13035) );
  XNOR2_X1 U14759 ( .A(n14301), .B(n14008), .ZN(n14149) );
  XNOR2_X1 U14760 ( .A(n14295), .B(n14007), .ZN(n13430) );
  NAND2_X1 U14761 ( .A1(n14295), .A2(n14007), .ZN(n13036) );
  XNOR2_X1 U14762 ( .A(n14290), .B(n14006), .ZN(n13428) );
  NAND2_X1 U14763 ( .A1(n14290), .A2(n14006), .ZN(n13037) );
  NAND2_X1 U14764 ( .A1(n14285), .A2(n14090), .ZN(n13401) );
  NAND2_X1 U14765 ( .A1(n14278), .A2(n14005), .ZN(n13039) );
  XNOR2_X1 U14766 ( .A(n14271), .B(n14044), .ZN(n13433) );
  OR2_X1 U14767 ( .A1(n14337), .A2(n13040), .ZN(n13041) );
  NAND2_X1 U14768 ( .A1(n13042), .A2(n13041), .ZN(n14239) );
  NAND2_X1 U14769 ( .A1(n14239), .A2(n14238), .ZN(n14237) );
  INV_X1 U14770 ( .A(n14013), .ZN(n13043) );
  OR2_X1 U14771 ( .A1(n14332), .A2(n13043), .ZN(n13044) );
  NAND2_X1 U14772 ( .A1(n14237), .A2(n13044), .ZN(n14212) );
  NAND2_X1 U14773 ( .A1(n14327), .A2(n14190), .ZN(n13045) );
  NAND2_X1 U14774 ( .A1(n14212), .A2(n13045), .ZN(n13047) );
  OR2_X1 U14775 ( .A1(n14327), .A2(n14190), .ZN(n13046) );
  INV_X1 U14776 ( .A(n14011), .ZN(n13049) );
  NOR2_X1 U14777 ( .A1(n14317), .A2(n13049), .ZN(n13048) );
  NAND2_X1 U14778 ( .A1(n14317), .A2(n13049), .ZN(n13050) );
  INV_X1 U14779 ( .A(n14010), .ZN(n14192) );
  AND2_X1 U14780 ( .A1(n14314), .A2(n14192), .ZN(n13051) );
  INV_X1 U14781 ( .A(n14009), .ZN(n14144) );
  NOR2_X1 U14782 ( .A1(n14309), .A2(n14144), .ZN(n13052) );
  INV_X1 U14783 ( .A(n14309), .ZN(n14172) );
  NAND2_X1 U14784 ( .A1(n14152), .A2(n14008), .ZN(n13053) );
  NAND2_X1 U14785 ( .A1(n14147), .A2(n13053), .ZN(n14128) );
  NAND2_X1 U14786 ( .A1(n14295), .A2(n14145), .ZN(n13054) );
  OR2_X1 U14787 ( .A1(n14295), .A2(n14145), .ZN(n13055) );
  INV_X1 U14788 ( .A(n14006), .ZN(n14100) );
  NAND2_X1 U14789 ( .A1(n14290), .A2(n14100), .ZN(n13057) );
  NAND2_X1 U14790 ( .A1(n14108), .A2(n14090), .ZN(n13058) );
  OR2_X1 U14791 ( .A1(n14108), .A2(n14090), .ZN(n13059) );
  XNOR2_X1 U14792 ( .A(n14278), .B(n14005), .ZN(n14087) );
  NAND2_X1 U14793 ( .A1(n14278), .A2(n14101), .ZN(n13060) );
  INV_X1 U14794 ( .A(n13433), .ZN(n14042) );
  OAI22_X1 U14795 ( .A1(n13889), .A2(n14191), .B1(n14101), .B2(n14189), .ZN(
        n13061) );
  INV_X1 U14796 ( .A(n13061), .ZN(n13062) );
  INV_X1 U14797 ( .A(n14332), .ZN(n14232) );
  OR2_X1 U14798 ( .A1(n14327), .A2(n14229), .ZN(n14216) );
  INV_X1 U14799 ( .A(n14314), .ZN(n14185) );
  OR2_X2 U14800 ( .A1(n14102), .A2(n14278), .ZN(n14082) );
  NAND2_X1 U14801 ( .A1(n14082), .A2(n14271), .ZN(n13064) );
  NAND2_X1 U14802 ( .A1(n14075), .A2(n13064), .ZN(n14273) );
  AOI22_X1 U14803 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(n16156), .B1(n13887), 
        .B2(n16146), .ZN(n13066) );
  NAND2_X1 U14804 ( .A1(n14271), .A2(n16147), .ZN(n13065) );
  OAI211_X1 U14805 ( .C1(n14273), .C2(n14206), .A(n13066), .B(n13065), .ZN(
        n13067) );
  AOI21_X1 U14806 ( .B1(n13063), .B2(n16151), .A(n13067), .ZN(n13068) );
  OAI21_X1 U14807 ( .B1(n14276), .B2(n16156), .A(n13068), .ZN(P2_U3238) );
  XNOR2_X1 U14808 ( .A(n13070), .B(n13069), .ZN(n13071) );
  OAI22_X1 U14809 ( .A1(n15012), .A2(n14531), .B1(n14587), .B2(n15916), .ZN(
        n13075) );
  AOI21_X1 U14810 ( .B1(n15042), .B2(n14885), .A(n14872), .ZN(n15043) );
  NOR2_X1 U14811 ( .A1(n14383), .A2(n15933), .ZN(n13079) );
  OAI22_X1 U14812 ( .A1(n15942), .A2(n13077), .B1(n14536), .B2(n15931), .ZN(
        n13078) );
  AOI211_X1 U14813 ( .C1(n15043), .C2(n14958), .A(n13079), .B(n13078), .ZN(
        n13081) );
  NAND2_X1 U14814 ( .A1(n15041), .A2(n15941), .ZN(n13080) );
  OAI211_X1 U14815 ( .C1(n15045), .C2(n14997), .A(n13081), .B(n13080), .ZN(
        P1_U3266) );
  XNOR2_X1 U14816 ( .A(n13807), .B(n13119), .ZN(n13088) );
  INV_X1 U14817 ( .A(n13084), .ZN(n13085) );
  NAND2_X1 U14818 ( .A1(n13085), .A2(n13573), .ZN(n13086) );
  NAND2_X1 U14819 ( .A1(n13087), .A2(n13086), .ZN(n13512) );
  XNOR2_X1 U14820 ( .A(n13088), .B(n13734), .ZN(n13513) );
  XNOR2_X1 U14821 ( .A(n13544), .B(n13119), .ZN(n13089) );
  XNOR2_X1 U14822 ( .A(n13089), .B(n13745), .ZN(n13545) );
  INV_X1 U14823 ( .A(n13089), .ZN(n13090) );
  XNOR2_X1 U14824 ( .A(n13860), .B(n13119), .ZN(n13091) );
  XNOR2_X1 U14825 ( .A(n13091), .B(n13735), .ZN(n13483) );
  NAND2_X1 U14826 ( .A1(n13484), .A2(n13483), .ZN(n13093) );
  NAND2_X1 U14827 ( .A1(n13091), .A2(n13707), .ZN(n13092) );
  XNOR2_X1 U14828 ( .A(n13532), .B(n13119), .ZN(n13094) );
  NAND2_X1 U14829 ( .A1(n13094), .A2(n13721), .ZN(n13095) );
  OAI21_X1 U14830 ( .B1(n13094), .B2(n13721), .A(n13095), .ZN(n13529) );
  INV_X1 U14831 ( .A(n13096), .ZN(n13098) );
  MUX2_X1 U14832 ( .A(n13098), .B(n13097), .S(n13119), .Z(n13492) );
  INV_X1 U14833 ( .A(n13099), .ZN(n13100) );
  MUX2_X1 U14834 ( .A(n7208), .B(n13100), .S(n11350), .Z(n13491) );
  XNOR2_X1 U14835 ( .A(n13539), .B(n13119), .ZN(n13101) );
  INV_X1 U14836 ( .A(n13101), .ZN(n13102) );
  NOR2_X1 U14837 ( .A1(n13103), .A2(n13102), .ZN(n13104) );
  XNOR2_X1 U14838 ( .A(n13474), .B(n13119), .ZN(n13105) );
  XNOR2_X1 U14839 ( .A(n13107), .B(n13105), .ZN(n13475) );
  NAND2_X1 U14840 ( .A1(n13475), .A2(n13676), .ZN(n13109) );
  INV_X1 U14841 ( .A(n13105), .ZN(n13106) );
  OR2_X1 U14842 ( .A1(n13107), .A2(n13106), .ZN(n13108) );
  NAND2_X1 U14843 ( .A1(n13109), .A2(n13108), .ZN(n13519) );
  XNOR2_X1 U14844 ( .A(n13522), .B(n13119), .ZN(n13110) );
  XNOR2_X1 U14845 ( .A(n13110), .B(n13665), .ZN(n13520) );
  NAND2_X1 U14846 ( .A1(n13519), .A2(n13520), .ZN(n13112) );
  NAND2_X1 U14847 ( .A1(n13110), .A2(n13504), .ZN(n13111) );
  NAND2_X1 U14848 ( .A1(n13112), .A2(n13111), .ZN(n13501) );
  XNOR2_X1 U14849 ( .A(n13505), .B(n13119), .ZN(n13113) );
  XNOR2_X1 U14850 ( .A(n13113), .B(n13569), .ZN(n13502) );
  NAND2_X1 U14851 ( .A1(n13113), .A2(n13656), .ZN(n13114) );
  XNOR2_X1 U14852 ( .A(n13560), .B(n13119), .ZN(n13116) );
  XNOR2_X1 U14853 ( .A(n13116), .B(n13637), .ZN(n13556) );
  XNOR2_X1 U14854 ( .A(n13117), .B(n13119), .ZN(n13118) );
  XNOR2_X1 U14855 ( .A(n13118), .B(n13568), .ZN(n13466) );
  AOI22_X1 U14856 ( .A1(n13467), .A2(n13466), .B1(n13627), .B2(n13118), .ZN(
        n13121) );
  XNOR2_X1 U14857 ( .A(n13608), .B(n13119), .ZN(n13120) );
  XNOR2_X1 U14858 ( .A(n13121), .B(n13120), .ZN(n13127) );
  AOI22_X1 U14859 ( .A1(n13568), .A2(n13549), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13122) );
  OAI21_X1 U14860 ( .B1(n13610), .B2(n13551), .A(n13122), .ZN(n13125) );
  NOR2_X1 U14861 ( .A1(n13828), .A2(n13561), .ZN(n13124) );
  AOI211_X1 U14862 ( .C1(n13613), .C2(n13564), .A(n13125), .B(n13124), .ZN(
        n13126) );
  OAI21_X1 U14863 ( .B1(n13127), .B2(n13566), .A(n13126), .ZN(P3_U3160) );
  INV_X1 U14864 ( .A(n13351), .ZN(n13465) );
  OAI222_X1 U14865 ( .A1(P1_U3086), .A2(n8517), .B1(n15160), .B2(n13465), .C1(
        n13128), .C2(n15157), .ZN(P1_U3325) );
  INV_X1 U14866 ( .A(n13129), .ZN(n13130) );
  OAI222_X1 U14867 ( .A1(n13132), .A2(P3_U3151), .B1(n13131), .B2(n13130), 
        .C1(n15283), .C2(n13880), .ZN(P3_U3268) );
  INV_X1 U14868 ( .A(n13138), .ZN(n13133) );
  NAND2_X1 U14869 ( .A1(n13133), .A2(n13365), .ZN(n13142) );
  NAND2_X1 U14870 ( .A1(n13135), .A2(n13393), .ZN(n13134) );
  NAND2_X1 U14871 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  NAND3_X1 U14872 ( .A1(n13142), .A2(n13141), .A3(n13140), .ZN(n13153) );
  NAND2_X1 U14873 ( .A1(n13144), .A2(n13393), .ZN(n13145) );
  NAND2_X1 U14874 ( .A1(n13146), .A2(n13145), .ZN(n13154) );
  NAND2_X1 U14875 ( .A1(n13153), .A2(n13154), .ZN(n13150) );
  NAND2_X1 U14876 ( .A1(n13144), .A2(n13365), .ZN(n13148) );
  NAND2_X1 U14877 ( .A1(n13143), .A2(n13393), .ZN(n13147) );
  NAND2_X1 U14878 ( .A1(n13148), .A2(n13147), .ZN(n13149) );
  NAND2_X1 U14879 ( .A1(n13150), .A2(n13149), .ZN(n13159) );
  NAND2_X1 U14880 ( .A1(n14248), .A2(n13393), .ZN(n13151) );
  NAND2_X1 U14881 ( .A1(n13152), .A2(n13151), .ZN(n13160) );
  NAND2_X1 U14882 ( .A1(n13160), .A2(n13161), .ZN(n13158) );
  INV_X1 U14883 ( .A(n13153), .ZN(n13156) );
  NAND2_X1 U14884 ( .A1(n13156), .A2(n13155), .ZN(n13157) );
  NAND3_X1 U14885 ( .A1(n13159), .A2(n13158), .A3(n13157), .ZN(n13165) );
  INV_X1 U14886 ( .A(n13160), .ZN(n13163) );
  INV_X1 U14887 ( .A(n13161), .ZN(n13162) );
  NAND2_X1 U14888 ( .A1(n13163), .A2(n13162), .ZN(n13164) );
  NAND2_X1 U14889 ( .A1(n13165), .A2(n13164), .ZN(n13171) );
  NAND2_X1 U14890 ( .A1(n14026), .A2(n13393), .ZN(n13167) );
  NAND2_X1 U14891 ( .A1(n13168), .A2(n13365), .ZN(n13166) );
  NAND2_X1 U14892 ( .A1(n13167), .A2(n13166), .ZN(n13172) );
  AOI22_X1 U14893 ( .A1(n13365), .A2(n14026), .B1(n13168), .B2(n13393), .ZN(
        n13169) );
  INV_X1 U14894 ( .A(n13169), .ZN(n13170) );
  INV_X1 U14895 ( .A(n13172), .ZN(n13173) );
  NAND2_X1 U14896 ( .A1(n13176), .A2(n13393), .ZN(n13175) );
  NAND2_X1 U14897 ( .A1(n14025), .A2(n13365), .ZN(n13174) );
  NAND2_X1 U14898 ( .A1(n13176), .A2(n13365), .ZN(n13177) );
  OAI21_X1 U14899 ( .B1(n13178), .B2(n13365), .A(n13177), .ZN(n13179) );
  NAND2_X1 U14900 ( .A1(n13182), .A2(n13365), .ZN(n13181) );
  NAND2_X1 U14901 ( .A1(n14024), .A2(n13340), .ZN(n13180) );
  NAND2_X1 U14902 ( .A1(n13181), .A2(n13180), .ZN(n13185) );
  AOI22_X1 U14903 ( .A1(n13182), .A2(n13340), .B1(n13365), .B2(n14024), .ZN(
        n13183) );
  AOI21_X1 U14904 ( .B1(n13186), .B2(n13185), .A(n13183), .ZN(n13184) );
  INV_X1 U14905 ( .A(n13184), .ZN(n13187) );
  NAND2_X1 U14906 ( .A1(n16043), .A2(n13340), .ZN(n13189) );
  NAND2_X1 U14907 ( .A1(n14023), .A2(n13365), .ZN(n13188) );
  NAND2_X1 U14908 ( .A1(n13189), .A2(n13188), .ZN(n13191) );
  AOI22_X1 U14909 ( .A1(n16043), .A2(n13365), .B1(n14023), .B2(n13340), .ZN(
        n13190) );
  NAND2_X1 U14910 ( .A1(n13195), .A2(n13365), .ZN(n13194) );
  NAND2_X1 U14911 ( .A1(n14022), .A2(n13340), .ZN(n13193) );
  NAND2_X1 U14912 ( .A1(n13195), .A2(n13340), .ZN(n13196) );
  OAI21_X1 U14913 ( .B1(n13197), .B2(n13393), .A(n13196), .ZN(n13198) );
  NAND2_X1 U14914 ( .A1(n13202), .A2(n13340), .ZN(n13201) );
  NAND2_X1 U14915 ( .A1(n14021), .A2(n13365), .ZN(n13200) );
  AOI22_X1 U14916 ( .A1(n13202), .A2(n13365), .B1(n14021), .B2(n13340), .ZN(
        n13203) );
  INV_X1 U14917 ( .A(n13203), .ZN(n13204) );
  NAND2_X1 U14918 ( .A1(n13205), .A2(n13204), .ZN(n13207) );
  NAND2_X1 U14919 ( .A1(n7268), .A2(n7204), .ZN(n13206) );
  NAND2_X1 U14920 ( .A1(n13210), .A2(n13365), .ZN(n13209) );
  NAND2_X1 U14921 ( .A1(n14020), .A2(n13340), .ZN(n13208) );
  NAND2_X1 U14922 ( .A1(n13210), .A2(n13340), .ZN(n13211) );
  OAI21_X1 U14923 ( .B1(n13212), .B2(n13393), .A(n13211), .ZN(n13213) );
  NAND2_X1 U14924 ( .A1(n13216), .A2(n13340), .ZN(n13215) );
  NAND2_X1 U14925 ( .A1(n14019), .A2(n13365), .ZN(n13214) );
  NAND2_X1 U14926 ( .A1(n13215), .A2(n13214), .ZN(n13220) );
  AOI22_X1 U14927 ( .A1(n13216), .A2(n13365), .B1(n14019), .B2(n13340), .ZN(
        n13217) );
  INV_X1 U14928 ( .A(n13217), .ZN(n13218) );
  NAND2_X1 U14929 ( .A1(n13219), .A2(n13218), .ZN(n13221) );
  NAND2_X1 U14930 ( .A1(n13224), .A2(n13365), .ZN(n13223) );
  NAND2_X1 U14931 ( .A1(n14018), .A2(n13340), .ZN(n13222) );
  NAND2_X1 U14932 ( .A1(n13223), .A2(n13222), .ZN(n13230) );
  NAND2_X1 U14933 ( .A1(n13224), .A2(n13340), .ZN(n13225) );
  NAND2_X1 U14934 ( .A1(n13228), .A2(n13227), .ZN(n13234) );
  INV_X1 U14935 ( .A(n13229), .ZN(n13232) );
  INV_X1 U14936 ( .A(n13230), .ZN(n13231) );
  NAND2_X1 U14937 ( .A1(n13232), .A2(n13231), .ZN(n13233) );
  NAND2_X1 U14938 ( .A1(n13237), .A2(n13340), .ZN(n13236) );
  NAND2_X1 U14939 ( .A1(n14017), .A2(n13365), .ZN(n13235) );
  NAND2_X1 U14940 ( .A1(n13236), .A2(n13235), .ZN(n13240) );
  AOI22_X1 U14941 ( .A1(n13237), .A2(n13365), .B1(n14017), .B2(n13340), .ZN(
        n13238) );
  INV_X1 U14942 ( .A(n13238), .ZN(n13239) );
  INV_X1 U14943 ( .A(n13240), .ZN(n13241) );
  NAND2_X1 U14944 ( .A1(n16148), .A2(n13365), .ZN(n13243) );
  NAND2_X1 U14945 ( .A1(n13244), .A2(n13340), .ZN(n13242) );
  NAND2_X1 U14946 ( .A1(n13243), .A2(n13242), .ZN(n13246) );
  AOI22_X1 U14947 ( .A1(n16148), .A2(n13340), .B1(n13365), .B2(n13244), .ZN(
        n13245) );
  NAND2_X1 U14948 ( .A1(n13249), .A2(n13340), .ZN(n13248) );
  NAND2_X1 U14949 ( .A1(n14016), .A2(n13365), .ZN(n13247) );
  NAND2_X1 U14950 ( .A1(n13248), .A2(n13247), .ZN(n13253) );
  NAND2_X1 U14951 ( .A1(n13249), .A2(n13365), .ZN(n13250) );
  OAI21_X1 U14952 ( .B1(n13251), .B2(n13365), .A(n13250), .ZN(n13252) );
  NAND2_X1 U14953 ( .A1(n14342), .A2(n13365), .ZN(n13256) );
  NAND2_X1 U14954 ( .A1(n14015), .A2(n13340), .ZN(n13255) );
  NAND2_X1 U14955 ( .A1(n13256), .A2(n13255), .ZN(n13258) );
  AOI22_X1 U14956 ( .A1(n14342), .A2(n13340), .B1(n13365), .B2(n14015), .ZN(
        n13257) );
  NAND2_X1 U14957 ( .A1(n14337), .A2(n13340), .ZN(n13261) );
  NAND2_X1 U14958 ( .A1(n14014), .A2(n13365), .ZN(n13260) );
  NAND2_X1 U14959 ( .A1(n14337), .A2(n13365), .ZN(n13263) );
  NAND2_X1 U14960 ( .A1(n14014), .A2(n13340), .ZN(n13262) );
  NAND2_X1 U14961 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  NAND2_X1 U14962 ( .A1(n14332), .A2(n13365), .ZN(n13266) );
  NAND2_X1 U14963 ( .A1(n14013), .A2(n13340), .ZN(n13265) );
  NAND2_X1 U14964 ( .A1(n13266), .A2(n13265), .ZN(n13270) );
  NAND2_X1 U14965 ( .A1(n13271), .A2(n13270), .ZN(n13269) );
  AOI22_X1 U14966 ( .A1(n14332), .A2(n13340), .B1(n13365), .B2(n14013), .ZN(
        n13267) );
  NAND2_X1 U14967 ( .A1(n14327), .A2(n13340), .ZN(n13274) );
  NAND2_X1 U14968 ( .A1(n14012), .A2(n13365), .ZN(n13273) );
  NAND2_X1 U14969 ( .A1(n13274), .A2(n13273), .ZN(n13277) );
  NAND2_X1 U14970 ( .A1(n14327), .A2(n13365), .ZN(n13275) );
  OAI21_X1 U14971 ( .B1(n14190), .B2(n13365), .A(n13275), .ZN(n13276) );
  NAND2_X1 U14972 ( .A1(n14317), .A2(n13365), .ZN(n13280) );
  NAND2_X1 U14973 ( .A1(n14011), .A2(n13340), .ZN(n13279) );
  NAND2_X1 U14974 ( .A1(n13280), .A2(n13279), .ZN(n13284) );
  AOI22_X1 U14975 ( .A1(n14317), .A2(n13340), .B1(n13365), .B2(n14011), .ZN(
        n13281) );
  NAND2_X1 U14976 ( .A1(n13283), .A2(n13282), .ZN(n13286) );
  NAND2_X1 U14977 ( .A1(n14314), .A2(n13340), .ZN(n13288) );
  NAND2_X1 U14978 ( .A1(n14010), .A2(n13365), .ZN(n13287) );
  NAND2_X1 U14979 ( .A1(n14314), .A2(n13365), .ZN(n13289) );
  OAI21_X1 U14980 ( .B1(n14192), .B2(n13365), .A(n13289), .ZN(n13290) );
  NAND2_X1 U14981 ( .A1(n14309), .A2(n13365), .ZN(n13292) );
  NAND2_X1 U14982 ( .A1(n14009), .A2(n13340), .ZN(n13291) );
  NAND2_X1 U14983 ( .A1(n13292), .A2(n13291), .ZN(n13294) );
  AOI22_X1 U14984 ( .A1(n14309), .A2(n13340), .B1(n13365), .B2(n14009), .ZN(
        n13293) );
  AOI21_X1 U14985 ( .B1(n13295), .B2(n13294), .A(n13293), .ZN(n13296) );
  NAND2_X1 U14986 ( .A1(n14301), .A2(n13340), .ZN(n13298) );
  NAND2_X1 U14987 ( .A1(n14008), .A2(n13365), .ZN(n13297) );
  NAND2_X1 U14988 ( .A1(n13298), .A2(n13297), .ZN(n13301) );
  AOI22_X1 U14989 ( .A1(n14301), .A2(n13365), .B1(n14008), .B2(n13340), .ZN(
        n13299) );
  INV_X1 U14990 ( .A(n13299), .ZN(n13300) );
  INV_X1 U14991 ( .A(n13301), .ZN(n13302) );
  AND2_X1 U14992 ( .A1(n14007), .A2(n13340), .ZN(n13303) );
  AOI21_X1 U14993 ( .B1(n14295), .B2(n13365), .A(n13303), .ZN(n13309) );
  INV_X1 U14994 ( .A(n13309), .ZN(n13304) );
  NAND2_X1 U14995 ( .A1(n13308), .A2(n13304), .ZN(n13307) );
  NAND2_X1 U14996 ( .A1(n14295), .A2(n13340), .ZN(n13305) );
  OAI21_X1 U14997 ( .B1(n14145), .B2(n13393), .A(n13305), .ZN(n13306) );
  NAND2_X1 U14998 ( .A1(n13307), .A2(n13306), .ZN(n13312) );
  INV_X1 U14999 ( .A(n13308), .ZN(n13310) );
  NAND2_X1 U15000 ( .A1(n13310), .A2(n13309), .ZN(n13311) );
  NAND2_X1 U15001 ( .A1(n14290), .A2(n13340), .ZN(n13314) );
  NAND2_X1 U15002 ( .A1(n14006), .A2(n13365), .ZN(n13313) );
  AOI22_X1 U15003 ( .A1(n14290), .A2(n13365), .B1(n14006), .B2(n13340), .ZN(
        n13315) );
  INV_X1 U15004 ( .A(n13315), .ZN(n13316) );
  NAND2_X1 U15005 ( .A1(n14364), .A2(n13350), .ZN(n13318) );
  NAND2_X1 U15006 ( .A1(n10741), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13317) );
  INV_X1 U15007 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U15008 ( .A1(n10552), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U15009 ( .A1(n13357), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n13319) );
  OAI211_X1 U15010 ( .C1(n10553), .C2(n13321), .A(n13320), .B(n13319), .ZN(
        n14003) );
  XNOR2_X1 U15011 ( .A(n14032), .B(n14003), .ZN(n13436) );
  NAND2_X1 U15012 ( .A1(n14369), .A2(n13350), .ZN(n13323) );
  NAND2_X1 U15013 ( .A1(n10535), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13322) );
  AND2_X1 U15014 ( .A1(n14004), .A2(n13340), .ZN(n13324) );
  AOI21_X1 U15015 ( .B1(n14260), .B2(n13365), .A(n13324), .ZN(n13369) );
  NAND2_X1 U15016 ( .A1(n14260), .A2(n13340), .ZN(n13326) );
  NAND2_X1 U15017 ( .A1(n14004), .A2(n13365), .ZN(n13325) );
  NAND2_X1 U15018 ( .A1(n13326), .A2(n13325), .ZN(n13368) );
  NAND2_X1 U15019 ( .A1(n13369), .A2(n13368), .ZN(n13375) );
  AND2_X1 U15020 ( .A1(n14054), .A2(n13340), .ZN(n13327) );
  AOI21_X1 U15021 ( .B1(n14267), .B2(n13365), .A(n13327), .ZN(n13374) );
  NAND2_X1 U15022 ( .A1(n14267), .A2(n13340), .ZN(n13329) );
  NAND2_X1 U15023 ( .A1(n14054), .A2(n13365), .ZN(n13328) );
  NAND2_X1 U15024 ( .A1(n13329), .A2(n13328), .ZN(n13373) );
  NAND2_X1 U15025 ( .A1(n13374), .A2(n13373), .ZN(n13330) );
  AND2_X1 U15026 ( .A1(n13375), .A2(n13330), .ZN(n13331) );
  AND2_X1 U15027 ( .A1(n13436), .A2(n13331), .ZN(n13345) );
  AND2_X1 U15028 ( .A1(n14092), .A2(n13340), .ZN(n13332) );
  AOI21_X1 U15029 ( .B1(n14271), .B2(n13365), .A(n13332), .ZN(n13347) );
  NAND2_X1 U15030 ( .A1(n14271), .A2(n13340), .ZN(n13334) );
  NAND2_X1 U15031 ( .A1(n14092), .A2(n13365), .ZN(n13333) );
  NAND2_X1 U15032 ( .A1(n13334), .A2(n13333), .ZN(n13346) );
  NAND2_X1 U15033 ( .A1(n13347), .A2(n13346), .ZN(n13335) );
  AND2_X1 U15034 ( .A1(n13345), .A2(n13335), .ZN(n13342) );
  AND2_X1 U15035 ( .A1(n14005), .A2(n13340), .ZN(n13336) );
  AOI21_X1 U15036 ( .B1(n14278), .B2(n13365), .A(n13336), .ZN(n13344) );
  NAND2_X1 U15037 ( .A1(n14278), .A2(n13340), .ZN(n13338) );
  NAND2_X1 U15038 ( .A1(n14005), .A2(n13365), .ZN(n13337) );
  NAND2_X1 U15039 ( .A1(n13338), .A2(n13337), .ZN(n13343) );
  NAND2_X1 U15040 ( .A1(n13344), .A2(n13343), .ZN(n13339) );
  AOI22_X1 U15041 ( .A1(n14285), .A2(n13365), .B1(n14090), .B2(n13340), .ZN(
        n13384) );
  OAI22_X1 U15042 ( .A1(n14108), .A2(n13365), .B1(n14118), .B2(n13393), .ZN(
        n13383) );
  AND2_X1 U15043 ( .A1(n13384), .A2(n13383), .ZN(n13341) );
  INV_X1 U15044 ( .A(n13345), .ZN(n13381) );
  INV_X1 U15045 ( .A(n13346), .ZN(n13349) );
  INV_X1 U15046 ( .A(n13347), .ZN(n13348) );
  NAND2_X1 U15047 ( .A1(n13349), .A2(n13348), .ZN(n13380) );
  NAND2_X1 U15048 ( .A1(n13351), .A2(n13350), .ZN(n13353) );
  NAND2_X1 U15049 ( .A1(n10741), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13352) );
  INV_X1 U15050 ( .A(n13354), .ZN(n13355) );
  MUX2_X1 U15051 ( .A(n14003), .B(n13355), .S(n13399), .Z(n13362) );
  NAND2_X1 U15052 ( .A1(n13356), .A2(n13445), .ZN(n13361) );
  INV_X1 U15053 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13360) );
  NAND2_X1 U15054 ( .A1(n10552), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n13359) );
  NAND2_X1 U15055 ( .A1(n13357), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n13358) );
  OAI211_X1 U15056 ( .C1(n10553), .C2(n13360), .A(n13359), .B(n13358), .ZN(
        n14048) );
  OAI21_X1 U15057 ( .B1(n13362), .B2(n13361), .A(n14048), .ZN(n13363) );
  INV_X1 U15058 ( .A(n13363), .ZN(n13364) );
  AOI21_X1 U15059 ( .B1(n14035), .B2(n13365), .A(n13364), .ZN(n13390) );
  NAND2_X1 U15060 ( .A1(n14035), .A2(n13340), .ZN(n13367) );
  NAND2_X1 U15061 ( .A1(n14048), .A2(n13365), .ZN(n13366) );
  NAND2_X1 U15062 ( .A1(n13367), .A2(n13366), .ZN(n13389) );
  OAI22_X1 U15063 ( .A1(n13390), .A2(n13389), .B1(n13369), .B2(n13368), .ZN(
        n13372) );
  NAND2_X1 U15064 ( .A1(n14032), .A2(n13340), .ZN(n13370) );
  NAND2_X1 U15065 ( .A1(n14003), .A2(n13365), .ZN(n13395) );
  OAI211_X1 U15066 ( .C1(n14032), .C2(n14003), .A(n13370), .B(n13395), .ZN(
        n13371) );
  NAND2_X1 U15067 ( .A1(n13372), .A2(n13371), .ZN(n13379) );
  INV_X1 U15068 ( .A(n13373), .ZN(n13377) );
  INV_X1 U15069 ( .A(n13374), .ZN(n13376) );
  NAND4_X1 U15070 ( .A1(n13436), .A2(n13377), .A3(n13376), .A4(n13375), .ZN(
        n13378) );
  OAI211_X1 U15071 ( .C1(n13381), .C2(n13380), .A(n13379), .B(n13378), .ZN(
        n13382) );
  AOI21_X1 U15072 ( .B1(n13388), .B2(n13387), .A(n13386), .ZN(n13398) );
  INV_X1 U15073 ( .A(n13389), .ZN(n13392) );
  INV_X1 U15074 ( .A(n13390), .ZN(n13391) );
  NOR2_X1 U15075 ( .A1(n13392), .A2(n13391), .ZN(n13397) );
  INV_X1 U15076 ( .A(n14003), .ZN(n14031) );
  NAND2_X1 U15077 ( .A1(n14031), .A2(n13393), .ZN(n13394) );
  MUX2_X1 U15078 ( .A(n13395), .B(n13394), .S(n14032), .Z(n13396) );
  INV_X1 U15079 ( .A(n13447), .ZN(n13400) );
  NAND2_X1 U15080 ( .A1(n13402), .A2(n13401), .ZN(n14099) );
  NAND4_X1 U15081 ( .A1(n13404), .A2(n15898), .A3(n13403), .A4(n13442), .ZN(
        n13406) );
  NOR2_X1 U15082 ( .A1(n13406), .A2(n13405), .ZN(n13409) );
  NAND4_X1 U15083 ( .A1(n13410), .A2(n13409), .A3(n13408), .A4(n13407), .ZN(
        n13411) );
  NOR3_X1 U15084 ( .A1(n13413), .A2(n13412), .A3(n13411), .ZN(n13416) );
  NAND4_X1 U15085 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13418) );
  NOR2_X1 U15086 ( .A1(n13419), .A2(n13418), .ZN(n13422) );
  NAND4_X1 U15087 ( .A1(n13423), .A2(n13422), .A3(n13421), .A4(n13420), .ZN(
        n13424) );
  NOR2_X1 U15088 ( .A1(n13425), .A2(n13424), .ZN(n13426) );
  AND4_X1 U15089 ( .A1(n14194), .A2(n13426), .A3(n14211), .A4(n14238), .ZN(
        n13427) );
  XNOR2_X1 U15090 ( .A(n14314), .B(n14010), .ZN(n14177) );
  XNOR2_X1 U15091 ( .A(n14309), .B(n14009), .ZN(n14163) );
  AND4_X1 U15092 ( .A1(n13428), .A2(n13427), .A3(n14177), .A4(n14163), .ZN(
        n13429) );
  AND2_X1 U15093 ( .A1(n14099), .A2(n13429), .ZN(n13431) );
  NAND4_X1 U15094 ( .A1(n14087), .A2(n13431), .A3(n13430), .A4(n14149), .ZN(
        n13432) );
  NOR3_X1 U15095 ( .A1(n14072), .A2(n13433), .A3(n13432), .ZN(n13435) );
  XNOR2_X1 U15096 ( .A(n14035), .B(n14048), .ZN(n13434) );
  XNOR2_X1 U15097 ( .A(n14260), .B(n14004), .ZN(n14056) );
  OAI21_X1 U15098 ( .B1(n10435), .B2(n13442), .A(n10458), .ZN(n13444) );
  NAND2_X1 U15099 ( .A1(n13444), .A2(n13443), .ZN(n13449) );
  INV_X1 U15100 ( .A(n13444), .ZN(n13446) );
  NAND2_X1 U15101 ( .A1(n13446), .A2(n13445), .ZN(n13448) );
  MUX2_X1 U15102 ( .A(n13449), .B(n13448), .S(n13447), .Z(n13450) );
  INV_X1 U15103 ( .A(n13450), .ZN(n13451) );
  AOI21_X1 U15104 ( .B1(n13453), .B2(n13452), .A(n13451), .ZN(n13459) );
  NOR4_X1 U15105 ( .A1(n15406), .A2(n10950), .A3(n13455), .A4(n13454), .ZN(
        n13457) );
  OAI21_X1 U15106 ( .B1(n13458), .B2(n10435), .A(P2_B_REG_SCAN_IN), .ZN(n13456) );
  OAI22_X1 U15107 ( .A1(n13459), .A2(n13458), .B1(n13457), .B2(n13456), .ZN(
        P2_U3328) );
  INV_X1 U15108 ( .A(n13460), .ZN(n13461) );
  OAI222_X1 U15109 ( .A1(P3_U3151), .A2(n9078), .B1(n13880), .B2(n15281), .C1(
        n13131), .C2(n13461), .ZN(P3_U3265) );
  INV_X1 U15110 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13463) );
  OAI222_X1 U15111 ( .A1(n14378), .A2(n13465), .B1(P2_U3088), .B2(n13464), 
        .C1(n13463), .C2(n14370), .ZN(P2_U3297) );
  XNOR2_X1 U15112 ( .A(n13467), .B(n13466), .ZN(n13468) );
  NAND2_X1 U15113 ( .A1(n13468), .A2(n13476), .ZN(n13473) );
  AOI22_X1 U15114 ( .A1(n13637), .A2(n13549), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13469) );
  OAI21_X1 U15115 ( .B1(n13470), .B2(n13551), .A(n13469), .ZN(n13471) );
  AOI21_X1 U15116 ( .B1(n13619), .B2(n13564), .A(n13471), .ZN(n13472) );
  OAI211_X1 U15117 ( .C1(n13768), .C2(n13561), .A(n13473), .B(n13472), .ZN(
        P3_U3154) );
  XNOR2_X1 U15118 ( .A(n13475), .B(n13676), .ZN(n13477) );
  NAND2_X1 U15119 ( .A1(n13477), .A2(n13476), .ZN(n13482) );
  OAI22_X1 U15120 ( .A1(n13504), .A2(n13551), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13478), .ZN(n13480) );
  NOR2_X1 U15121 ( .A1(n13496), .A2(n13559), .ZN(n13479) );
  AOI211_X1 U15122 ( .C1(n13668), .C2(n13564), .A(n13480), .B(n13479), .ZN(
        n13481) );
  OAI211_X1 U15123 ( .C1(n13844), .C2(n13561), .A(n13482), .B(n13481), .ZN(
        P3_U3156) );
  XNOR2_X1 U15124 ( .A(n13484), .B(n13483), .ZN(n13490) );
  NAND2_X1 U15125 ( .A1(n13687), .A2(n13557), .ZN(n13486) );
  OAI211_X1 U15126 ( .C1(n13745), .C2(n13559), .A(n13486), .B(n13485), .ZN(
        n13488) );
  NOR2_X1 U15127 ( .A1(n13860), .A2(n13561), .ZN(n13487) );
  AOI211_X1 U15128 ( .C1(n13724), .C2(n13564), .A(n13488), .B(n13487), .ZN(
        n13489) );
  OAI21_X1 U15129 ( .B1(n13490), .B2(n13566), .A(n13489), .ZN(P3_U3159) );
  NAND2_X1 U15130 ( .A1(n8307), .A2(n13492), .ZN(n13493) );
  XNOR2_X1 U15131 ( .A(n13494), .B(n13493), .ZN(n13500) );
  AOI22_X1 U15132 ( .A1(n13687), .A2(n13549), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13495) );
  OAI21_X1 U15133 ( .B1(n13496), .B2(n13551), .A(n13495), .ZN(n13498) );
  INV_X1 U15134 ( .A(n13697), .ZN(n13852) );
  NOR2_X1 U15135 ( .A1(n13852), .A2(n13561), .ZN(n13497) );
  AOI211_X1 U15136 ( .C1(n13695), .C2(n13564), .A(n13498), .B(n13497), .ZN(
        n13499) );
  OAI21_X1 U15137 ( .B1(n13500), .B2(n13566), .A(n13499), .ZN(P3_U3163) );
  XOR2_X1 U15138 ( .A(n13502), .B(n13501), .Z(n13509) );
  AOI22_X1 U15139 ( .A1(n13557), .A2(n13637), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13503) );
  OAI21_X1 U15140 ( .B1(n13504), .B2(n13559), .A(n13503), .ZN(n13507) );
  NOR2_X1 U15141 ( .A1(n13836), .A2(n13561), .ZN(n13506) );
  AOI211_X1 U15142 ( .C1(n13644), .C2(n13564), .A(n13507), .B(n13506), .ZN(
        n13508) );
  OAI21_X1 U15143 ( .B1(n13509), .B2(n13566), .A(n13508), .ZN(P3_U3165) );
  INV_X1 U15144 ( .A(n13510), .ZN(n13511) );
  AOI21_X1 U15145 ( .B1(n13513), .B2(n13512), .A(n13511), .ZN(n13518) );
  NOR2_X1 U15146 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9392), .ZN(n15819) );
  AOI21_X1 U15147 ( .B1(n13571), .B2(n13557), .A(n15819), .ZN(n13514) );
  OAI21_X1 U15148 ( .B1(n13746), .B2(n13559), .A(n13514), .ZN(n13516) );
  INV_X1 U15149 ( .A(n13807), .ZN(n13755) );
  NOR2_X1 U15150 ( .A1(n13755), .A2(n13561), .ZN(n13515) );
  AOI211_X1 U15151 ( .C1(n13752), .C2(n13564), .A(n13516), .B(n13515), .ZN(
        n13517) );
  OAI21_X1 U15152 ( .B1(n13518), .B2(n13566), .A(n13517), .ZN(P3_U3168) );
  XOR2_X1 U15153 ( .A(n13520), .B(n13519), .Z(n13526) );
  AOI22_X1 U15154 ( .A1(n13569), .A2(n13557), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13521) );
  OAI21_X1 U15155 ( .B1(n13676), .B2(n13559), .A(n13521), .ZN(n13524) );
  NOR2_X1 U15156 ( .A1(n13840), .A2(n13561), .ZN(n13523) );
  AOI211_X1 U15157 ( .C1(n13657), .C2(n13564), .A(n13524), .B(n13523), .ZN(
        n13525) );
  OAI21_X1 U15158 ( .B1(n13526), .B2(n13566), .A(n13525), .ZN(P3_U3169) );
  INV_X1 U15159 ( .A(n13527), .ZN(n13528) );
  AOI21_X1 U15160 ( .B1(n13530), .B2(n13529), .A(n13528), .ZN(n13536) );
  AOI22_X1 U15161 ( .A1(n13707), .A2(n13549), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13531) );
  OAI21_X1 U15162 ( .B1(n13675), .B2(n13551), .A(n13531), .ZN(n13534) );
  NOR2_X1 U15163 ( .A1(n13856), .A2(n13561), .ZN(n13533) );
  AOI211_X1 U15164 ( .C1(n13712), .C2(n13564), .A(n13534), .B(n13533), .ZN(
        n13535) );
  OAI21_X1 U15165 ( .B1(n13536), .B2(n13566), .A(n13535), .ZN(P3_U3173) );
  XNOR2_X1 U15166 ( .A(n13537), .B(n13688), .ZN(n13543) );
  AOI22_X1 U15167 ( .A1(n13709), .A2(n13549), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13538) );
  OAI21_X1 U15168 ( .B1(n13676), .B2(n13551), .A(n13538), .ZN(n13541) );
  NOR2_X1 U15169 ( .A1(n13848), .A2(n13561), .ZN(n13540) );
  AOI211_X1 U15170 ( .C1(n13679), .C2(n13564), .A(n13541), .B(n13540), .ZN(
        n13542) );
  OAI21_X1 U15171 ( .B1(n13543), .B2(n13566), .A(n13542), .ZN(P3_U3175) );
  INV_X1 U15172 ( .A(n13544), .ZN(n13865) );
  AOI21_X1 U15173 ( .B1(n13546), .B2(n13545), .A(n13566), .ZN(n13548) );
  NAND2_X1 U15174 ( .A1(n13548), .A2(n13547), .ZN(n13554) );
  NAND2_X1 U15175 ( .A1(n13572), .A2(n13549), .ZN(n13550) );
  NAND2_X1 U15176 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n15849)
         );
  OAI211_X1 U15177 ( .C1(n13735), .C2(n13551), .A(n13550), .B(n15849), .ZN(
        n13552) );
  AOI21_X1 U15178 ( .B1(n13739), .B2(n13564), .A(n13552), .ZN(n13553) );
  OAI211_X1 U15179 ( .C1(n13865), .C2(n13561), .A(n13554), .B(n13553), .ZN(
        P3_U3178) );
  XOR2_X1 U15180 ( .A(n13556), .B(n13555), .Z(n13567) );
  AOI22_X1 U15181 ( .A1(n13568), .A2(n13557), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13558) );
  OAI21_X1 U15182 ( .B1(n13656), .B2(n13559), .A(n13558), .ZN(n13563) );
  NOR2_X1 U15183 ( .A1(n13832), .A2(n13561), .ZN(n13562) );
  AOI211_X1 U15184 ( .C1(n13630), .C2(n13564), .A(n13563), .B(n13562), .ZN(
        n13565) );
  OAI21_X1 U15185 ( .B1(n13567), .B2(n13566), .A(n13565), .ZN(P3_U3180) );
  MUX2_X1 U15186 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n9881), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15187 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13568), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15188 ( .A(n13637), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13589), .Z(
        P3_U3517) );
  MUX2_X1 U15189 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13569), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15190 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13665), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15191 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13570), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15192 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13688), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15193 ( .A(n13709), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13589), .Z(
        P3_U3512) );
  MUX2_X1 U15194 ( .A(n13687), .B(P3_DATAO_REG_20__SCAN_IN), .S(n13589), .Z(
        P3_U3511) );
  MUX2_X1 U15195 ( .A(n13707), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13589), .Z(
        P3_U3510) );
  MUX2_X1 U15196 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13571), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15197 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13572), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15198 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13573), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15199 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13574), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15200 ( .A(n13575), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13589), .Z(
        P3_U3505) );
  MUX2_X1 U15201 ( .A(n13576), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13589), .Z(
        P3_U3504) );
  MUX2_X1 U15202 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13577), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15203 ( .A(n13578), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13589), .Z(
        P3_U3502) );
  MUX2_X1 U15204 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13579), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15205 ( .A(n13580), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13589), .Z(
        P3_U3500) );
  MUX2_X1 U15206 ( .A(n13581), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13589), .Z(
        P3_U3499) );
  MUX2_X1 U15207 ( .A(n13582), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13589), .Z(
        P3_U3498) );
  MUX2_X1 U15208 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13583), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15209 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13584), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15210 ( .A(n13585), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13589), .Z(
        P3_U3495) );
  MUX2_X1 U15211 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13586), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15212 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13587), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15213 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13588), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15214 ( .A(n13590), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13589), .Z(
        P3_U3491) );
  NOR2_X1 U15215 ( .A1(n13593), .A2(n13592), .ZN(n13819) );
  NOR2_X1 U15216 ( .A1(n15967), .A2(n13594), .ZN(n13603) );
  NOR3_X1 U15217 ( .A1(n13819), .A2(n7188), .A3(n13603), .ZN(n13598) );
  NOR2_X1 U15218 ( .A1(n13715), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13595) );
  OAI22_X1 U15219 ( .A1(n13821), .A2(n13754), .B1(n13598), .B2(n13595), .ZN(
        P3_U3202) );
  NOR2_X1 U15220 ( .A1(n13715), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13597) );
  OAI22_X1 U15221 ( .A1(n13824), .A2(n13754), .B1(n13598), .B2(n13597), .ZN(
        P3_U3203) );
  INV_X1 U15222 ( .A(n13599), .ZN(n13606) );
  NAND2_X1 U15223 ( .A1(n13600), .A2(n13715), .ZN(n13605) );
  NOR2_X1 U15224 ( .A1(n13601), .A2(n13754), .ZN(n13602) );
  AOI211_X1 U15225 ( .C1(n7188), .C2(P3_REG2_REG_29__SCAN_IN), .A(n13603), .B(
        n13602), .ZN(n13604) );
  OAI211_X1 U15226 ( .C1(n13606), .C2(n13717), .A(n13605), .B(n13604), .ZN(
        P3_U3204) );
  XNOR2_X1 U15227 ( .A(n13607), .B(n13608), .ZN(n13762) );
  INV_X1 U15228 ( .A(n13762), .ZN(n13617) );
  OAI22_X1 U15229 ( .A1(n13627), .A2(n15960), .B1(n13610), .B2(n15962), .ZN(
        n13611) );
  INV_X1 U15230 ( .A(n13611), .ZN(n13612) );
  AOI22_X1 U15231 ( .A1(n7188), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n15909), 
        .B2(n13613), .ZN(n13614) );
  OAI21_X1 U15232 ( .B1(n13828), .B2(n13754), .A(n13614), .ZN(n13615) );
  AOI21_X1 U15233 ( .B1(n13763), .B2(n13715), .A(n13615), .ZN(n13616) );
  OAI21_X1 U15234 ( .B1(n13617), .B2(n13717), .A(n13616), .ZN(P3_U3205) );
  INV_X1 U15235 ( .A(n13618), .ZN(n13624) );
  AOI22_X1 U15236 ( .A1(n7188), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n15909), 
        .B2(n13619), .ZN(n13620) );
  OAI21_X1 U15237 ( .B1(n13768), .B2(n13754), .A(n13620), .ZN(n13621) );
  AOI21_X1 U15238 ( .B1(n13622), .B2(n13715), .A(n13621), .ZN(n13623) );
  OAI21_X1 U15239 ( .B1(n13717), .B2(n13624), .A(n13623), .ZN(P3_U3206) );
  XOR2_X1 U15240 ( .A(n13625), .B(n13628), .Z(n13626) );
  OAI222_X1 U15241 ( .A1(n15962), .A2(n13627), .B1(n15960), .B2(n13656), .C1(
        n13626), .C2(n15959), .ZN(n13769) );
  INV_X1 U15242 ( .A(n13769), .ZN(n13634) );
  XOR2_X1 U15243 ( .A(n13629), .B(n13628), .Z(n13770) );
  AOI22_X1 U15244 ( .A1(n7188), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n15909), 
        .B2(n13630), .ZN(n13631) );
  OAI21_X1 U15245 ( .B1(n13832), .B2(n13754), .A(n13631), .ZN(n13632) );
  AOI21_X1 U15246 ( .B1(n13770), .B2(n13757), .A(n13632), .ZN(n13633) );
  OAI21_X1 U15247 ( .B1(n13634), .B2(n7188), .A(n13633), .ZN(P3_U3207) );
  XNOR2_X1 U15248 ( .A(n13636), .B(n13635), .ZN(n13643) );
  AOI22_X1 U15249 ( .A1(n13665), .A2(n13708), .B1(n9880), .B2(n13637), .ZN(
        n13642) );
  OAI211_X1 U15250 ( .C1(n13640), .C2(n13639), .A(n13638), .B(n13705), .ZN(
        n13641) );
  OAI211_X1 U15251 ( .C1(n13643), .C2(n13694), .A(n13642), .B(n13641), .ZN(
        n13773) );
  INV_X1 U15252 ( .A(n13773), .ZN(n13649) );
  INV_X1 U15253 ( .A(n13643), .ZN(n13774) );
  AOI22_X1 U15254 ( .A1(n7188), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15909), 
        .B2(n13644), .ZN(n13645) );
  OAI21_X1 U15255 ( .B1(n13836), .B2(n13754), .A(n13645), .ZN(n13646) );
  AOI21_X1 U15256 ( .B1(n13774), .B2(n13647), .A(n13646), .ZN(n13648) );
  OAI21_X1 U15257 ( .B1(n13649), .B2(n7188), .A(n13648), .ZN(P3_U3208) );
  XOR2_X1 U15258 ( .A(n13650), .B(n13654), .Z(n13778) );
  INV_X1 U15259 ( .A(n13778), .ZN(n13661) );
  INV_X1 U15260 ( .A(n13651), .ZN(n13652) );
  AOI21_X1 U15261 ( .B1(n13654), .B2(n13653), .A(n13652), .ZN(n13655) );
  OAI222_X1 U15262 ( .A1(n15962), .A2(n13656), .B1(n15960), .B2(n13676), .C1(
        n15959), .C2(n13655), .ZN(n13777) );
  AOI22_X1 U15263 ( .A1(n7188), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15909), 
        .B2(n13657), .ZN(n13658) );
  OAI21_X1 U15264 ( .B1(n13840), .B2(n13754), .A(n13658), .ZN(n13659) );
  AOI21_X1 U15265 ( .B1(n13777), .B2(n13715), .A(n13659), .ZN(n13660) );
  OAI21_X1 U15266 ( .B1(n13661), .B2(n13717), .A(n13660), .ZN(P3_U3209) );
  XOR2_X1 U15267 ( .A(n13662), .B(n13663), .Z(n13782) );
  INV_X1 U15268 ( .A(n13782), .ZN(n13672) );
  OAI211_X1 U15269 ( .C1(n7246), .C2(n7458), .A(n13705), .B(n13664), .ZN(
        n13667) );
  AOI22_X1 U15270 ( .A1(n13688), .A2(n13708), .B1(n9880), .B2(n13665), .ZN(
        n13666) );
  NAND2_X1 U15271 ( .A1(n13667), .A2(n13666), .ZN(n13781) );
  AOI22_X1 U15272 ( .A1(n7188), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15909), 
        .B2(n13668), .ZN(n13669) );
  OAI21_X1 U15273 ( .B1(n13844), .B2(n13754), .A(n13669), .ZN(n13670) );
  AOI21_X1 U15274 ( .B1(n13781), .B2(n13715), .A(n13670), .ZN(n13671) );
  OAI21_X1 U15275 ( .B1(n13672), .B2(n13717), .A(n13671), .ZN(P3_U3210) );
  XNOR2_X1 U15276 ( .A(n13673), .B(n13678), .ZN(n13674) );
  OAI222_X1 U15277 ( .A1(n15962), .A2(n13676), .B1(n15960), .B2(n13675), .C1(
        n15959), .C2(n13674), .ZN(n13785) );
  INV_X1 U15278 ( .A(n13785), .ZN(n13683) );
  XOR2_X1 U15279 ( .A(n13678), .B(n13677), .Z(n13786) );
  AOI22_X1 U15280 ( .A1(n13679), .A2(n15909), .B1(n7188), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n13680) );
  OAI21_X1 U15281 ( .B1(n13848), .B2(n13754), .A(n13680), .ZN(n13681) );
  AOI21_X1 U15282 ( .B1(n13786), .B2(n13757), .A(n13681), .ZN(n13682) );
  OAI21_X1 U15283 ( .B1(n13683), .B2(n7188), .A(n13682), .ZN(P3_U3211) );
  OR2_X1 U15284 ( .A1(n13684), .A2(n13689), .ZN(n13685) );
  NAND2_X1 U15285 ( .A1(n13686), .A2(n13685), .ZN(n13789) );
  AOI22_X1 U15286 ( .A1(n13688), .A2(n9880), .B1(n13708), .B2(n13687), .ZN(
        n13693) );
  XNOR2_X1 U15287 ( .A(n13690), .B(n13689), .ZN(n13691) );
  NAND2_X1 U15288 ( .A1(n13691), .A2(n13705), .ZN(n13692) );
  OAI211_X1 U15289 ( .C1(n13789), .C2(n13694), .A(n13693), .B(n13692), .ZN(
        n13790) );
  AOI22_X1 U15290 ( .A1(n7188), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13695), 
        .B2(n15909), .ZN(n13699) );
  NAND2_X1 U15291 ( .A1(n13697), .A2(n13696), .ZN(n13698) );
  OAI211_X1 U15292 ( .C1(n13789), .C2(n13700), .A(n13699), .B(n13698), .ZN(
        n13701) );
  AOI21_X1 U15293 ( .B1(n13790), .B2(n13715), .A(n13701), .ZN(n13702) );
  INV_X1 U15294 ( .A(n13702), .ZN(P3_U3212) );
  XOR2_X1 U15295 ( .A(n13704), .B(n13703), .Z(n13795) );
  INV_X1 U15296 ( .A(n13795), .ZN(n13718) );
  OAI211_X1 U15297 ( .C1(n7312), .C2(n7903), .A(n13706), .B(n13705), .ZN(
        n13711) );
  AOI22_X1 U15298 ( .A1(n13709), .A2(n9880), .B1(n13708), .B2(n13707), .ZN(
        n13710) );
  NAND2_X1 U15299 ( .A1(n13711), .A2(n13710), .ZN(n13794) );
  AOI22_X1 U15300 ( .A1(n7188), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15909), 
        .B2(n13712), .ZN(n13713) );
  OAI21_X1 U15301 ( .B1(n13856), .B2(n13754), .A(n13713), .ZN(n13714) );
  AOI21_X1 U15302 ( .B1(n13794), .B2(n13715), .A(n13714), .ZN(n13716) );
  OAI21_X1 U15303 ( .B1(n13718), .B2(n13717), .A(n13716), .ZN(P3_U3213) );
  XNOR2_X1 U15304 ( .A(n13719), .B(n13722), .ZN(n13720) );
  OAI222_X1 U15305 ( .A1(n15962), .A2(n13721), .B1(n15960), .B2(n13745), .C1(
        n15959), .C2(n13720), .ZN(n13798) );
  INV_X1 U15306 ( .A(n13798), .ZN(n13728) );
  XNOR2_X1 U15307 ( .A(n13723), .B(n13722), .ZN(n13799) );
  AOI22_X1 U15308 ( .A1(n7188), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15909), 
        .B2(n13724), .ZN(n13725) );
  OAI21_X1 U15309 ( .B1(n13860), .B2(n13754), .A(n13725), .ZN(n13726) );
  AOI21_X1 U15310 ( .B1(n13799), .B2(n13757), .A(n13726), .ZN(n13727) );
  OAI21_X1 U15311 ( .B1(n13728), .B2(n7188), .A(n13727), .ZN(P3_U3214) );
  AOI21_X1 U15312 ( .B1(n13729), .B2(n13731), .A(n13730), .ZN(n13732) );
  NOR2_X1 U15313 ( .A1(n7307), .A2(n13732), .ZN(n13733) );
  OAI222_X1 U15314 ( .A1(n15962), .A2(n13735), .B1(n15960), .B2(n13734), .C1(
        n15959), .C2(n13733), .ZN(n13802) );
  INV_X1 U15315 ( .A(n13802), .ZN(n13743) );
  OAI21_X1 U15316 ( .B1(n13738), .B2(n13737), .A(n13736), .ZN(n13803) );
  AOI22_X1 U15317 ( .A1(n7188), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15909), 
        .B2(n13739), .ZN(n13740) );
  OAI21_X1 U15318 ( .B1(n13865), .B2(n13754), .A(n13740), .ZN(n13741) );
  AOI21_X1 U15319 ( .B1(n13803), .B2(n13757), .A(n13741), .ZN(n13742) );
  OAI21_X1 U15320 ( .B1(n13743), .B2(n7188), .A(n13742), .ZN(P3_U3215) );
  AOI21_X1 U15321 ( .B1(n13744), .B2(n13750), .A(n15959), .ZN(n13748) );
  OAI22_X1 U15322 ( .A1(n13746), .A2(n15960), .B1(n13745), .B2(n15962), .ZN(
        n13747) );
  AOI21_X1 U15323 ( .B1(n13748), .B2(n13729), .A(n13747), .ZN(n13809) );
  OAI21_X1 U15324 ( .B1(n13751), .B2(n13750), .A(n13749), .ZN(n13808) );
  AOI22_X1 U15325 ( .A1(n7188), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15909), 
        .B2(n13752), .ZN(n13753) );
  OAI21_X1 U15326 ( .B1(n13755), .B2(n13754), .A(n13753), .ZN(n13756) );
  AOI21_X1 U15327 ( .B1(n13808), .B2(n13757), .A(n13756), .ZN(n13758) );
  OAI21_X1 U15328 ( .B1(n13809), .B2(n7188), .A(n13758), .ZN(P3_U3216) );
  NAND2_X1 U15329 ( .A1(n13819), .A2(n16165), .ZN(n13760) );
  NAND2_X1 U15330 ( .A1(n9674), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13759) );
  OAI211_X1 U15331 ( .C1(n13821), .C2(n13806), .A(n13760), .B(n13759), .ZN(
        P3_U3490) );
  NAND2_X1 U15332 ( .A1(n9674), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13761) );
  OAI211_X1 U15333 ( .C1(n13824), .C2(n13806), .A(n13761), .B(n13760), .ZN(
        P3_U3489) );
  INV_X1 U15334 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13764) );
  INV_X1 U15335 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13766) );
  MUX2_X1 U15336 ( .A(n13766), .B(n13765), .S(n16165), .Z(n13767) );
  OAI21_X1 U15337 ( .B1(n13768), .B2(n13806), .A(n13767), .ZN(P3_U3486) );
  INV_X1 U15338 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13771) );
  AOI21_X1 U15339 ( .B1(n16160), .B2(n13770), .A(n13769), .ZN(n13829) );
  MUX2_X1 U15340 ( .A(n13771), .B(n13829), .S(n16165), .Z(n13772) );
  OAI21_X1 U15341 ( .B1(n13832), .B2(n13806), .A(n13772), .ZN(P3_U3485) );
  INV_X1 U15342 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13775) );
  AOI21_X1 U15343 ( .B1(n16103), .B2(n13774), .A(n13773), .ZN(n13833) );
  MUX2_X1 U15344 ( .A(n13775), .B(n13833), .S(n16165), .Z(n13776) );
  OAI21_X1 U15345 ( .B1(n13836), .B2(n13806), .A(n13776), .ZN(P3_U3484) );
  INV_X1 U15346 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13779) );
  AOI21_X1 U15347 ( .B1(n16160), .B2(n13778), .A(n13777), .ZN(n13837) );
  MUX2_X1 U15348 ( .A(n13779), .B(n13837), .S(n16165), .Z(n13780) );
  OAI21_X1 U15349 ( .B1(n13840), .B2(n13806), .A(n13780), .ZN(P3_U3483) );
  INV_X1 U15350 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13783) );
  AOI21_X1 U15351 ( .B1(n13782), .B2(n16160), .A(n13781), .ZN(n13841) );
  MUX2_X1 U15352 ( .A(n13783), .B(n13841), .S(n16165), .Z(n13784) );
  OAI21_X1 U15353 ( .B1(n13844), .B2(n13806), .A(n13784), .ZN(P3_U3482) );
  INV_X1 U15354 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13787) );
  AOI21_X1 U15355 ( .B1(n16160), .B2(n13786), .A(n13785), .ZN(n13845) );
  MUX2_X1 U15356 ( .A(n13787), .B(n13845), .S(n16165), .Z(n13788) );
  OAI21_X1 U15357 ( .B1(n13848), .B2(n13806), .A(n13788), .ZN(P3_U3481) );
  INV_X1 U15358 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13792) );
  INV_X1 U15359 ( .A(n13789), .ZN(n13791) );
  AOI21_X1 U15360 ( .B1(n16103), .B2(n13791), .A(n13790), .ZN(n13849) );
  MUX2_X1 U15361 ( .A(n13792), .B(n13849), .S(n16165), .Z(n13793) );
  OAI21_X1 U15362 ( .B1(n13852), .B2(n13806), .A(n13793), .ZN(P3_U3480) );
  INV_X1 U15363 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13796) );
  AOI21_X1 U15364 ( .B1(n13795), .B2(n16160), .A(n13794), .ZN(n13853) );
  MUX2_X1 U15365 ( .A(n13796), .B(n13853), .S(n16165), .Z(n13797) );
  OAI21_X1 U15366 ( .B1(n13856), .B2(n13806), .A(n13797), .ZN(P3_U3479) );
  INV_X1 U15367 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13800) );
  AOI21_X1 U15368 ( .B1(n13799), .B2(n16160), .A(n13798), .ZN(n13857) );
  MUX2_X1 U15369 ( .A(n13800), .B(n13857), .S(n16165), .Z(n13801) );
  OAI21_X1 U15370 ( .B1(n13806), .B2(n13860), .A(n13801), .ZN(P3_U3478) );
  INV_X1 U15371 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13804) );
  AOI21_X1 U15372 ( .B1(n16160), .B2(n13803), .A(n13802), .ZN(n13861) );
  MUX2_X1 U15373 ( .A(n13804), .B(n13861), .S(n16165), .Z(n13805) );
  OAI21_X1 U15374 ( .B1(n13865), .B2(n13806), .A(n13805), .ZN(P3_U3477) );
  AOI22_X1 U15375 ( .A1(n13808), .A2(n16160), .B1(n16107), .B2(n13807), .ZN(
        n13810) );
  NAND2_X1 U15376 ( .A1(n13810), .A2(n13809), .ZN(n13866) );
  MUX2_X1 U15377 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13866), .S(n16165), .Z(
        P3_U3476) );
  AOI22_X1 U15378 ( .A1(n13812), .A2(n16160), .B1(n16107), .B2(n13811), .ZN(
        n13813) );
  NAND2_X1 U15379 ( .A1(n13814), .A2(n13813), .ZN(n13867) );
  MUX2_X1 U15380 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13867), .S(n16165), .Z(
        P3_U3475) );
  AOI22_X1 U15381 ( .A1(n13816), .A2(n16160), .B1(n16107), .B2(n13815), .ZN(
        n13817) );
  NAND2_X1 U15382 ( .A1(n13818), .A2(n13817), .ZN(n13868) );
  MUX2_X1 U15383 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13868), .S(n16165), .Z(
        P3_U3474) );
  NAND2_X1 U15384 ( .A1(n13819), .A2(n16169), .ZN(n13822) );
  NAND2_X1 U15385 ( .A1(n16166), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13820) );
  OAI211_X1 U15386 ( .C1(n13821), .C2(n13864), .A(n13822), .B(n13820), .ZN(
        P3_U3458) );
  NAND2_X1 U15387 ( .A1(n16166), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13823) );
  OAI211_X1 U15388 ( .C1(n13824), .C2(n13864), .A(n13823), .B(n13822), .ZN(
        P3_U3457) );
  INV_X1 U15389 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13826) );
  OAI21_X1 U15390 ( .B1(n13828), .B2(n13864), .A(n13827), .ZN(P3_U3455) );
  INV_X1 U15391 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13830) );
  MUX2_X1 U15392 ( .A(n13830), .B(n13829), .S(n16169), .Z(n13831) );
  OAI21_X1 U15393 ( .B1(n13832), .B2(n13864), .A(n13831), .ZN(P3_U3453) );
  INV_X1 U15394 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13834) );
  MUX2_X1 U15395 ( .A(n13834), .B(n13833), .S(n16169), .Z(n13835) );
  OAI21_X1 U15396 ( .B1(n13836), .B2(n13864), .A(n13835), .ZN(P3_U3452) );
  INV_X1 U15397 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13838) );
  MUX2_X1 U15398 ( .A(n13838), .B(n13837), .S(n16169), .Z(n13839) );
  OAI21_X1 U15399 ( .B1(n13840), .B2(n13864), .A(n13839), .ZN(P3_U3451) );
  INV_X1 U15400 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13842) );
  MUX2_X1 U15401 ( .A(n13842), .B(n13841), .S(n16169), .Z(n13843) );
  OAI21_X1 U15402 ( .B1(n13844), .B2(n13864), .A(n13843), .ZN(P3_U3450) );
  MUX2_X1 U15403 ( .A(n13846), .B(n13845), .S(n16169), .Z(n13847) );
  OAI21_X1 U15404 ( .B1(n13848), .B2(n13864), .A(n13847), .ZN(P3_U3449) );
  INV_X1 U15405 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13850) );
  MUX2_X1 U15406 ( .A(n13850), .B(n13849), .S(n16169), .Z(n13851) );
  OAI21_X1 U15407 ( .B1(n13852), .B2(n13864), .A(n13851), .ZN(P3_U3448) );
  INV_X1 U15408 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13854) );
  MUX2_X1 U15409 ( .A(n13854), .B(n13853), .S(n16169), .Z(n13855) );
  OAI21_X1 U15410 ( .B1(n13856), .B2(n13864), .A(n13855), .ZN(P3_U3447) );
  INV_X1 U15411 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13858) );
  MUX2_X1 U15412 ( .A(n13858), .B(n13857), .S(n16169), .Z(n13859) );
  OAI21_X1 U15413 ( .B1(n13864), .B2(n13860), .A(n13859), .ZN(P3_U3446) );
  INV_X1 U15414 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13862) );
  MUX2_X1 U15415 ( .A(n13862), .B(n13861), .S(n16169), .Z(n13863) );
  OAI21_X1 U15416 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(P3_U3444) );
  MUX2_X1 U15417 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13866), .S(n16169), .Z(
        P3_U3441) );
  MUX2_X1 U15418 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13867), .S(n16169), .Z(
        P3_U3438) );
  MUX2_X1 U15419 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13868), .S(n16169), .Z(
        P3_U3435) );
  MUX2_X1 U15420 ( .A(P3_D_REG_1__SCAN_IN), .B(n13869), .S(n13870), .Z(
        P3_U3377) );
  MUX2_X1 U15421 ( .A(P3_D_REG_0__SCAN_IN), .B(n13871), .S(n13870), .Z(
        P3_U3376) );
  NAND3_X1 U15422 ( .A1(n13872), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13874) );
  OAI22_X1 U15423 ( .A1(n9076), .A2(n13874), .B1(n13873), .B2(n13880), .ZN(
        n13875) );
  AOI21_X1 U15424 ( .B1(n13877), .B2(n13876), .A(n13875), .ZN(n13878) );
  INV_X1 U15425 ( .A(n13878), .ZN(P3_U3264) );
  INV_X1 U15426 ( .A(n13879), .ZN(n13882) );
  OAI222_X1 U15427 ( .A1(n13131), .A2(n13882), .B1(n13881), .B2(P3_U3151), 
        .C1(n15277), .C2(n13880), .ZN(P3_U3266) );
  MUX2_X1 U15428 ( .A(n13884), .B(n13883), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3294) );
  XNOR2_X1 U15429 ( .A(n13885), .B(n13886), .ZN(n13893) );
  NOR2_X1 U15430 ( .A1(n14101), .A2(n13992), .ZN(n13891) );
  AOI22_X1 U15431 ( .A1(n13887), .A2(n13994), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13888) );
  OAI21_X1 U15432 ( .B1(n13889), .B2(n13996), .A(n13888), .ZN(n13890) );
  AOI211_X1 U15433 ( .C1(n14271), .C2(n13999), .A(n13891), .B(n13890), .ZN(
        n13892) );
  OAI21_X1 U15434 ( .B1(n13893), .B2(n14001), .A(n13892), .ZN(P2_U3186) );
  INV_X1 U15435 ( .A(n14008), .ZN(n13894) );
  OAI22_X1 U15436 ( .A1(n14100), .A2(n14191), .B1(n13894), .B2(n14189), .ZN(
        n14129) );
  INV_X1 U15437 ( .A(n14129), .ZN(n13896) );
  AOI22_X1 U15438 ( .A1(n13994), .A2(n14136), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13895) );
  OAI21_X1 U15439 ( .B1(n13896), .B2(n13984), .A(n13895), .ZN(n13900) );
  NOR3_X1 U15440 ( .A1(n13898), .A2(n14145), .A3(n13897), .ZN(n13899) );
  AOI211_X1 U15441 ( .C1(n14295), .C2(n13999), .A(n13900), .B(n13899), .ZN(
        n13901) );
  OAI21_X1 U15442 ( .B1(n13902), .B2(n14001), .A(n13901), .ZN(P2_U3188) );
  XNOR2_X1 U15443 ( .A(n13904), .B(n13903), .ZN(n13910) );
  NOR2_X1 U15444 ( .A1(n13992), .A2(n14190), .ZN(n13908) );
  NAND2_X1 U15445 ( .A1(n13994), .A2(n14203), .ZN(n13906) );
  OAI211_X1 U15446 ( .C1(n13996), .C2(n14192), .A(n13906), .B(n13905), .ZN(
        n13907) );
  AOI211_X1 U15447 ( .C1(n14317), .C2(n13999), .A(n13908), .B(n13907), .ZN(
        n13909) );
  OAI21_X1 U15448 ( .B1(n13910), .B2(n14001), .A(n13909), .ZN(P2_U3191) );
  XNOR2_X1 U15449 ( .A(n13912), .B(n13911), .ZN(n13918) );
  AND2_X1 U15450 ( .A1(n14010), .A2(n14089), .ZN(n13913) );
  AOI21_X1 U15451 ( .B1(n14008), .B2(n14091), .A(n13913), .ZN(n14165) );
  INV_X1 U15452 ( .A(n13914), .ZN(n14169) );
  AOI22_X1 U15453 ( .A1(n13994), .A2(n14169), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13915) );
  OAI21_X1 U15454 ( .B1(n14165), .B2(n13984), .A(n13915), .ZN(n13916) );
  AOI21_X1 U15455 ( .B1(n14309), .B2(n13999), .A(n13916), .ZN(n13917) );
  OAI21_X1 U15456 ( .B1(n13918), .B2(n14001), .A(n13917), .ZN(P2_U3195) );
  XNOR2_X1 U15457 ( .A(n13919), .B(n13920), .ZN(n13925) );
  NOR2_X1 U15458 ( .A1(n13992), .A2(n14100), .ZN(n13923) );
  AOI22_X1 U15459 ( .A1(n14105), .A2(n13994), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13921) );
  OAI21_X1 U15460 ( .B1(n14101), .B2(n13996), .A(n13921), .ZN(n13922) );
  AOI211_X1 U15461 ( .C1(n14285), .C2(n13999), .A(n13923), .B(n13922), .ZN(
        n13924) );
  OAI21_X1 U15462 ( .B1(n13925), .B2(n14001), .A(n13924), .ZN(P2_U3197) );
  OAI21_X1 U15463 ( .B1(n13928), .B2(n13927), .A(n13926), .ZN(n13929) );
  NAND2_X1 U15464 ( .A1(n13929), .A2(n13940), .ZN(n13936) );
  NOR2_X1 U15465 ( .A1(n13931), .A2(n13930), .ZN(n13934) );
  NOR2_X1 U15466 ( .A1(n13984), .A2(n13932), .ZN(n13933) );
  AOI211_X1 U15467 ( .C1(P2_REG3_REG_16__SCAN_IN), .C2(P2_U3088), .A(n13934), 
        .B(n13933), .ZN(n13935) );
  OAI211_X1 U15468 ( .C1(n7762), .C2(n13978), .A(n13936), .B(n13935), .ZN(
        P2_U3198) );
  OAI21_X1 U15469 ( .B1(n13939), .B2(n13938), .A(n13937), .ZN(n13941) );
  NAND2_X1 U15470 ( .A1(n13941), .A2(n13940), .ZN(n13947) );
  INV_X1 U15471 ( .A(n14233), .ZN(n13945) );
  AND2_X1 U15472 ( .A1(n14014), .A2(n14089), .ZN(n13942) );
  AOI21_X1 U15473 ( .B1(n14012), .B2(n14091), .A(n13942), .ZN(n14240) );
  NOR2_X1 U15474 ( .A1(n13984), .A2(n14240), .ZN(n13943) );
  AOI211_X1 U15475 ( .C1(n13994), .C2(n13945), .A(n13944), .B(n13943), .ZN(
        n13946) );
  OAI211_X1 U15476 ( .C1(n14232), .C2(n13978), .A(n13947), .B(n13946), .ZN(
        P2_U3200) );
  AOI21_X1 U15477 ( .B1(n13949), .B2(n13948), .A(n14001), .ZN(n13951) );
  NAND2_X1 U15478 ( .A1(n13951), .A2(n13950), .ZN(n13957) );
  INV_X1 U15479 ( .A(n13952), .ZN(n14123) );
  AOI22_X1 U15480 ( .A1(n14123), .A2(n13994), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13953) );
  OAI21_X1 U15481 ( .B1(n14118), .B2(n13996), .A(n13953), .ZN(n13954) );
  AOI21_X1 U15482 ( .B1(n13955), .B2(n14007), .A(n13954), .ZN(n13956) );
  OAI211_X1 U15483 ( .C1(n7765), .C2(n13978), .A(n13957), .B(n13956), .ZN(
        P2_U3201) );
  OAI21_X1 U15484 ( .B1(n13960), .B2(n13959), .A(n13958), .ZN(n13961) );
  INV_X1 U15485 ( .A(n13961), .ZN(n13967) );
  AND2_X1 U15486 ( .A1(n14011), .A2(n14089), .ZN(n13962) );
  AOI21_X1 U15487 ( .B1(n14009), .B2(n14091), .A(n13962), .ZN(n14178) );
  INV_X1 U15488 ( .A(n13963), .ZN(n14182) );
  AOI22_X1 U15489 ( .A1(n13994), .A2(n14182), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13964) );
  OAI21_X1 U15490 ( .B1(n13984), .B2(n14178), .A(n13964), .ZN(n13965) );
  AOI21_X1 U15491 ( .B1(n14314), .B2(n13999), .A(n13965), .ZN(n13966) );
  OAI21_X1 U15492 ( .B1(n13967), .B2(n14001), .A(n13966), .ZN(P2_U3205) );
  NAND2_X1 U15493 ( .A1(n13968), .A2(n14008), .ZN(n13972) );
  OR2_X1 U15494 ( .A1(n14001), .A2(n13969), .ZN(n13971) );
  MUX2_X1 U15495 ( .A(n13972), .B(n13971), .S(n13970), .Z(n13977) );
  AOI22_X1 U15496 ( .A1(n13994), .A2(n14155), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13973) );
  OAI21_X1 U15497 ( .B1(n13992), .B2(n14144), .A(n13973), .ZN(n13974) );
  AOI21_X1 U15498 ( .B1(n13975), .B2(n14007), .A(n13974), .ZN(n13976) );
  OAI211_X1 U15499 ( .C1(n14152), .C2(n13978), .A(n13977), .B(n13976), .ZN(
        P2_U3207) );
  XNOR2_X1 U15500 ( .A(n13980), .B(n13979), .ZN(n13987) );
  AND2_X1 U15501 ( .A1(n14013), .A2(n14089), .ZN(n13981) );
  AOI21_X1 U15502 ( .B1(n14011), .B2(n14091), .A(n13981), .ZN(n14213) );
  INV_X1 U15503 ( .A(n13982), .ZN(n14218) );
  AOI22_X1 U15504 ( .A1(n13994), .A2(n14218), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13983) );
  OAI21_X1 U15505 ( .B1(n13984), .B2(n14213), .A(n13983), .ZN(n13985) );
  AOI21_X1 U15506 ( .B1(n14327), .B2(n13999), .A(n13985), .ZN(n13986) );
  OAI21_X1 U15507 ( .B1(n13987), .B2(n14001), .A(n13986), .ZN(P2_U3210) );
  INV_X1 U15508 ( .A(n13989), .ZN(n13990) );
  AOI21_X1 U15509 ( .B1(n13991), .B2(n13988), .A(n13990), .ZN(n14002) );
  NOR2_X1 U15510 ( .A1(n14118), .A2(n13992), .ZN(n13998) );
  INV_X1 U15511 ( .A(n13993), .ZN(n14084) );
  AOI22_X1 U15512 ( .A1(n14084), .A2(n13994), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13995) );
  OAI21_X1 U15513 ( .B1(n14044), .B2(n13996), .A(n13995), .ZN(n13997) );
  AOI211_X1 U15514 ( .C1(n14278), .C2(n13999), .A(n13998), .B(n13997), .ZN(
        n14000) );
  OAI21_X1 U15515 ( .B1(n14002), .B2(n14001), .A(n14000), .ZN(P2_U3212) );
  MUX2_X1 U15516 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n14003), .S(n15405), .Z(
        P2_U3562) );
  MUX2_X1 U15517 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n14048), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15518 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n14004), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15519 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n14054), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15520 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n14092), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15521 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n14005), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15522 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n14090), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15523 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n14006), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15524 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n14007), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15525 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14008), .S(n15405), .Z(
        P2_U3553) );
  MUX2_X1 U15526 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n14009), .S(n15405), .Z(
        P2_U3552) );
  MUX2_X1 U15527 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n14010), .S(n15405), .Z(
        P2_U3551) );
  MUX2_X1 U15528 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n14011), .S(n15405), .Z(
        P2_U3550) );
  MUX2_X1 U15529 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n14012), .S(n15405), .Z(
        P2_U3549) );
  MUX2_X1 U15530 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n14013), .S(n15405), .Z(
        P2_U3548) );
  MUX2_X1 U15531 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n14014), .S(n15405), .Z(
        P2_U3547) );
  MUX2_X1 U15532 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n14015), .S(n15405), .Z(
        P2_U3546) );
  MUX2_X1 U15533 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n14016), .S(n15405), .Z(
        P2_U3545) );
  MUX2_X1 U15534 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n14017), .S(n15405), .Z(
        P2_U3543) );
  MUX2_X1 U15535 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n14018), .S(n15405), .Z(
        P2_U3542) );
  MUX2_X1 U15536 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n14019), .S(n15405), .Z(
        P2_U3541) );
  MUX2_X1 U15537 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n14020), .S(n15405), .Z(
        P2_U3540) );
  MUX2_X1 U15538 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n14021), .S(n15405), .Z(
        P2_U3539) );
  MUX2_X1 U15539 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n14022), .S(n15405), .Z(
        P2_U3538) );
  MUX2_X1 U15540 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n14023), .S(n15405), .Z(
        P2_U3537) );
  MUX2_X1 U15541 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n14024), .S(n15405), .Z(
        P2_U3536) );
  MUX2_X1 U15542 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n14025), .S(n15405), .Z(
        P2_U3535) );
  MUX2_X1 U15543 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n14026), .S(n15405), .Z(
        P2_U3534) );
  MUX2_X1 U15544 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n14027), .S(n15405), .Z(
        P2_U3533) );
  MUX2_X1 U15545 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13144), .S(n15405), .Z(
        P2_U3532) );
  INV_X1 U15546 ( .A(n14260), .ZN(n14061) );
  XNOR2_X1 U15547 ( .A(n14036), .B(n14032), .ZN(n14028) );
  NAND2_X1 U15548 ( .A1(n14028), .A2(n14302), .ZN(n14254) );
  NAND2_X1 U15549 ( .A1(n14029), .A2(P2_B_REG_SCAN_IN), .ZN(n14030) );
  NAND2_X1 U15550 ( .A1(n14091), .A2(n14030), .ZN(n14050) );
  OR2_X1 U15551 ( .A1(n14031), .A2(n14050), .ZN(n14256) );
  NOR2_X1 U15552 ( .A1(n16156), .A2(n14256), .ZN(n14040) );
  INV_X1 U15553 ( .A(n14032), .ZN(n14255) );
  NOR2_X1 U15554 ( .A1(n14255), .A2(n14231), .ZN(n14033) );
  AOI211_X1 U15555 ( .C1(n16156), .C2(P2_REG2_REG_31__SCAN_IN), .A(n14040), 
        .B(n14033), .ZN(n14034) );
  OAI21_X1 U15556 ( .B1(n16045), .B2(n14254), .A(n14034), .ZN(P2_U3234) );
  INV_X1 U15557 ( .A(n14060), .ZN(n14038) );
  OAI211_X1 U15558 ( .C1(n14258), .C2(n14038), .A(n14037), .B(n14302), .ZN(
        n14257) );
  NOR2_X1 U15559 ( .A1(n14258), .A2(n14231), .ZN(n14039) );
  AOI211_X1 U15560 ( .C1(n16156), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14040), 
        .B(n14039), .ZN(n14041) );
  OAI21_X1 U15561 ( .B1(n16045), .B2(n14257), .A(n14041), .ZN(P2_U3235) );
  NAND2_X1 U15562 ( .A1(n14069), .A2(n14045), .ZN(n14047) );
  INV_X1 U15563 ( .A(n14056), .ZN(n14046) );
  XNOR2_X1 U15564 ( .A(n14047), .B(n14046), .ZN(n14053) );
  INV_X1 U15565 ( .A(n14048), .ZN(n14051) );
  NAND2_X1 U15566 ( .A1(n14054), .A2(n14089), .ZN(n14049) );
  OAI21_X1 U15567 ( .B1(n14051), .B2(n14050), .A(n14049), .ZN(n14052) );
  NAND2_X1 U15568 ( .A1(n14071), .A2(n14055), .ZN(n14057) );
  XNOR2_X1 U15569 ( .A(n14057), .B(n14046), .ZN(n14259) );
  NAND2_X1 U15570 ( .A1(n14259), .A2(n14151), .ZN(n14065) );
  INV_X1 U15571 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n14058) );
  OAI22_X1 U15572 ( .A1(n14059), .A2(n16038), .B1(n14058), .B2(n16041), .ZN(
        n14063) );
  OAI211_X1 U15573 ( .C1(n14074), .C2(n14061), .A(n14302), .B(n14060), .ZN(
        n14261) );
  NOR2_X1 U15574 ( .A1(n14261), .A2(n16045), .ZN(n14062) );
  AOI211_X1 U15575 ( .C1(n16147), .C2(n14260), .A(n14063), .B(n14062), .ZN(
        n14064) );
  OAI211_X1 U15576 ( .C1(n14263), .C2(n16156), .A(n14065), .B(n14064), .ZN(
        P2_U3236) );
  AOI21_X1 U15577 ( .B1(n14066), .B2(n14072), .A(n14214), .ZN(n14070) );
  INV_X1 U15578 ( .A(n14067), .ZN(n14068) );
  AOI21_X1 U15579 ( .B1(n14070), .B2(n14069), .A(n14068), .ZN(n14269) );
  OAI21_X1 U15580 ( .B1(n14073), .B2(n14072), .A(n14071), .ZN(n14265) );
  NAND2_X1 U15581 ( .A1(n14265), .A2(n14151), .ZN(n14080) );
  AOI211_X1 U15582 ( .C1(n14267), .C2(n14075), .A(n14319), .B(n14074), .ZN(
        n14266) );
  AOI22_X1 U15583 ( .A1(n14076), .A2(n16146), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n16156), .ZN(n14077) );
  OAI21_X1 U15584 ( .B1(n7758), .B2(n14231), .A(n14077), .ZN(n14078) );
  AOI21_X1 U15585 ( .B1(n14266), .B2(n16150), .A(n14078), .ZN(n14079) );
  OAI211_X1 U15586 ( .C1(n16156), .C2(n14269), .A(n14080), .B(n14079), .ZN(
        P2_U3237) );
  XNOR2_X1 U15587 ( .A(n14081), .B(n14087), .ZN(n14282) );
  INV_X1 U15588 ( .A(n14082), .ZN(n14083) );
  AOI21_X1 U15589 ( .B1(n14278), .B2(n14102), .A(n14083), .ZN(n14279) );
  INV_X1 U15590 ( .A(n14278), .ZN(n14086) );
  AOI22_X1 U15591 ( .A1(n16156), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n14084), 
        .B2(n16146), .ZN(n14085) );
  OAI21_X1 U15592 ( .B1(n14086), .B2(n14231), .A(n14085), .ZN(n14095) );
  XNOR2_X1 U15593 ( .A(n14088), .B(n14087), .ZN(n14093) );
  AOI222_X1 U15594 ( .A1(n14236), .A2(n14093), .B1(n14092), .B2(n14091), .C1(
        n14090), .C2(n14089), .ZN(n14281) );
  NOR2_X1 U15595 ( .A1(n14281), .A2(n16156), .ZN(n14094) );
  AOI211_X1 U15596 ( .C1(n14159), .C2(n14279), .A(n14095), .B(n14094), .ZN(
        n14096) );
  OAI21_X1 U15597 ( .B1(n14244), .B2(n14282), .A(n14096), .ZN(P2_U3239) );
  XOR2_X1 U15598 ( .A(n14099), .B(n14097), .Z(n14287) );
  INV_X1 U15599 ( .A(n14122), .ZN(n14104) );
  INV_X1 U15600 ( .A(n14102), .ZN(n14103) );
  AOI211_X1 U15601 ( .C1(n14285), .C2(n14104), .A(n14319), .B(n14103), .ZN(
        n14284) );
  NAND2_X1 U15602 ( .A1(n14284), .A2(n16150), .ZN(n14107) );
  AOI22_X1 U15603 ( .A1(n16156), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n14105), 
        .B2(n16146), .ZN(n14106) );
  OAI211_X1 U15604 ( .C1(n14108), .C2(n14231), .A(n14107), .B(n14106), .ZN(
        n14109) );
  AOI21_X1 U15605 ( .B1(n14283), .B2(n16041), .A(n14109), .ZN(n14110) );
  OAI21_X1 U15606 ( .B1(n14287), .B2(n14244), .A(n14110), .ZN(P2_U3240) );
  OR2_X1 U15607 ( .A1(n14111), .A2(n14114), .ZN(n14112) );
  NAND2_X1 U15608 ( .A1(n14115), .A2(n14114), .ZN(n14116) );
  AOI21_X1 U15609 ( .B1(n14117), .B2(n14116), .A(n14214), .ZN(n14120) );
  OAI22_X1 U15610 ( .A1(n14118), .A2(n14191), .B1(n14145), .B2(n14189), .ZN(
        n14119) );
  AOI211_X1 U15611 ( .C1(n14288), .C2(n14121), .A(n14120), .B(n14119), .ZN(
        n14292) );
  AOI211_X1 U15612 ( .C1(n14290), .C2(n14134), .A(n14319), .B(n14122), .ZN(
        n14289) );
  NAND2_X1 U15613 ( .A1(n14289), .A2(n16150), .ZN(n14125) );
  AOI22_X1 U15614 ( .A1(n16156), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n14123), 
        .B2(n16146), .ZN(n14124) );
  OAI211_X1 U15615 ( .C1(n7765), .C2(n14231), .A(n14125), .B(n14124), .ZN(
        n14126) );
  AOI21_X1 U15616 ( .B1(n14288), .B2(n16151), .A(n14126), .ZN(n14127) );
  OAI21_X1 U15617 ( .B1(n14292), .B2(n16156), .A(n14127), .ZN(P2_U3241) );
  XNOR2_X1 U15618 ( .A(n14128), .B(n14132), .ZN(n14130) );
  AOI21_X1 U15619 ( .B1(n14130), .B2(n14236), .A(n14129), .ZN(n14297) );
  OAI21_X1 U15620 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(n14298) );
  INV_X1 U15621 ( .A(n14298), .ZN(n14141) );
  INV_X1 U15622 ( .A(n14295), .ZN(n14139) );
  AOI21_X1 U15623 ( .B1(n14154), .B2(n14295), .A(n14319), .ZN(n14135) );
  AND2_X1 U15624 ( .A1(n14135), .A2(n14134), .ZN(n14294) );
  NAND2_X1 U15625 ( .A1(n14294), .A2(n16150), .ZN(n14138) );
  AOI22_X1 U15626 ( .A1(n16156), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14136), 
        .B2(n16146), .ZN(n14137) );
  OAI211_X1 U15627 ( .C1(n14139), .C2(n14231), .A(n14138), .B(n14137), .ZN(
        n14140) );
  AOI21_X1 U15628 ( .B1(n14141), .B2(n14151), .A(n14140), .ZN(n14142) );
  OAI21_X1 U15629 ( .B1(n16156), .B2(n14297), .A(n14142), .ZN(P2_U3242) );
  AOI21_X1 U15630 ( .B1(n14143), .B2(n8058), .A(n14214), .ZN(n14148) );
  OAI22_X1 U15631 ( .A1(n14145), .A2(n14191), .B1(n14144), .B2(n14189), .ZN(
        n14146) );
  AOI21_X1 U15632 ( .B1(n14148), .B2(n14147), .A(n14146), .ZN(n14305) );
  NAND2_X1 U15633 ( .A1(n14150), .A2(n14149), .ZN(n14299) );
  NAND3_X1 U15634 ( .A1(n14300), .A2(n14299), .A3(n14151), .ZN(n14161) );
  OR2_X1 U15635 ( .A1(n14167), .A2(n14152), .ZN(n14153) );
  AND2_X1 U15636 ( .A1(n14154), .A2(n14153), .ZN(n14303) );
  NAND2_X1 U15637 ( .A1(n14301), .A2(n16147), .ZN(n14157) );
  AOI22_X1 U15638 ( .A1(n16156), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14155), 
        .B2(n16146), .ZN(n14156) );
  NAND2_X1 U15639 ( .A1(n14157), .A2(n14156), .ZN(n14158) );
  AOI21_X1 U15640 ( .B1(n14303), .B2(n14159), .A(n14158), .ZN(n14160) );
  OAI211_X1 U15641 ( .C1(n16156), .C2(n14305), .A(n14161), .B(n14160), .ZN(
        P2_U3243) );
  XOR2_X1 U15642 ( .A(n14163), .B(n14162), .Z(n14311) );
  XNOR2_X1 U15643 ( .A(n14164), .B(n14163), .ZN(n14166) );
  OAI21_X1 U15644 ( .B1(n14166), .B2(n14214), .A(n14165), .ZN(n14307) );
  INV_X1 U15645 ( .A(n14180), .ZN(n14168) );
  AOI211_X1 U15646 ( .C1(n14309), .C2(n14168), .A(n14319), .B(n14167), .ZN(
        n14308) );
  NAND2_X1 U15647 ( .A1(n14308), .A2(n16150), .ZN(n14171) );
  AOI22_X1 U15648 ( .A1(n16156), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14169), 
        .B2(n16146), .ZN(n14170) );
  OAI211_X1 U15649 ( .C1(n14172), .C2(n14231), .A(n14171), .B(n14170), .ZN(
        n14173) );
  AOI21_X1 U15650 ( .B1(n16041), .B2(n14307), .A(n14173), .ZN(n14174) );
  OAI21_X1 U15651 ( .B1(n14311), .B2(n14244), .A(n14174), .ZN(P2_U3244) );
  XOR2_X1 U15652 ( .A(n14177), .B(n14175), .Z(n14316) );
  XOR2_X1 U15653 ( .A(n14177), .B(n14176), .Z(n14179) );
  OAI21_X1 U15654 ( .B1(n14179), .B2(n14214), .A(n14178), .ZN(n14312) );
  INV_X1 U15655 ( .A(n14201), .ZN(n14181) );
  AOI211_X1 U15656 ( .C1(n14314), .C2(n14181), .A(n14319), .B(n14180), .ZN(
        n14313) );
  NAND2_X1 U15657 ( .A1(n14313), .A2(n16150), .ZN(n14184) );
  AOI22_X1 U15658 ( .A1(n16156), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14182), 
        .B2(n16146), .ZN(n14183) );
  OAI211_X1 U15659 ( .C1(n14185), .C2(n14231), .A(n14184), .B(n14183), .ZN(
        n14186) );
  AOI21_X1 U15660 ( .B1(n14312), .B2(n16041), .A(n14186), .ZN(n14187) );
  OAI21_X1 U15661 ( .B1(n14316), .B2(n14244), .A(n14187), .ZN(P2_U3245) );
  XOR2_X1 U15662 ( .A(n14194), .B(n14188), .Z(n14200) );
  OAI22_X1 U15663 ( .A1(n14192), .A2(n14191), .B1(n14190), .B2(n14189), .ZN(
        n14199) );
  NAND2_X1 U15664 ( .A1(n14193), .A2(n14194), .ZN(n14195) );
  NAND2_X1 U15665 ( .A1(n14196), .A2(n14195), .ZN(n14324) );
  NOR2_X1 U15666 ( .A1(n14324), .A2(n14197), .ZN(n14198) );
  AOI211_X1 U15667 ( .C1(n14200), .C2(n14236), .A(n14199), .B(n14198), .ZN(
        n14323) );
  INV_X1 U15668 ( .A(n14324), .ZN(n14208) );
  AND2_X1 U15669 ( .A1(n14317), .A2(n14216), .ZN(n14202) );
  OR2_X1 U15670 ( .A1(n14202), .A2(n14201), .ZN(n14320) );
  AOI22_X1 U15671 ( .A1(n16156), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14203), 
        .B2(n16146), .ZN(n14205) );
  NAND2_X1 U15672 ( .A1(n14317), .A2(n16147), .ZN(n14204) );
  OAI211_X1 U15673 ( .C1(n14320), .C2(n14206), .A(n14205), .B(n14204), .ZN(
        n14207) );
  AOI21_X1 U15674 ( .B1(n14208), .B2(n16151), .A(n14207), .ZN(n14209) );
  OAI21_X1 U15675 ( .B1(n14323), .B2(n16156), .A(n14209), .ZN(P2_U3246) );
  XNOR2_X1 U15676 ( .A(n14210), .B(n14211), .ZN(n14329) );
  XNOR2_X1 U15677 ( .A(n14212), .B(n14211), .ZN(n14215) );
  OAI21_X1 U15678 ( .B1(n14215), .B2(n14214), .A(n14213), .ZN(n14325) );
  INV_X1 U15679 ( .A(n14327), .ZN(n14221) );
  INV_X1 U15680 ( .A(n14216), .ZN(n14217) );
  AOI211_X1 U15681 ( .C1(n14327), .C2(n14229), .A(n14319), .B(n14217), .ZN(
        n14326) );
  NAND2_X1 U15682 ( .A1(n14326), .A2(n16150), .ZN(n14220) );
  AOI22_X1 U15683 ( .A1(n16156), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14218), 
        .B2(n16146), .ZN(n14219) );
  OAI211_X1 U15684 ( .C1(n14221), .C2(n14231), .A(n14220), .B(n14219), .ZN(
        n14222) );
  AOI21_X1 U15685 ( .B1(n16041), .B2(n14325), .A(n14222), .ZN(n14223) );
  OAI21_X1 U15686 ( .B1(n14244), .B2(n14329), .A(n14223), .ZN(P2_U3247) );
  OAI21_X1 U15687 ( .B1(n14226), .B2(n14225), .A(n14224), .ZN(n14227) );
  INV_X1 U15688 ( .A(n14227), .ZN(n14334) );
  INV_X1 U15689 ( .A(n14229), .ZN(n14230) );
  AOI211_X1 U15690 ( .C1(n14332), .C2(n7764), .A(n14319), .B(n14230), .ZN(
        n14331) );
  NOR2_X1 U15691 ( .A1(n14232), .A2(n14231), .ZN(n14235) );
  OAI22_X1 U15692 ( .A1(n16041), .A2(n12414), .B1(n14233), .B2(n16038), .ZN(
        n14234) );
  AOI211_X1 U15693 ( .C1(n14331), .C2(n16150), .A(n14235), .B(n14234), .ZN(
        n14243) );
  OAI211_X1 U15694 ( .C1(n14239), .C2(n14238), .A(n14237), .B(n14236), .ZN(
        n14241) );
  NAND2_X1 U15695 ( .A1(n14241), .A2(n14240), .ZN(n14330) );
  NAND2_X1 U15696 ( .A1(n14330), .A2(n16041), .ZN(n14242) );
  OAI211_X1 U15697 ( .C1(n14334), .C2(n14244), .A(n14243), .B(n14242), .ZN(
        P2_U3248) );
  OAI22_X1 U15698 ( .A1(n16045), .A2(n14246), .B1(n14245), .B2(n16038), .ZN(
        n14247) );
  AOI21_X1 U15699 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n16156), .A(n14247), .ZN(
        n14253) );
  AOI22_X1 U15700 ( .A1(n16151), .A2(n14249), .B1(n16147), .B2(n14248), .ZN(
        n14252) );
  NAND2_X1 U15701 ( .A1(n16041), .A2(n14250), .ZN(n14251) );
  NAND3_X1 U15702 ( .A1(n14253), .A2(n14252), .A3(n14251), .ZN(P2_U3263) );
  OAI211_X1 U15703 ( .C1(n14255), .C2(n16182), .A(n14254), .B(n14256), .ZN(
        n14347) );
  MUX2_X1 U15704 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14347), .S(n16189), .Z(
        P2_U3530) );
  OAI211_X1 U15705 ( .C1(n14258), .C2(n16182), .A(n14257), .B(n14256), .ZN(
        n14348) );
  MUX2_X1 U15706 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14348), .S(n16189), .Z(
        P2_U3529) );
  NAND2_X1 U15707 ( .A1(n14259), .A2(n16186), .ZN(n14264) );
  NAND2_X1 U15708 ( .A1(n14260), .A2(n14343), .ZN(n14262) );
  NAND2_X1 U15709 ( .A1(n14264), .A2(n8415), .ZN(n14349) );
  MUX2_X1 U15710 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14349), .S(n16189), .Z(
        P2_U3528) );
  INV_X1 U15711 ( .A(n14265), .ZN(n14270) );
  AOI21_X1 U15712 ( .B1(n14343), .B2(n14267), .A(n14266), .ZN(n14268) );
  OAI211_X1 U15713 ( .C1(n14270), .C2(n14346), .A(n14269), .B(n14268), .ZN(
        n14350) );
  MUX2_X1 U15714 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14350), .S(n16189), .Z(
        P2_U3527) );
  INV_X1 U15715 ( .A(n14271), .ZN(n14272) );
  OAI22_X1 U15716 ( .A1(n14273), .A2(n14319), .B1(n14272), .B2(n16182), .ZN(
        n14274) );
  INV_X1 U15717 ( .A(n14274), .ZN(n14275) );
  OAI211_X1 U15718 ( .C1(n15897), .C2(n14277), .A(n14276), .B(n14275), .ZN(
        n14351) );
  MUX2_X1 U15719 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14351), .S(n16189), .Z(
        P2_U3526) );
  AOI22_X1 U15720 ( .A1(n14279), .A2(n14302), .B1(n14343), .B2(n14278), .ZN(
        n14280) );
  OAI211_X1 U15721 ( .C1(n14282), .C2(n14346), .A(n14281), .B(n14280), .ZN(
        n14352) );
  MUX2_X1 U15722 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14352), .S(n16189), .Z(
        P2_U3525) );
  AOI211_X1 U15723 ( .C1(n14343), .C2(n14285), .A(n14284), .B(n14283), .ZN(
        n14286) );
  OAI21_X1 U15724 ( .B1(n14346), .B2(n14287), .A(n14286), .ZN(n14353) );
  MUX2_X1 U15725 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14353), .S(n16189), .Z(
        P2_U3524) );
  INV_X1 U15726 ( .A(n14288), .ZN(n14293) );
  AOI21_X1 U15727 ( .B1(n14343), .B2(n14290), .A(n14289), .ZN(n14291) );
  OAI211_X1 U15728 ( .C1(n15897), .C2(n14293), .A(n14292), .B(n14291), .ZN(
        n14354) );
  MUX2_X1 U15729 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14354), .S(n16189), .Z(
        P2_U3523) );
  AOI21_X1 U15730 ( .B1(n14343), .B2(n14295), .A(n14294), .ZN(n14296) );
  OAI211_X1 U15731 ( .C1(n14298), .C2(n14346), .A(n14297), .B(n14296), .ZN(
        n14355) );
  MUX2_X1 U15732 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14355), .S(n16189), .Z(
        P2_U3522) );
  NAND3_X1 U15733 ( .A1(n14300), .A2(n16186), .A3(n14299), .ZN(n14306) );
  AOI22_X1 U15734 ( .A1(n14303), .A2(n14302), .B1(n14343), .B2(n14301), .ZN(
        n14304) );
  NAND3_X1 U15735 ( .A1(n14306), .A2(n14305), .A3(n14304), .ZN(n14356) );
  MUX2_X1 U15736 ( .A(n14356), .B(P2_REG1_REG_22__SCAN_IN), .S(n16188), .Z(
        P2_U3521) );
  AOI211_X1 U15737 ( .C1(n14343), .C2(n14309), .A(n14308), .B(n14307), .ZN(
        n14310) );
  OAI21_X1 U15738 ( .B1(n14311), .B2(n14346), .A(n14310), .ZN(n14357) );
  MUX2_X1 U15739 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14357), .S(n16189), .Z(
        P2_U3520) );
  AOI211_X1 U15740 ( .C1(n14343), .C2(n14314), .A(n14313), .B(n14312), .ZN(
        n14315) );
  OAI21_X1 U15741 ( .B1(n14346), .B2(n14316), .A(n14315), .ZN(n14358) );
  MUX2_X1 U15742 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14358), .S(n16189), .Z(
        P2_U3519) );
  INV_X1 U15743 ( .A(n14317), .ZN(n14318) );
  OAI22_X1 U15744 ( .A1(n14320), .A2(n14319), .B1(n14318), .B2(n16182), .ZN(
        n14321) );
  INV_X1 U15745 ( .A(n14321), .ZN(n14322) );
  OAI211_X1 U15746 ( .C1(n15897), .C2(n14324), .A(n14323), .B(n14322), .ZN(
        n14359) );
  MUX2_X1 U15747 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14359), .S(n16189), .Z(
        P2_U3518) );
  AOI211_X1 U15748 ( .C1(n14343), .C2(n14327), .A(n14326), .B(n14325), .ZN(
        n14328) );
  OAI21_X1 U15749 ( .B1(n14346), .B2(n14329), .A(n14328), .ZN(n14360) );
  MUX2_X1 U15750 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14360), .S(n16189), .Z(
        P2_U3517) );
  AOI211_X1 U15751 ( .C1(n14343), .C2(n14332), .A(n14331), .B(n14330), .ZN(
        n14333) );
  OAI21_X1 U15752 ( .B1(n14334), .B2(n14346), .A(n14333), .ZN(n14361) );
  MUX2_X1 U15753 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14361), .S(n16189), .Z(
        P2_U3516) );
  AOI211_X1 U15754 ( .C1(n14343), .C2(n14337), .A(n14336), .B(n14335), .ZN(
        n14338) );
  OAI21_X1 U15755 ( .B1(n14339), .B2(n14346), .A(n14338), .ZN(n14362) );
  MUX2_X1 U15756 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14362), .S(n16189), .Z(
        P2_U3515) );
  AOI211_X1 U15757 ( .C1(n14343), .C2(n14342), .A(n14341), .B(n14340), .ZN(
        n14344) );
  OAI21_X1 U15758 ( .B1(n14346), .B2(n14345), .A(n14344), .ZN(n14363) );
  MUX2_X1 U15759 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14363), .S(n16189), .Z(
        P2_U3514) );
  MUX2_X1 U15760 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14347), .S(n16192), .Z(
        P2_U3498) );
  MUX2_X1 U15761 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14348), .S(n16192), .Z(
        P2_U3497) );
  MUX2_X1 U15762 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14349), .S(n16192), .Z(
        P2_U3496) );
  MUX2_X1 U15763 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14350), .S(n16192), .Z(
        P2_U3495) );
  MUX2_X1 U15764 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14351), .S(n16192), .Z(
        P2_U3494) );
  MUX2_X1 U15765 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14352), .S(n16192), .Z(
        P2_U3493) );
  MUX2_X1 U15766 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14353), .S(n16192), .Z(
        P2_U3492) );
  MUX2_X1 U15767 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14354), .S(n16192), .Z(
        P2_U3491) );
  MUX2_X1 U15768 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14355), .S(n16192), .Z(
        P2_U3490) );
  MUX2_X1 U15769 ( .A(n14356), .B(P2_REG0_REG_22__SCAN_IN), .S(n16190), .Z(
        P2_U3489) );
  MUX2_X1 U15770 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14357), .S(n16192), .Z(
        P2_U3488) );
  MUX2_X1 U15771 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14358), .S(n16192), .Z(
        P2_U3487) );
  MUX2_X1 U15772 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14359), .S(n16192), .Z(
        P2_U3486) );
  MUX2_X1 U15773 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14360), .S(n16192), .Z(
        P2_U3484) );
  MUX2_X1 U15774 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14361), .S(n16192), .Z(
        P2_U3481) );
  MUX2_X1 U15775 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14362), .S(n16192), .Z(
        P2_U3478) );
  MUX2_X1 U15776 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14363), .S(n16192), .Z(
        P2_U3475) );
  INV_X1 U15777 ( .A(n14364), .ZN(n15153) );
  INV_X1 U15778 ( .A(n14365), .ZN(n14366) );
  NOR4_X1 U15779 ( .A1(n14366), .A2(P2_IR_REG_30__SCAN_IN), .A3(n10415), .A4(
        P2_U3088), .ZN(n14367) );
  AOI21_X1 U15780 ( .B1(n14376), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14367), 
        .ZN(n14368) );
  OAI21_X1 U15781 ( .B1(n15153), .B2(n14378), .A(n14368), .ZN(P2_U3296) );
  INV_X1 U15782 ( .A(n14369), .ZN(n15155) );
  OAI222_X1 U15783 ( .A1(n14378), .A2(n15155), .B1(P2_U3088), .B2(n14372), 
        .C1(n14371), .C2(n14370), .ZN(P2_U3298) );
  INV_X1 U15784 ( .A(n14374), .ZN(n15159) );
  AOI21_X1 U15785 ( .B1(n14376), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14375), 
        .ZN(n14377) );
  OAI21_X1 U15786 ( .B1(n15159), .B2(n14378), .A(n14377), .ZN(P2_U3299) );
  INV_X1 U15787 ( .A(n14379), .ZN(n14380) );
  MUX2_X1 U15788 ( .A(n14380), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OR2_X1 U15789 ( .A1(n14383), .A2(n14588), .ZN(n14382) );
  NAND2_X1 U15790 ( .A1(n14480), .A2(n14745), .ZN(n14381) );
  NAND2_X1 U15791 ( .A1(n14382), .A2(n14381), .ZN(n14581) );
  OAI22_X1 U15792 ( .A1(n14383), .A2(n14585), .B1(n14595), .B2(n14588), .ZN(
        n14384) );
  XNOR2_X1 U15793 ( .A(n14384), .B(n14589), .ZN(n14580) );
  XOR2_X1 U15794 ( .A(n14581), .B(n14580), .Z(n14584) );
  NOR2_X1 U15795 ( .A1(n14586), .A2(n14385), .ZN(n14386) );
  AOI21_X1 U15796 ( .B1(n14387), .B2(n14533), .A(n14386), .ZN(n14410) );
  INV_X1 U15797 ( .A(n14410), .ZN(n14413) );
  NAND2_X1 U15798 ( .A1(n14387), .A2(n14526), .ZN(n14389) );
  NAND2_X1 U15799 ( .A1(n14533), .A2(n14758), .ZN(n14388) );
  NAND2_X1 U15800 ( .A1(n14389), .A2(n14388), .ZN(n14390) );
  XNOR2_X1 U15801 ( .A(n14390), .B(n14529), .ZN(n14411) );
  INV_X1 U15802 ( .A(n14411), .ZN(n14412) );
  NAND2_X1 U15803 ( .A1(n14661), .A2(n14526), .ZN(n14395) );
  NAND2_X1 U15804 ( .A1(n11917), .A2(n14761), .ZN(n14394) );
  NAND2_X1 U15805 ( .A1(n14395), .A2(n14394), .ZN(n14396) );
  XNOR2_X1 U15806 ( .A(n14396), .B(n14529), .ZN(n14653) );
  NOR2_X1 U15807 ( .A1(n14586), .A2(n14397), .ZN(n14398) );
  AOI21_X1 U15808 ( .B1(n14661), .B2(n14533), .A(n14398), .ZN(n14399) );
  NAND2_X1 U15809 ( .A1(n14653), .A2(n14399), .ZN(n14401) );
  INV_X1 U15810 ( .A(n14653), .ZN(n14400) );
  INV_X1 U15811 ( .A(n14399), .ZN(n14652) );
  AOI22_X1 U15812 ( .A1(n14560), .A2(n14526), .B1(n14533), .B2(n14760), .ZN(
        n14402) );
  XNOR2_X1 U15813 ( .A(n14402), .B(n14589), .ZN(n14404) );
  NOR2_X1 U15814 ( .A1(n14586), .A2(n14696), .ZN(n14403) );
  AOI21_X1 U15815 ( .B1(n14560), .B2(n14533), .A(n14403), .ZN(n14405) );
  XNOR2_X1 U15816 ( .A(n14404), .B(n14405), .ZN(n14554) );
  OAI22_X1 U15817 ( .A1(n14407), .A2(n14585), .B1(n14615), .B2(n14588), .ZN(
        n14406) );
  XNOR2_X1 U15818 ( .A(n14406), .B(n14589), .ZN(n14409) );
  OAI22_X1 U15819 ( .A1(n14407), .A2(n14588), .B1(n14615), .B2(n14586), .ZN(
        n14408) );
  XNOR2_X1 U15820 ( .A(n14409), .B(n14408), .ZN(n14695) );
  NOR2_X1 U15821 ( .A1(n14409), .A2(n14408), .ZN(n14611) );
  XNOR2_X1 U15822 ( .A(n14411), .B(n14410), .ZN(n14610) );
  AOI22_X1 U15823 ( .A1(n14679), .A2(n14533), .B1(n14480), .B2(n14757), .ZN(
        n14418) );
  NAND2_X1 U15824 ( .A1(n14679), .A2(n14526), .ZN(n14415) );
  NAND2_X1 U15825 ( .A1(n11917), .A2(n14757), .ZN(n14414) );
  NAND2_X1 U15826 ( .A1(n14415), .A2(n14414), .ZN(n14416) );
  XNOR2_X1 U15827 ( .A(n14416), .B(n14589), .ZN(n14417) );
  XOR2_X1 U15828 ( .A(n14418), .B(n14417), .Z(n14672) );
  NAND2_X1 U15829 ( .A1(n16177), .A2(n14526), .ZN(n14420) );
  NAND2_X1 U15830 ( .A1(n11917), .A2(n14756), .ZN(n14419) );
  NAND2_X1 U15831 ( .A1(n14420), .A2(n14419), .ZN(n14421) );
  XNOR2_X1 U15832 ( .A(n14421), .B(n14529), .ZN(n14425) );
  NOR2_X1 U15833 ( .A1(n14586), .A2(n14422), .ZN(n14423) );
  AOI21_X1 U15834 ( .B1(n16177), .B2(n14533), .A(n14423), .ZN(n14424) );
  NAND2_X1 U15835 ( .A1(n14425), .A2(n14424), .ZN(n14426) );
  OAI21_X1 U15836 ( .B1(n14425), .B2(n14424), .A(n14426), .ZN(n16173) );
  NAND2_X1 U15837 ( .A1(n14738), .A2(n14526), .ZN(n14428) );
  NAND2_X1 U15838 ( .A1(n11917), .A2(n14755), .ZN(n14427) );
  NAND2_X1 U15839 ( .A1(n14428), .A2(n14427), .ZN(n14429) );
  XNOR2_X1 U15840 ( .A(n14429), .B(n14589), .ZN(n14434) );
  OAI22_X1 U15842 ( .A1(n14431), .A2(n14588), .B1(n14430), .B2(n14586), .ZN(
        n14731) );
  INV_X1 U15843 ( .A(n14432), .ZN(n14433) );
  NAND2_X1 U15844 ( .A1(n16199), .A2(n14526), .ZN(n14436) );
  NAND2_X1 U15845 ( .A1(n11917), .A2(n14754), .ZN(n14435) );
  NAND2_X1 U15846 ( .A1(n14436), .A2(n14435), .ZN(n14437) );
  XNOR2_X1 U15847 ( .A(n14437), .B(n14529), .ZN(n14441) );
  INV_X1 U15848 ( .A(n14441), .ZN(n14443) );
  NOR2_X1 U15849 ( .A1(n14586), .A2(n14438), .ZN(n14439) );
  AOI21_X1 U15850 ( .B1(n16199), .B2(n14533), .A(n14439), .ZN(n14440) );
  INV_X1 U15851 ( .A(n14440), .ZN(n14442) );
  AND2_X1 U15852 ( .A1(n14441), .A2(n14440), .ZN(n14444) );
  AOI21_X1 U15853 ( .B1(n14443), .B2(n14442), .A(n14444), .ZN(n16194) );
  INV_X1 U15854 ( .A(n14444), .ZN(n14634) );
  NAND2_X1 U15855 ( .A1(n14449), .A2(n14526), .ZN(n14446) );
  NAND2_X1 U15856 ( .A1(n14753), .A2(n14533), .ZN(n14445) );
  NAND2_X1 U15857 ( .A1(n14446), .A2(n14445), .ZN(n14447) );
  XNOR2_X1 U15858 ( .A(n14447), .B(n14529), .ZN(n14450) );
  NOR2_X1 U15859 ( .A1(n14586), .A2(n15013), .ZN(n14448) );
  AOI21_X1 U15860 ( .B1(n14449), .B2(n14533), .A(n14448), .ZN(n14451) );
  NAND2_X1 U15861 ( .A1(n14450), .A2(n14451), .ZN(n14455) );
  INV_X1 U15862 ( .A(n14450), .ZN(n14453) );
  INV_X1 U15863 ( .A(n14451), .ZN(n14452) );
  NAND2_X1 U15864 ( .A1(n14453), .A2(n14452), .ZN(n14454) );
  NAND2_X1 U15865 ( .A1(n14455), .A2(n14454), .ZN(n14633) );
  INV_X1 U15866 ( .A(n14455), .ZN(n14708) );
  NAND2_X1 U15867 ( .A1(n15025), .A2(n14526), .ZN(n14457) );
  NAND2_X1 U15868 ( .A1(n14752), .A2(n14533), .ZN(n14456) );
  NAND2_X1 U15869 ( .A1(n14457), .A2(n14456), .ZN(n14458) );
  XNOR2_X1 U15870 ( .A(n14458), .B(n14529), .ZN(n14460) );
  AND2_X1 U15871 ( .A1(n14480), .A2(n14752), .ZN(n14459) );
  AOI21_X1 U15872 ( .B1(n15025), .B2(n14533), .A(n14459), .ZN(n14461) );
  NAND2_X1 U15873 ( .A1(n14460), .A2(n14461), .ZN(n14465) );
  INV_X1 U15874 ( .A(n14460), .ZN(n14463) );
  INV_X1 U15875 ( .A(n14461), .ZN(n14462) );
  NAND2_X1 U15876 ( .A1(n14463), .A2(n14462), .ZN(n14464) );
  AND2_X1 U15877 ( .A1(n14465), .A2(n14464), .ZN(n14707) );
  NAND2_X1 U15878 ( .A1(n15105), .A2(n14526), .ZN(n14467) );
  NAND2_X1 U15879 ( .A1(n14751), .A2(n14533), .ZN(n14466) );
  NAND2_X1 U15880 ( .A1(n14467), .A2(n14466), .ZN(n14468) );
  XNOR2_X1 U15881 ( .A(n14468), .B(n14589), .ZN(n14469) );
  AOI22_X1 U15882 ( .A1(n15105), .A2(n14533), .B1(n14480), .B2(n14751), .ZN(
        n14470) );
  XNOR2_X1 U15883 ( .A(n14469), .B(n14470), .ZN(n14573) );
  INV_X1 U15884 ( .A(n14469), .ZN(n14471) );
  NAND2_X1 U15885 ( .A1(n14471), .A2(n14470), .ZN(n14665) );
  NAND2_X1 U15886 ( .A1(n15099), .A2(n14526), .ZN(n14473) );
  NAND2_X1 U15887 ( .A1(n14750), .A2(n14533), .ZN(n14472) );
  NAND2_X1 U15888 ( .A1(n14473), .A2(n14472), .ZN(n14474) );
  XNOR2_X1 U15889 ( .A(n14474), .B(n14589), .ZN(n14484) );
  AND2_X1 U15890 ( .A1(n14750), .A2(n14480), .ZN(n14475) );
  AOI21_X1 U15891 ( .B1(n15099), .B2(n14533), .A(n14475), .ZN(n14482) );
  XNOR2_X1 U15892 ( .A(n14484), .B(n14482), .ZN(n14664) );
  NAND2_X1 U15893 ( .A1(n15086), .A2(n14526), .ZN(n14478) );
  NAND2_X1 U15894 ( .A1(n14749), .A2(n14533), .ZN(n14477) );
  NAND2_X1 U15895 ( .A1(n14478), .A2(n14477), .ZN(n14479) );
  XNOR2_X1 U15896 ( .A(n14479), .B(n14589), .ZN(n14488) );
  AND2_X1 U15897 ( .A1(n14749), .A2(n14480), .ZN(n14481) );
  AOI21_X1 U15898 ( .B1(n15086), .B2(n14533), .A(n14481), .ZN(n14486) );
  XNOR2_X1 U15899 ( .A(n14488), .B(n14486), .ZN(n14602) );
  INV_X1 U15900 ( .A(n14482), .ZN(n14483) );
  NAND2_X1 U15901 ( .A1(n14484), .A2(n14483), .ZN(n14603) );
  INV_X1 U15902 ( .A(n14486), .ZN(n14487) );
  NOR2_X1 U15903 ( .A1(n14586), .A2(n14490), .ZN(n14491) );
  AOI21_X1 U15904 ( .B1(n15077), .B2(n14533), .A(n14491), .ZN(n14501) );
  NAND2_X1 U15905 ( .A1(n15077), .A2(n14526), .ZN(n14493) );
  NAND2_X1 U15906 ( .A1(n11917), .A2(n14748), .ZN(n14492) );
  NAND2_X1 U15907 ( .A1(n14493), .A2(n14492), .ZN(n14494) );
  XNOR2_X1 U15908 ( .A(n14494), .B(n14589), .ZN(n14503) );
  XOR2_X1 U15909 ( .A(n14501), .B(n14503), .Z(n14684) );
  NAND2_X1 U15910 ( .A1(n15073), .A2(n14526), .ZN(n14496) );
  NAND2_X1 U15911 ( .A1(n11917), .A2(n14912), .ZN(n14495) );
  NAND2_X1 U15912 ( .A1(n14496), .A2(n14495), .ZN(n14497) );
  XNOR2_X1 U15913 ( .A(n14497), .B(n14529), .ZN(n14500) );
  NOR2_X1 U15914 ( .A1(n14586), .A2(n14686), .ZN(n14498) );
  AOI21_X1 U15915 ( .B1(n15073), .B2(n14533), .A(n14498), .ZN(n14499) );
  NAND2_X1 U15916 ( .A1(n14500), .A2(n14499), .ZN(n14646) );
  OAI21_X1 U15917 ( .B1(n14500), .B2(n14499), .A(n14646), .ZN(n14547) );
  INV_X1 U15918 ( .A(n14501), .ZN(n14502) );
  AND2_X1 U15919 ( .A1(n14503), .A2(n14502), .ZN(n14548) );
  NOR2_X1 U15920 ( .A1(n14547), .A2(n14548), .ZN(n14504) );
  NAND2_X1 U15921 ( .A1(n15063), .A2(n14526), .ZN(n14506) );
  NAND2_X1 U15922 ( .A1(n11917), .A2(n14747), .ZN(n14505) );
  NAND2_X1 U15923 ( .A1(n14506), .A2(n14505), .ZN(n14507) );
  XNOR2_X1 U15924 ( .A(n14507), .B(n14529), .ZN(n14510) );
  NOR2_X1 U15925 ( .A1(n14586), .A2(n14508), .ZN(n14509) );
  AOI21_X1 U15926 ( .B1(n15063), .B2(n14533), .A(n14509), .ZN(n14511) );
  NAND2_X1 U15927 ( .A1(n14510), .A2(n14511), .ZN(n14515) );
  INV_X1 U15928 ( .A(n14510), .ZN(n14513) );
  INV_X1 U15929 ( .A(n14511), .ZN(n14512) );
  NAND2_X1 U15930 ( .A1(n14513), .A2(n14512), .ZN(n14514) );
  AND2_X1 U15931 ( .A1(n14515), .A2(n14514), .ZN(n14644) );
  OAI22_X1 U15932 ( .A1(n14517), .A2(n14588), .B1(n14516), .B2(n14586), .ZN(
        n14522) );
  NAND2_X1 U15933 ( .A1(n15055), .A2(n14526), .ZN(n14519) );
  NAND2_X1 U15934 ( .A1(n14533), .A2(n14913), .ZN(n14518) );
  NAND2_X1 U15935 ( .A1(n14519), .A2(n14518), .ZN(n14520) );
  XNOR2_X1 U15936 ( .A(n14520), .B(n14589), .ZN(n14521) );
  XOR2_X1 U15937 ( .A(n14522), .B(n14521), .Z(n14623) );
  NAND2_X1 U15938 ( .A1(n14622), .A2(n14623), .ZN(n14621) );
  INV_X1 U15939 ( .A(n14521), .ZN(n14524) );
  INV_X1 U15940 ( .A(n14522), .ZN(n14523) );
  NAND2_X1 U15941 ( .A1(n14524), .A2(n14523), .ZN(n14525) );
  NAND2_X1 U15942 ( .A1(n15047), .A2(n14526), .ZN(n14528) );
  NAND2_X1 U15943 ( .A1(n11917), .A2(n14746), .ZN(n14527) );
  NAND2_X1 U15944 ( .A1(n14528), .A2(n14527), .ZN(n14530) );
  XNOR2_X1 U15945 ( .A(n14530), .B(n14529), .ZN(n14535) );
  NOR2_X1 U15946 ( .A1(n14586), .A2(n14531), .ZN(n14532) );
  AOI21_X1 U15947 ( .B1(n15047), .B2(n14533), .A(n14532), .ZN(n14534) );
  OR2_X1 U15948 ( .A1(n14535), .A2(n14534), .ZN(n14720) );
  NAND2_X1 U15949 ( .A1(n14535), .A2(n14534), .ZN(n14723) );
  NOR2_X1 U15950 ( .A1(n16203), .A2(n14536), .ZN(n14540) );
  AOI22_X1 U15951 ( .A1(n14714), .A2(n14746), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14537) );
  OAI21_X1 U15952 ( .B1(n14587), .B2(n14538), .A(n14537), .ZN(n14539) );
  AOI211_X1 U15953 ( .C1(n15042), .C2(n7185), .A(n14540), .B(n14539), .ZN(
        n14541) );
  OAI21_X1 U15954 ( .B1(n14542), .B2(n14740), .A(n14541), .ZN(P1_U3214) );
  NAND2_X1 U15955 ( .A1(n14914), .A2(n14747), .ZN(n14544) );
  NAND2_X1 U15956 ( .A1(n15925), .A2(n14748), .ZN(n14543) );
  NAND2_X1 U15957 ( .A1(n14544), .A2(n14543), .ZN(n15072) );
  AOI22_X1 U15958 ( .A1(n16197), .A2(n15072), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14545) );
  OAI21_X1 U15959 ( .B1(n14935), .B2(n16203), .A(n14545), .ZN(n14552) );
  INV_X1 U15960 ( .A(n14546), .ZN(n14682) );
  OAI21_X1 U15961 ( .B1(n14682), .B2(n14548), .A(n14547), .ZN(n14550) );
  AOI21_X1 U15962 ( .B1(n14550), .B2(n14549), .A(n14740), .ZN(n14551) );
  AOI211_X1 U15963 ( .C1(n15073), .C2(n7185), .A(n14552), .B(n14551), .ZN(
        n14553) );
  INV_X1 U15964 ( .A(n14553), .ZN(P1_U3216) );
  XNOR2_X1 U15965 ( .A(n14555), .B(n14554), .ZN(n14562) );
  AOI22_X1 U15966 ( .A1(n16197), .A2(n14556), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14557) );
  OAI21_X1 U15967 ( .B1(n14558), .B2(n16203), .A(n14557), .ZN(n14559) );
  AOI21_X1 U15968 ( .B1(n14560), .B2(n7185), .A(n14559), .ZN(n14561) );
  OAI21_X1 U15969 ( .B1(n14562), .B2(n14740), .A(n14561), .ZN(P1_U3217) );
  OAI211_X1 U15970 ( .C1(n14565), .C2(n14564), .A(n14563), .B(n16195), .ZN(
        n14570) );
  AOI22_X1 U15971 ( .A1(n7185), .A2(n14566), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n14569) );
  AOI22_X1 U15972 ( .A1(n14699), .A2(n14766), .B1(n14714), .B2(n14768), .ZN(
        n14568) );
  INV_X1 U15973 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14783) );
  NAND2_X1 U15974 ( .A1(n14690), .A2(n14783), .ZN(n14567) );
  NAND4_X1 U15975 ( .A1(n14570), .A2(n14569), .A3(n14568), .A4(n14567), .ZN(
        P1_U3218) );
  OAI21_X1 U15976 ( .B1(n14573), .B2(n14572), .A(n14571), .ZN(n14574) );
  NAND2_X1 U15977 ( .A1(n14574), .A2(n16195), .ZN(n14579) );
  INV_X1 U15978 ( .A(n14575), .ZN(n14994) );
  AND2_X1 U15979 ( .A1(n14752), .A2(n15925), .ZN(n14576) );
  AOI21_X1 U15980 ( .B1(n14750), .B2(n14914), .A(n14576), .ZN(n15103) );
  NAND2_X1 U15981 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14837)
         );
  OAI21_X1 U15982 ( .B1(n15103), .B2(n14711), .A(n14837), .ZN(n14577) );
  AOI21_X1 U15983 ( .B1(n14994), .B2(n14690), .A(n14577), .ZN(n14578) );
  OAI211_X1 U15984 ( .C1(n8878), .C2(n14717), .A(n14579), .B(n14578), .ZN(
        P1_U3219) );
  INV_X1 U15985 ( .A(n14580), .ZN(n14583) );
  INV_X1 U15986 ( .A(n14581), .ZN(n14582) );
  OAI22_X1 U15987 ( .A1(n15036), .A2(n14585), .B1(n14587), .B2(n14588), .ZN(
        n14592) );
  OAI22_X1 U15988 ( .A1(n15036), .A2(n14588), .B1(n14587), .B2(n14586), .ZN(
        n14590) );
  XNOR2_X1 U15989 ( .A(n14590), .B(n14589), .ZN(n14591) );
  XOR2_X1 U15990 ( .A(n14592), .B(n14591), .Z(n14593) );
  OAI22_X1 U15991 ( .A1(n15012), .A2(n14595), .B1(n14594), .B2(n15916), .ZN(
        n14869) );
  AOI22_X1 U15992 ( .A1(n16197), .A2(n14869), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14596) );
  OAI21_X1 U15993 ( .B1(n14876), .B2(n16203), .A(n14596), .ZN(n14597) );
  AOI21_X1 U15994 ( .B1(n14878), .B2(n7185), .A(n14597), .ZN(n14598) );
  OAI21_X1 U15995 ( .B1(n14599), .B2(n14740), .A(n14598), .ZN(P1_U3220) );
  INV_X1 U15996 ( .A(n14600), .ZN(n14605) );
  AOI21_X1 U15997 ( .B1(n14601), .B2(n14603), .A(n14602), .ZN(n14604) );
  OAI21_X1 U15998 ( .B1(n14605), .B2(n14604), .A(n16195), .ZN(n14609) );
  AOI22_X1 U15999 ( .A1(n14750), .A2(n15925), .B1(n14914), .B2(n14748), .ZN(
        n15088) );
  INV_X1 U16000 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14606) );
  OAI22_X1 U16001 ( .A1(n15088), .A2(n14711), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14606), .ZN(n14607) );
  AOI21_X1 U16002 ( .B1(n14965), .B2(n14690), .A(n14607), .ZN(n14608) );
  OAI211_X1 U16003 ( .C1(n14967), .C2(n14717), .A(n14609), .B(n14608), .ZN(
        P1_U3223) );
  OAI21_X1 U16004 ( .B1(n14693), .B2(n14611), .A(n14610), .ZN(n14612) );
  NAND3_X1 U16005 ( .A1(n7384), .A2(n16195), .A3(n14612), .ZN(n14619) );
  NOR2_X1 U16006 ( .A1(n16203), .A2(n14613), .ZN(n14617) );
  OAI21_X1 U16007 ( .B1(n14697), .B2(n14615), .A(n14614), .ZN(n14616) );
  AOI211_X1 U16008 ( .C1(n14699), .C2(n14757), .A(n14617), .B(n14616), .ZN(
        n14618) );
  OAI211_X1 U16009 ( .C1(n14620), .C2(n14717), .A(n14619), .B(n14618), .ZN(
        P1_U3224) );
  OAI21_X1 U16010 ( .B1(n14623), .B2(n14622), .A(n14621), .ZN(n14624) );
  INV_X1 U16011 ( .A(n14624), .ZN(n14630) );
  NAND2_X1 U16012 ( .A1(n14914), .A2(n14746), .ZN(n14626) );
  NAND2_X1 U16013 ( .A1(n15925), .A2(n14747), .ZN(n14625) );
  NAND2_X1 U16014 ( .A1(n14626), .A2(n14625), .ZN(n15054) );
  AOI22_X1 U16015 ( .A1(n16197), .A2(n15054), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14627) );
  OAI21_X1 U16016 ( .B1(n14904), .B2(n16203), .A(n14627), .ZN(n14628) );
  AOI21_X1 U16017 ( .B1(n15055), .B2(n7185), .A(n14628), .ZN(n14629) );
  OAI21_X1 U16018 ( .B1(n14630), .B2(n14740), .A(n14629), .ZN(P1_U3225) );
  AND3_X1 U16019 ( .A1(n14632), .A2(n14634), .A3(n14633), .ZN(n14635) );
  OAI21_X1 U16020 ( .B1(n14631), .B2(n14635), .A(n16195), .ZN(n14641) );
  NOR2_X1 U16021 ( .A1(n16203), .A2(n14636), .ZN(n14637) );
  AOI211_X1 U16022 ( .C1(n16197), .C2(n14639), .A(n14638), .B(n14637), .ZN(
        n14640) );
  OAI211_X1 U16023 ( .C1(n15121), .C2(n14717), .A(n14641), .B(n14640), .ZN(
        P1_U3228) );
  AOI22_X1 U16024 ( .A1(n14714), .A2(n14912), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14643) );
  NAND2_X1 U16025 ( .A1(n14699), .A2(n14913), .ZN(n14642) );
  OAI211_X1 U16026 ( .C1(n16203), .C2(n14923), .A(n14643), .B(n14642), .ZN(
        n14650) );
  INV_X1 U16027 ( .A(n14644), .ZN(n14645) );
  NAND3_X1 U16028 ( .A1(n14549), .A2(n14646), .A3(n14645), .ZN(n14647) );
  AOI21_X1 U16029 ( .B1(n14648), .B2(n14647), .A(n14740), .ZN(n14649) );
  AOI211_X1 U16030 ( .C1(n15063), .C2(n7185), .A(n14650), .B(n14649), .ZN(
        n14651) );
  INV_X1 U16031 ( .A(n14651), .ZN(P1_U3229) );
  XNOR2_X1 U16032 ( .A(n14653), .B(n14652), .ZN(n14654) );
  XNOR2_X1 U16033 ( .A(n7342), .B(n14654), .ZN(n14663) );
  OAI21_X1 U16034 ( .B1(n14697), .B2(n14656), .A(n14655), .ZN(n14657) );
  AOI21_X1 U16035 ( .B1(n14699), .B2(n14760), .A(n14657), .ZN(n14658) );
  OAI21_X1 U16036 ( .B1(n14659), .B2(n16203), .A(n14658), .ZN(n14660) );
  AOI21_X1 U16037 ( .B1(n14661), .B2(n7185), .A(n14660), .ZN(n14662) );
  OAI21_X1 U16038 ( .B1(n14663), .B2(n14740), .A(n14662), .ZN(P1_U3231) );
  NAND2_X1 U16039 ( .A1(n14601), .A2(n16195), .ZN(n14671) );
  AOI21_X1 U16040 ( .B1(n14571), .B2(n14665), .A(n14664), .ZN(n14670) );
  OAI22_X1 U16041 ( .A1(n14666), .A2(n15916), .B1(n8877), .B2(n15012), .ZN(
        n15098) );
  AOI22_X1 U16042 ( .A1(n15098), .A2(n16197), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14667) );
  OAI21_X1 U16043 ( .B1(n14980), .B2(n16203), .A(n14667), .ZN(n14668) );
  AOI21_X1 U16044 ( .B1(n15099), .B2(n7185), .A(n14668), .ZN(n14669) );
  OAI21_X1 U16045 ( .B1(n14671), .B2(n14670), .A(n14669), .ZN(P1_U3233) );
  XNOR2_X1 U16046 ( .A(n14673), .B(n14672), .ZN(n14681) );
  NAND2_X1 U16047 ( .A1(n16197), .A2(n14674), .ZN(n14675) );
  OAI211_X1 U16048 ( .C1(n16203), .C2(n14677), .A(n14676), .B(n14675), .ZN(
        n14678) );
  AOI21_X1 U16049 ( .B1(n14679), .B2(n7185), .A(n14678), .ZN(n14680) );
  OAI21_X1 U16050 ( .B1(n14681), .B2(n14740), .A(n14680), .ZN(P1_U3234) );
  AOI211_X1 U16051 ( .C1(n14684), .C2(n14683), .A(n14740), .B(n14682), .ZN(
        n14685) );
  INV_X1 U16052 ( .A(n14685), .ZN(n14692) );
  NOR2_X1 U16053 ( .A1(n15916), .A2(n14686), .ZN(n14687) );
  AOI21_X1 U16054 ( .B1(n14749), .B2(n15925), .A(n14687), .ZN(n15078) );
  OAI22_X1 U16055 ( .A1(n15078), .A2(n14711), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14688), .ZN(n14689) );
  AOI21_X1 U16056 ( .B1(n14948), .B2(n14690), .A(n14689), .ZN(n14691) );
  OAI211_X1 U16057 ( .C1(n14717), .C2(n14952), .A(n14692), .B(n14691), .ZN(
        P1_U3235) );
  AOI21_X1 U16058 ( .B1(n14695), .B2(n14694), .A(n14693), .ZN(n14705) );
  NAND2_X1 U16059 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14797)
         );
  OAI21_X1 U16060 ( .B1(n14697), .B2(n14696), .A(n14797), .ZN(n14698) );
  AOI21_X1 U16061 ( .B1(n14699), .B2(n14758), .A(n14698), .ZN(n14700) );
  OAI21_X1 U16062 ( .B1(n14701), .B2(n16203), .A(n14700), .ZN(n14702) );
  AOI21_X1 U16063 ( .B1(n14703), .B2(n7185), .A(n14702), .ZN(n14704) );
  OAI21_X1 U16064 ( .B1(n14705), .B2(n14740), .A(n14704), .ZN(P1_U3236) );
  INV_X1 U16065 ( .A(n14706), .ZN(n14710) );
  NOR3_X1 U16066 ( .A1(n14631), .A2(n14708), .A3(n14707), .ZN(n14709) );
  OAI21_X1 U16067 ( .B1(n14710), .B2(n14709), .A(n16195), .ZN(n14716) );
  NOR2_X1 U16068 ( .A1(n16203), .A2(n15019), .ZN(n14713) );
  NAND2_X1 U16069 ( .A1(n14751), .A2(n14914), .ZN(n15011) );
  NAND2_X1 U16070 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14818)
         );
  OAI21_X1 U16071 ( .B1(n14711), .B2(n15011), .A(n14818), .ZN(n14712) );
  AOI211_X1 U16072 ( .C1(n14714), .C2(n14753), .A(n14713), .B(n14712), .ZN(
        n14715) );
  OAI211_X1 U16073 ( .C1(n8857), .C2(n14717), .A(n14716), .B(n14715), .ZN(
        P1_U3238) );
  INV_X1 U16074 ( .A(n14718), .ZN(n14724) );
  INV_X1 U16075 ( .A(n14719), .ZN(n14722) );
  NAND2_X1 U16076 ( .A1(n14720), .A2(n14723), .ZN(n14721) );
  AOI22_X1 U16077 ( .A1(n14724), .A2(n14723), .B1(n14722), .B2(n14721), .ZN(
        n14730) );
  NAND2_X1 U16078 ( .A1(n14914), .A2(n14745), .ZN(n14726) );
  NAND2_X1 U16079 ( .A1(n15925), .A2(n14913), .ZN(n14725) );
  NAND2_X1 U16080 ( .A1(n14726), .A2(n14725), .ZN(n15046) );
  AOI22_X1 U16081 ( .A1(n16197), .A2(n15046), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14727) );
  OAI21_X1 U16082 ( .B1(n14888), .B2(n16203), .A(n14727), .ZN(n14728) );
  AOI21_X1 U16083 ( .B1(n15047), .B2(n7185), .A(n14728), .ZN(n14729) );
  OAI21_X1 U16084 ( .B1(n14730), .B2(n14740), .A(n14729), .ZN(P1_U3240) );
  XNOR2_X1 U16085 ( .A(n14732), .B(n14731), .ZN(n14741) );
  NAND2_X1 U16086 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15541)
         );
  NAND2_X1 U16087 ( .A1(n16197), .A2(n14733), .ZN(n14734) );
  OAI211_X1 U16088 ( .C1(n16203), .C2(n14735), .A(n15541), .B(n14734), .ZN(
        n14736) );
  AOI21_X1 U16089 ( .B1(n14738), .B2(n7185), .A(n14736), .ZN(n14739) );
  OAI21_X1 U16090 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(P1_U3241) );
  MUX2_X1 U16091 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14840), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16092 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14742), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16093 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14743), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16094 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14744), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16095 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14745), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16096 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14746), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16097 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14913), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16098 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14747), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16099 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14912), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16100 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14748), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16101 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14749), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16102 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14750), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16103 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14751), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16104 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14752), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16105 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14753), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16106 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14754), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16107 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14755), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16108 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14756), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16109 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14757), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16110 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14758), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16111 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14759), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16112 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14760), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16113 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14761), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16114 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14762), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16115 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14763), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16116 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14764), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16117 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14765), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16118 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14766), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16119 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14767), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16120 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14768), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16121 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14769), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16122 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15924), .S(P1_U4016), .Z(
        P1_U3560) );
  AND2_X1 U16123 ( .A1(n15398), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n14771) );
  OAI211_X1 U16124 ( .C1(n14772), .C2(n14771), .A(n15539), .B(n14770), .ZN(
        n14780) );
  AOI22_X1 U16125 ( .A1(n15526), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14779) );
  NAND2_X1 U16126 ( .A1(n15862), .A2(n14773), .ZN(n14778) );
  OAI211_X1 U16127 ( .C1(n14776), .C2(n14775), .A(n15869), .B(n14774), .ZN(
        n14777) );
  NAND4_X1 U16128 ( .A1(n14780), .A2(n14779), .A3(n14778), .A4(n14777), .ZN(
        P1_U3244) );
  OAI211_X1 U16129 ( .C1(n14782), .C2(n14781), .A(n15539), .B(n15856), .ZN(
        n14792) );
  NOR2_X1 U16130 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14783), .ZN(n14784) );
  AOI21_X1 U16131 ( .B1(n15526), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14784), .ZN(
        n14791) );
  NAND2_X1 U16132 ( .A1(n15862), .A2(n15393), .ZN(n14790) );
  MUX2_X1 U16133 ( .A(n11152), .B(P1_REG2_REG_3__SCAN_IN), .S(n15393), .Z(
        n14787) );
  NAND3_X1 U16134 ( .A1(n14787), .A2(n14786), .A3(n14785), .ZN(n14788) );
  NAND3_X1 U16135 ( .A1(n15869), .A2(n15865), .A3(n14788), .ZN(n14789) );
  NAND4_X1 U16136 ( .A1(n14792), .A2(n14791), .A3(n14790), .A4(n14789), .ZN(
        P1_U3246) );
  OAI21_X1 U16137 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(n14796) );
  NAND2_X1 U16138 ( .A1(n14796), .A2(n15539), .ZN(n14809) );
  INV_X1 U16139 ( .A(n14797), .ZN(n14798) );
  AOI21_X1 U16140 ( .B1(n15526), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n14798), 
        .ZN(n14808) );
  INV_X1 U16141 ( .A(n14799), .ZN(n14804) );
  NAND3_X1 U16142 ( .A1(n14802), .A2(n14801), .A3(n14800), .ZN(n14803) );
  NAND3_X1 U16143 ( .A1(n15869), .A2(n14804), .A3(n14803), .ZN(n14807) );
  NAND2_X1 U16144 ( .A1(n15862), .A2(n14805), .ZN(n14806) );
  NAND4_X1 U16145 ( .A1(n14809), .A2(n14808), .A3(n14807), .A4(n14806), .ZN(
        P1_U3254) );
  OAI21_X1 U16146 ( .B1(n14812), .B2(n14811), .A(n14810), .ZN(n14827) );
  XNOR2_X1 U16147 ( .A(n14827), .B(n14826), .ZN(n14828) );
  XNOR2_X1 U16148 ( .A(n14828), .B(n15020), .ZN(n14822) );
  AND2_X1 U16149 ( .A1(n14817), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14824) );
  INV_X1 U16150 ( .A(n14824), .ZN(n14816) );
  OAI211_X1 U16151 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14817), .A(n14816), 
        .B(n15539), .ZN(n14821) );
  OAI21_X1 U16152 ( .B1(n15876), .B2(n10398), .A(n14818), .ZN(n14819) );
  AOI21_X1 U16153 ( .B1(n14826), .B2(n15862), .A(n14819), .ZN(n14820) );
  OAI211_X1 U16154 ( .C1(n14822), .C2(n15536), .A(n14821), .B(n14820), .ZN(
        P1_U3261) );
  NOR2_X1 U16155 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  XNOR2_X1 U16156 ( .A(n14825), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14833) );
  NAND2_X1 U16157 ( .A1(n14827), .A2(n14826), .ZN(n14830) );
  OR2_X1 U16158 ( .A1(n14828), .A2(n15020), .ZN(n14829) );
  NAND2_X1 U16159 ( .A1(n14830), .A2(n14829), .ZN(n14831) );
  XOR2_X1 U16160 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14831), .Z(n14832) );
  AOI22_X1 U16161 ( .A1(n14833), .A2(n15539), .B1(n15869), .B2(n14832), .ZN(
        n14836) );
  INV_X1 U16162 ( .A(n14832), .ZN(n14834) );
  NAND2_X1 U16163 ( .A1(n14845), .A2(n15035), .ZN(n14844) );
  XOR2_X1 U16164 ( .A(n10245), .B(n14844), .Z(n14838) );
  NAND2_X1 U16165 ( .A1(n14838), .A2(n16012), .ZN(n15031) );
  AND2_X1 U16166 ( .A1(n14840), .A2(n14839), .ZN(n14841) );
  NAND2_X1 U16167 ( .A1(n14914), .A2(n14841), .ZN(n15033) );
  NOR2_X1 U16168 ( .A1(n14997), .A2(n15033), .ZN(n14847) );
  INV_X1 U16169 ( .A(n10245), .ZN(n15032) );
  NOR2_X1 U16170 ( .A1(n15032), .A2(n15933), .ZN(n14842) );
  AOI211_X1 U16171 ( .C1(n15894), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14847), 
        .B(n14842), .ZN(n14843) );
  OAI21_X1 U16172 ( .B1(n14880), .B2(n15031), .A(n14843), .ZN(P1_U3263) );
  OAI211_X1 U16173 ( .C1(n14845), .C2(n15035), .A(n16012), .B(n14844), .ZN(
        n15034) );
  AND2_X1 U16174 ( .A1(n15894), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14846) );
  NOR2_X1 U16175 ( .A1(n14847), .A2(n14846), .ZN(n14850) );
  NAND2_X1 U16176 ( .A1(n14848), .A2(n15026), .ZN(n14849) );
  OAI211_X1 U16177 ( .C1(n15034), .C2(n14880), .A(n14850), .B(n14849), .ZN(
        P1_U3264) );
  OAI22_X1 U16178 ( .A1(n14853), .A2(n14852), .B1(n14851), .B2(n15931), .ZN(
        n14856) );
  NOR2_X1 U16179 ( .A1(n14997), .A2(n14854), .ZN(n14855) );
  AOI211_X1 U16180 ( .C1(n15894), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14856), 
        .B(n14855), .ZN(n14857) );
  OAI21_X1 U16181 ( .B1(n14858), .B2(n15933), .A(n14857), .ZN(n14859) );
  AOI21_X1 U16182 ( .B1(n14861), .B2(n14860), .A(n14859), .ZN(n14864) );
  NAND2_X1 U16183 ( .A1(n14862), .A2(n15001), .ZN(n14863) );
  OAI211_X1 U16184 ( .C1(n14865), .C2(n15003), .A(n14864), .B(n14863), .ZN(
        P1_U3356) );
  AOI211_X1 U16185 ( .C1(n14868), .C2(n14867), .A(n16134), .B(n14866), .ZN(
        n14870) );
  OAI21_X1 U16186 ( .B1(n14872), .B2(n15036), .A(n16012), .ZN(n14873) );
  NAND2_X1 U16187 ( .A1(n14997), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14875) );
  OAI21_X1 U16188 ( .B1(n15931), .B2(n14876), .A(n14875), .ZN(n14877) );
  AOI21_X1 U16189 ( .B1(n14878), .B2(n15026), .A(n14877), .ZN(n14879) );
  OAI21_X1 U16190 ( .B1(n15038), .B2(n14880), .A(n14879), .ZN(n14881) );
  AOI21_X1 U16191 ( .B1(n15040), .B2(n15001), .A(n14881), .ZN(n14882) );
  OAI21_X1 U16192 ( .B1(n8416), .B2(n14997), .A(n14882), .ZN(P1_U3265) );
  XOR2_X1 U16193 ( .A(n7285), .B(n14884), .Z(n15053) );
  XOR2_X1 U16194 ( .A(n14884), .B(n14883), .Z(n15051) );
  OAI21_X1 U16195 ( .B1(n7775), .B2(n14886), .A(n14885), .ZN(n15049) );
  NOR2_X1 U16196 ( .A1(n15942), .A2(n14887), .ZN(n14891) );
  INV_X1 U16197 ( .A(n15046), .ZN(n14889) );
  OAI22_X1 U16198 ( .A1(n14997), .A2(n14889), .B1(n14888), .B2(n15931), .ZN(
        n14890) );
  AOI211_X1 U16199 ( .C1(n15047), .C2(n15026), .A(n14891), .B(n14890), .ZN(
        n14892) );
  OAI21_X1 U16200 ( .B1(n15049), .B2(n15936), .A(n14892), .ZN(n14893) );
  AOI21_X1 U16201 ( .B1(n15051), .B2(n15001), .A(n14893), .ZN(n14894) );
  OAI21_X1 U16202 ( .B1(n15053), .B2(n15003), .A(n14894), .ZN(P1_U3267) );
  AOI21_X1 U16203 ( .B1(n14898), .B2(n14896), .A(n14895), .ZN(n15061) );
  OAI21_X1 U16204 ( .B1(n14899), .B2(n14898), .A(n14897), .ZN(n14900) );
  INV_X1 U16205 ( .A(n14900), .ZN(n15059) );
  NAND2_X1 U16206 ( .A1(n14919), .A2(n15055), .ZN(n14901) );
  NAND2_X1 U16207 ( .A1(n14902), .A2(n14901), .ZN(n15057) );
  NOR2_X1 U16208 ( .A1(n15942), .A2(n14903), .ZN(n14907) );
  INV_X1 U16209 ( .A(n15054), .ZN(n14905) );
  OAI22_X1 U16210 ( .A1(n14997), .A2(n14905), .B1(n14904), .B2(n15931), .ZN(
        n14906) );
  AOI211_X1 U16211 ( .C1(n15055), .C2(n15026), .A(n14907), .B(n14906), .ZN(
        n14908) );
  OAI21_X1 U16212 ( .B1(n15057), .B2(n15936), .A(n14908), .ZN(n14909) );
  AOI21_X1 U16213 ( .B1(n15059), .B2(n15001), .A(n14909), .ZN(n14910) );
  OAI21_X1 U16214 ( .B1(n15061), .B2(n15003), .A(n14910), .ZN(P1_U3268) );
  AOI21_X1 U16215 ( .B1(n14916), .B2(n14911), .A(n7247), .ZN(n15067) );
  AOI22_X1 U16216 ( .A1(n14914), .A2(n14913), .B1(n15925), .B2(n14912), .ZN(
        n14918) );
  OAI211_X1 U16217 ( .C1(n7296), .C2(n14916), .A(n14915), .B(n16019), .ZN(
        n14917) );
  OAI211_X1 U16218 ( .C1(n15067), .C2(n15927), .A(n14918), .B(n14917), .ZN(
        n15062) );
  NAND2_X1 U16219 ( .A1(n15062), .A2(n15942), .ZN(n14928) );
  INV_X1 U16220 ( .A(n15069), .ZN(n14921) );
  INV_X1 U16221 ( .A(n14919), .ZN(n14920) );
  AOI21_X1 U16222 ( .B1(n15063), .B2(n14921), .A(n14920), .ZN(n15064) );
  NOR2_X1 U16223 ( .A1(n14922), .A2(n15933), .ZN(n14926) );
  OAI22_X1 U16224 ( .A1(n15942), .A2(n14924), .B1(n14923), .B2(n15931), .ZN(
        n14925) );
  AOI211_X1 U16225 ( .C1(n15064), .C2(n14958), .A(n14926), .B(n14925), .ZN(
        n14927) );
  OAI211_X1 U16226 ( .C1(n15067), .C2(n15029), .A(n14928), .B(n14927), .ZN(
        P1_U3269) );
  AOI21_X1 U16227 ( .B1(n14930), .B2(n14932), .A(n14929), .ZN(n15076) );
  OAI21_X1 U16228 ( .B1(n14933), .B2(n14932), .A(n14931), .ZN(n14934) );
  INV_X1 U16229 ( .A(n14934), .ZN(n15068) );
  NAND2_X1 U16230 ( .A1(n15068), .A2(n15001), .ZN(n14943) );
  INV_X1 U16231 ( .A(n14935), .ZN(n14936) );
  AOI22_X1 U16232 ( .A1(n15942), .A2(n15072), .B1(n14936), .B2(n15887), .ZN(
        n14937) );
  OAI21_X1 U16233 ( .B1(n14938), .B2(n15942), .A(n14937), .ZN(n14941) );
  NOR2_X1 U16234 ( .A1(n14939), .A2(n14947), .ZN(n15070) );
  NOR3_X1 U16235 ( .A1(n15070), .A2(n15069), .A3(n15936), .ZN(n14940) );
  AOI211_X1 U16236 ( .C1(n15026), .C2(n15073), .A(n14941), .B(n14940), .ZN(
        n14942) );
  OAI211_X1 U16237 ( .C1(n15076), .C2(n15003), .A(n14943), .B(n14942), .ZN(
        P1_U3270) );
  XNOR2_X1 U16238 ( .A(n14944), .B(n14945), .ZN(n15085) );
  AND2_X1 U16239 ( .A1(n15077), .A2(n7225), .ZN(n14946) );
  NOR2_X1 U16240 ( .A1(n14947), .A2(n14946), .ZN(n15083) );
  INV_X1 U16241 ( .A(n14948), .ZN(n14949) );
  OAI22_X1 U16242 ( .A1(n15078), .A2(n14997), .B1(n14949), .B2(n15931), .ZN(
        n14950) );
  AOI21_X1 U16243 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(n14997), .A(n14950), 
        .ZN(n14951) );
  OAI21_X1 U16244 ( .B1(n14952), .B2(n15933), .A(n14951), .ZN(n14957) );
  AOI21_X1 U16245 ( .B1(n14955), .B2(n14954), .A(n14953), .ZN(n15080) );
  NOR2_X1 U16246 ( .A1(n15080), .A2(n14974), .ZN(n14956) );
  AOI211_X1 U16247 ( .C1(n15083), .C2(n14958), .A(n14957), .B(n14956), .ZN(
        n14959) );
  OAI21_X1 U16248 ( .B1(n15085), .B2(n15003), .A(n14959), .ZN(P1_U3271) );
  XNOR2_X1 U16249 ( .A(n14961), .B(n14960), .ZN(n15093) );
  XNOR2_X1 U16250 ( .A(n14962), .B(n14963), .ZN(n15091) );
  INV_X1 U16251 ( .A(n14964), .ZN(n15095) );
  OAI21_X1 U16252 ( .B1(n15095), .B2(n14967), .A(n7225), .ZN(n15089) );
  INV_X1 U16253 ( .A(n14965), .ZN(n14966) );
  OAI22_X1 U16254 ( .A1(n15088), .A2(n15894), .B1(n14966), .B2(n15931), .ZN(
        n14969) );
  NOR2_X1 U16255 ( .A1(n14967), .A2(n15933), .ZN(n14968) );
  AOI211_X1 U16256 ( .C1(n15894), .C2(P1_REG2_REG_21__SCAN_IN), .A(n14969), 
        .B(n14968), .ZN(n14970) );
  OAI21_X1 U16257 ( .B1(n15089), .B2(n15936), .A(n14970), .ZN(n14971) );
  AOI21_X1 U16258 ( .B1(n15091), .B2(n14972), .A(n14971), .ZN(n14973) );
  OAI21_X1 U16259 ( .B1(n15093), .B2(n14974), .A(n14973), .ZN(P1_U3272) );
  OAI21_X1 U16260 ( .B1(n14976), .B2(n14979), .A(n14975), .ZN(n15102) );
  AOI21_X1 U16261 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n15094) );
  NAND2_X1 U16262 ( .A1(n15094), .A2(n15001), .ZN(n14988) );
  INV_X1 U16263 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14983) );
  INV_X1 U16264 ( .A(n14980), .ZN(n14981) );
  AOI22_X1 U16265 ( .A1(n15098), .A2(n15942), .B1(n14981), .B2(n15887), .ZN(
        n14982) );
  OAI21_X1 U16266 ( .B1(n14983), .B2(n15942), .A(n14982), .ZN(n14986) );
  NOR2_X1 U16267 ( .A1(n14992), .A2(n14984), .ZN(n15096) );
  NOR3_X1 U16268 ( .A1(n15096), .A2(n15095), .A3(n15936), .ZN(n14985) );
  AOI211_X1 U16269 ( .C1(n15026), .C2(n15099), .A(n14986), .B(n14985), .ZN(
        n14987) );
  OAI211_X1 U16270 ( .C1(n15102), .C2(n15003), .A(n14988), .B(n14987), .ZN(
        P1_U3273) );
  XNOR2_X1 U16271 ( .A(n7330), .B(n14990), .ZN(n15111) );
  OAI21_X1 U16272 ( .B1(n14991), .B2(n14990), .A(n14989), .ZN(n15109) );
  AND2_X1 U16273 ( .A1(n15105), .A2(n15022), .ZN(n14993) );
  OR2_X1 U16274 ( .A1(n14993), .A2(n14992), .ZN(n15107) );
  NAND2_X1 U16275 ( .A1(n15887), .A2(n14994), .ZN(n14996) );
  NAND2_X1 U16276 ( .A1(n14997), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n14995) );
  OAI211_X1 U16277 ( .C1(n15103), .C2(n14997), .A(n14996), .B(n14995), .ZN(
        n14998) );
  AOI21_X1 U16278 ( .B1(n15105), .B2(n15026), .A(n14998), .ZN(n14999) );
  OAI21_X1 U16279 ( .B1(n15107), .B2(n15936), .A(n14999), .ZN(n15000) );
  AOI21_X1 U16280 ( .B1(n15109), .B2(n15001), .A(n15000), .ZN(n15002) );
  OAI21_X1 U16281 ( .B1(n15111), .B2(n15003), .A(n15002), .ZN(P1_U3274) );
  NAND2_X1 U16282 ( .A1(n15005), .A2(n15004), .ZN(n15006) );
  NAND2_X1 U16283 ( .A1(n15007), .A2(n15006), .ZN(n15112) );
  INV_X1 U16284 ( .A(n15112), .ZN(n15030) );
  NAND2_X1 U16285 ( .A1(n15112), .A2(n15877), .ZN(n15018) );
  INV_X1 U16286 ( .A(n15008), .ZN(n15016) );
  AOI21_X1 U16287 ( .B1(n15010), .B2(n15009), .A(n16134), .ZN(n15015) );
  OAI21_X1 U16288 ( .B1(n15013), .B2(n15012), .A(n15011), .ZN(n15014) );
  AOI21_X1 U16289 ( .B1(n15016), .B2(n15015), .A(n15014), .ZN(n15017) );
  NAND2_X1 U16290 ( .A1(n15018), .A2(n15017), .ZN(n15115) );
  NAND2_X1 U16291 ( .A1(n15115), .A2(n15942), .ZN(n15028) );
  OAI22_X1 U16292 ( .A1(n15942), .A2(n15020), .B1(n15019), .B2(n15931), .ZN(
        n15024) );
  NAND2_X1 U16293 ( .A1(n15025), .A2(n15118), .ZN(n15021) );
  NAND2_X1 U16294 ( .A1(n15022), .A2(n15021), .ZN(n15113) );
  NOR2_X1 U16295 ( .A1(n15113), .A2(n15936), .ZN(n15023) );
  AOI211_X1 U16296 ( .C1(n15026), .C2(n15025), .A(n15024), .B(n15023), .ZN(
        n15027) );
  OAI211_X1 U16297 ( .C1(n15030), .C2(n15029), .A(n15028), .B(n15027), .ZN(
        P1_U3275) );
  OAI211_X1 U16298 ( .C1(n15032), .C2(n16133), .A(n15031), .B(n15033), .ZN(
        n15133) );
  MUX2_X1 U16299 ( .A(n15133), .B(P1_REG1_REG_31__SCAN_IN), .S(n16140), .Z(
        P1_U3559) );
  OAI211_X1 U16300 ( .C1(n15035), .C2(n16133), .A(n15034), .B(n15033), .ZN(
        n15134) );
  MUX2_X1 U16301 ( .A(n15134), .B(P1_REG1_REG_30__SCAN_IN), .S(n16140), .Z(
        P1_U3558) );
  NAND2_X1 U16302 ( .A1(n14878), .A2(n16009), .ZN(n15037) );
  MUX2_X1 U16303 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15136), .S(n16141), .Z(
        P1_U3556) );
  AOI22_X1 U16304 ( .A1(n15043), .A2(n16012), .B1(n15042), .B2(n15126), .ZN(
        n15044) );
  MUX2_X1 U16305 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15137), .S(n16141), .Z(
        P1_U3555) );
  AOI21_X1 U16306 ( .B1(n15047), .B2(n15126), .A(n15046), .ZN(n15048) );
  OAI21_X1 U16307 ( .B1(n15049), .B2(n16077), .A(n15048), .ZN(n15050) );
  AOI21_X1 U16308 ( .B1(n15051), .B2(n16139), .A(n15050), .ZN(n15052) );
  OAI21_X1 U16309 ( .B1(n16134), .B2(n15053), .A(n15052), .ZN(n15138) );
  MUX2_X1 U16310 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15138), .S(n16141), .Z(
        P1_U3554) );
  AOI21_X1 U16311 ( .B1(n15055), .B2(n15126), .A(n15054), .ZN(n15056) );
  OAI21_X1 U16312 ( .B1(n15057), .B2(n16077), .A(n15056), .ZN(n15058) );
  AOI21_X1 U16313 ( .B1(n15059), .B2(n16139), .A(n15058), .ZN(n15060) );
  OAI21_X1 U16314 ( .B1(n16134), .B2(n15061), .A(n15060), .ZN(n15139) );
  MUX2_X1 U16315 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15139), .S(n16141), .Z(
        P1_U3553) );
  INV_X1 U16316 ( .A(n15062), .ZN(n15066) );
  AOI22_X1 U16317 ( .A1(n15064), .A2(n16012), .B1(n15063), .B2(n15126), .ZN(
        n15065) );
  OAI211_X1 U16318 ( .C1(n15067), .C2(n15881), .A(n15066), .B(n15065), .ZN(
        n15140) );
  MUX2_X1 U16319 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15140), .S(n16141), .Z(
        P1_U3552) );
  NAND2_X1 U16320 ( .A1(n15068), .A2(n16139), .ZN(n15075) );
  NOR3_X1 U16321 ( .A1(n15070), .A2(n15069), .A3(n16077), .ZN(n15071) );
  AOI211_X1 U16322 ( .C1(n15073), .C2(n16009), .A(n15072), .B(n15071), .ZN(
        n15074) );
  OAI211_X1 U16323 ( .C1(n16134), .C2(n15076), .A(n15075), .B(n15074), .ZN(
        n15141) );
  MUX2_X1 U16324 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15141), .S(n16141), .Z(
        P1_U3551) );
  NAND2_X1 U16325 ( .A1(n15077), .A2(n16009), .ZN(n15079) );
  NAND2_X1 U16326 ( .A1(n15079), .A2(n15078), .ZN(n15082) );
  NOR2_X1 U16327 ( .A1(n15080), .A2(n16015), .ZN(n15081) );
  AOI211_X1 U16328 ( .C1(n16012), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        n15084) );
  OAI21_X1 U16329 ( .B1(n16134), .B2(n15085), .A(n15084), .ZN(n15142) );
  MUX2_X1 U16330 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15142), .S(n16141), .Z(
        P1_U3550) );
  NAND2_X1 U16331 ( .A1(n15086), .A2(n15126), .ZN(n15087) );
  OAI211_X1 U16332 ( .C1(n15089), .C2(n16077), .A(n15088), .B(n15087), .ZN(
        n15090) );
  AOI21_X1 U16333 ( .B1(n15091), .B2(n16019), .A(n15090), .ZN(n15092) );
  OAI21_X1 U16334 ( .B1(n15093), .B2(n16015), .A(n15092), .ZN(n15143) );
  MUX2_X1 U16335 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15143), .S(n16141), .Z(
        P1_U3549) );
  NAND2_X1 U16336 ( .A1(n15094), .A2(n16139), .ZN(n15101) );
  NOR3_X1 U16337 ( .A1(n15096), .A2(n15095), .A3(n16077), .ZN(n15097) );
  AOI211_X1 U16338 ( .C1(n15099), .C2(n15126), .A(n15098), .B(n15097), .ZN(
        n15100) );
  OAI211_X1 U16339 ( .C1(n16134), .C2(n15102), .A(n15101), .B(n15100), .ZN(
        n15144) );
  MUX2_X1 U16340 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15144), .S(n16141), .Z(
        P1_U3548) );
  INV_X1 U16341 ( .A(n15103), .ZN(n15104) );
  AOI21_X1 U16342 ( .B1(n15105), .B2(n15126), .A(n15104), .ZN(n15106) );
  OAI21_X1 U16343 ( .B1(n15107), .B2(n16077), .A(n15106), .ZN(n15108) );
  AOI21_X1 U16344 ( .B1(n15109), .B2(n16139), .A(n15108), .ZN(n15110) );
  OAI21_X1 U16345 ( .B1(n15111), .B2(n16134), .A(n15110), .ZN(n15145) );
  MUX2_X1 U16346 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15145), .S(n16141), .Z(
        P1_U3547) );
  AND2_X1 U16347 ( .A1(n15112), .A2(n7680), .ZN(n15116) );
  OAI22_X1 U16348 ( .A1(n15113), .A2(n16077), .B1(n8857), .B2(n16133), .ZN(
        n15114) );
  MUX2_X1 U16349 ( .A(n15146), .B(P1_REG1_REG_18__SCAN_IN), .S(n16140), .Z(
        P1_U3546) );
  NAND3_X1 U16350 ( .A1(n15118), .A2(n16012), .A3(n15117), .ZN(n15120) );
  OAI211_X1 U16351 ( .C1(n15121), .C2(n16133), .A(n15120), .B(n15119), .ZN(
        n15122) );
  AOI21_X1 U16352 ( .B1(n15123), .B2(n16019), .A(n15122), .ZN(n15124) );
  OAI21_X1 U16353 ( .B1(n15125), .B2(n16015), .A(n15124), .ZN(n15147) );
  MUX2_X1 U16354 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15147), .S(n16141), .Z(
        P1_U3545) );
  AOI21_X1 U16355 ( .B1(n16199), .B2(n15126), .A(n16198), .ZN(n15127) );
  OAI21_X1 U16356 ( .B1(n15128), .B2(n16077), .A(n15127), .ZN(n15129) );
  AOI21_X1 U16357 ( .B1(n15130), .B2(n16139), .A(n15129), .ZN(n15131) );
  OAI21_X1 U16358 ( .B1(n16134), .B2(n15132), .A(n15131), .ZN(n15148) );
  MUX2_X1 U16359 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15148), .S(n16141), .Z(
        P1_U3544) );
  MUX2_X1 U16360 ( .A(n15133), .B(P1_REG0_REG_31__SCAN_IN), .S(n16142), .Z(
        P1_U3527) );
  MUX2_X1 U16361 ( .A(n15134), .B(P1_REG0_REG_30__SCAN_IN), .S(n16142), .Z(
        P1_U3526) );
  MUX2_X1 U16362 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15136), .S(n15984), .Z(
        P1_U3524) );
  MUX2_X1 U16363 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15137), .S(n15984), .Z(
        P1_U3523) );
  MUX2_X1 U16364 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15138), .S(n15984), .Z(
        P1_U3522) );
  MUX2_X1 U16365 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15139), .S(n15984), .Z(
        P1_U3521) );
  MUX2_X1 U16366 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15140), .S(n15984), .Z(
        P1_U3520) );
  MUX2_X1 U16367 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15141), .S(n15984), .Z(
        P1_U3519) );
  MUX2_X1 U16368 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15142), .S(n15984), .Z(
        P1_U3518) );
  MUX2_X1 U16369 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15143), .S(n15984), .Z(
        P1_U3517) );
  MUX2_X1 U16370 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15144), .S(n15984), .Z(
        P1_U3516) );
  MUX2_X1 U16371 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15145), .S(n15984), .Z(
        P1_U3515) );
  MUX2_X1 U16372 ( .A(n15146), .B(P1_REG0_REG_18__SCAN_IN), .S(n16142), .Z(
        P1_U3513) );
  MUX2_X1 U16373 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15147), .S(n15984), .Z(
        P1_U3510) );
  MUX2_X1 U16374 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15148), .S(n15984), .Z(
        P1_U3507) );
  MUX2_X1 U16375 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15149), .S(n15984), .Z(
        P1_U3504) );
  MUX2_X1 U16376 ( .A(n15150), .B(P1_D_REG_1__SCAN_IN), .S(n15400), .Z(
        P1_U3446) );
  NOR4_X1 U16377 ( .A1(n7575), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n7791), .ZN(n15151) );
  AOI21_X1 U16378 ( .B1(n15392), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15151), 
        .ZN(n15152) );
  OAI21_X1 U16379 ( .B1(n15153), .B2(n15160), .A(n15152), .ZN(P1_U3324) );
  OAI222_X1 U16380 ( .A1(P1_U3086), .A2(n15156), .B1(n15160), .B2(n15155), 
        .C1(n15154), .C2(n15157), .ZN(P1_U3326) );
  OAI222_X1 U16381 ( .A1(P1_U3086), .A2(n15161), .B1(n15160), .B2(n15159), 
        .C1(n15158), .C2(n15157), .ZN(P1_U3327) );
  MUX2_X1 U16382 ( .A(n15163), .B(n15162), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  AOI22_X1 U16383 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_62), .B1(n15165), .B2(keyinput_61), .ZN(n15164) );
  OAI221_X1 U16384 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_62), .C1(
        n15165), .C2(keyinput_61), .A(n15164), .ZN(n15391) );
  INV_X1 U16385 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15261) );
  INV_X1 U16386 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15968) );
  OAI22_X1 U16387 ( .A1(n15261), .A2(keyinput_60), .B1(n15968), .B2(
        keyinput_59), .ZN(n15166) );
  AOI221_X1 U16388 ( .B1(n15261), .B2(keyinput_60), .C1(keyinput_59), .C2(
        n15968), .A(n15166), .ZN(n15390) );
  INV_X1 U16389 ( .A(keyinput_58), .ZN(n15259) );
  INV_X1 U16390 ( .A(keyinput_57), .ZN(n15257) );
  INV_X1 U16391 ( .A(keyinput_56), .ZN(n15255) );
  INV_X1 U16392 ( .A(keyinput_55), .ZN(n15253) );
  INV_X1 U16393 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15619) );
  INV_X1 U16394 ( .A(keyinput_54), .ZN(n15251) );
  INV_X1 U16395 ( .A(keyinput_47), .ZN(n15240) );
  INV_X1 U16396 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15354) );
  INV_X1 U16397 ( .A(keyinput_40), .ZN(n15228) );
  INV_X1 U16398 ( .A(keyinput_39), .ZN(n15226) );
  INV_X1 U16399 ( .A(keyinput_38), .ZN(n15224) );
  INV_X1 U16400 ( .A(keyinput_37), .ZN(n15222) );
  XNOR2_X1 U16401 ( .A(SI_3_), .B(keyinput_29), .ZN(n15220) );
  OAI22_X1 U16402 ( .A1(SI_7_), .A2(keyinput_25), .B1(keyinput_27), .B2(SI_5_), 
        .ZN(n15167) );
  AOI221_X1 U16403 ( .B1(SI_7_), .B2(keyinput_25), .C1(SI_5_), .C2(keyinput_27), .A(n15167), .ZN(n15210) );
  OAI22_X1 U16404 ( .A1(SI_6_), .A2(keyinput_26), .B1(keyinput_28), .B2(SI_4_), 
        .ZN(n15168) );
  AOI221_X1 U16405 ( .B1(SI_6_), .B2(keyinput_26), .C1(SI_4_), .C2(keyinput_28), .A(n15168), .ZN(n15209) );
  OAI22_X1 U16406 ( .A1(n15170), .A2(keyinput_22), .B1(keyinput_23), .B2(SI_9_), .ZN(n15169) );
  AOI221_X1 U16407 ( .B1(n15170), .B2(keyinput_22), .C1(SI_9_), .C2(
        keyinput_23), .A(n15169), .ZN(n15206) );
  INV_X1 U16408 ( .A(keyinput_21), .ZN(n15204) );
  INV_X1 U16409 ( .A(SI_23_), .ZN(n15172) );
  OAI22_X1 U16410 ( .A1(n15172), .A2(keyinput_9), .B1(keyinput_10), .B2(SI_22_), .ZN(n15171) );
  AOI221_X1 U16411 ( .B1(n15172), .B2(keyinput_9), .C1(SI_22_), .C2(
        keyinput_10), .A(n15171), .ZN(n15187) );
  INV_X1 U16412 ( .A(keyinput_8), .ZN(n15185) );
  INV_X1 U16413 ( .A(keyinput_7), .ZN(n15183) );
  INV_X1 U16414 ( .A(keyinput_2), .ZN(n15175) );
  OAI22_X1 U16415 ( .A1(SI_31_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        P3_WR_REG_SCAN_IN), .ZN(n15173) );
  AOI221_X1 U16416 ( .B1(SI_31_), .B2(keyinput_1), .C1(P3_WR_REG_SCAN_IN), 
        .C2(keyinput_0), .A(n15173), .ZN(n15174) );
  AOI221_X1 U16417 ( .B1(SI_30_), .B2(keyinput_2), .C1(n15281), .C2(n15175), 
        .A(n15174), .ZN(n15181) );
  AOI22_X1 U16418 ( .A1(n15177), .A2(keyinput_4), .B1(n15277), .B2(keyinput_3), 
        .ZN(n15176) );
  OAI221_X1 U16419 ( .B1(n15177), .B2(keyinput_4), .C1(n15277), .C2(keyinput_3), .A(n15176), .ZN(n15180) );
  OAI22_X1 U16420 ( .A1(n15283), .A2(keyinput_5), .B1(keyinput_6), .B2(SI_26_), 
        .ZN(n15178) );
  AOI221_X1 U16421 ( .B1(n15283), .B2(keyinput_5), .C1(SI_26_), .C2(keyinput_6), .A(n15178), .ZN(n15179) );
  OAI21_X1 U16422 ( .B1(n15181), .B2(n15180), .A(n15179), .ZN(n15182) );
  OAI221_X1 U16423 ( .B1(SI_25_), .B2(keyinput_7), .C1(n15290), .C2(n15183), 
        .A(n15182), .ZN(n15184) );
  OAI221_X1 U16424 ( .B1(SI_24_), .B2(n15185), .C1(n15293), .C2(keyinput_8), 
        .A(n15184), .ZN(n15186) );
  OAI211_X1 U16425 ( .C1(n15189), .C2(keyinput_11), .A(n15187), .B(n15186), 
        .ZN(n15188) );
  AOI21_X1 U16426 ( .B1(n15189), .B2(keyinput_11), .A(n15188), .ZN(n15190) );
  AOI21_X1 U16427 ( .B1(SI_20_), .B2(keyinput_12), .A(n15190), .ZN(n15194) );
  AOI22_X1 U16428 ( .A1(SI_18_), .A2(keyinput_14), .B1(n15192), .B2(
        keyinput_13), .ZN(n15191) );
  OAI221_X1 U16429 ( .B1(SI_18_), .B2(keyinput_14), .C1(n15192), .C2(
        keyinput_13), .A(n15191), .ZN(n15193) );
  AOI221_X1 U16430 ( .B1(SI_20_), .B2(n15194), .C1(keyinput_12), .C2(n15194), 
        .A(n15193), .ZN(n15202) );
  AOI22_X1 U16431 ( .A1(n15196), .A2(keyinput_16), .B1(n15275), .B2(
        keyinput_15), .ZN(n15195) );
  OAI221_X1 U16432 ( .B1(n15196), .B2(keyinput_16), .C1(n15275), .C2(
        keyinput_15), .A(n15195), .ZN(n15201) );
  OAI22_X1 U16433 ( .A1(SI_15_), .A2(keyinput_17), .B1(SI_12_), .B2(
        keyinput_20), .ZN(n15197) );
  AOI221_X1 U16434 ( .B1(SI_15_), .B2(keyinput_17), .C1(keyinput_20), .C2(
        SI_12_), .A(n15197), .ZN(n15200) );
  OAI22_X1 U16435 ( .A1(SI_14_), .A2(keyinput_18), .B1(SI_13_), .B2(
        keyinput_19), .ZN(n15198) );
  AOI221_X1 U16436 ( .B1(SI_14_), .B2(keyinput_18), .C1(keyinput_19), .C2(
        SI_13_), .A(n15198), .ZN(n15199) );
  OAI211_X1 U16437 ( .C1(n15202), .C2(n15201), .A(n15200), .B(n15199), .ZN(
        n15203) );
  OAI221_X1 U16438 ( .B1(SI_11_), .B2(keyinput_21), .C1(n15313), .C2(n15204), 
        .A(n15203), .ZN(n15205) );
  AOI22_X1 U16439 ( .A1(keyinput_24), .A2(n15320), .B1(n15206), .B2(n15205), 
        .ZN(n15207) );
  OAI21_X1 U16440 ( .B1(n15320), .B2(keyinput_24), .A(n15207), .ZN(n15208) );
  NAND3_X1 U16441 ( .A1(n15210), .A2(n15209), .A3(n15208), .ZN(n15219) );
  AOI22_X1 U16442 ( .A1(SI_2_), .A2(keyinput_30), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(keyinput_36), .ZN(n15211) );
  OAI221_X1 U16443 ( .B1(SI_2_), .B2(keyinput_30), .C1(P3_REG3_REG_27__SCAN_IN), .C2(keyinput_36), .A(n15211), .ZN(n15218) );
  INV_X1 U16444 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15852) );
  AOI22_X1 U16445 ( .A1(P3_U3151), .A2(keyinput_34), .B1(keyinput_33), .B2(
        n15852), .ZN(n15212) );
  OAI221_X1 U16446 ( .B1(P3_U3151), .B2(keyinput_34), .C1(n15852), .C2(
        keyinput_33), .A(n15212), .ZN(n15215) );
  INV_X1 U16447 ( .A(SI_1_), .ZN(n15266) );
  AOI22_X1 U16448 ( .A1(SI_0_), .A2(keyinput_32), .B1(n15266), .B2(keyinput_31), .ZN(n15213) );
  OAI221_X1 U16449 ( .B1(SI_0_), .B2(keyinput_32), .C1(n15266), .C2(
        keyinput_31), .A(n15213), .ZN(n15214) );
  AOI211_X1 U16450 ( .C1(keyinput_35), .C2(P3_REG3_REG_7__SCAN_IN), .A(n15215), 
        .B(n15214), .ZN(n15216) );
  OAI21_X1 U16451 ( .B1(keyinput_35), .B2(P3_REG3_REG_7__SCAN_IN), .A(n15216), 
        .ZN(n15217) );
  AOI211_X1 U16452 ( .C1(n15220), .C2(n15219), .A(n15218), .B(n15217), .ZN(
        n15221) );
  AOI221_X1 U16453 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(
        n15335), .C2(n15222), .A(n15221), .ZN(n15223) );
  AOI221_X1 U16454 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        n13478), .C2(n15224), .A(n15223), .ZN(n15225) );
  AOI221_X1 U16455 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(n15226), .C1(n15339), 
        .C2(keyinput_39), .A(n15225), .ZN(n15227) );
  AOI221_X1 U16456 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(n15343), .C2(n15228), .A(n15227), .ZN(n15238) );
  AOI22_X1 U16457 ( .A1(n15230), .A2(keyinput_46), .B1(n15348), .B2(
        keyinput_45), .ZN(n15229) );
  OAI221_X1 U16458 ( .B1(n15230), .B2(keyinput_46), .C1(n15348), .C2(
        keyinput_45), .A(n15229), .ZN(n15237) );
  INV_X1 U16459 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15232) );
  AOI22_X1 U16460 ( .A1(n15232), .A2(keyinput_41), .B1(keyinput_43), .B2(
        n15346), .ZN(n15231) );
  OAI221_X1 U16461 ( .B1(n15232), .B2(keyinput_41), .C1(n15346), .C2(
        keyinput_43), .A(n15231), .ZN(n15236) );
  INV_X1 U16462 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U16463 ( .A1(n9570), .A2(keyinput_42), .B1(keyinput_44), .B2(n15234), .ZN(n15233) );
  OAI221_X1 U16464 ( .B1(n9570), .B2(keyinput_42), .C1(n15234), .C2(
        keyinput_44), .A(n15233), .ZN(n15235) );
  NOR4_X1 U16465 ( .A1(n15238), .A2(n15237), .A3(n15236), .A4(n15235), .ZN(
        n15239) );
  AOI221_X1 U16466 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n15240), .C1(n15354), 
        .C2(keyinput_47), .A(n15239), .ZN(n15244) );
  OAI22_X1 U16467 ( .A1(n9392), .A2(keyinput_50), .B1(n9158), .B2(keyinput_49), 
        .ZN(n15241) );
  AOI221_X1 U16468 ( .B1(n9392), .B2(keyinput_50), .C1(keyinput_49), .C2(n9158), .A(n15241), .ZN(n15242) );
  OAI21_X1 U16469 ( .B1(keyinput_48), .B2(P3_REG3_REG_16__SCAN_IN), .A(n15242), 
        .ZN(n15243) );
  AOI211_X1 U16470 ( .C1(keyinput_48), .C2(P3_REG3_REG_16__SCAN_IN), .A(n15244), .B(n15243), .ZN(n15248) );
  AOI22_X1 U16471 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(keyinput_52), .B1(n15246), 
        .B2(keyinput_51), .ZN(n15245) );
  OAI221_X1 U16472 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .C1(n15246), .C2(keyinput_51), .A(n15245), .ZN(n15247) );
  AOI211_X1 U16473 ( .C1(P3_REG3_REG_9__SCAN_IN), .C2(keyinput_53), .A(n15248), 
        .B(n15247), .ZN(n15249) );
  OAI21_X1 U16474 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .A(n15249), 
        .ZN(n15250) );
  OAI221_X1 U16475 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .C1(n15619), .C2(n15251), .A(n15250), .ZN(n15252) );
  OAI221_X1 U16476 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(
        n15369), .C2(n15253), .A(n15252), .ZN(n15254) );
  OAI221_X1 U16477 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(n15255), .C1(n9318), 
        .C2(keyinput_56), .A(n15254), .ZN(n15256) );
  OAI221_X1 U16478 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .C1(
        n15374), .C2(n15257), .A(n15256), .ZN(n15258) );
  OAI221_X1 U16479 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .C1(
        n15377), .C2(n15259), .A(n15258), .ZN(n15389) );
  INV_X1 U16480 ( .A(keyinput_127), .ZN(n15382) );
  OAI22_X1 U16481 ( .A1(n15261), .A2(keyinput_124), .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .ZN(n15260) );
  AOI221_X1 U16482 ( .B1(n15261), .B2(keyinput_124), .C1(keyinput_123), .C2(
        P3_REG3_REG_2__SCAN_IN), .A(n15260), .ZN(n15381) );
  INV_X1 U16483 ( .A(keyinput_122), .ZN(n15376) );
  INV_X1 U16484 ( .A(keyinput_121), .ZN(n15373) );
  INV_X1 U16485 ( .A(keyinput_120), .ZN(n15371) );
  INV_X1 U16486 ( .A(keyinput_119), .ZN(n15368) );
  INV_X1 U16487 ( .A(keyinput_118), .ZN(n15366) );
  INV_X1 U16488 ( .A(keyinput_111), .ZN(n15355) );
  INV_X1 U16489 ( .A(keyinput_104), .ZN(n15342) );
  INV_X1 U16490 ( .A(keyinput_103), .ZN(n15340) );
  INV_X1 U16491 ( .A(keyinput_102), .ZN(n15337) );
  INV_X1 U16492 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15264) );
  OAI22_X1 U16493 ( .A1(n15264), .A2(keyinput_100), .B1(n15263), .B2(
        keyinput_99), .ZN(n15262) );
  AOI221_X1 U16494 ( .B1(n15264), .B2(keyinput_100), .C1(keyinput_99), .C2(
        n15263), .A(n15262), .ZN(n15273) );
  OAI22_X1 U16495 ( .A1(n15266), .A2(keyinput_95), .B1(keyinput_98), .B2(
        P3_STATE_REG_SCAN_IN), .ZN(n15265) );
  AOI221_X1 U16496 ( .B1(n15266), .B2(keyinput_95), .C1(P3_STATE_REG_SCAN_IN), 
        .C2(keyinput_98), .A(n15265), .ZN(n15272) );
  XNOR2_X1 U16497 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_97), .ZN(n15271) );
  XOR2_X1 U16498 ( .A(SI_2_), .B(keyinput_94), .Z(n15269) );
  INV_X1 U16499 ( .A(SI_0_), .ZN(n15267) );
  XNOR2_X1 U16500 ( .A(keyinput_96), .B(n15267), .ZN(n15268) );
  NOR2_X1 U16501 ( .A1(n15269), .A2(n15268), .ZN(n15270) );
  NAND4_X1 U16502 ( .A1(n15273), .A2(n15272), .A3(n15271), .A4(n15270), .ZN(
        n15333) );
  INV_X1 U16503 ( .A(keyinput_93), .ZN(n15330) );
  INV_X1 U16504 ( .A(keyinput_85), .ZN(n15314) );
  OAI22_X1 U16505 ( .A1(n15275), .A2(keyinput_79), .B1(SI_16_), .B2(
        keyinput_80), .ZN(n15274) );
  AOI221_X1 U16506 ( .B1(n15275), .B2(keyinput_79), .C1(keyinput_80), .C2(
        SI_16_), .A(n15274), .ZN(n15311) );
  XOR2_X1 U16507 ( .A(SI_20_), .B(keyinput_76), .Z(n15302) );
  INV_X1 U16508 ( .A(keyinput_72), .ZN(n15292) );
  INV_X1 U16509 ( .A(keyinput_71), .ZN(n15289) );
  OAI22_X1 U16510 ( .A1(n15277), .A2(keyinput_67), .B1(SI_28_), .B2(
        keyinput_68), .ZN(n15276) );
  AOI221_X1 U16511 ( .B1(n15277), .B2(keyinput_67), .C1(keyinput_68), .C2(
        SI_28_), .A(n15276), .ZN(n15287) );
  INV_X1 U16512 ( .A(keyinput_66), .ZN(n15280) );
  AOI22_X1 U16513 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n15278) );
  OAI221_X1 U16514 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n15278), .ZN(n15279) );
  OAI221_X1 U16515 ( .B1(SI_30_), .B2(keyinput_66), .C1(n15281), .C2(n15280), 
        .A(n15279), .ZN(n15286) );
  AOI22_X1 U16516 ( .A1(n15284), .A2(keyinput_70), .B1(n15283), .B2(
        keyinput_69), .ZN(n15282) );
  OAI221_X1 U16517 ( .B1(n15284), .B2(keyinput_70), .C1(n15283), .C2(
        keyinput_69), .A(n15282), .ZN(n15285) );
  AOI21_X1 U16518 ( .B1(n15287), .B2(n15286), .A(n15285), .ZN(n15288) );
  AOI221_X1 U16519 ( .B1(SI_25_), .B2(keyinput_71), .C1(n15290), .C2(n15289), 
        .A(n15288), .ZN(n15291) );
  AOI221_X1 U16520 ( .B1(SI_24_), .B2(keyinput_72), .C1(n15293), .C2(n15292), 
        .A(n15291), .ZN(n15298) );
  OAI22_X1 U16521 ( .A1(n15295), .A2(keyinput_74), .B1(keyinput_73), .B2(
        SI_23_), .ZN(n15294) );
  AOI221_X1 U16522 ( .B1(n15295), .B2(keyinput_74), .C1(SI_23_), .C2(
        keyinput_73), .A(n15294), .ZN(n15296) );
  OAI21_X1 U16523 ( .B1(keyinput_75), .B2(SI_21_), .A(n15296), .ZN(n15297) );
  AOI211_X1 U16524 ( .C1(keyinput_75), .C2(SI_21_), .A(n15298), .B(n15297), 
        .ZN(n15301) );
  OAI22_X1 U16525 ( .A1(SI_19_), .A2(keyinput_77), .B1(keyinput_78), .B2(
        SI_18_), .ZN(n15299) );
  AOI221_X1 U16526 ( .B1(SI_19_), .B2(keyinput_77), .C1(SI_18_), .C2(
        keyinput_78), .A(n15299), .ZN(n15300) );
  OAI21_X1 U16527 ( .B1(n15302), .B2(n15301), .A(n15300), .ZN(n15310) );
  AOI22_X1 U16528 ( .A1(n15305), .A2(keyinput_81), .B1(keyinput_83), .B2(
        n15304), .ZN(n15303) );
  OAI221_X1 U16529 ( .B1(n15305), .B2(keyinput_81), .C1(n15304), .C2(
        keyinput_83), .A(n15303), .ZN(n15309) );
  AOI22_X1 U16530 ( .A1(SI_14_), .A2(keyinput_82), .B1(n15307), .B2(
        keyinput_84), .ZN(n15306) );
  OAI221_X1 U16531 ( .B1(SI_14_), .B2(keyinput_82), .C1(n15307), .C2(
        keyinput_84), .A(n15306), .ZN(n15308) );
  AOI211_X1 U16532 ( .C1(n15311), .C2(n15310), .A(n15309), .B(n15308), .ZN(
        n15312) );
  AOI221_X1 U16533 ( .B1(SI_11_), .B2(n15314), .C1(n15313), .C2(keyinput_85), 
        .A(n15312), .ZN(n15318) );
  XOR2_X1 U16534 ( .A(SI_10_), .B(keyinput_86), .Z(n15316) );
  XNOR2_X1 U16535 ( .A(SI_9_), .B(keyinput_87), .ZN(n15315) );
  NAND2_X1 U16536 ( .A1(n15316), .A2(n15315), .ZN(n15317) );
  OAI22_X1 U16537 ( .A1(n15318), .A2(n15317), .B1(keyinput_88), .B2(n15320), 
        .ZN(n15319) );
  AOI21_X1 U16538 ( .B1(keyinput_88), .B2(n15320), .A(n15319), .ZN(n15328) );
  AOI22_X1 U16539 ( .A1(n15323), .A2(keyinput_92), .B1(n15322), .B2(
        keyinput_89), .ZN(n15321) );
  OAI221_X1 U16540 ( .B1(n15323), .B2(keyinput_92), .C1(n15322), .C2(
        keyinput_89), .A(n15321), .ZN(n15327) );
  AOI22_X1 U16541 ( .A1(SI_6_), .A2(keyinput_90), .B1(n15325), .B2(keyinput_91), .ZN(n15324) );
  OAI221_X1 U16542 ( .B1(SI_6_), .B2(keyinput_90), .C1(n15325), .C2(
        keyinput_91), .A(n15324), .ZN(n15326) );
  NOR3_X1 U16543 ( .A1(n15328), .A2(n15327), .A3(n15326), .ZN(n15329) );
  AOI221_X1 U16544 ( .B1(SI_3_), .B2(keyinput_93), .C1(n15331), .C2(n15330), 
        .A(n15329), .ZN(n15332) );
  OAI22_X1 U16545 ( .A1(keyinput_101), .A2(n15335), .B1(n15333), .B2(n15332), 
        .ZN(n15334) );
  AOI21_X1 U16546 ( .B1(keyinput_101), .B2(n15335), .A(n15334), .ZN(n15336) );
  AOI221_X1 U16547 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(n15337), .C1(n13478), 
        .C2(keyinput_102), .A(n15336), .ZN(n15338) );
  AOI221_X1 U16548 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(n15340), .C1(n15339), 
        .C2(keyinput_103), .A(n15338), .ZN(n15341) );
  AOI221_X1 U16549 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .C1(
        n15343), .C2(n15342), .A(n15341), .ZN(n15352) );
  AOI22_X1 U16550 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_108), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .ZN(n15344) );
  OAI221_X1 U16551 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_108), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_110), .A(n15344), .ZN(n15351)
         );
  AOI22_X1 U16552 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_105), .B1(
        n15346), .B2(keyinput_107), .ZN(n15345) );
  OAI221_X1 U16553 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .C1(
        n15346), .C2(keyinput_107), .A(n15345), .ZN(n15350) );
  AOI22_X1 U16554 ( .A1(n15348), .A2(keyinput_109), .B1(n9570), .B2(
        keyinput_106), .ZN(n15347) );
  OAI221_X1 U16555 ( .B1(n15348), .B2(keyinput_109), .C1(n9570), .C2(
        keyinput_106), .A(n15347), .ZN(n15349) );
  NOR4_X1 U16556 ( .A1(n15352), .A2(n15351), .A3(n15350), .A4(n15349), .ZN(
        n15353) );
  AOI221_X1 U16557 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n15355), .C1(n15354), 
        .C2(keyinput_111), .A(n15353), .ZN(n15360) );
  OAI22_X1 U16558 ( .A1(n15357), .A2(keyinput_112), .B1(keyinput_113), .B2(
        P3_REG3_REG_5__SCAN_IN), .ZN(n15356) );
  AOI221_X1 U16559 ( .B1(n15357), .B2(keyinput_112), .C1(
        P3_REG3_REG_5__SCAN_IN), .C2(keyinput_113), .A(n15356), .ZN(n15358) );
  OAI21_X1 U16560 ( .B1(keyinput_114), .B2(P3_REG3_REG_17__SCAN_IN), .A(n15358), .ZN(n15359) );
  AOI211_X1 U16561 ( .C1(keyinput_114), .C2(P3_REG3_REG_17__SCAN_IN), .A(
        n15360), .B(n15359), .ZN(n15363) );
  AOI22_X1 U16562 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_115), .B1(n9231), .B2(keyinput_117), .ZN(n15361) );
  OAI221_X1 U16563 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(
        n9231), .C2(keyinput_117), .A(n15361), .ZN(n15362) );
  AOI211_X1 U16564 ( .C1(P3_REG3_REG_4__SCAN_IN), .C2(keyinput_116), .A(n15363), .B(n15362), .ZN(n15364) );
  OAI21_X1 U16565 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(keyinput_116), .A(n15364), 
        .ZN(n15365) );
  OAI221_X1 U16566 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15366), .C1(n15619), 
        .C2(keyinput_118), .A(n15365), .ZN(n15367) );
  OAI221_X1 U16567 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        n15369), .C2(n15368), .A(n15367), .ZN(n15370) );
  OAI221_X1 U16568 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_120), .C1(
        n9318), .C2(n15371), .A(n15370), .ZN(n15372) );
  OAI221_X1 U16569 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .C1(
        n15374), .C2(n15373), .A(n15372), .ZN(n15375) );
  OAI221_X1 U16570 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        n15377), .C2(n15376), .A(n15375), .ZN(n15380) );
  AOI22_X1 U16571 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_125), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_126), .ZN(n15378) );
  OAI221_X1 U16572 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_126), .A(n15378), .ZN(n15379)
         );
  AOI21_X1 U16573 ( .B1(n15381), .B2(n15380), .A(n15379), .ZN(n15385) );
  OAI211_X1 U16574 ( .C1(n15382), .C2(n15385), .A(P3_REG3_REG_15__SCAN_IN), 
        .B(keyinput_63), .ZN(n15387) );
  INV_X1 U16575 ( .A(keyinput_63), .ZN(n15383) );
  OAI211_X1 U16576 ( .C1(n15385), .C2(keyinput_127), .A(n15384), .B(n15383), 
        .ZN(n15386) );
  NAND2_X1 U16577 ( .A1(n15387), .A2(n15386), .ZN(n15388) );
  OAI221_X1 U16578 ( .B1(n15391), .B2(n15390), .C1(n15391), .C2(n15389), .A(
        n15388), .ZN(n15397) );
  AOI222_X1 U16579 ( .A1(n15395), .A2(n15394), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15393), .C1(P2_DATAO_REG_3__SCAN_IN), .C2(n15392), .ZN(n15396) );
  XOR2_X1 U16580 ( .A(n15397), .B(n15396), .Z(P1_U3352) );
  MUX2_X1 U16581 ( .A(n15399), .B(n15398), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  AND2_X1 U16582 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15400), .ZN(P1_U3323) );
  AND2_X1 U16583 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15400), .ZN(P1_U3322) );
  AND2_X1 U16584 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15400), .ZN(P1_U3321) );
  AND2_X1 U16585 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15400), .ZN(P1_U3320) );
  AND2_X1 U16586 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15400), .ZN(P1_U3319) );
  AND2_X1 U16587 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15400), .ZN(P1_U3318) );
  AND2_X1 U16588 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15400), .ZN(P1_U3317) );
  AND2_X1 U16589 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15400), .ZN(P1_U3316) );
  AND2_X1 U16590 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15400), .ZN(P1_U3315) );
  AND2_X1 U16591 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15400), .ZN(P1_U3314) );
  AND2_X1 U16592 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15400), .ZN(P1_U3313) );
  AND2_X1 U16593 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15400), .ZN(P1_U3312) );
  AND2_X1 U16594 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15400), .ZN(P1_U3311) );
  AND2_X1 U16595 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15400), .ZN(P1_U3310) );
  AND2_X1 U16596 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15400), .ZN(P1_U3309) );
  AND2_X1 U16597 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15400), .ZN(P1_U3308) );
  AND2_X1 U16598 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15400), .ZN(P1_U3307) );
  AND2_X1 U16599 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15400), .ZN(P1_U3306) );
  AND2_X1 U16600 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15400), .ZN(P1_U3305) );
  AND2_X1 U16601 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15400), .ZN(P1_U3304) );
  AND2_X1 U16602 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15400), .ZN(P1_U3303) );
  AND2_X1 U16603 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15400), .ZN(P1_U3302) );
  AND2_X1 U16604 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15400), .ZN(P1_U3301) );
  AND2_X1 U16605 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15400), .ZN(P1_U3300) );
  AND2_X1 U16606 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15400), .ZN(P1_U3299) );
  AND2_X1 U16607 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15400), .ZN(P1_U3298) );
  AND2_X1 U16608 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15400), .ZN(P1_U3297) );
  AND2_X1 U16609 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15400), .ZN(P1_U3296) );
  AND2_X1 U16610 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15400), .ZN(P1_U3295) );
  AND2_X1 U16611 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15400), .ZN(P1_U3294) );
  AOI21_X1 U16612 ( .B1(n15402), .B2(n15406), .A(n15401), .ZN(P2_U3417) );
  AND2_X1 U16613 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15404), .ZN(P2_U3295) );
  AND2_X1 U16614 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15404), .ZN(P2_U3294) );
  AND2_X1 U16615 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15404), .ZN(P2_U3293) );
  AND2_X1 U16616 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15404), .ZN(P2_U3292) );
  AND2_X1 U16617 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15404), .ZN(P2_U3291) );
  AND2_X1 U16618 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15404), .ZN(P2_U3290) );
  AND2_X1 U16619 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15404), .ZN(P2_U3289) );
  AND2_X1 U16620 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15404), .ZN(P2_U3288) );
  AND2_X1 U16621 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15404), .ZN(P2_U3287) );
  AND2_X1 U16622 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15404), .ZN(P2_U3286) );
  AND2_X1 U16623 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15404), .ZN(P2_U3285) );
  AND2_X1 U16624 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15404), .ZN(P2_U3284) );
  AND2_X1 U16625 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15404), .ZN(P2_U3283) );
  AND2_X1 U16626 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15404), .ZN(P2_U3282) );
  AND2_X1 U16627 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15404), .ZN(P2_U3281) );
  AND2_X1 U16628 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15404), .ZN(P2_U3280) );
  AND2_X1 U16629 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15404), .ZN(P2_U3279) );
  AND2_X1 U16630 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15404), .ZN(P2_U3278) );
  AND2_X1 U16631 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15404), .ZN(P2_U3277) );
  AND2_X1 U16632 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15404), .ZN(P2_U3276) );
  AND2_X1 U16633 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15404), .ZN(P2_U3275) );
  AND2_X1 U16634 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15404), .ZN(P2_U3274) );
  AND2_X1 U16635 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15404), .ZN(P2_U3273) );
  AND2_X1 U16636 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15404), .ZN(P2_U3272) );
  AND2_X1 U16637 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15404), .ZN(P2_U3271) );
  AND2_X1 U16638 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15404), .ZN(P2_U3270) );
  AND2_X1 U16639 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15404), .ZN(P2_U3269) );
  AND2_X1 U16640 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15404), .ZN(P2_U3268) );
  AND2_X1 U16641 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15404), .ZN(P2_U3267) );
  AND2_X1 U16642 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15404), .ZN(P2_U3266) );
  NOR2_X1 U16643 ( .A1(n15502), .A2(n15405), .ZN(P2_U3087) );
  NOR2_X1 U16644 ( .A1(P3_U3897), .A2(n15832), .ZN(P3_U3150) );
  AOI22_X1 U16645 ( .A1(n15409), .A2(n15408), .B1(n15407), .B2(n15406), .ZN(
        P2_U3416) );
  AOI22_X1 U16646 ( .A1(n15502), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15424) );
  NAND2_X1 U16647 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15415) );
  INV_X1 U16648 ( .A(n15410), .ZN(n15414) );
  INV_X1 U16649 ( .A(n15411), .ZN(n15413) );
  AOI211_X1 U16650 ( .C1(n15415), .C2(n15414), .A(n15413), .B(n15412), .ZN(
        n15416) );
  AOI21_X1 U16651 ( .B1(n15452), .B2(n15417), .A(n15416), .ZN(n15423) );
  INV_X1 U16652 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15901) );
  NOR2_X1 U16653 ( .A1(n15418), .A2(n15901), .ZN(n15421) );
  OAI211_X1 U16654 ( .C1(n15421), .C2(n15420), .A(n15494), .B(n15419), .ZN(
        n15422) );
  NAND3_X1 U16655 ( .A1(n15424), .A2(n15423), .A3(n15422), .ZN(P2_U3215) );
  AOI22_X1 U16656 ( .A1(n15502), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15436) );
  OAI211_X1 U16657 ( .C1(n15427), .C2(n15426), .A(n15512), .B(n15425), .ZN(
        n15428) );
  OAI21_X1 U16658 ( .B1(n15468), .B2(n15429), .A(n15428), .ZN(n15430) );
  INV_X1 U16659 ( .A(n15430), .ZN(n15435) );
  OAI211_X1 U16660 ( .C1(n15433), .C2(n15432), .A(n15494), .B(n15431), .ZN(
        n15434) );
  NAND3_X1 U16661 ( .A1(n15436), .A2(n15435), .A3(n15434), .ZN(P2_U3216) );
  INV_X1 U16662 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15442) );
  OAI211_X1 U16663 ( .C1(n15439), .C2(n15438), .A(n15512), .B(n15437), .ZN(
        n15440) );
  OAI21_X1 U16664 ( .B1(n15442), .B2(n15441), .A(n15440), .ZN(n15443) );
  AOI21_X1 U16665 ( .B1(n15444), .B2(n15504), .A(n15443), .ZN(n15451) );
  AOI211_X1 U16666 ( .C1(n15447), .C2(n15446), .A(n15445), .B(n15508), .ZN(
        n15448) );
  INV_X1 U16667 ( .A(n15448), .ZN(n15449) );
  NAND3_X1 U16668 ( .A1(n15451), .A2(n15450), .A3(n15449), .ZN(P2_U3218) );
  INV_X1 U16669 ( .A(n15452), .ZN(n15454) );
  OAI21_X1 U16670 ( .B1(n15454), .B2(n15453), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15455) );
  OAI21_X1 U16671 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15455), .ZN(n15466) );
  NOR2_X1 U16672 ( .A1(n15457), .A2(n15456), .ZN(n15458) );
  XNOR2_X1 U16673 ( .A(n15459), .B(n15458), .ZN(n15460) );
  AOI22_X1 U16674 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n15502), .B1(n15512), 
        .B2(n15460), .ZN(n15465) );
  OAI211_X1 U16675 ( .C1(n15463), .C2(n15462), .A(n15461), .B(n15494), .ZN(
        n15464) );
  NAND3_X1 U16676 ( .A1(n15466), .A2(n15465), .A3(n15464), .ZN(P2_U3228) );
  NOR2_X1 U16677 ( .A1(n15468), .A2(n15467), .ZN(n15469) );
  AOI211_X1 U16678 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n15502), .A(n15470), 
        .B(n15469), .ZN(n15477) );
  OAI211_X1 U16679 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15472), .A(n15512), 
        .B(n15471), .ZN(n15476) );
  OAI211_X1 U16680 ( .C1(n15474), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15494), 
        .B(n15473), .ZN(n15475) );
  NAND3_X1 U16681 ( .A1(n15477), .A2(n15476), .A3(n15475), .ZN(P2_U3229) );
  AOI22_X1 U16682 ( .A1(n15502), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n15488) );
  OAI211_X1 U16683 ( .C1(n15480), .C2(n15479), .A(n15512), .B(n15478), .ZN(
        n15487) );
  NAND2_X1 U16684 ( .A1(n15504), .A2(n15481), .ZN(n15486) );
  OAI211_X1 U16685 ( .C1(n15484), .C2(n15483), .A(n15494), .B(n15482), .ZN(
        n15485) );
  NAND4_X1 U16686 ( .A1(n15488), .A2(n15487), .A3(n15486), .A4(n15485), .ZN(
        P2_U3230) );
  AOI22_X1 U16687 ( .A1(n15489), .A2(n15504), .B1(P2_ADDR_REG_13__SCAN_IN), 
        .B2(n15502), .ZN(n15501) );
  NAND2_X1 U16688 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n15500)
         );
  AOI21_X1 U16689 ( .B1(n15492), .B2(n15491), .A(n15490), .ZN(n15493) );
  NAND2_X1 U16690 ( .A1(n15512), .A2(n15493), .ZN(n15499) );
  OAI211_X1 U16691 ( .C1(n15497), .C2(n15496), .A(n15495), .B(n15494), .ZN(
        n15498) );
  NAND4_X1 U16692 ( .A1(n15501), .A2(n15500), .A3(n15499), .A4(n15498), .ZN(
        P2_U3227) );
  AOI22_X1 U16693 ( .A1(n15504), .A2(n15503), .B1(n15502), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n15517) );
  AOI21_X1 U16694 ( .B1(n15507), .B2(n15506), .A(n15505), .ZN(n15509) );
  OR2_X1 U16695 ( .A1(n15509), .A2(n15508), .ZN(n15515) );
  XNOR2_X1 U16696 ( .A(n15511), .B(n15510), .ZN(n15513) );
  NAND2_X1 U16697 ( .A1(n15513), .A2(n15512), .ZN(n15514) );
  NAND4_X1 U16698 ( .A1(n15517), .A2(n15516), .A3(n15515), .A4(n15514), .ZN(
        P2_U3226) );
  NOR2_X1 U16699 ( .A1(n15518), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15520) );
  OR2_X1 U16700 ( .A1(n15519), .A2(n15520), .ZN(n15523) );
  INV_X1 U16701 ( .A(n15520), .ZN(n15522) );
  MUX2_X1 U16702 ( .A(n15523), .B(n15522), .S(n15521), .Z(n15525) );
  NAND2_X1 U16703 ( .A1(n15525), .A2(n15524), .ZN(n15528) );
  AOI22_X1 U16704 ( .A1(n15526), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15527) );
  OAI21_X1 U16705 ( .B1(n15529), .B2(n15528), .A(n15527), .ZN(P1_U3243) );
  OAI21_X1 U16706 ( .B1(n15531), .B2(n8798), .A(n15530), .ZN(n15540) );
  AOI21_X1 U16707 ( .B1(n15533), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15532), 
        .ZN(n15537) );
  OAI22_X1 U16708 ( .A1(n15537), .A2(n15536), .B1(n15535), .B2(n15534), .ZN(
        n15538) );
  AOI21_X1 U16709 ( .B1(n15540), .B2(n15539), .A(n15538), .ZN(n15542) );
  OAI211_X1 U16710 ( .C1(n15543), .C2(n15876), .A(n15542), .B(n15541), .ZN(
        P1_U3258) );
  XOR2_X1 U16711 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15544), .Z(SUB_1596_U53) );
  OAI21_X1 U16712 ( .B1(n15547), .B2(n15546), .A(n15545), .ZN(n15548) );
  XNOR2_X1 U16713 ( .A(n15548), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  OAI21_X1 U16714 ( .B1(n15551), .B2(n15550), .A(n15549), .ZN(SUB_1596_U60) );
  AOI21_X1 U16715 ( .B1(n15554), .B2(n15553), .A(n15552), .ZN(SUB_1596_U59) );
  AOI21_X1 U16716 ( .B1(n15557), .B2(n15556), .A(n15555), .ZN(SUB_1596_U58) );
  AOI21_X1 U16717 ( .B1(n15560), .B2(n15559), .A(n15558), .ZN(SUB_1596_U56) );
  AOI21_X1 U16718 ( .B1(n15563), .B2(n15562), .A(n15561), .ZN(SUB_1596_U55) );
  AOI21_X1 U16719 ( .B1(n15566), .B2(n15565), .A(n15564), .ZN(n15567) );
  XOR2_X1 U16720 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n15567), .Z(SUB_1596_U54) );
  AOI21_X1 U16721 ( .B1(n15570), .B2(n15569), .A(n15568), .ZN(n15571) );
  XOR2_X1 U16722 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n15571), .Z(SUB_1596_U70)
         );
  AOI21_X1 U16723 ( .B1(n15574), .B2(n15573), .A(n15572), .ZN(n15575) );
  XOR2_X1 U16724 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15575), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16725 ( .B1(n15578), .B2(n15577), .A(n15576), .ZN(SUB_1596_U68) );
  OAI21_X1 U16726 ( .B1(n15581), .B2(n15580), .A(n15579), .ZN(n15582) );
  XNOR2_X1 U16727 ( .A(n15582), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16728 ( .B1(n15585), .B2(n15584), .A(n15583), .ZN(n15586) );
  XNOR2_X1 U16729 ( .A(n15586), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16730 ( .A1(n15591), .A2(n15590), .B1(n15591), .B2(n15589), .C1(
        n15588), .C2(n15587), .ZN(SUB_1596_U65) );
  OAI222_X1 U16731 ( .A1(n15596), .A2(n15595), .B1(n15596), .B2(n15594), .C1(
        n15593), .C2(n15592), .ZN(SUB_1596_U64) );
  AOI21_X1 U16732 ( .B1(n15599), .B2(n15598), .A(n15597), .ZN(SUB_1596_U63) );
  AOI21_X1 U16733 ( .B1(n15604), .B2(n15603), .A(n15602), .ZN(n15605) );
  XOR2_X1 U16734 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n15605), .Z(SUB_1596_U57) );
  AOI21_X1 U16735 ( .B1(n15608), .B2(n15607), .A(n15606), .ZN(SUB_1596_U5) );
  AOI22_X1 U16736 ( .A1(n15845), .A2(n15609), .B1(n15832), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n15618) );
  OR2_X1 U16737 ( .A1(n15844), .A2(n15806), .ZN(n15614) );
  INV_X1 U16738 ( .A(n15610), .ZN(n15611) );
  NAND2_X1 U16739 ( .A1(n15614), .A2(n15611), .ZN(n15612) );
  MUX2_X1 U16740 ( .A(n15612), .B(n15822), .S(P3_IR_REG_0__SCAN_IN), .Z(n15616) );
  OAI21_X1 U16741 ( .B1(n15614), .B2(n15845), .A(n15613), .ZN(n15615) );
  AND2_X1 U16742 ( .A1(n15616), .A2(n15615), .ZN(n15617) );
  OAI211_X1 U16743 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n15619), .A(n15618), .B(
        n15617), .ZN(P3_U3182) );
  AOI21_X1 U16744 ( .B1(n15622), .B2(n15621), .A(n15620), .ZN(n15637) );
  INV_X1 U16745 ( .A(n15623), .ZN(n15624) );
  NAND3_X1 U16746 ( .A1(n15626), .A2(n15625), .A3(n15624), .ZN(n15627) );
  AOI21_X1 U16747 ( .B1(n15645), .B2(n15627), .A(n15840), .ZN(n15632) );
  AOI21_X1 U16748 ( .B1(n15832), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n15628), .ZN(
        n15629) );
  OAI21_X1 U16749 ( .B1(n15822), .B2(n15630), .A(n15629), .ZN(n15631) );
  NOR2_X1 U16750 ( .A1(n15632), .A2(n15631), .ZN(n15636) );
  XNOR2_X1 U16751 ( .A(n15633), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n15634) );
  NAND2_X1 U16752 ( .A1(n15844), .A2(n15634), .ZN(n15635) );
  OAI211_X1 U16753 ( .C1(n15637), .C2(n15830), .A(n15636), .B(n15635), .ZN(
        P3_U3185) );
  AOI21_X1 U16754 ( .B1(n15639), .B2(n7349), .A(n15638), .ZN(n15657) );
  INV_X1 U16755 ( .A(n15832), .ZN(n15772) );
  INV_X1 U16756 ( .A(n15640), .ZN(n15641) );
  OAI21_X1 U16757 ( .B1(n15772), .B2(n10303), .A(n15641), .ZN(n15649) );
  INV_X1 U16758 ( .A(n15642), .ZN(n15643) );
  NAND3_X1 U16759 ( .A1(n15645), .A2(n15644), .A3(n15643), .ZN(n15646) );
  AOI21_X1 U16760 ( .B1(n15647), .B2(n15646), .A(n15840), .ZN(n15648) );
  AOI211_X1 U16761 ( .C1(n15834), .C2(n15650), .A(n15649), .B(n15648), .ZN(
        n15656) );
  AND2_X1 U16762 ( .A1(n15652), .A2(n15651), .ZN(n15653) );
  OAI21_X1 U16763 ( .B1(n15654), .B2(n15653), .A(n15844), .ZN(n15655) );
  OAI211_X1 U16764 ( .C1(n15657), .C2(n15830), .A(n15656), .B(n15655), .ZN(
        P3_U3186) );
  AOI21_X1 U16765 ( .B1(n15660), .B2(n15659), .A(n15658), .ZN(n15674) );
  OAI21_X1 U16766 ( .B1(n15663), .B2(n15662), .A(n15661), .ZN(n15665) );
  AOI22_X1 U16767 ( .A1(n15665), .A2(n15806), .B1(n15664), .B2(n15834), .ZN(
        n15666) );
  INV_X1 U16768 ( .A(n15666), .ZN(n15667) );
  AOI211_X1 U16769 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n15832), .A(n15668), .B(
        n15667), .ZN(n15673) );
  OAI21_X1 U16770 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n15670), .A(n15669), .ZN(
        n15671) );
  NAND2_X1 U16771 ( .A1(n15671), .A2(n15844), .ZN(n15672) );
  OAI211_X1 U16772 ( .C1(n15674), .C2(n15830), .A(n15673), .B(n15672), .ZN(
        P3_U3187) );
  AOI21_X1 U16773 ( .B1(n15677), .B2(n15676), .A(n15675), .ZN(n15693) );
  INV_X1 U16774 ( .A(n15678), .ZN(n15680) );
  NAND2_X1 U16775 ( .A1(n15680), .A2(n15679), .ZN(n15681) );
  XNOR2_X1 U16776 ( .A(n15682), .B(n15681), .ZN(n15684) );
  OAI22_X1 U16777 ( .A1(n15684), .A2(n15840), .B1(n15683), .B2(n15822), .ZN(
        n15685) );
  AOI211_X1 U16778 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n15832), .A(n15686), .B(
        n15685), .ZN(n15692) );
  OAI21_X1 U16779 ( .B1(n15689), .B2(n15688), .A(n15687), .ZN(n15690) );
  NAND2_X1 U16780 ( .A1(n15690), .A2(n15844), .ZN(n15691) );
  OAI211_X1 U16781 ( .C1(n15693), .C2(n15830), .A(n15692), .B(n15691), .ZN(
        P3_U3188) );
  AOI21_X1 U16782 ( .B1(n7338), .B2(n15695), .A(n15694), .ZN(n15709) );
  OAI21_X1 U16783 ( .B1(n15698), .B2(n15697), .A(n15696), .ZN(n15699) );
  AND2_X1 U16784 ( .A1(n15699), .A2(n15844), .ZN(n15700) );
  AOI211_X1 U16785 ( .C1(P3_ADDR_REG_10__SCAN_IN), .C2(n15832), .A(n15701), 
        .B(n15700), .ZN(n15708) );
  OAI21_X1 U16786 ( .B1(n15704), .B2(n15703), .A(n15702), .ZN(n15706) );
  AOI22_X1 U16787 ( .A1(n15706), .A2(n15806), .B1(n15705), .B2(n15834), .ZN(
        n15707) );
  OAI211_X1 U16788 ( .C1(n15709), .C2(n15830), .A(n15708), .B(n15707), .ZN(
        P3_U3192) );
  AOI21_X1 U16789 ( .B1(n15712), .B2(n15711), .A(n15710), .ZN(n15725) );
  XNOR2_X1 U16790 ( .A(n15714), .B(n15713), .ZN(n15723) );
  OAI21_X1 U16791 ( .B1(n15716), .B2(P3_REG1_REG_11__SCAN_IN), .A(n15715), 
        .ZN(n15717) );
  NAND2_X1 U16792 ( .A1(n15717), .A2(n15844), .ZN(n15720) );
  AOI21_X1 U16793 ( .B1(n15832), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n15718), 
        .ZN(n15719) );
  OAI211_X1 U16794 ( .C1(n15822), .C2(n15721), .A(n15720), .B(n15719), .ZN(
        n15722) );
  AOI21_X1 U16795 ( .B1(n15806), .B2(n15723), .A(n15722), .ZN(n15724) );
  OAI21_X1 U16796 ( .B1(n15725), .B2(n15830), .A(n15724), .ZN(P3_U3193) );
  AOI21_X1 U16797 ( .B1(n15728), .B2(n15727), .A(n15726), .ZN(n15744) );
  XNOR2_X1 U16798 ( .A(n15730), .B(n15729), .ZN(n15741) );
  OAI21_X1 U16799 ( .B1(n15733), .B2(n15732), .A(n15731), .ZN(n15734) );
  NAND2_X1 U16800 ( .A1(n15734), .A2(n15844), .ZN(n15740) );
  AOI21_X1 U16801 ( .B1(n15832), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n15735), 
        .ZN(n15736) );
  OAI21_X1 U16802 ( .B1(n15822), .B2(n15737), .A(n15736), .ZN(n15738) );
  INV_X1 U16803 ( .A(n15738), .ZN(n15739) );
  OAI211_X1 U16804 ( .C1(n15741), .C2(n15840), .A(n15740), .B(n15739), .ZN(
        n15742) );
  INV_X1 U16805 ( .A(n15742), .ZN(n15743) );
  OAI21_X1 U16806 ( .B1(n15744), .B2(n15830), .A(n15743), .ZN(P3_U3194) );
  AOI22_X1 U16807 ( .A1(n15834), .A2(n15745), .B1(n15832), .B2(
        P3_ADDR_REG_13__SCAN_IN), .ZN(n15760) );
  OAI21_X1 U16808 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15747), .A(n15746), 
        .ZN(n15752) );
  OAI21_X1 U16809 ( .B1(n15750), .B2(n15749), .A(n15748), .ZN(n15751) );
  AOI22_X1 U16810 ( .A1(n15752), .A2(n15844), .B1(n15806), .B2(n15751), .ZN(
        n15759) );
  INV_X1 U16811 ( .A(n15753), .ZN(n15758) );
  OAI221_X1 U16812 ( .B1(n15756), .B2(n15755), .C1(n15756), .C2(n15754), .A(
        n15845), .ZN(n15757) );
  NAND4_X1 U16813 ( .A1(n15760), .A2(n15759), .A3(n15758), .A4(n15757), .ZN(
        P3_U3195) );
  INV_X1 U16814 ( .A(n15761), .ZN(n15762) );
  AOI21_X1 U16815 ( .B1(n15764), .B2(n15763), .A(n15762), .ZN(n15781) );
  OAI21_X1 U16816 ( .B1(n15767), .B2(n15766), .A(n15765), .ZN(n15779) );
  INV_X1 U16817 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15773) );
  NAND2_X1 U16818 ( .A1(n15834), .A2(n15768), .ZN(n15771) );
  INV_X1 U16819 ( .A(n15769), .ZN(n15770) );
  OAI211_X1 U16820 ( .C1(n15773), .C2(n15772), .A(n15771), .B(n15770), .ZN(
        n15778) );
  AOI211_X1 U16821 ( .C1(n15776), .C2(n15775), .A(n15840), .B(n15774), .ZN(
        n15777) );
  AOI211_X1 U16822 ( .C1(n15844), .C2(n15779), .A(n15778), .B(n15777), .ZN(
        n15780) );
  OAI21_X1 U16823 ( .B1(n15781), .B2(n15830), .A(n15780), .ZN(P3_U3196) );
  AOI21_X1 U16824 ( .B1(n15784), .B2(n15783), .A(n15782), .ZN(n15797) );
  OAI21_X1 U16825 ( .B1(n15786), .B2(P3_REG1_REG_15__SCAN_IN), .A(n15785), 
        .ZN(n15795) );
  AOI21_X1 U16826 ( .B1(n15832), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n15787), 
        .ZN(n15788) );
  OAI21_X1 U16827 ( .B1(n15822), .B2(n15789), .A(n15788), .ZN(n15794) );
  AOI211_X1 U16828 ( .C1(n15792), .C2(n15791), .A(n15840), .B(n15790), .ZN(
        n15793) );
  AOI211_X1 U16829 ( .C1(n15844), .C2(n15795), .A(n15794), .B(n15793), .ZN(
        n15796) );
  OAI21_X1 U16830 ( .B1(n15797), .B2(n15830), .A(n15796), .ZN(P3_U3197) );
  AOI22_X1 U16831 ( .A1(n15834), .A2(n15798), .B1(n15832), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n15813) );
  OAI21_X1 U16832 ( .B1(n15801), .B2(n15800), .A(n15799), .ZN(n15807) );
  OAI21_X1 U16833 ( .B1(n15804), .B2(n15803), .A(n15802), .ZN(n15805) );
  AOI22_X1 U16834 ( .A1(n15807), .A2(n15806), .B1(n15844), .B2(n15805), .ZN(
        n15812) );
  OAI221_X1 U16835 ( .B1(n7232), .B2(n15809), .C1(n7232), .C2(n15808), .A(
        n15845), .ZN(n15810) );
  NAND4_X1 U16836 ( .A1(n15813), .A2(n15812), .A3(n15811), .A4(n15810), .ZN(
        P3_U3198) );
  AOI21_X1 U16837 ( .B1(n15816), .B2(n15815), .A(n15814), .ZN(n15831) );
  OAI21_X1 U16838 ( .B1(n15818), .B2(P3_REG1_REG_17__SCAN_IN), .A(n15817), 
        .ZN(n15828) );
  AOI21_X1 U16839 ( .B1(n15832), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n15819), 
        .ZN(n15820) );
  OAI21_X1 U16840 ( .B1(n15822), .B2(n15821), .A(n15820), .ZN(n15827) );
  AOI211_X1 U16841 ( .C1(n15825), .C2(n15824), .A(n15840), .B(n15823), .ZN(
        n15826) );
  AOI211_X1 U16842 ( .C1(n15844), .C2(n15828), .A(n15827), .B(n15826), .ZN(
        n15829) );
  OAI21_X1 U16843 ( .B1(n15831), .B2(n15830), .A(n15829), .ZN(P3_U3199) );
  AOI22_X1 U16844 ( .A1(n15834), .A2(n15833), .B1(n15832), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n15851) );
  XNOR2_X1 U16845 ( .A(n15836), .B(n15835), .ZN(n15843) );
  AOI21_X1 U16846 ( .B1(n15839), .B2(n15838), .A(n15837), .ZN(n15841) );
  NOR2_X1 U16847 ( .A1(n15841), .A2(n15840), .ZN(n15842) );
  AOI21_X1 U16848 ( .B1(n15844), .B2(n15843), .A(n15842), .ZN(n15850) );
  OAI221_X1 U16849 ( .B1(n7233), .B2(n15847), .C1(n7233), .C2(n15846), .A(
        n15845), .ZN(n15848) );
  NAND4_X1 U16850 ( .A1(n15851), .A2(n15850), .A3(n15849), .A4(n15848), .ZN(
        P3_U3200) );
  INV_X1 U16851 ( .A(P2_RD_REG_SCAN_IN), .ZN(n15853) );
  OAI221_X1 U16852 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n15853), .C2(n7802), .A(n15852), .ZN(U29) );
  AND3_X1 U16853 ( .A1(n15856), .A2(n15855), .A3(n15854), .ZN(n15857) );
  NOR3_X1 U16854 ( .A1(n15859), .A2(n15858), .A3(n15857), .ZN(n15860) );
  AOI21_X1 U16855 ( .B1(n15862), .B2(n15861), .A(n15860), .ZN(n15871) );
  MUX2_X1 U16856 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11155), .S(n15863), .Z(
        n15866) );
  NAND3_X1 U16857 ( .A1(n15866), .A2(n15865), .A3(n15864), .ZN(n15867) );
  NAND3_X1 U16858 ( .A1(n15869), .A2(n15868), .A3(n15867), .ZN(n15870) );
  AND3_X1 U16859 ( .A1(n15872), .A2(n15871), .A3(n15870), .ZN(n15874) );
  OAI211_X1 U16860 ( .C1(n15876), .C2(n15875), .A(n15874), .B(n15873), .ZN(
        P1_U3247) );
  INV_X1 U16861 ( .A(n15882), .ZN(n15890) );
  OAI21_X1 U16862 ( .B1(n15877), .B2(n16019), .A(n15890), .ZN(n15879) );
  AND2_X1 U16863 ( .A1(n15879), .A2(n15878), .ZN(n15893) );
  INV_X1 U16864 ( .A(n15893), .ZN(n15884) );
  OAI22_X1 U16865 ( .A1(n15882), .A2(n15881), .B1(n15888), .B2(n15880), .ZN(
        n15883) );
  NOR2_X1 U16866 ( .A1(n15884), .A2(n15883), .ZN(n15886) );
  AOI22_X1 U16867 ( .A1(n16141), .A2(n15886), .B1(n15885), .B2(n16140), .ZN(
        P1_U3528) );
  AOI22_X1 U16868 ( .A1(n15984), .A2(n15886), .B1(n8556), .B2(n16142), .ZN(
        P1_U3459) );
  AOI22_X1 U16869 ( .A1(n15887), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n15894), .ZN(n15892) );
  AOI21_X1 U16870 ( .B1(n15936), .B2(n15933), .A(n15888), .ZN(n15889) );
  AOI21_X1 U16871 ( .B1(n15941), .B2(n15890), .A(n15889), .ZN(n15891) );
  OAI211_X1 U16872 ( .C1(n15894), .C2(n15893), .A(n15892), .B(n15891), .ZN(
        P1_U3293) );
  OAI22_X1 U16873 ( .A1(n15898), .A2(n15897), .B1(n15896), .B2(n15895), .ZN(
        n15899) );
  NOR2_X1 U16874 ( .A1(n15900), .A2(n15899), .ZN(n15902) );
  AOI22_X1 U16875 ( .A1(n16189), .A2(n15902), .B1(n15901), .B2(n16188), .ZN(
        P2_U3499) );
  AOI22_X1 U16876 ( .A1(n16192), .A2(n15902), .B1(n10522), .B2(n16190), .ZN(
        P2_U3430) );
  AND3_X1 U16877 ( .A1(n15904), .A2(n15974), .A3(n15903), .ZN(n15907) );
  INV_X1 U16878 ( .A(n15905), .ZN(n15906) );
  AOI211_X1 U16879 ( .C1(n15966), .C2(n15908), .A(n15907), .B(n15906), .ZN(
        n15911) );
  AOI22_X1 U16880 ( .A1(P3_REG2_REG_1__SCAN_IN), .A2(n7188), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(n15909), .ZN(n15910) );
  OAI21_X1 U16881 ( .B1(n7188), .B2(n15911), .A(n15910), .ZN(P3_U3232) );
  INV_X1 U16882 ( .A(n15912), .ZN(n15913) );
  XOR2_X1 U16883 ( .A(n15913), .B(n15920), .Z(n15928) );
  INV_X1 U16884 ( .A(n15928), .ZN(n15940) );
  XNOR2_X1 U16885 ( .A(n15917), .B(n15914), .ZN(n15935) );
  NOR2_X1 U16886 ( .A1(n15916), .A2(n7694), .ZN(n15939) );
  INV_X1 U16887 ( .A(n15939), .ZN(n15919) );
  NAND2_X1 U16888 ( .A1(n16009), .A2(n15917), .ZN(n15918) );
  OAI211_X1 U16889 ( .C1(n16077), .C2(n15935), .A(n15919), .B(n15918), .ZN(
        n15929) );
  AOI211_X1 U16890 ( .C1(n15922), .C2(n10207), .A(n16134), .B(n15921), .ZN(
        n15923) );
  AOI21_X1 U16891 ( .B1(n15925), .B2(n15924), .A(n15923), .ZN(n15926) );
  OAI21_X1 U16892 ( .B1(n15928), .B2(n15927), .A(n15926), .ZN(n15943) );
  AOI211_X1 U16893 ( .C1(n7680), .C2(n15940), .A(n15929), .B(n15943), .ZN(
        n15930) );
  AOI22_X1 U16894 ( .A1(n16141), .A2(n15930), .B1(n11140), .B2(n16140), .ZN(
        P1_U3529) );
  AOI22_X1 U16895 ( .A1(n15984), .A2(n15930), .B1(n8546), .B2(n16142), .ZN(
        P1_U3462) );
  INV_X1 U16896 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n15932) );
  OAI22_X1 U16897 ( .A1(n15942), .A2(n11148), .B1(n15932), .B2(n15931), .ZN(
        n15938) );
  OAI22_X1 U16898 ( .A1(n15936), .A2(n15935), .B1(n15934), .B2(n15933), .ZN(
        n15937) );
  AOI211_X1 U16899 ( .C1(n15939), .C2(n15942), .A(n15938), .B(n15937), .ZN(
        n15945) );
  AOI22_X1 U16900 ( .A1(n15943), .A2(n15942), .B1(n15941), .B2(n15940), .ZN(
        n15944) );
  NAND2_X1 U16901 ( .A1(n15945), .A2(n15944), .ZN(P1_U3292) );
  INV_X1 U16902 ( .A(n15946), .ZN(n15952) );
  OAI21_X1 U16903 ( .B1(n15948), .B2(n16182), .A(n15947), .ZN(n15951) );
  INV_X1 U16904 ( .A(n15949), .ZN(n15950) );
  AOI211_X1 U16905 ( .C1(n16121), .C2(n15952), .A(n15951), .B(n15950), .ZN(
        n15953) );
  AOI22_X1 U16906 ( .A1(n16189), .A2(n15953), .B1(n11058), .B2(n16188), .ZN(
        P2_U3500) );
  AOI22_X1 U16907 ( .A1(n16192), .A2(n15953), .B1(n10530), .B2(n16190), .ZN(
        P2_U3433) );
  OAI21_X1 U16908 ( .B1(n15955), .B2(n15957), .A(n15954), .ZN(n15973) );
  NOR2_X1 U16909 ( .A1(n15970), .A2(n16157), .ZN(n15963) );
  XNOR2_X1 U16910 ( .A(n15956), .B(n15957), .ZN(n15958) );
  OAI222_X1 U16911 ( .A1(n15962), .A2(n15961), .B1(n15960), .B2(n11228), .C1(
        n15959), .C2(n15958), .ZN(n15971) );
  AOI211_X1 U16912 ( .C1(n16160), .C2(n15973), .A(n15963), .B(n15971), .ZN(
        n15965) );
  AOI22_X1 U16913 ( .A1(n16165), .A2(n15965), .B1(n9973), .B2(n9674), .ZN(
        P3_U3461) );
  INV_X1 U16914 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15964) );
  AOI22_X1 U16915 ( .A1(n16169), .A2(n15965), .B1(n15964), .B2(n16166), .ZN(
        P3_U3396) );
  INV_X1 U16916 ( .A(n15966), .ZN(n15969) );
  OAI22_X1 U16917 ( .A1(n15970), .A2(n15969), .B1(n15968), .B2(n15967), .ZN(
        n15972) );
  AOI211_X1 U16918 ( .C1(n15974), .C2(n15973), .A(n15972), .B(n15971), .ZN(
        n15975) );
  AOI22_X1 U16919 ( .A1(n7188), .A2(n9974), .B1(n15975), .B2(n13715), .ZN(
        P3_U3231) );
  INV_X1 U16920 ( .A(n15976), .ZN(n15982) );
  OAI22_X1 U16921 ( .A1(n15978), .A2(n16133), .B1(n16077), .B2(n15977), .ZN(
        n15981) );
  INV_X1 U16922 ( .A(n15979), .ZN(n15980) );
  AOI211_X1 U16923 ( .C1(n15982), .C2(n16139), .A(n15981), .B(n15980), .ZN(
        n15983) );
  AOI22_X1 U16924 ( .A1(n16141), .A2(n15983), .B1(n11141), .B2(n16140), .ZN(
        P1_U3530) );
  AOI22_X1 U16925 ( .A1(n15984), .A2(n15983), .B1(n8566), .B2(n16142), .ZN(
        P1_U3465) );
  INV_X1 U16926 ( .A(n15988), .ZN(n15990) );
  INV_X1 U16927 ( .A(n16103), .ZN(n16055) );
  AOI21_X1 U16928 ( .B1(n15986), .B2(n16107), .A(n15985), .ZN(n15987) );
  OAI21_X1 U16929 ( .B1(n15988), .B2(n16055), .A(n15987), .ZN(n15989) );
  AOI21_X1 U16930 ( .B1(n15990), .B2(n16057), .A(n15989), .ZN(n15992) );
  AOI22_X1 U16931 ( .A1(n16165), .A2(n15992), .B1(n9979), .B2(n9674), .ZN(
        P3_U3462) );
  INV_X1 U16932 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15991) );
  AOI22_X1 U16933 ( .A1(n16169), .A2(n15992), .B1(n15991), .B2(n16166), .ZN(
        P3_U3399) );
  INV_X1 U16934 ( .A(n15993), .ZN(n15998) );
  OAI21_X1 U16935 ( .B1(n15995), .B2(n16182), .A(n15994), .ZN(n15997) );
  AOI211_X1 U16936 ( .C1(n16121), .C2(n15998), .A(n15997), .B(n15996), .ZN(
        n15999) );
  AOI22_X1 U16937 ( .A1(n16189), .A2(n15999), .B1(n10513), .B2(n16188), .ZN(
        P2_U3502) );
  AOI22_X1 U16938 ( .A1(n16192), .A2(n15999), .B1(n10512), .B2(n16190), .ZN(
        P2_U3439) );
  INV_X1 U16939 ( .A(n16003), .ZN(n16005) );
  AOI21_X1 U16940 ( .B1(n16001), .B2(n16107), .A(n16000), .ZN(n16002) );
  OAI21_X1 U16941 ( .B1(n16055), .B2(n16003), .A(n16002), .ZN(n16004) );
  AOI21_X1 U16942 ( .B1(n16005), .B2(n16057), .A(n16004), .ZN(n16007) );
  AOI22_X1 U16943 ( .A1(n16165), .A2(n16007), .B1(n9985), .B2(n9674), .ZN(
        P3_U3463) );
  INV_X1 U16944 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n16006) );
  AOI22_X1 U16945 ( .A1(n16169), .A2(n16007), .B1(n16006), .B2(n16166), .ZN(
        P3_U3402) );
  AND2_X1 U16946 ( .A1(n16009), .A2(n16008), .ZN(n16011) );
  AOI211_X1 U16947 ( .C1(n16013), .C2(n16012), .A(n16011), .B(n16010), .ZN(
        n16014) );
  OAI21_X1 U16948 ( .B1(n16016), .B2(n16015), .A(n16014), .ZN(n16017) );
  AOI21_X1 U16949 ( .B1(n16019), .B2(n16018), .A(n16017), .ZN(n16020) );
  AOI22_X1 U16950 ( .A1(n16141), .A2(n16020), .B1(n11142), .B2(n16140), .ZN(
        P1_U3532) );
  AOI22_X1 U16951 ( .A1(n15984), .A2(n16020), .B1(n8610), .B2(n16142), .ZN(
        P1_U3471) );
  INV_X1 U16952 ( .A(n16024), .ZN(n16026) );
  AOI21_X1 U16953 ( .B1(n16022), .B2(n16107), .A(n16021), .ZN(n16023) );
  OAI21_X1 U16954 ( .B1(n16055), .B2(n16024), .A(n16023), .ZN(n16025) );
  AOI21_X1 U16955 ( .B1(n16026), .B2(n16057), .A(n16025), .ZN(n16029) );
  INV_X1 U16956 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n16027) );
  AOI22_X1 U16957 ( .A1(n16165), .A2(n16029), .B1(n16027), .B2(n9674), .ZN(
        P3_U3464) );
  INV_X1 U16958 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n16028) );
  AOI22_X1 U16959 ( .A1(n16169), .A2(n16029), .B1(n16028), .B2(n16166), .ZN(
        P3_U3405) );
  INV_X1 U16960 ( .A(n16030), .ZN(n16034) );
  OAI21_X1 U16961 ( .B1(n16032), .B2(n16157), .A(n16031), .ZN(n16033) );
  AOI21_X1 U16962 ( .B1(n16034), .B2(n16160), .A(n16033), .ZN(n16036) );
  AOI22_X1 U16963 ( .A1(n16165), .A2(n16036), .B1(n9995), .B2(n9674), .ZN(
        P3_U3465) );
  INV_X1 U16964 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n16035) );
  AOI22_X1 U16965 ( .A1(n16169), .A2(n16036), .B1(n16035), .B2(n16166), .ZN(
        P3_U3408) );
  INV_X1 U16966 ( .A(n16037), .ZN(n16046) );
  OAI22_X1 U16967 ( .A1(n16041), .A2(n16040), .B1(n16039), .B2(n16038), .ZN(
        n16042) );
  AOI21_X1 U16968 ( .B1(n16147), .B2(n16043), .A(n16042), .ZN(n16044) );
  OAI21_X1 U16969 ( .B1(n16046), .B2(n16045), .A(n16044), .ZN(n16047) );
  AOI21_X1 U16970 ( .B1(n16151), .B2(n16048), .A(n16047), .ZN(n16049) );
  OAI21_X1 U16971 ( .B1(n16156), .B2(n16050), .A(n16049), .ZN(P2_U3259) );
  INV_X1 U16972 ( .A(n16054), .ZN(n16058) );
  AOI21_X1 U16973 ( .B1(n16052), .B2(n16107), .A(n16051), .ZN(n16053) );
  OAI21_X1 U16974 ( .B1(n16055), .B2(n16054), .A(n16053), .ZN(n16056) );
  AOI21_X1 U16975 ( .B1(n16058), .B2(n16057), .A(n16056), .ZN(n16061) );
  INV_X1 U16976 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n16059) );
  AOI22_X1 U16977 ( .A1(n16165), .A2(n16061), .B1(n16059), .B2(n9674), .ZN(
        P3_U3466) );
  INV_X1 U16978 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n16060) );
  AOI22_X1 U16979 ( .A1(n16169), .A2(n16061), .B1(n16060), .B2(n16166), .ZN(
        P3_U3411) );
  OAI21_X1 U16980 ( .B1(n16063), .B2(n16182), .A(n16062), .ZN(n16065) );
  AOI211_X1 U16981 ( .C1(n16121), .C2(n16066), .A(n16065), .B(n16064), .ZN(
        n16068) );
  AOI22_X1 U16982 ( .A1(n16189), .A2(n16068), .B1(n11068), .B2(n16188), .ZN(
        P2_U3506) );
  INV_X1 U16983 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n16067) );
  AOI22_X1 U16984 ( .A1(n16192), .A2(n16068), .B1(n16067), .B2(n16190), .ZN(
        P2_U3451) );
  NOR2_X1 U16985 ( .A1(n16069), .A2(n16157), .ZN(n16071) );
  AOI211_X1 U16986 ( .C1(n16160), .C2(n16072), .A(n16071), .B(n16070), .ZN(
        n16075) );
  AOI22_X1 U16987 ( .A1(n16165), .A2(n16075), .B1(n16073), .B2(n9674), .ZN(
        P3_U3467) );
  INV_X1 U16988 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U16989 ( .A1(n16169), .A2(n16075), .B1(n16074), .B2(n16166), .ZN(
        P3_U3414) );
  OAI22_X1 U16990 ( .A1(n16078), .A2(n16077), .B1(n8318), .B2(n16133), .ZN(
        n16080) );
  AOI211_X1 U16991 ( .C1(n7680), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        n16082) );
  AOI22_X1 U16992 ( .A1(n16141), .A2(n16082), .B1(n11291), .B2(n16140), .ZN(
        P1_U3536) );
  AOI22_X1 U16993 ( .A1(n15984), .A2(n16082), .B1(n8675), .B2(n16142), .ZN(
        P1_U3483) );
  INV_X1 U16994 ( .A(n16083), .ZN(n16087) );
  NOR2_X1 U16995 ( .A1(n16084), .A2(n16157), .ZN(n16086) );
  AOI211_X1 U16996 ( .C1(n16087), .C2(n16103), .A(n16086), .B(n16085), .ZN(
        n16090) );
  INV_X1 U16997 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n16088) );
  AOI22_X1 U16998 ( .A1(n16165), .A2(n16090), .B1(n16088), .B2(n9674), .ZN(
        P3_U3468) );
  INV_X1 U16999 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16089) );
  AOI22_X1 U17000 ( .A1(n16169), .A2(n16090), .B1(n16089), .B2(n16166), .ZN(
        P3_U3417) );
  INV_X1 U17001 ( .A(n16091), .ZN(n16095) );
  OAI21_X1 U17002 ( .B1(n7756), .B2(n16182), .A(n16092), .ZN(n16094) );
  AOI211_X1 U17003 ( .C1(n16121), .C2(n16095), .A(n16094), .B(n16093), .ZN(
        n16097) );
  AOI22_X1 U17004 ( .A1(n16189), .A2(n16097), .B1(n10478), .B2(n16188), .ZN(
        P2_U3508) );
  INV_X1 U17005 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n16096) );
  AOI22_X1 U17006 ( .A1(n16192), .A2(n16097), .B1(n16096), .B2(n16190), .ZN(
        P2_U3457) );
  INV_X1 U17007 ( .A(n16098), .ZN(n16102) );
  NOR2_X1 U17008 ( .A1(n16099), .A2(n16157), .ZN(n16101) );
  AOI211_X1 U17009 ( .C1(n16103), .C2(n16102), .A(n16101), .B(n16100), .ZN(
        n16106) );
  AOI22_X1 U17010 ( .A1(n16165), .A2(n16106), .B1(n16104), .B2(n9674), .ZN(
        P3_U3469) );
  INV_X1 U17011 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n16105) );
  AOI22_X1 U17012 ( .A1(n16169), .A2(n16106), .B1(n16105), .B2(n16166), .ZN(
        P3_U3420) );
  AOI22_X1 U17013 ( .A1(n16109), .A2(n16160), .B1(n16108), .B2(n16107), .ZN(
        n16111) );
  AND2_X1 U17014 ( .A1(n16111), .A2(n16110), .ZN(n16114) );
  INV_X1 U17015 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n16112) );
  AOI22_X1 U17016 ( .A1(n16165), .A2(n16114), .B1(n16112), .B2(n9674), .ZN(
        P3_U3470) );
  INV_X1 U17017 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16113) );
  AOI22_X1 U17018 ( .A1(n16169), .A2(n16114), .B1(n16113), .B2(n16166), .ZN(
        P3_U3423) );
  INV_X1 U17019 ( .A(n16115), .ZN(n16120) );
  OAI21_X1 U17020 ( .B1(n16117), .B2(n16182), .A(n16116), .ZN(n16119) );
  AOI211_X1 U17021 ( .C1(n16121), .C2(n16120), .A(n16119), .B(n16118), .ZN(
        n16123) );
  AOI22_X1 U17022 ( .A1(n16189), .A2(n16123), .B1(n11279), .B2(n16188), .ZN(
        P2_U3510) );
  INV_X1 U17023 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n16122) );
  AOI22_X1 U17024 ( .A1(n16192), .A2(n16123), .B1(n16122), .B2(n16190), .ZN(
        P2_U3463) );
  NOR2_X1 U17025 ( .A1(n16124), .A2(n16157), .ZN(n16126) );
  AOI211_X1 U17026 ( .C1(n16160), .C2(n16127), .A(n16126), .B(n16125), .ZN(
        n16130) );
  INV_X1 U17027 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n16128) );
  AOI22_X1 U17028 ( .A1(n16165), .A2(n16130), .B1(n16128), .B2(n9674), .ZN(
        P3_U3472) );
  INV_X1 U17029 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n16129) );
  AOI22_X1 U17030 ( .A1(n16169), .A2(n16130), .B1(n16129), .B2(n16166), .ZN(
        P3_U3429) );
  OAI211_X1 U17031 ( .C1(n8322), .C2(n16133), .A(n16132), .B(n16131), .ZN(
        n16137) );
  NOR2_X1 U17032 ( .A1(n16135), .A2(n16134), .ZN(n16136) );
  AOI211_X1 U17033 ( .C1(n16139), .C2(n16138), .A(n16137), .B(n16136), .ZN(
        n16143) );
  AOI22_X1 U17034 ( .A1(n16141), .A2(n16143), .B1(n11810), .B2(n16140), .ZN(
        P1_U3541) );
  AOI22_X1 U17035 ( .A1(n15984), .A2(n16143), .B1(n8764), .B2(n16142), .ZN(
        P1_U3498) );
  INV_X1 U17036 ( .A(n16144), .ZN(n16145) );
  AOI222_X1 U17037 ( .A1(n16148), .A2(n16147), .B1(P2_REG2_REG_13__SCAN_IN), 
        .B2(n16156), .C1(n16146), .C2(n16145), .ZN(n16154) );
  AOI22_X1 U17038 ( .A1(n16152), .A2(n16151), .B1(n16150), .B2(n16149), .ZN(
        n16153) );
  OAI211_X1 U17039 ( .C1(n16156), .C2(n16155), .A(n16154), .B(n16153), .ZN(
        P2_U3252) );
  NOR2_X1 U17040 ( .A1(n16158), .A2(n16157), .ZN(n16159) );
  AOI21_X1 U17041 ( .B1(n16161), .B2(n16160), .A(n16159), .ZN(n16162) );
  AND2_X1 U17042 ( .A1(n16163), .A2(n16162), .ZN(n16168) );
  AOI22_X1 U17043 ( .A1(n16165), .A2(n16168), .B1(n16164), .B2(n9674), .ZN(
        P3_U3473) );
  INV_X1 U17044 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n16167) );
  AOI22_X1 U17045 ( .A1(n16169), .A2(n16168), .B1(n16167), .B2(n16166), .ZN(
        P3_U3432) );
  INV_X1 U17046 ( .A(n16170), .ZN(n16171) );
  AOI21_X1 U17047 ( .B1(n16173), .B2(n16172), .A(n16171), .ZN(n16174) );
  INV_X1 U17048 ( .A(n16174), .ZN(n16175) );
  AOI222_X1 U17049 ( .A1(n7185), .A2(n16177), .B1(n16176), .B2(n16197), .C1(
        n16175), .C2(n16195), .ZN(n16179) );
  OAI211_X1 U17050 ( .C1(n16203), .C2(n16180), .A(n16179), .B(n16178), .ZN(
        P1_U3215) );
  OAI21_X1 U17051 ( .B1(n16183), .B2(n16182), .A(n16181), .ZN(n16185) );
  AOI211_X1 U17052 ( .C1(n16187), .C2(n16186), .A(n16185), .B(n16184), .ZN(
        n16191) );
  AOI22_X1 U17053 ( .A1(n16189), .A2(n16191), .B1(n12425), .B2(n16188), .ZN(
        P2_U3513) );
  AOI22_X1 U17054 ( .A1(n16192), .A2(n16191), .B1(n10666), .B2(n16190), .ZN(
        P2_U3472) );
  OAI21_X1 U17055 ( .B1(n16194), .B2(n16193), .A(n14632), .ZN(n16196) );
  AOI222_X1 U17056 ( .A1(n7185), .A2(n16199), .B1(n16198), .B2(n16197), .C1(
        n16196), .C2(n16195), .ZN(n16201) );
  OAI211_X1 U17057 ( .C1(n16203), .C2(n16202), .A(n16201), .B(n16200), .ZN(
        P1_U3226) );
  AOI21_X1 U17058 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16204) );
  OAI21_X1 U17059 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16204), 
        .ZN(U28) );
  CLKBUF_X1 U7300 ( .A(n9138), .Z(n9601) );
  CLKBUF_X1 U7302 ( .A(n10416), .Z(n10447) );
  XNOR2_X1 U7336 ( .A(n14432), .B(n14434), .ZN(n14732) );
  CLKBUF_X2 U9052 ( .A(n9598), .Z(n7187) );
  CLKBUF_X1 U15841 ( .A(n10040), .Z(n15162) );
endmodule

