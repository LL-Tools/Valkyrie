

module b22_C_AntiSAT_k_256_9 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617;

  INV_X4 U7390 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  BUF_X1 U7391 ( .A(n10208), .Z(n13459) );
  CLKBUF_X2 U7392 ( .A(n11811), .Z(n12322) );
  BUF_X1 U7393 ( .A(n7865), .Z(n6644) );
  INV_X1 U7394 ( .A(n9601), .ZN(n11490) );
  BUF_X2 U7395 ( .A(n11619), .Z(n6652) );
  AOI21_X1 U7396 ( .B1(n12032), .B2(n8779), .A(n8778), .ZN(n9949) );
  NAND4_X2 U7397 ( .A1(n8341), .A2(n8340), .A3(n6683), .A4(n8339), .ZN(n9350)
         );
  OAI21_X1 U7398 ( .B1(n9446), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9445) );
  AND2_X1 U7399 ( .A1(n11486), .A2(n7033), .ZN(n11488) );
  INV_X1 U7400 ( .A(n11693), .ZN(n11699) );
  OR2_X1 U7401 ( .A1(n11586), .A2(n11585), .ZN(n11670) );
  OAI22_X1 U7402 ( .A1(n11083), .A2(n8117), .B1(n11230), .B2(n14535), .ZN(
        n11150) );
  NAND2_X1 U7403 ( .A1(n9645), .A2(n11759), .ZN(n9850) );
  AND2_X1 U7404 ( .A1(n9601), .A2(n9468), .ZN(n11619) );
  INV_X1 U7405 ( .A(n9850), .ZN(n11995) );
  INV_X1 U7406 ( .A(n10936), .ZN(n10208) );
  INV_X1 U7407 ( .A(n7741), .ZN(n12467) );
  NAND2_X1 U7408 ( .A1(n8116), .A2(n8115), .ZN(n11083) );
  INV_X1 U7409 ( .A(n8911), .ZN(n15124) );
  NAND2_X1 U7410 ( .A1(n9580), .A2(n11757), .ZN(n11759) );
  NAND2_X1 U7411 ( .A1(n8772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U7412 ( .A1(n10563), .A2(n10562), .ZN(n10651) );
  MUX2_X1 U7413 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13694), .S(n9601), .Z(n13654)
         );
  NOR2_X1 U7414 ( .A1(n11212), .A2(n10966), .ZN(n7514) );
  NAND2_X1 U7415 ( .A1(n8411), .A2(n8410), .ZN(n12052) );
  NAND2_X1 U7416 ( .A1(n14173), .A2(n8634), .ZN(n14150) );
  INV_X1 U7417 ( .A(n11968), .ZN(n9017) );
  CLKBUF_X3 U7418 ( .A(n8235), .Z(n6643) );
  INV_X1 U7419 ( .A(n14114), .ZN(n8775) );
  AND2_X1 U7420 ( .A1(n8222), .A2(n8230), .ZN(n6642) );
  INV_X2 U7421 ( .A(n6655), .ZN(n11692) );
  NAND2_X2 U7422 ( .A1(n14174), .A2(n8633), .ZN(n14173) );
  INV_X1 U7423 ( .A(n6883), .ZN(n7078) );
  OAI21_X1 U7424 ( .B1(n9055), .B2(P2_IR_REG_27__SCAN_IN), .A(n6674), .ZN(
        n7055) );
  NAND2_X1 U7425 ( .A1(n8890), .A2(n8891), .ZN(n9055) );
  NAND2_X2 U7426 ( .A1(n11780), .A2(n7492), .ZN(n7491) );
  NAND2_X2 U7427 ( .A1(n11249), .A2(n11248), .ZN(n11780) );
  AND2_X1 U7428 ( .A1(n7705), .A2(n7704), .ZN(n7865) );
  XNOR2_X2 U7429 ( .A(n7701), .B(n7700), .ZN(n7706) );
  INV_X1 U7430 ( .A(n11324), .ZN(n13179) );
  AND3_X2 U7431 ( .A1(n9564), .A2(n9565), .A3(n9563), .ZN(n11324) );
  XNOR2_X2 U7432 ( .A(n7670), .B(n7669), .ZN(n11319) );
  OAI21_X2 U7433 ( .B1(n13203), .B2(n7339), .A(n7337), .ZN(n13170) );
  NAND2_X2 U7434 ( .A1(n11971), .A2(n11970), .ZN(n13203) );
  NAND2_X1 U7435 ( .A1(n13161), .A2(n7304), .ZN(n7306) );
  INV_X1 U7436 ( .A(n11323), .ZN(n11337) );
  NAND4_X2 U7437 ( .A1(n9467), .A2(n7407), .A3(n7408), .A4(n7406), .ZN(n11331)
         );
  MUX2_X2 U7438 ( .A(n7676), .B(n7675), .S(P1_ADDR_REG_19__SCAN_IN), .Z(n8235)
         );
  INV_X1 U7439 ( .A(n9468), .ZN(n9560) );
  BUF_X4 U7440 ( .A(n7865), .Z(n6645) );
  NAND2_X2 U7441 ( .A1(n7514), .A2(n9017), .ZN(n9225) );
  OAI22_X2 U7442 ( .A1(n11386), .A2(n7424), .B1(n7423), .B2(n11387), .ZN(
        n11395) );
  NOR2_X2 U7443 ( .A1(n10132), .A2(n10131), .ZN(n10136) );
  NOR2_X2 U7444 ( .A1(n9854), .A2(n9853), .ZN(n10132) );
  XNOR2_X2 U7445 ( .A(n7495), .B(n7494), .ZN(n13812) );
  NAND2_X2 U7446 ( .A1(n7491), .A2(n6739), .ZN(n7495) );
  OAI21_X2 U7447 ( .B1(n8624), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8625) );
  XNOR2_X2 U7448 ( .A(n8774), .B(n8773), .ZN(n12025) );
  INV_X1 U7449 ( .A(n6642), .ZN(n6646) );
  INV_X4 U7450 ( .A(n6642), .ZN(n6647) );
  OAI21_X2 U7451 ( .B1(n10990), .B2(n12234), .A(n8576), .ZN(n11096) );
  AOI21_X1 U7452 ( .B1(n11719), .B2(n11718), .A(n11717), .ZN(n11761) );
  OAI22_X1 U7453 ( .A1(n11488), .A2(n11487), .B1(n11486), .B2(n7033), .ZN(
        n11503) );
  OAI21_X1 U7454 ( .B1(n7430), .B2(n11429), .A(n7431), .ZN(n11440) );
  OR2_X1 U7455 ( .A1(n11428), .A2(n7432), .ZN(n7430) );
  NAND2_X1 U7456 ( .A1(n10434), .A2(n7510), .ZN(n7509) );
  INV_X4 U7457 ( .A(n11692), .ZN(n11693) );
  CLKBUF_X3 U7458 ( .A(n9850), .Z(n12012) );
  INV_X4 U7459 ( .A(n11380), .ZN(n11716) );
  AND2_X1 U7460 ( .A1(n8370), .A2(n6713), .ZN(n14714) );
  INV_X1 U7461 ( .A(n7719), .ZN(n7741) );
  NAND2_X1 U7462 ( .A1(n12267), .A2(n13683), .ZN(n9466) );
  CLKBUF_X2 U7463 ( .A(n8381), .Z(n8626) );
  BUF_X2 U7464 ( .A(n9580), .Z(n6656) );
  CLKBUF_X2 U7465 ( .A(n8819), .Z(n6650) );
  CLKBUF_X2 U7466 ( .A(n8819), .Z(n6651) );
  NAND2_X1 U7467 ( .A1(n8222), .A2(n8221), .ZN(n8819) );
  AOI21_X1 U7468 ( .B1(n14006), .B2(n14144), .A(n14005), .ZN(n14202) );
  NAND2_X1 U7469 ( .A1(n13263), .A2(n7326), .ZN(n13148) );
  MUX2_X1 U7470 ( .A(n15375), .B(n13078), .S(n15197), .Z(n13079) );
  NOR2_X1 U7471 ( .A1(n14007), .A2(n8749), .ZN(n8760) );
  NOR2_X1 U7472 ( .A1(n14008), .A2(n14009), .ZN(n14007) );
  NAND2_X1 U7473 ( .A1(n14020), .A2(n6826), .ZN(n14008) );
  OAI21_X1 U7474 ( .B1(n11951), .B2(n13372), .A(n13521), .ZN(n13368) );
  OAI21_X1 U7475 ( .B1(n11789), .B2(n7479), .A(n7478), .ZN(n7476) );
  OR2_X1 U7476 ( .A1(n11990), .A2(n11989), .ZN(n7562) );
  NAND2_X1 U7477 ( .A1(n10838), .A2(n10837), .ZN(n10842) );
  NAND2_X1 U7478 ( .A1(n8661), .A2(n8660), .ZN(n14303) );
  NAND2_X1 U7479 ( .A1(n7509), .A2(n6762), .ZN(n10838) );
  INV_X1 U7480 ( .A(n12703), .ZN(n12412) );
  OR2_X1 U7481 ( .A1(n11016), .A2(n11738), .ZN(n11166) );
  OR2_X1 U7482 ( .A1(n8289), .A2(n15493), .ZN(n7403) );
  NAND2_X2 U7483 ( .A1(n11065), .A2(n11064), .ZN(n13637) );
  NAND2_X1 U7484 ( .A1(n10935), .A2(n10934), .ZN(n13643) );
  NAND2_X1 U7485 ( .A1(n8550), .A2(n8549), .ZN(n14584) );
  NOR2_X1 U7486 ( .A1(n7024), .A2(n7023), .ZN(n7022) );
  OR2_X1 U7487 ( .A1(n7823), .A2(n10788), .ZN(n7001) );
  XNOR2_X1 U7488 ( .A(n6840), .B(n8564), .ZN(n11062) );
  AOI21_X1 U7489 ( .B1(n8562), .B2(n8561), .A(n8560), .ZN(n6840) );
  NAND2_X1 U7490 ( .A1(n7373), .A2(n7372), .ZN(n8599) );
  NAND2_X1 U7491 ( .A1(n10751), .A2(n10750), .ZN(n14558) );
  NAND2_X1 U7492 ( .A1(n9388), .A2(n9387), .ZN(n9805) );
  AND2_X1 U7493 ( .A1(n11958), .A2(n9381), .ZN(n9388) );
  NAND2_X1 U7494 ( .A1(n8277), .A2(n8276), .ZN(n8559) );
  NAND2_X1 U7495 ( .A1(n10518), .A2(n10517), .ZN(n14918) );
  NAND2_X1 U7496 ( .A1(n10266), .A2(n10265), .ZN(n11417) );
  NAND2_X1 U7497 ( .A1(n10204), .A2(n10203), .ZN(n11411) );
  NAND2_X1 U7498 ( .A1(n7385), .A2(n7383), .ZN(n8499) );
  NAND2_X1 U7499 ( .A1(n8428), .A2(n8427), .ZN(n12056) );
  INV_X2 U7500 ( .A(n15144), .ZN(n15146) );
  NAND2_X1 U7501 ( .A1(n8262), .A2(n8261), .ZN(n8467) );
  XNOR2_X1 U7502 ( .A(n8454), .B(n8453), .ZN(n10201) );
  INV_X1 U7503 ( .A(n9731), .ZN(n12212) );
  NAND2_X1 U7504 ( .A1(n9668), .A2(n9667), .ZN(n14874) );
  AND2_X1 U7505 ( .A1(n12565), .A2(n12571), .ZN(n12500) );
  AND2_X1 U7506 ( .A1(n12549), .A2(n12550), .ZN(n12507) );
  AND2_X1 U7507 ( .A1(n9604), .A2(n9603), .ZN(n11354) );
  NAND4_X1 U7509 ( .A1(n7716), .A2(n7715), .A3(n7714), .A4(n7713), .ZN(n15125)
         );
  BUF_X1 U7510 ( .A(n8356), .Z(n12034) );
  AND2_X1 U7511 ( .A1(n13839), .A2(n14714), .ZN(n12039) );
  NOR2_X1 U7512 ( .A1(n13839), .A2(n14714), .ZN(n12038) );
  NAND4_X1 U7513 ( .A1(n9623), .A2(n9622), .A3(n9621), .A4(n9620), .ZN(n13299)
         );
  INV_X2 U7514 ( .A(n11836), .ZN(n12323) );
  INV_X2 U7515 ( .A(n9657), .ZN(n10936) );
  NOR2_X1 U7516 ( .A1(n11834), .A2(n14176), .ZN(n11811) );
  INV_X2 U7517 ( .A(n7741), .ZN(n8138) );
  INV_X1 U7518 ( .A(n11836), .ZN(n6648) );
  NAND2_X1 U7519 ( .A1(n8777), .A2(n9995), .ZN(n12032) );
  NAND2_X1 U7520 ( .A1(n11756), .A2(n11690), .ZN(n13521) );
  NAND4_X1 U7521 ( .A1(n9578), .A2(n9577), .A3(n9576), .A4(n9575), .ZN(n11346)
         );
  AND2_X1 U7522 ( .A1(n11750), .A2(n9569), .ZN(n13653) );
  CLKBUF_X3 U7523 ( .A(n9605), .Z(n11658) );
  AND2_X1 U7524 ( .A1(n9225), .A2(n9962), .ZN(n9345) );
  NAND2_X2 U7525 ( .A1(n9491), .A2(n9560), .ZN(n8089) );
  AND2_X1 U7526 ( .A1(n7706), .A2(n13144), .ZN(n7719) );
  INV_X1 U7527 ( .A(n7706), .ZN(n7705) );
  INV_X1 U7528 ( .A(n13838), .ZN(n6649) );
  INV_X2 U7529 ( .A(n9466), .ZN(n11686) );
  NAND4_X2 U7530 ( .A1(n8361), .A2(n8360), .A3(n8359), .A4(n8358), .ZN(n13839)
         );
  INV_X1 U7531 ( .A(n9581), .ZN(n9569) );
  NAND4_X2 U7532 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), .ZN(n13841)
         );
  INV_X2 U7533 ( .A(n12693), .ZN(n12758) );
  NAND2_X1 U7534 ( .A1(n8767), .A2(n8772), .ZN(n12206) );
  NAND2_X1 U7535 ( .A1(n9456), .A2(n13683), .ZN(n11689) );
  INV_X1 U7536 ( .A(n12025), .ZN(n14335) );
  NAND2_X2 U7537 ( .A1(n11319), .A2(n9517), .ZN(n9491) );
  NAND2_X1 U7538 ( .A1(n8833), .A2(n8832), .ZN(n11968) );
  NAND2_X1 U7539 ( .A1(n13138), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7701) );
  XNOR2_X1 U7540 ( .A(n7703), .B(P3_IR_REG_29__SCAN_IN), .ZN(n7704) );
  XNOR2_X1 U7541 ( .A(n9447), .B(P2_IR_REG_19__SCAN_IN), .ZN(n11748) );
  MUX2_X1 U7542 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9046), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n9048) );
  NAND2_X1 U7543 ( .A1(n8837), .A2(n8836), .ZN(n11212) );
  INV_X1 U7544 ( .A(n10649), .ZN(n12205) );
  MUX2_X1 U7545 ( .A(n8764), .B(P1_IR_REG_31__SCAN_IN), .S(n8765), .Z(n8767)
         );
  OR2_X1 U7546 ( .A1(n6646), .A2(n9999), .ZN(n8340) );
  NAND2_X2 U7547 ( .A1(n8220), .A2(n8230), .ZN(n12179) );
  XNOR2_X1 U7548 ( .A(n8839), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U7549 ( .A1(n8837), .A2(n8828), .ZN(n8833) );
  NAND2_X1 U7550 ( .A1(n8771), .A2(n8770), .ZN(n10649) );
  OR2_X1 U7551 ( .A1(n7702), .A2(n7699), .ZN(n13138) );
  MUX2_X1 U7552 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9449), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n9451) );
  OAI21_X1 U7553 ( .B1(n7702), .B2(P3_IR_REG_28__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7703) );
  OR2_X1 U7554 ( .A1(n9053), .A2(n9689), .ZN(n9046) );
  NAND2_X1 U7555 ( .A1(n8841), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8839) );
  INV_X1 U7556 ( .A(n8221), .ZN(n8230) );
  OR2_X1 U7557 ( .A1(n8834), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n8837) );
  AND2_X2 U7558 ( .A1(n8220), .A2(n8221), .ZN(n12178) );
  NAND2_X1 U7559 ( .A1(n7593), .A2(n7118), .ZN(n7702) );
  XNOR2_X1 U7560 ( .A(n9057), .B(n9056), .ZN(n13691) );
  NAND2_X2 U7561 ( .A1(n9560), .A2(P1_U3086), .ZN(n14330) );
  NOR2_X1 U7562 ( .A1(n8831), .A2(n8830), .ZN(n8832) );
  OR2_X1 U7563 ( .A1(n8763), .A2(n8762), .ZN(n8768) );
  NAND2_X2 U7564 ( .A1(n6643), .A2(P3_U3151), .ZN(n12350) );
  NOR2_X1 U7565 ( .A1(n8825), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n8838) );
  OR2_X1 U7566 ( .A1(n8217), .A2(n8317), .ZN(n8219) );
  NOR2_X1 U7567 ( .A1(n7121), .A2(n6738), .ZN(n7120) );
  AND2_X1 U7568 ( .A1(n8894), .A2(n8889), .ZN(n8890) );
  AND2_X2 U7569 ( .A1(n9043), .A2(n8879), .ZN(n8891) );
  NOR2_X1 U7570 ( .A1(n8888), .A2(n8887), .ZN(n8894) );
  AND2_X1 U7571 ( .A1(n8761), .A2(n6764), .ZN(n8212) );
  NAND2_X1 U7572 ( .A1(n7054), .A2(n9689), .ZN(n7053) );
  AND4_X1 U7573 ( .A1(n7884), .A2(n15471), .A3(n7580), .A4(n7857), .ZN(n7581)
         );
  AND3_X1 U7574 ( .A1(n8210), .A2(n8209), .A3(n8579), .ZN(n8761) );
  AND4_X1 U7575 ( .A1(n8875), .A2(n8874), .A3(n8873), .A4(n8872), .ZN(n8876)
         );
  AND3_X1 U7576 ( .A1(n8204), .A2(n8203), .A3(n8500), .ZN(n8208) );
  AND2_X1 U7577 ( .A1(n8955), .A2(n8956), .ZN(n8965) );
  INV_X1 U7578 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7130) );
  NOR2_X1 U7579 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n8213) );
  NOR2_X1 U7580 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n8214) );
  NOR2_X1 U7581 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7577) );
  NOR2_X1 U7582 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8881) );
  NOR2_X1 U7583 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8209) );
  NOR2_X1 U7584 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n8210) );
  INV_X4 U7585 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7586 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9444) );
  NOR2_X1 U7587 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n8201) );
  NOR2_X1 U7588 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8202) );
  INV_X1 U7589 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7674) );
  NOR2_X1 U7590 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8203) );
  INV_X1 U7591 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7794) );
  INV_X4 U7592 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7593 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n8830) );
  INV_X1 U7594 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8886) );
  INV_X1 U7595 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8902) );
  INV_X1 U7596 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8765) );
  INV_X1 U7597 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7857) );
  NOR2_X1 U7598 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8874) );
  NOR2_X1 U7599 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n8875) );
  INV_X1 U7600 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9188) );
  NOR2_X1 U7601 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8955) );
  INV_X1 U7602 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9757) );
  INV_X1 U7603 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9334) );
  OAI21_X2 U7604 ( .B1(n12864), .B2(n7007), .A(n7004), .ZN(n12838) );
  NAND2_X2 U7605 ( .A1(n12531), .A2(n12532), .ZN(n12854) );
  NAND2_X1 U7606 ( .A1(n6823), .A2(n9373), .ZN(n9356) );
  OR2_X1 U7607 ( .A1(n9350), .A2(n14708), .ZN(n8779) );
  OAI222_X1 U7608 ( .A1(n14330), .A2(n14327), .B1(P1_U3086), .B2(n8221), .C1(
        n14326), .C2(n14332), .ZN(P1_U3326) );
  OR2_X1 U7609 ( .A1(n12822), .A2(n12802), .ZN(n12671) );
  NOR2_X1 U7610 ( .A1(n11834), .A2(n14176), .ZN(n6653) );
  INV_X1 U7611 ( .A(n9657), .ZN(n6654) );
  BUF_X4 U7612 ( .A(n11598), .Z(n6655) );
  INV_X1 U7613 ( .A(n11716), .ZN(n11598) );
  XNOR2_X1 U7614 ( .A(n9445), .B(n9444), .ZN(n9580) );
  NOR2_X4 U7615 ( .A1(n14110), .A2(n14119), .ZN(n14113) );
  INV_X1 U7616 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7122) );
  INV_X1 U7617 ( .A(n7266), .ZN(n7123) );
  AND3_X1 U7618 ( .A1(n6956), .A2(n6709), .A3(n7579), .ZN(n6955) );
  AND2_X1 U7619 ( .A1(n7265), .A2(n7591), .ZN(n6956) );
  AND2_X1 U7620 ( .A1(n7581), .A2(n7762), .ZN(n6957) );
  NAND2_X1 U7621 ( .A1(n11976), .A2(n11977), .ZN(n7345) );
  INV_X1 U7622 ( .A(n13683), .ZN(n9452) );
  NAND2_X1 U7623 ( .A1(n9601), .A2(n9560), .ZN(n9592) );
  INV_X1 U7624 ( .A(n8324), .ZN(n8381) );
  NAND2_X1 U7625 ( .A1(n7706), .A2(n7704), .ZN(n7919) );
  NAND2_X1 U7626 ( .A1(n7760), .A2(n7614), .ZN(n6927) );
  NOR2_X2 U7627 ( .A1(n13978), .A2(n13985), .ZN(n13980) );
  AOI21_X1 U7628 ( .B1(n7558), .B2(n7556), .A(n6711), .ZN(n7555) );
  MUX2_X1 U7629 ( .A(n12036), .B(n12035), .S(n12034), .Z(n12037) );
  NAND2_X1 U7630 ( .A1(n7413), .A2(n7412), .ZN(n7411) );
  NOR2_X1 U7631 ( .A1(n6703), .A2(n7415), .ZN(n7413) );
  NAND2_X1 U7632 ( .A1(n6865), .A2(n7434), .ZN(n12142) );
  OR2_X1 U7633 ( .A1(n11522), .A2(n11521), .ZN(n7029) );
  INV_X1 U7634 ( .A(n7419), .ZN(n7421) );
  INV_X1 U7635 ( .A(n10854), .ZN(n7323) );
  INV_X1 U7636 ( .A(n8622), .ZN(n6982) );
  NAND2_X1 U7637 ( .A1(n11893), .A2(n12656), .ZN(n7243) );
  NAND2_X1 U7638 ( .A1(n13134), .A2(n8904), .ZN(n8906) );
  OR2_X1 U7639 ( .A1(n15011), .A2(n7133), .ZN(n6851) );
  NAND2_X1 U7640 ( .A1(n7134), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U7641 ( .A1(n10704), .A2(n7134), .ZN(n7132) );
  NOR2_X1 U7642 ( .A1(n12816), .A2(n12666), .ZN(n6999) );
  AND2_X1 U7643 ( .A1(n7098), .A2(n6759), .ZN(n7097) );
  INV_X1 U7644 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n15471) );
  NOR2_X1 U7645 ( .A1(n13389), .A2(n13567), .ZN(n7058) );
  NAND2_X1 U7646 ( .A1(n10777), .A2(n10776), .ZN(n7295) );
  INV_X1 U7647 ( .A(n10776), .ZN(n7298) );
  AND2_X1 U7648 ( .A1(n7181), .A2(n11734), .ZN(n7180) );
  NAND2_X1 U7649 ( .A1(n7183), .A2(n10519), .ZN(n7181) );
  INV_X1 U7650 ( .A(n10519), .ZN(n7182) );
  OR2_X1 U7651 ( .A1(n14887), .A2(n11399), .ZN(n7199) );
  INV_X1 U7652 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8884) );
  AND4_X1 U7653 ( .A1(n8878), .A2(n9188), .A3(n9334), .A4(n8877), .ZN(n8879)
         );
  INV_X1 U7654 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8877) );
  AND2_X1 U7655 ( .A1(n14083), .A2(n8806), .ZN(n7370) );
  INV_X1 U7656 ( .A(n7544), .ZN(n7541) );
  NAND2_X1 U7657 ( .A1(n7544), .A2(n7545), .ZN(n7542) );
  NAND2_X1 U7658 ( .A1(n7393), .A2(n7391), .ZN(n11680) );
  AOI21_X1 U7659 ( .B1(n11612), .B2(n7392), .A(n6816), .ZN(n7391) );
  NAND2_X1 U7660 ( .A1(n8735), .A2(n7389), .ZN(n7393) );
  INV_X1 U7661 ( .A(n7395), .ZN(n7392) );
  NAND2_X1 U7662 ( .A1(n8314), .A2(n6974), .ZN(n6976) );
  INV_X1 U7663 ( .A(n8712), .ZN(n6974) );
  INV_X1 U7664 ( .A(n8312), .ZN(n8313) );
  NAND2_X1 U7665 ( .A1(n10812), .A2(n8304), .ZN(n8683) );
  NAND2_X1 U7666 ( .A1(n8599), .A2(n8598), .ZN(n8288) );
  AOI21_X1 U7667 ( .B1(n7386), .B2(n7388), .A(n7384), .ZN(n7383) );
  INV_X1 U7668 ( .A(n8268), .ZN(n7384) );
  AOI21_X1 U7669 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15009), .A(n14351), .ZN(
        n14408) );
  AND2_X1 U7670 ( .A1(n14423), .A2(n6903), .ZN(n6902) );
  NAND3_X1 U7671 ( .A1(n9888), .A2(n8924), .A3(n8921), .ZN(n10152) );
  XNOR2_X1 U7672 ( .A(n7672), .B(n7671), .ZN(n9517) );
  NAND2_X1 U7673 ( .A1(n7003), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U7674 ( .A1(n15043), .A2(n12725), .ZN(n15044) );
  OR2_X1 U7675 ( .A1(n13080), .A2(n12354), .ZN(n7570) );
  NAND2_X1 U7676 ( .A1(n12822), .A2(n12802), .ZN(n12797) );
  AOI21_X1 U7677 ( .B1(n7006), .B2(n8128), .A(n7005), .ZN(n7004) );
  INV_X1 U7678 ( .A(n12532), .ZN(n7005) );
  AND2_X1 U7679 ( .A1(n12603), .A2(n12596), .ZN(n7010) );
  AND4_X1 U7680 ( .A1(n7745), .A2(n7744), .A3(n7743), .A4(n7742), .ZN(n15111)
         );
  INV_X1 U7681 ( .A(n8089), .ZN(n12480) );
  NAND2_X1 U7682 ( .A1(n8192), .A2(n10250), .ZN(n15182) );
  AND2_X1 U7683 ( .A1(n8934), .A2(n8183), .ZN(n12690) );
  NAND2_X1 U7684 ( .A1(n8155), .A2(n11043), .ZN(n7270) );
  AND2_X1 U7685 ( .A1(n7120), .A2(n7671), .ZN(n7118) );
  XNOR2_X1 U7686 ( .A(n8149), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U7687 ( .A1(n8148), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U7688 ( .A1(n7641), .A2(n7640), .ZN(n7995) );
  OAI21_X1 U7689 ( .B1(n7149), .B2(n6918), .A(n6916), .ZN(n7641) );
  AND2_X1 U7690 ( .A1(n6917), .A2(n7172), .ZN(n6916) );
  NAND2_X1 U7691 ( .A1(n7149), .A2(n6919), .ZN(n7637) );
  NAND2_X1 U7692 ( .A1(n6927), .A2(n7616), .ZN(n7777) );
  NOR2_X1 U7693 ( .A1(n7611), .A2(n7170), .ZN(n7169) );
  INV_X1 U7694 ( .A(n7609), .ZN(n7170) );
  NAND2_X1 U7695 ( .A1(n7345), .A2(n13202), .ZN(n7342) );
  NAND2_X1 U7696 ( .A1(n7343), .A2(n7345), .ZN(n7340) );
  INV_X1 U7697 ( .A(n11974), .ZN(n7344) );
  OR2_X1 U7698 ( .A1(n11494), .A2(n11493), .ZN(n11529) );
  AOI21_X1 U7699 ( .B1(n7310), .B2(n7311), .A(n7308), .ZN(n7307) );
  INV_X1 U7700 ( .A(n11200), .ZN(n7308) );
  NAND2_X1 U7701 ( .A1(n11558), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n11576) );
  AND4_X1 U7702 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11930) );
  AND2_X1 U7703 ( .A1(n9456), .A2(n9452), .ZN(n9605) );
  NOR2_X1 U7704 ( .A1(n13358), .A2(n13365), .ZN(n13359) );
  NAND2_X1 U7705 ( .A1(n13682), .A2(n6652), .ZN(n6960) );
  INV_X1 U7706 ( .A(n7058), .ZN(n13377) );
  NAND2_X1 U7707 ( .A1(n7058), .A2(n7057), .ZN(n13358) );
  NAND2_X1 U7708 ( .A1(n13504), .A2(n11911), .ZN(n13495) );
  AOI21_X1 U7709 ( .B1(n7273), .B2(n7275), .A(n6790), .ZN(n6945) );
  AOI21_X1 U7710 ( .B1(n7209), .B2(n7207), .A(n6756), .ZN(n7206) );
  NAND2_X1 U7711 ( .A1(n11934), .A2(n7215), .ZN(n7210) );
  NAND2_X1 U7712 ( .A1(n11908), .A2(n6665), .ZN(n13535) );
  OR2_X1 U7713 ( .A1(n11182), .A2(n11181), .ZN(n11184) );
  OAI21_X1 U7714 ( .B1(n7272), .B2(n6933), .A(n6931), .ZN(n10350) );
  AND2_X1 U7715 ( .A1(n6932), .A2(n10277), .ZN(n6931) );
  OR2_X1 U7716 ( .A1(n7271), .A2(n6933), .ZN(n6932) );
  INV_X1 U7717 ( .A(n10262), .ZN(n6933) );
  INV_X1 U7718 ( .A(n13562), .ZN(n7228) );
  NAND2_X1 U7719 ( .A1(n14098), .A2(n7528), .ZN(n14076) );
  NOR2_X1 U7720 ( .A1(n14083), .A2(n7529), .ZN(n7528) );
  INV_X1 U7721 ( .A(n8696), .ZN(n7529) );
  INV_X1 U7722 ( .A(n8597), .ZN(n7559) );
  OAI21_X1 U7723 ( .B1(n10640), .B2(n7547), .A(n7546), .ZN(n10990) );
  INV_X1 U7724 ( .A(n7548), .ZN(n7547) );
  AOI21_X1 U7725 ( .B1(n7548), .B2(n12228), .A(n6726), .ZN(n7546) );
  AOI21_X1 U7726 ( .B1(n10019), .B2(n7521), .A(n6734), .ZN(n7520) );
  INV_X1 U7727 ( .A(n8450), .ZN(n7521) );
  NAND2_X1 U7728 ( .A1(n10050), .A2(n8435), .ZN(n9906) );
  INV_X1 U7729 ( .A(n8404), .ZN(n7527) );
  INV_X1 U7730 ( .A(n9957), .ZN(n7079) );
  NAND2_X1 U7731 ( .A1(n8754), .A2(n8753), .ZN(n13992) );
  NAND2_X1 U7732 ( .A1(n8588), .A2(n8587), .ZN(n14276) );
  INV_X2 U7733 ( .A(n8369), .ZN(n12195) );
  AND2_X1 U7734 ( .A1(n8206), .A2(n8205), .ZN(n8207) );
  INV_X1 U7735 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8211) );
  OR2_X1 U7736 ( .A1(n8698), .A2(n8697), .ZN(n8700) );
  OR2_X1 U7737 ( .A1(n8640), .A2(n8639), .ZN(n8657) );
  AND2_X1 U7738 ( .A1(P3_U3897), .A2(n11319), .ZN(n15096) );
  INV_X1 U7739 ( .A(n13541), .ZN(n13284) );
  NAND2_X1 U7740 ( .A1(n11353), .A2(n6693), .ZN(n11361) );
  NOR2_X1 U7741 ( .A1(n12040), .A2(n12212), .ZN(n7438) );
  OR2_X1 U7742 ( .A1(n12055), .A2(n12053), .ZN(n7473) );
  NOR2_X1 U7743 ( .A1(n11385), .A2(n11388), .ZN(n7424) );
  INV_X1 U7744 ( .A(n11385), .ZN(n7423) );
  INV_X1 U7745 ( .A(n11394), .ZN(n7032) );
  NAND3_X1 U7746 ( .A1(n7445), .A2(n7444), .A3(n12065), .ZN(n7443) );
  INV_X1 U7747 ( .A(n12063), .ZN(n7446) );
  INV_X1 U7748 ( .A(n12068), .ZN(n6882) );
  OAI22_X1 U7749 ( .A1(n12073), .A2(n6864), .B1(n12074), .B2(n6863), .ZN(
        n12077) );
  NOR2_X1 U7750 ( .A1(n12075), .A2(n12072), .ZN(n6864) );
  INV_X1 U7751 ( .A(n12072), .ZN(n6863) );
  NAND2_X1 U7752 ( .A1(n7451), .A2(n7450), .ZN(n12073) );
  AND2_X1 U7753 ( .A1(n7026), .A2(n7025), .ZN(n7024) );
  NOR2_X1 U7754 ( .A1(n11413), .A2(n11412), .ZN(n7023) );
  INV_X1 U7755 ( .A(n6774), .ZN(n7026) );
  AND2_X1 U7756 ( .A1(n11412), .A2(n11413), .ZN(n7433) );
  NOR2_X1 U7757 ( .A1(n12118), .A2(n6875), .ZN(n6874) );
  NAND2_X1 U7758 ( .A1(n6877), .A2(n14168), .ZN(n6875) );
  INV_X1 U7759 ( .A(n11446), .ZN(n7429) );
  NAND2_X1 U7760 ( .A1(n11434), .A2(n6720), .ZN(n7431) );
  NAND2_X1 U7761 ( .A1(n11439), .A2(n6721), .ZN(n7017) );
  AND2_X1 U7762 ( .A1(n7019), .A2(n11438), .ZN(n7018) );
  INV_X1 U7763 ( .A(n11479), .ZN(n7414) );
  NAND2_X1 U7764 ( .A1(n6659), .A2(n7410), .ZN(n7409) );
  AOI21_X1 U7765 ( .B1(n12142), .B2(n12141), .A(n12139), .ZN(n12140) );
  OR2_X1 U7766 ( .A1(n12147), .A2(n12148), .ZN(n7462) );
  NAND2_X1 U7767 ( .A1(n12150), .A2(n12151), .ZN(n7461) );
  INV_X1 U7768 ( .A(n12150), .ZN(n7465) );
  AOI22_X1 U7769 ( .A1(n11508), .A2(n11507), .B1(n11506), .B2(n11505), .ZN(
        n11519) );
  INV_X1 U7770 ( .A(n6893), .ZN(n14340) );
  INV_X1 U7771 ( .A(n10705), .ZN(n7134) );
  NOR2_X1 U7772 ( .A1(n8031), .A2(n6924), .ZN(n6923) );
  INV_X1 U7773 ( .A(n7646), .ZN(n6924) );
  INV_X1 U7774 ( .A(n8019), .ZN(n6921) );
  INV_X1 U7775 ( .A(n7626), .ZN(n7148) );
  INV_X1 U7776 ( .A(n7147), .ZN(n7146) );
  OAI21_X1 U7777 ( .B1(n7148), .B2(n7625), .A(n7888), .ZN(n7147) );
  NAND2_X1 U7778 ( .A1(n6964), .A2(n6963), .ZN(n6962) );
  INV_X1 U7779 ( .A(n11679), .ZN(n6963) );
  INV_X1 U7780 ( .A(n11678), .ZN(n6964) );
  NAND2_X1 U7781 ( .A1(n7405), .A2(n7404), .ZN(n8312) );
  AOI21_X1 U7782 ( .B1(n6680), .B2(n8697), .A(n6805), .ZN(n7404) );
  AOI21_X1 U7783 ( .B1(n8284), .B2(n8278), .A(n7376), .ZN(n7375) );
  INV_X1 U7784 ( .A(n8577), .ZN(n7376) );
  INV_X1 U7785 ( .A(n8284), .ZN(n7377) );
  INV_X1 U7786 ( .A(n8235), .ZN(n8237) );
  INV_X1 U7787 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7673) );
  INV_X1 U7788 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6929) );
  INV_X1 U7789 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15391) );
  INV_X1 U7790 ( .A(n12448), .ZN(n7238) );
  AND3_X1 U7791 ( .A1(n7739), .A2(n7738), .A3(n7737), .ZN(n8915) );
  OR2_X1 U7792 ( .A1(n7882), .A2(SI_2_), .ZN(n7739) );
  AOI21_X1 U7793 ( .B1(n14959), .B2(n14960), .A(n6705), .ZN(n10379) );
  NAND2_X1 U7794 ( .A1(n14972), .A2(n6985), .ZN(n10688) );
  OR2_X1 U7795 ( .A1(n10389), .A2(n15205), .ZN(n6985) );
  NAND2_X1 U7796 ( .A1(n6993), .A2(n6992), .ZN(n10692) );
  OR2_X1 U7797 ( .A1(n15000), .A2(n15208), .ZN(n6992) );
  NAND2_X1 U7798 ( .A1(n14994), .A2(n14995), .ZN(n6993) );
  NAND2_X1 U7799 ( .A1(n15048), .A2(n6986), .ZN(n12779) );
  NAND2_X1 U7800 ( .A1(n15051), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6986) );
  INV_X1 U7801 ( .A(n6999), .ZN(n6998) );
  INV_X1 U7802 ( .A(n12854), .ZN(n7008) );
  AND2_X1 U7803 ( .A1(n6758), .A2(n12499), .ZN(n7106) );
  INV_X1 U7804 ( .A(n7111), .ZN(n7110) );
  NAND2_X1 U7805 ( .A1(n12917), .A2(n7112), .ZN(n7111) );
  INV_X1 U7806 ( .A(n7564), .ZN(n7112) );
  OR2_X1 U7807 ( .A1(n11869), .A2(n12918), .ZN(n12625) );
  NAND2_X1 U7808 ( .A1(n12505), .A2(n7115), .ZN(n8110) );
  INV_X1 U7809 ( .A(n10917), .ZN(n7115) );
  NAND2_X1 U7810 ( .A1(n15116), .A2(n8102), .ZN(n10503) );
  INV_X1 U7811 ( .A(n10049), .ZN(n8191) );
  INV_X1 U7812 ( .A(n10250), .ZN(n12535) );
  NAND2_X1 U7813 ( .A1(n7667), .A2(n7267), .ZN(n7266) );
  INV_X1 U7814 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7267) );
  INV_X1 U7815 ( .A(n7121), .ZN(n7119) );
  INV_X1 U7816 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7589) );
  INV_X1 U7817 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7265) );
  OR2_X1 U7818 ( .A1(n6919), .A2(n6918), .ZN(n6917) );
  AND2_X1 U7819 ( .A1(n10941), .A2(n7318), .ZN(n7317) );
  NAND2_X1 U7820 ( .A1(n7322), .A2(n7320), .ZN(n7318) );
  OR2_X1 U7821 ( .A1(n10943), .A2(n10948), .ZN(n10940) );
  NAND2_X1 U7822 ( .A1(n7317), .A2(n7319), .ZN(n7315) );
  INV_X1 U7823 ( .A(n7320), .ZN(n7319) );
  NAND2_X1 U7824 ( .A1(n7323), .A2(n6811), .ZN(n7320) );
  INV_X1 U7825 ( .A(n10209), .ZN(n7334) );
  OR2_X1 U7826 ( .A1(n11698), .A2(n13354), .ZN(n11713) );
  AND2_X1 U7827 ( .A1(n11602), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U7828 ( .A1(n11919), .A2(n7289), .ZN(n7288) );
  INV_X1 U7829 ( .A(n11918), .ZN(n7289) );
  NAND2_X1 U7830 ( .A1(n6668), .A2(n6937), .ZN(n6935) );
  AND2_X1 U7831 ( .A1(n11917), .A2(n11941), .ZN(n7220) );
  NOR2_X1 U7832 ( .A1(n13588), .A2(n13596), .ZN(n7068) );
  NOR2_X1 U7833 ( .A1(n7188), .A2(n13467), .ZN(n7187) );
  NOR2_X1 U7834 ( .A1(n6690), .A2(n7189), .ZN(n7188) );
  INV_X1 U7835 ( .A(n11939), .ZN(n7189) );
  INV_X1 U7836 ( .A(n7209), .ZN(n7208) );
  NOR2_X1 U7837 ( .A1(n11935), .A2(n7216), .ZN(n7215) );
  INV_X1 U7838 ( .A(n11932), .ZN(n7216) );
  AND2_X1 U7839 ( .A1(n10753), .A2(n11012), .ZN(n7201) );
  NAND2_X1 U7840 ( .A1(n6745), .A2(n10355), .ZN(n7183) );
  NOR2_X1 U7841 ( .A1(n14918), .A2(n11424), .ZN(n7074) );
  NOR2_X1 U7842 ( .A1(n7193), .A2(n11732), .ZN(n7191) );
  INV_X1 U7843 ( .A(n7197), .ZN(n7193) );
  INV_X1 U7844 ( .A(n7199), .ZN(n7195) );
  AND2_X1 U7845 ( .A1(n11732), .A2(n10261), .ZN(n7271) );
  AND2_X1 U7846 ( .A1(n9616), .A2(n9597), .ZN(n11722) );
  NAND2_X1 U7847 ( .A1(n9582), .A2(n13349), .ZN(n9645) );
  XNOR2_X1 U7848 ( .A(n9581), .B(n11759), .ZN(n9582) );
  INV_X1 U7849 ( .A(n10367), .ZN(n10368) );
  OR2_X1 U7850 ( .A1(n10296), .A2(n11417), .ZN(n10367) );
  INV_X1 U7851 ( .A(n13742), .ZN(n7481) );
  NAND2_X1 U7852 ( .A1(n12174), .A2(n7470), .ZN(n7469) );
  NAND2_X1 U7853 ( .A1(n6871), .A2(n6672), .ZN(n6870) );
  OR2_X1 U7854 ( .A1(n6661), .A2(n6768), .ZN(n6871) );
  OR2_X1 U7855 ( .A1(n6661), .A2(n12176), .ZN(n6868) );
  INV_X1 U7856 ( .A(n12125), .ZN(n7364) );
  INV_X1 U7857 ( .A(n8797), .ZN(n7358) );
  NOR2_X1 U7858 ( .A1(n14584), .A2(n7087), .ZN(n7086) );
  INV_X1 U7859 ( .A(n7088), .ZN(n7087) );
  NOR2_X1 U7860 ( .A1(n12082), .A2(n12092), .ZN(n7088) );
  NAND2_X1 U7861 ( .A1(n14022), .A2(n14021), .ZN(n14020) );
  INV_X1 U7862 ( .A(n7370), .ZN(n7369) );
  AND2_X1 U7863 ( .A1(n8807), .A2(n7368), .ZN(n7367) );
  NAND2_X1 U7864 ( .A1(n7370), .A2(n8694), .ZN(n7368) );
  NOR2_X1 U7865 ( .A1(n8751), .A2(n7400), .ZN(n7399) );
  INV_X1 U7866 ( .A(n8734), .ZN(n7400) );
  NAND2_X1 U7867 ( .A1(n7397), .A2(n7396), .ZN(n7395) );
  INV_X1 U7868 ( .A(n8750), .ZN(n7397) );
  NAND2_X1 U7869 ( .A1(n6681), .A2(n6795), .ZN(n6984) );
  INV_X1 U7870 ( .A(n8583), .ZN(n8585) );
  INV_X1 U7871 ( .A(n7381), .ZN(n7380) );
  INV_X1 U7872 ( .A(n8251), .ZN(n7382) );
  INV_X1 U7873 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14379) );
  INV_X1 U7874 ( .A(n6894), .ZN(n14344) );
  XNOR2_X1 U7875 ( .A(n14344), .B(n9716), .ZN(n14392) );
  OAI22_X1 U7876 ( .A1(n14397), .A2(n14347), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14989), .ZN(n14348) );
  INV_X1 U7877 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U7878 ( .A1(n11295), .A2(n11303), .ZN(n7252) );
  NAND2_X1 U7879 ( .A1(n10152), .A2(n8925), .ZN(n10341) );
  NAND2_X1 U7880 ( .A1(n7255), .A2(n7254), .ZN(n10737) );
  AND2_X1 U7881 ( .A1(n10605), .A2(n10606), .ZN(n7254) );
  OAI21_X1 U7882 ( .B1(n12425), .B2(n7258), .A(n7256), .ZN(n11883) );
  AOI21_X1 U7883 ( .B1(n7259), .B2(n7257), .A(n6792), .ZN(n7256) );
  INV_X1 U7884 ( .A(n7259), .ZN(n7258) );
  INV_X1 U7885 ( .A(n12424), .ZN(n7257) );
  INV_X1 U7886 ( .A(n12710), .ZN(n11028) );
  INV_X1 U7887 ( .A(n11884), .ZN(n7234) );
  AND2_X1 U7888 ( .A1(n7243), .A2(n11890), .ZN(n7242) );
  INV_X1 U7889 ( .A(n7252), .ZN(n7251) );
  INV_X1 U7890 ( .A(n7250), .ZN(n7249) );
  OAI21_X1 U7891 ( .B1(n7253), .B2(n7251), .A(n11307), .ZN(n7250) );
  NAND2_X1 U7892 ( .A1(n13137), .A2(n7130), .ZN(n7129) );
  NOR2_X1 U7893 ( .A1(n9703), .A2(n6862), .ZN(n14958) );
  AND2_X1 U7894 ( .A1(n9704), .A2(n6995), .ZN(n6862) );
  OAI21_X1 U7895 ( .B1(n9710), .B2(n9709), .A(n6994), .ZN(n14959) );
  NAND2_X1 U7896 ( .A1(n9707), .A2(n6995), .ZN(n6994) );
  NOR2_X1 U7897 ( .A1(n14957), .A2(n14958), .ZN(n14956) );
  NAND2_X1 U7898 ( .A1(n14974), .A2(n14973), .ZN(n14972) );
  OAI21_X1 U7899 ( .B1(n10374), .B2(n7137), .A(n7135), .ZN(n14969) );
  NAND2_X1 U7900 ( .A1(n7138), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U7901 ( .A1(n10375), .A2(n7138), .ZN(n7135) );
  INV_X1 U7902 ( .A(n7136), .ZN(n14971) );
  OAI21_X1 U7903 ( .B1(n10374), .B2(n10486), .A(n10373), .ZN(n7136) );
  XNOR2_X1 U7904 ( .A(n10688), .B(n10698), .ZN(n10383) );
  NOR2_X1 U7905 ( .A1(n14969), .A2(n7139), .ZN(n10697) );
  NOR2_X1 U7906 ( .A1(n10389), .A2(n10376), .ZN(n7139) );
  NOR2_X1 U7907 ( .A1(n12741), .A2(n6954), .ZN(n15038) );
  AND2_X1 U7908 ( .A1(n12742), .A2(n12774), .ZN(n6954) );
  OR2_X1 U7909 ( .A1(n15027), .A2(n12724), .ZN(n15043) );
  NAND2_X1 U7910 ( .A1(n15050), .A2(n15049), .ZN(n15048) );
  NOR2_X1 U7911 ( .A1(n15038), .A2(n15037), .ZN(n15036) );
  XNOR2_X1 U7912 ( .A(n12779), .B(n12749), .ZN(n15068) );
  NAND2_X1 U7913 ( .A1(n6852), .A2(n12753), .ZN(n12731) );
  OAI21_X1 U7914 ( .B1(n15066), .B2(n15065), .A(n6853), .ZN(n6852) );
  NAND2_X1 U7915 ( .A1(n6858), .A2(n6682), .ZN(n6857) );
  NAND2_X1 U7916 ( .A1(n12733), .A2(n6856), .ZN(n6855) );
  OR2_X1 U7917 ( .A1(n14463), .A2(n14464), .ZN(n6861) );
  OAI22_X1 U7918 ( .A1(n14505), .A2(n7140), .B1(n6686), .B2(n14521), .ZN(
        n14523) );
  OR2_X1 U7919 ( .A1(n14521), .A2(n15481), .ZN(n7140) );
  NAND2_X1 U7920 ( .A1(n8135), .A2(n8134), .ZN(n12805) );
  NAND2_X1 U7921 ( .A1(n12497), .A2(n12664), .ZN(n12832) );
  NAND2_X1 U7922 ( .A1(n12864), .A2(n12863), .ZN(n12866) );
  AOI21_X1 U7923 ( .B1(n12906), .B2(n12638), .A(n7014), .ZN(n7013) );
  AND2_X1 U7924 ( .A1(n12647), .A2(n12646), .ZN(n12881) );
  INV_X1 U7925 ( .A(n12640), .ZN(n12890) );
  NAND2_X1 U7926 ( .A1(n6704), .A2(n7101), .ZN(n7098) );
  NAND2_X1 U7927 ( .A1(n8121), .A2(n7102), .ZN(n7101) );
  INV_X1 U7928 ( .A(n7565), .ZN(n7102) );
  NAND2_X1 U7929 ( .A1(n6704), .A2(n7100), .ZN(n7099) );
  INV_X1 U7930 ( .A(n12599), .ZN(n7100) );
  AND2_X1 U7931 ( .A1(n12618), .A2(n12615), .ZN(n12965) );
  NAND2_X1 U7932 ( .A1(n11087), .A2(n12512), .ZN(n7011) );
  AND4_X1 U7933 ( .A1(n7914), .A2(n7913), .A3(n7912), .A4(n7911), .ZN(n11297)
         );
  AND2_X1 U7934 ( .A1(n12603), .A2(n12602), .ZN(n12599) );
  AND2_X1 U7935 ( .A1(n7891), .A2(n7890), .ZN(n11136) );
  AOI21_X1 U7936 ( .B1(n10719), .B2(n12568), .A(n8106), .ZN(n10981) );
  AND2_X1 U7937 ( .A1(n12559), .A2(n12563), .ZN(n12557) );
  AND3_X1 U7938 ( .A1(n7767), .A2(n7766), .A3(n7765), .ZN(n10252) );
  INV_X1 U7939 ( .A(n12987), .ZN(n15132) );
  AND2_X1 U7940 ( .A1(n8189), .A2(n8188), .ZN(n9936) );
  OAI21_X1 U7941 ( .B1(n11320), .B2(n8089), .A(n8090), .ZN(n8136) );
  OR2_X1 U7942 ( .A1(n7882), .A2(n7396), .ZN(n8090) );
  NAND2_X1 U7943 ( .A1(n7000), .A2(n12664), .ZN(n12812) );
  NAND2_X1 U7944 ( .A1(n8034), .A2(n8033), .ZN(n12651) );
  OR2_X1 U7945 ( .A1(n7882), .A2(SI_10_), .ZN(n7002) );
  AND3_X1 U7946 ( .A1(n7836), .A2(n7835), .A3(n7834), .ZN(n15183) );
  NAND2_X1 U7947 ( .A1(n7270), .A2(n8180), .ZN(n9271) );
  NAND2_X1 U7948 ( .A1(n7659), .A2(n7658), .ZN(n8088) );
  NAND2_X1 U7949 ( .A1(n8066), .A2(n7655), .ZN(n8078) );
  INV_X1 U7950 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8153) );
  INV_X1 U7951 ( .A(n7650), .ZN(n6926) );
  NAND2_X1 U7952 ( .A1(n7651), .A2(n7650), .ZN(n8042) );
  OAI21_X1 U7953 ( .B1(n7995), .B2(n7165), .A(n7161), .ZN(n8020) );
  AOI21_X1 U7954 ( .B1(n7164), .B2(n7163), .A(n7162), .ZN(n7161) );
  INV_X1 U7955 ( .A(n7644), .ZN(n7162) );
  INV_X1 U7956 ( .A(n7994), .ZN(n7163) );
  NAND2_X1 U7957 ( .A1(n8020), .A2(n8019), .ZN(n8018) );
  NAND2_X1 U7958 ( .A1(n7995), .A2(n7994), .ZN(n7167) );
  NAND2_X1 U7959 ( .A1(n7593), .A2(n7589), .ZN(n7666) );
  AND2_X1 U7960 ( .A1(n7762), .A2(n7265), .ZN(n6958) );
  INV_X1 U7961 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7585) );
  INV_X1 U7962 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7580) );
  AOI21_X1 U7963 ( .B1(n7635), .B2(n7152), .A(n6817), .ZN(n7151) );
  INV_X1 U7964 ( .A(n7634), .ZN(n7152) );
  NOR2_X1 U7965 ( .A1(n7953), .A2(n7965), .ZN(n7150) );
  OR2_X1 U7966 ( .A1(n7859), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U7967 ( .A1(n6906), .A2(n6908), .ZN(n7856) );
  AOI21_X1 U7968 ( .B1(n6911), .B2(n6909), .A(n6797), .ZN(n6908) );
  INV_X1 U7969 ( .A(n6691), .ZN(n6909) );
  AOI21_X1 U7970 ( .B1(n7159), .B2(n7158), .A(n6749), .ZN(n7157) );
  INV_X1 U7971 ( .A(n7620), .ZN(n7158) );
  NAND2_X1 U7972 ( .A1(n6914), .A2(n7160), .ZN(n7811) );
  INV_X1 U7973 ( .A(n7808), .ZN(n7160) );
  XNOR2_X1 U7974 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7798) );
  NAND2_X1 U7975 ( .A1(n7168), .A2(n6725), .ZN(n7760) );
  INV_X1 U7976 ( .A(n7757), .ZN(n7171) );
  INV_X1 U7977 ( .A(n10205), .ZN(n10206) );
  NOR2_X1 U7978 ( .A1(n11529), .A2(n11526), .ZN(n11544) );
  AOI21_X1 U7979 ( .B1(n11072), .B2(n11068), .A(n11197), .ZN(n7310) );
  INV_X1 U7980 ( .A(n11072), .ZN(n7311) );
  NOR2_X1 U7981 ( .A1(n11576), .A2(n13216), .ZN(n11590) );
  NAND2_X1 U7982 ( .A1(n6701), .A2(n7333), .ZN(n7332) );
  INV_X1 U7983 ( .A(n10332), .ZN(n7333) );
  OR2_X1 U7984 ( .A1(n10332), .A2(n10331), .ZN(n7331) );
  INV_X1 U7985 ( .A(n7332), .ZN(n7329) );
  NAND2_X1 U7986 ( .A1(n7330), .A2(n6701), .ZN(n10333) );
  INV_X1 U7987 ( .A(n10207), .ZN(n7330) );
  AOI21_X1 U7988 ( .B1(n7340), .B2(n7342), .A(n7338), .ZN(n7337) );
  INV_X1 U7989 ( .A(n13171), .ZN(n7338) );
  NOR2_X1 U7990 ( .A1(n9824), .A2(n9655), .ZN(n7304) );
  CLKBUF_X1 U7991 ( .A(n11070), .Z(n6837) );
  AND4_X1 U7992 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n13267) );
  AND2_X1 U7993 ( .A1(n11565), .A2(n11564), .ZN(n13237) );
  AND2_X1 U7994 ( .A1(n13475), .A2(n7064), .ZN(n13404) );
  AND2_X1 U7995 ( .A1(n7066), .A2(n7065), .ZN(n7064) );
  OAI21_X1 U7996 ( .B1(n11942), .B2(n7219), .A(n7217), .ZN(n13421) );
  INV_X1 U7997 ( .A(n7218), .ZN(n7217) );
  OAI21_X1 U7998 ( .B1(n7220), .B2(n7219), .A(n13417), .ZN(n7218) );
  INV_X1 U7999 ( .A(n13418), .ZN(n7219) );
  NAND2_X1 U8000 ( .A1(n11942), .A2(n7220), .ZN(n13432) );
  NAND2_X1 U8001 ( .A1(n6938), .A2(n6936), .ZN(n11916) );
  NAND2_X1 U8002 ( .A1(n11916), .A2(n6702), .ZN(n13428) );
  NAND2_X1 U8003 ( .A1(n13495), .A2(n6657), .ZN(n6938) );
  INV_X1 U8004 ( .A(n13282), .ZN(n13451) );
  AND2_X1 U8005 ( .A1(n6945), .A2(n13505), .ZN(n6943) );
  AND2_X1 U8006 ( .A1(n7213), .A2(n11936), .ZN(n7212) );
  OR2_X1 U8007 ( .A1(n11935), .A2(n7214), .ZN(n7213) );
  NAND2_X1 U8008 ( .A1(n11933), .A2(n11932), .ZN(n7214) );
  OAI21_X1 U8009 ( .B1(n11184), .B2(n7284), .A(n7282), .ZN(n11906) );
  INV_X1 U8010 ( .A(n7283), .ZN(n7282) );
  OAI21_X1 U8011 ( .B1(n6698), .B2(n7284), .A(n11275), .ZN(n7283) );
  INV_X1 U8012 ( .A(n7223), .ZN(n7222) );
  NOR2_X1 U8013 ( .A1(n11185), .A2(n11737), .ZN(n7285) );
  AND4_X1 U8014 ( .A1(n10773), .A2(n10772), .A3(n10771), .A4(n10770), .ZN(
        n11452) );
  NAND2_X1 U8015 ( .A1(n7225), .A2(n11740), .ZN(n11225) );
  OAI21_X1 U8016 ( .B1(n11010), .B2(n13290), .A(n11011), .ZN(n11182) );
  AOI21_X1 U8017 ( .B1(n7293), .B2(n7296), .A(n11445), .ZN(n7291) );
  NAND2_X1 U8018 ( .A1(n7177), .A2(n10748), .ZN(n7176) );
  NAND2_X1 U8019 ( .A1(n7180), .A2(n7182), .ZN(n7177) );
  NAND2_X1 U8020 ( .A1(n7175), .A2(n10753), .ZN(n14552) );
  INV_X1 U8021 ( .A(n10778), .ZN(n7300) );
  NAND2_X1 U8022 ( .A1(n10260), .A2(n10259), .ZN(n7272) );
  NAND2_X1 U8023 ( .A1(n7272), .A2(n7271), .ZN(n10290) );
  OAI21_X1 U8024 ( .B1(n9847), .B2(n11572), .A(n9849), .ZN(n11392) );
  XNOR2_X1 U8025 ( .A(n11392), .B(n13297), .ZN(n11727) );
  INV_X1 U8026 ( .A(n13298), .ZN(n11384) );
  INV_X1 U8027 ( .A(n13540), .ZN(n13650) );
  OR2_X1 U8028 ( .A1(n9592), .A2(n8959), .ZN(n9564) );
  XNOR2_X1 U8029 ( .A(n11323), .B(n13179), .ZN(n9570) );
  NAND2_X1 U8030 ( .A1(n9570), .A2(n9571), .ZN(n10226) );
  CLKBUF_X1 U8031 ( .A(n9645), .Z(n13647) );
  NAND2_X1 U8032 ( .A1(n11543), .A2(n11542), .ZN(n13601) );
  OR2_X1 U8033 ( .A1(n11541), .A2(n11572), .ZN(n11543) );
  AND2_X1 U8034 ( .A1(n13647), .A2(n13655), .ZN(n14890) );
  AND2_X1 U8035 ( .A1(n9420), .A2(n9421), .ZN(n14850) );
  NAND2_X1 U8036 ( .A1(n7425), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9448) );
  OR2_X1 U8037 ( .A1(n8897), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U8038 ( .A1(n6746), .A2(n7401), .ZN(n10812) );
  INV_X1 U8039 ( .A(n10810), .ZN(n8303) );
  CLKBUF_X1 U8040 ( .A(n9443), .Z(n8893) );
  OR2_X1 U8041 ( .A1(n8987), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9038) );
  AND2_X1 U8042 ( .A1(n13764), .A2(n12277), .ZN(n13703) );
  AOI22_X1 U8043 ( .A1(n9350), .A2(n6653), .B1(n9345), .B2(n12034), .ZN(n9351)
         );
  NOR2_X1 U8044 ( .A1(n8663), .A2(n8662), .ZN(n8671) );
  INV_X1 U8045 ( .A(n10841), .ZN(n7497) );
  INV_X1 U8046 ( .A(n9809), .ZN(n7503) );
  NOR2_X1 U8047 ( .A1(n14597), .A2(n7500), .ZN(n7499) );
  INV_X1 U8048 ( .A(n11118), .ZN(n7500) );
  NAND2_X1 U8049 ( .A1(n9354), .A2(n9353), .ZN(n9374) );
  OR2_X1 U8050 ( .A1(n8590), .A2(n8589), .ZN(n8616) );
  AND2_X1 U8051 ( .A1(n12257), .A2(n9219), .ZN(n9921) );
  INV_X1 U8052 ( .A(n12179), .ZN(n8718) );
  NAND2_X1 U8053 ( .A1(n8985), .A2(n7346), .ZN(n9001) );
  INV_X1 U8054 ( .A(n12240), .ZN(n14009) );
  NAND2_X1 U8055 ( .A1(n14113), .A2(n7089), .ZN(n14030) );
  NOR2_X1 U8056 ( .A1(n14032), .A2(n7091), .ZN(n7089) );
  AND2_X1 U8057 ( .A1(n14076), .A2(n8710), .ZN(n14071) );
  NAND2_X1 U8058 ( .A1(n14071), .A2(n14070), .ZN(n14069) );
  NAND2_X1 U8059 ( .A1(n14109), .A2(n7370), .ZN(n14054) );
  NAND2_X1 U8060 ( .A1(n8805), .A2(n14106), .ZN(n14109) );
  NAND2_X1 U8061 ( .A1(n7534), .A2(n7535), .ZN(n14127) );
  AOI21_X1 U8062 ( .B1(n7537), .B2(n7536), .A(n6736), .ZN(n7535) );
  INV_X1 U8063 ( .A(n14142), .ZN(n14133) );
  OR2_X1 U8064 ( .A1(n7366), .A2(n6658), .ZN(n14161) );
  INV_X1 U8065 ( .A(n13824), .ZN(n13745) );
  NAND2_X1 U8066 ( .A1(n11096), .A2(n12230), .ZN(n11095) );
  NAND2_X1 U8067 ( .A1(n10991), .A2(n6663), .ZN(n11093) );
  AND2_X1 U8068 ( .A1(n12102), .A2(n12103), .ZN(n12234) );
  AND2_X1 U8069 ( .A1(n12097), .A2(n12089), .ZN(n12209) );
  NOR2_X1 U8070 ( .A1(n12209), .A2(n7549), .ZN(n7548) );
  INV_X1 U8071 ( .A(n8544), .ZN(n7549) );
  OR2_X1 U8072 ( .A1(n9778), .A2(n7346), .ZN(n7349) );
  NAND2_X1 U8073 ( .A1(n10573), .A2(n8527), .ZN(n10640) );
  NAND2_X1 U8074 ( .A1(n10640), .A2(n10639), .ZN(n10638) );
  AOI21_X1 U8075 ( .B1(n12224), .B2(n8793), .A(n10418), .ZN(n7359) );
  OR2_X1 U8076 ( .A1(n12224), .A2(n7533), .ZN(n7532) );
  INV_X1 U8077 ( .A(n8497), .ZN(n7533) );
  OR2_X1 U8078 ( .A1(n10301), .A2(n12224), .ZN(n10302) );
  NAND2_X1 U8079 ( .A1(n10308), .A2(n12224), .ZN(n10307) );
  NAND2_X1 U8080 ( .A1(n7519), .A2(n7518), .ZN(n14653) );
  NAND2_X1 U8081 ( .A1(n9906), .A2(n9908), .ZN(n9905) );
  NAND2_X1 U8082 ( .A1(n7525), .A2(n7523), .ZN(n10050) );
  INV_X1 U8083 ( .A(n7524), .ZN(n7523) );
  OAI21_X1 U8084 ( .B1(n9747), .B2(n6685), .A(n12218), .ZN(n7524) );
  XNOR2_X1 U8085 ( .A(n12056), .B(n9910), .ZN(n12218) );
  AND2_X1 U8086 ( .A1(n7516), .A2(n8390), .ZN(n7515) );
  INV_X1 U8087 ( .A(n14176), .ZN(n14661) );
  INV_X1 U8088 ( .A(n14260), .ZN(n14079) );
  NAND2_X1 U8089 ( .A1(n12198), .A2(n12197), .ZN(n12202) );
  INV_X1 U8090 ( .A(n13821), .ZN(n14253) );
  NAND2_X1 U8091 ( .A1(n8628), .A2(n8627), .ZN(n14185) );
  NAND2_X1 U8092 ( .A1(n8615), .A2(n8614), .ZN(n11807) );
  AND2_X1 U8093 ( .A1(n9225), .A2(n9015), .ZN(n9924) );
  AND2_X1 U8094 ( .A1(n6662), .A2(n6887), .ZN(n6885) );
  NAND2_X1 U8095 ( .A1(n8732), .A2(n8731), .ZN(n8735) );
  AOI21_X1 U8096 ( .B1(n8288), .B2(n6979), .A(n6977), .ZN(n8658) );
  AND2_X1 U8097 ( .A1(n8299), .A2(n6789), .ZN(n6979) );
  NAND2_X1 U8098 ( .A1(n6806), .A2(n6978), .ZN(n6977) );
  OR2_X1 U8099 ( .A1(n8637), .A2(n10047), .ZN(n8655) );
  NAND2_X1 U8100 ( .A1(n8585), .A2(n8584), .ZN(n8600) );
  NAND2_X1 U8101 ( .A1(n7374), .A2(n8284), .ZN(n8578) );
  NAND2_X1 U8102 ( .A1(n8559), .A2(n8279), .ZN(n7374) );
  INV_X1 U8103 ( .A(n6968), .ZN(n8529) );
  AOI21_X1 U8104 ( .B1(n6973), .B2(n6971), .A(n6687), .ZN(n6968) );
  NAND2_X1 U8105 ( .A1(n8499), .A2(n8271), .ZN(n6973) );
  NAND2_X1 U8106 ( .A1(n8469), .A2(n8265), .ZN(n8488) );
  NAND2_X1 U8107 ( .A1(n8249), .A2(SI_5_), .ZN(n8251) );
  OAI21_X1 U8108 ( .B1(n8406), .B2(n7382), .A(n7380), .ZN(n8437) );
  NAND2_X1 U8109 ( .A1(n8394), .A2(n8248), .ZN(n8406) );
  NAND2_X1 U8110 ( .A1(n7047), .A2(n14400), .ZN(n14401) );
  NAND2_X1 U8111 ( .A1(n14441), .A2(n14440), .ZN(n7047) );
  INV_X1 U8112 ( .A(n6892), .ZN(n14410) );
  OAI21_X1 U8113 ( .B1(n14442), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6712), .ZN(
        n6892) );
  OAI21_X1 U8114 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14353), .A(n14352), .ZN(
        n14373) );
  AOI21_X1 U8115 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n15462), .A(n14357), .ZN(
        n14415) );
  OAI21_X1 U8116 ( .B1(n7039), .B2(n7038), .A(n7035), .ZN(n7043) );
  OAI21_X1 U8117 ( .B1(n14444), .B2(n14414), .A(n7041), .ZN(n7039) );
  NOR2_X1 U8118 ( .A1(n14449), .A2(n14429), .ZN(n14453) );
  AND3_X1 U8119 ( .A1(n8041), .A2(n8040), .A3(n8039), .ZN(n12650) );
  NAND2_X1 U8120 ( .A1(n9889), .A2(n8918), .ZN(n9888) );
  AND3_X1 U8121 ( .A1(n7843), .A2(n7842), .A3(n7841), .ZN(n15194) );
  XNOR2_X1 U8122 ( .A(n11883), .B(n11881), .ZN(n12430) );
  AND4_X1 U8123 ( .A1(n7774), .A2(n7773), .A3(n7772), .A4(n7771), .ZN(n10405)
         );
  INV_X1 U8124 ( .A(n13087), .ZN(n12457) );
  NAND2_X1 U8125 ( .A1(n8929), .A2(n12690), .ZN(n12459) );
  NAND2_X1 U8126 ( .A1(n8943), .A2(n8942), .ZN(n12451) );
  AOI21_X1 U8127 ( .B1(n12807), .B2(n6645), .A(n8096), .ZN(n12354) );
  AND3_X1 U8128 ( .A1(n8061), .A2(n8060), .A3(n8059), .ZN(n12656) );
  AND2_X1 U8129 ( .A1(n6951), .A2(n6950), .ZN(n9541) );
  NAND2_X1 U8130 ( .A1(n9519), .A2(n6952), .ZN(n6950) );
  NAND2_X1 U8131 ( .A1(n9520), .A2(n14949), .ZN(n6951) );
  OAI22_X1 U8132 ( .A1(n9541), .A2(n9540), .B1(n9539), .B2(n9543), .ZN(n9697)
         );
  OR2_X1 U8133 ( .A1(n10378), .A2(n10377), .ZN(n6854) );
  XNOR2_X1 U8134 ( .A(n10697), .B(n10698), .ZN(n10378) );
  INV_X1 U8135 ( .A(n15003), .ZN(n15087) );
  NOR2_X1 U8136 ( .A1(n14523), .A2(n7141), .ZN(n12736) );
  NOR2_X1 U8137 ( .A1(n14511), .A2(n12738), .ZN(n7141) );
  OAI21_X1 U8138 ( .B1(n6989), .B2(n15003), .A(n6988), .ZN(n6987) );
  INV_X1 U8139 ( .A(n12789), .ZN(n6988) );
  XNOR2_X1 U8140 ( .A(n6990), .B(n12788), .ZN(n6989) );
  INV_X1 U8141 ( .A(n11008), .ZN(n10926) );
  AND3_X1 U8142 ( .A1(n7786), .A2(n7785), .A3(n7784), .ZN(n15165) );
  AND3_X1 U8143 ( .A1(n7751), .A2(n7750), .A3(n7749), .ZN(n15155) );
  INV_X1 U8144 ( .A(n12998), .ZN(n14528) );
  NAND2_X1 U8145 ( .A1(n9941), .A2(n15108), .ZN(n15144) );
  NAND2_X1 U8146 ( .A1(n7918), .A2(n7917), .ZN(n13112) );
  AND2_X1 U8147 ( .A1(n8156), .A2(n7268), .ZN(n13134) );
  INV_X1 U8148 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7269) );
  INV_X1 U8149 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U8150 ( .A1(n7702), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7670) );
  XNOR2_X1 U8151 ( .A(n7584), .B(n7583), .ZN(n12769) );
  INV_X1 U8152 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7583) );
  OAI21_X1 U8153 ( .B1(n7942), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U8154 ( .A1(n10119), .A2(n10118), .ZN(n14887) );
  NAND2_X1 U8155 ( .A1(n10561), .A2(n10560), .ZN(n6841) );
  INV_X1 U8156 ( .A(n13493), .ZN(n13606) );
  NAND2_X1 U8157 ( .A1(n11263), .A2(n11262), .ZN(n13627) );
  NAND2_X1 U8158 ( .A1(n11510), .A2(n11509), .ZN(n13611) );
  OR2_X1 U8159 ( .A1(n12262), .A2(n11572), .ZN(n11510) );
  AND2_X1 U8160 ( .A1(n11537), .A2(n11536), .ZN(n13236) );
  NAND2_X1 U8161 ( .A1(n9463), .A2(n9462), .ZN(n13275) );
  INV_X1 U8162 ( .A(n13237), .ZN(n13469) );
  INV_X1 U8163 ( .A(n13236), .ZN(n13471) );
  OAI211_X1 U8164 ( .C1(n11218), .C2(n11551), .A(n10959), .B(n10958), .ZN(
        n13288) );
  NAND2_X1 U8165 ( .A1(n11685), .A2(n11684), .ZN(n13365) );
  XNOR2_X1 U8166 ( .A(n11924), .B(n11923), .ZN(n13565) );
  NAND2_X1 U8167 ( .A1(n13371), .A2(n11922), .ZN(n11924) );
  OR2_X1 U8168 ( .A1(n13368), .A2(n11955), .ZN(n7229) );
  AND2_X1 U8169 ( .A1(n11925), .A2(n13358), .ZN(n13563) );
  NAND2_X1 U8170 ( .A1(n11627), .A2(n11626), .ZN(n13567) );
  NAND2_X1 U8171 ( .A1(n13535), .A2(n11909), .ZN(n13518) );
  INV_X1 U8172 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12263) );
  XNOR2_X1 U8173 ( .A(n13695), .B(n13696), .ZN(n13697) );
  NAND2_X1 U8174 ( .A1(n13793), .A2(n12313), .ZN(n13695) );
  NAND2_X1 U8175 ( .A1(n10842), .A2(n10841), .ZN(n11119) );
  NAND2_X1 U8176 ( .A1(n8458), .A2(n8457), .ZN(n12067) );
  NAND2_X1 U8177 ( .A1(n8603), .A2(n8602), .ZN(n13761) );
  OR2_X1 U8178 ( .A1(n12262), .A2(n8369), .ZN(n8643) );
  NAND2_X1 U8179 ( .A1(n8505), .A2(n8504), .ZN(n14607) );
  AND2_X1 U8180 ( .A1(n7347), .A2(n6707), .ZN(n8370) );
  NAND4_X1 U8181 ( .A1(n8403), .A2(n8402), .A3(n8401), .A4(n8400), .ZN(n13837)
         );
  NAND2_X1 U8182 ( .A1(n12186), .A2(n12185), .ZN(n13985) );
  NAND2_X1 U8183 ( .A1(n7353), .A2(n7352), .ZN(n13987) );
  NAND2_X1 U8184 ( .A1(n13818), .A2(n14082), .ZN(n7352) );
  NAND2_X1 U8185 ( .A1(n8737), .A2(n8736), .ZN(n14200) );
  NAND2_X1 U8186 ( .A1(n14098), .A2(n8696), .ZN(n14078) );
  OR2_X1 U8187 ( .A1(n11573), .A2(n8369), .ZN(n8702) );
  NOR2_X1 U8188 ( .A1(n14204), .A2(n6830), .ZN(n14290) );
  NAND2_X1 U8189 ( .A1(n6832), .A2(n6831), .ZN(n6830) );
  INV_X1 U8190 ( .A(n14205), .ZN(n6831) );
  NAND2_X1 U8191 ( .A1(n14206), .A2(n14716), .ZN(n6832) );
  INV_X1 U8192 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10648) );
  XNOR2_X1 U8193 ( .A(n14410), .B(n7049), .ZN(n14443) );
  INV_X1 U8194 ( .A(n14411), .ZN(n7049) );
  NAND2_X1 U8195 ( .A1(n14626), .A2(n14625), .ZN(n14624) );
  NAND2_X1 U8196 ( .A1(n6890), .A2(n14624), .ZN(n14630) );
  OAI21_X1 U8197 ( .B1(n14626), .B2(n14625), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n6890) );
  NOR2_X1 U8198 ( .A1(n14630), .A2(n14631), .ZN(n14629) );
  XNOR2_X1 U8199 ( .A(n14453), .B(n14452), .ZN(n14451) );
  NAND2_X1 U8200 ( .A1(n11332), .A2(n11331), .ZN(n11330) );
  NAND2_X1 U8201 ( .A1(n13654), .A2(n11759), .ZN(n11329) );
  OR2_X1 U8202 ( .A1(n7475), .A2(n12054), .ZN(n7474) );
  INV_X1 U8203 ( .A(n11371), .ZN(n11372) );
  AND2_X1 U8204 ( .A1(n7452), .A2(n6880), .ZN(n6879) );
  NAND2_X1 U8205 ( .A1(n12068), .A2(n6881), .ZN(n6880) );
  OR2_X1 U8206 ( .A1(n12071), .A2(n7453), .ZN(n7450) );
  INV_X1 U8207 ( .A(n11420), .ZN(n7025) );
  NAND2_X1 U8208 ( .A1(n12084), .A2(n7458), .ZN(n7457) );
  OR2_X1 U8209 ( .A1(n12077), .A2(n12076), .ZN(n12081) );
  AND2_X1 U8210 ( .A1(n7459), .A2(n7456), .ZN(n7455) );
  NAND2_X1 U8211 ( .A1(n12083), .A2(n12085), .ZN(n7456) );
  NOR2_X1 U8212 ( .A1(n11434), .A2(n6720), .ZN(n7432) );
  NAND2_X1 U8213 ( .A1(n7021), .A2(n7020), .ZN(n11427) );
  OAI21_X1 U8214 ( .B1(n6752), .B2(n12123), .A(n14168), .ZN(n6872) );
  NAND2_X1 U8215 ( .A1(n12111), .A2(n6874), .ZN(n6873) );
  NAND2_X1 U8216 ( .A1(n7016), .A2(n7015), .ZN(n11455) );
  AOI21_X1 U8217 ( .B1(n6667), .B2(n7018), .A(n6755), .ZN(n7015) );
  NAND2_X1 U8218 ( .A1(n6703), .A2(n7415), .ZN(n7412) );
  NAND2_X1 U8219 ( .A1(n12136), .A2(n6867), .ZN(n6866) );
  INV_X1 U8220 ( .A(n12135), .ZN(n6867) );
  INV_X1 U8221 ( .A(n7412), .ZN(n7410) );
  INV_X1 U8222 ( .A(n12505), .ZN(n12590) );
  NAND2_X1 U8223 ( .A1(n7034), .A2(n6730), .ZN(n11486) );
  NAND2_X1 U8224 ( .A1(n7465), .A2(n7464), .ZN(n7463) );
  INV_X1 U8225 ( .A(n12151), .ZN(n7464) );
  NAND2_X1 U8226 ( .A1(n7028), .A2(n7027), .ZN(n7419) );
  NAND2_X1 U8227 ( .A1(n7422), .A2(n11540), .ZN(n7027) );
  INV_X1 U8228 ( .A(n11554), .ZN(n7417) );
  NAND2_X1 U8229 ( .A1(n12193), .A2(n7448), .ZN(n7447) );
  MUX2_X1 U8230 ( .A(n12666), .B(n12665), .S(n12672), .Z(n12667) );
  OR2_X1 U8231 ( .A1(n7986), .A2(n12913), .ZN(n7988) );
  NAND2_X1 U8232 ( .A1(n7009), .A2(n12571), .ZN(n7819) );
  OR2_X1 U8233 ( .A1(n11568), .A2(n11567), .ZN(n11569) );
  AND2_X1 U8234 ( .A1(n11568), .A2(n11567), .ZN(n11571) );
  NOR2_X1 U8235 ( .A1(n7281), .A2(n7280), .ZN(n7279) );
  INV_X1 U8236 ( .A(n10091), .ZN(n7280) );
  NAND2_X1 U8237 ( .A1(n10107), .A2(n10093), .ZN(n7277) );
  INV_X1 U8238 ( .A(n13752), .ZN(n7480) );
  INV_X1 U8239 ( .A(n12173), .ZN(n7470) );
  NAND2_X1 U8240 ( .A1(n12237), .A2(n7545), .ZN(n7543) );
  NAND2_X1 U8241 ( .A1(n14049), .A2(n14060), .ZN(n7544) );
  NOR2_X1 U8242 ( .A1(n7394), .A2(n7390), .ZN(n7389) );
  INV_X1 U8243 ( .A(n7399), .ZN(n7390) );
  INV_X1 U8244 ( .A(n11612), .ZN(n7394) );
  INV_X1 U8245 ( .A(n8639), .ZN(n8296) );
  NOR2_X1 U8246 ( .A1(n6687), .A2(n6967), .ZN(n6966) );
  INV_X1 U8247 ( .A(n8271), .ZN(n6967) );
  OR2_X1 U8248 ( .A1(n6971), .A2(n6687), .ZN(n6969) );
  INV_X1 U8249 ( .A(n7387), .ZN(n7386) );
  OAI21_X1 U8250 ( .B1(n8466), .B2(n7388), .A(n8267), .ZN(n7387) );
  INV_X1 U8251 ( .A(n8265), .ZN(n7388) );
  NOR2_X1 U8252 ( .A1(n14342), .A2(n14341), .ZN(n14343) );
  NOR2_X1 U8253 ( .A1(n14386), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n14342) );
  NOR2_X1 U8254 ( .A1(n9542), .A2(n7124), .ZN(n9702) );
  AND2_X1 U8255 ( .A1(n9543), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7124) );
  NAND2_X1 U8256 ( .A1(n15097), .A2(n12755), .ZN(n12756) );
  NAND2_X1 U8257 ( .A1(n15084), .A2(n12781), .ZN(n12782) );
  NOR2_X1 U8258 ( .A1(n14470), .A2(n12756), .ZN(n12757) );
  AND3_X1 U8259 ( .A1(n6857), .A2(n6855), .A3(n6822), .ZN(n12735) );
  INV_X1 U8260 ( .A(n12642), .ZN(n7014) );
  OR2_X1 U8261 ( .A1(n7863), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7876) );
  AND2_X1 U8262 ( .A1(n7819), .A2(n12557), .ZN(n10714) );
  NAND2_X1 U8263 ( .A1(n15171), .A2(n12714), .ZN(n12565) );
  NAND2_X1 U8264 ( .A1(n15139), .A2(n15126), .ZN(n15127) );
  NAND2_X1 U8265 ( .A1(n12719), .A2(n15124), .ZN(n12539) );
  INV_X1 U8266 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7668) );
  AOI21_X1 U8267 ( .B1(n6921), .B2(n6923), .A(n6821), .ZN(n6920) );
  INV_X1 U8268 ( .A(n6923), .ZN(n6922) );
  INV_X1 U8269 ( .A(n8005), .ZN(n7166) );
  INV_X1 U8270 ( .A(n7173), .ZN(n6918) );
  AND2_X1 U8271 ( .A1(n7915), .A2(n7639), .ZN(n7172) );
  AND2_X1 U8272 ( .A1(n7151), .A2(n6820), .ZN(n6919) );
  NOR2_X1 U8273 ( .A1(n7925), .A2(n7174), .ZN(n7173) );
  INV_X1 U8274 ( .A(n7636), .ZN(n7174) );
  NAND2_X1 U8275 ( .A1(n7144), .A2(n7143), .ZN(n7627) );
  AOI21_X1 U8276 ( .B1(n7146), .B2(n7148), .A(n6804), .ZN(n7143) );
  INV_X1 U8277 ( .A(n9850), .ZN(n7312) );
  NAND2_X1 U8278 ( .A1(n11696), .A2(n11697), .ZN(n11677) );
  INV_X1 U8279 ( .A(n11321), .ZN(n11322) );
  NAND2_X1 U8280 ( .A1(n11713), .A2(n11625), .ZN(n11747) );
  NAND2_X1 U8281 ( .A1(n9574), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7408) );
  INV_X1 U8282 ( .A(n13280), .ZN(n13266) );
  NOR2_X1 U8283 ( .A1(n13584), .A2(n7067), .ZN(n7066) );
  INV_X1 U8284 ( .A(n7068), .ZN(n7067) );
  INV_X1 U8285 ( .A(n11909), .ZN(n7275) );
  AND2_X1 U8286 ( .A1(n7212), .A2(n6770), .ZN(n7209) );
  INV_X1 U8287 ( .A(n7215), .ZN(n7207) );
  INV_X1 U8288 ( .A(n7285), .ZN(n7284) );
  OAI21_X1 U8289 ( .B1(n11740), .B2(n7224), .A(n11737), .ZN(n7223) );
  NOR2_X1 U8290 ( .A1(n10955), .A2(n10954), .ZN(n11075) );
  INV_X1 U8291 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U8292 ( .A1(n10275), .A2(n7198), .ZN(n7197) );
  INV_X1 U8293 ( .A(n10171), .ZN(n7198) );
  AND2_X1 U8294 ( .A1(n14881), .A2(n10445), .ZN(n10177) );
  INV_X1 U8295 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n15532) );
  NAND2_X1 U8296 ( .A1(n6809), .A2(n7056), .ZN(n10296) );
  INV_X1 U8297 ( .A(n7428), .ZN(n7427) );
  INV_X1 U8298 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U8299 ( .A1(n7054), .A2(n9056), .ZN(n7428) );
  NAND2_X1 U8300 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9049) );
  INV_X1 U8301 ( .A(n9806), .ZN(n7507) );
  INV_X1 U8302 ( .A(n11834), .ZN(n9346) );
  OR2_X1 U8303 ( .A1(n7481), .A2(n7480), .ZN(n7479) );
  OR2_X1 U8304 ( .A1(n7480), .A2(n11793), .ZN(n7478) );
  NOR2_X1 U8305 ( .A1(n14067), .A2(n14094), .ZN(n7093) );
  NAND2_X1 U8306 ( .A1(n6658), .A2(n8800), .ZN(n7363) );
  NOR2_X1 U8307 ( .A1(n14133), .A2(n7538), .ZN(n7537) );
  INV_X1 U8308 ( .A(n8653), .ZN(n7538) );
  NOR2_X1 U8309 ( .A1(n14175), .A2(n14185), .ZN(n7083) );
  NAND2_X1 U8310 ( .A1(n8621), .A2(n7553), .ZN(n7552) );
  INV_X1 U8311 ( .A(n7555), .ZN(n7553) );
  NOR2_X1 U8312 ( .A1(n6685), .A2(n7527), .ZN(n7526) );
  INV_X1 U8313 ( .A(n8372), .ZN(n7517) );
  NAND2_X1 U8314 ( .A1(n6649), .A2(n6883), .ZN(n12042) );
  NAND2_X1 U8315 ( .A1(n8775), .A2(n14335), .ZN(n12027) );
  NAND2_X1 U8316 ( .A1(n14136), .A2(n14234), .ZN(n14119) );
  NOR2_X1 U8317 ( .A1(n13815), .A2(n7085), .ZN(n7084) );
  INV_X1 U8318 ( .A(n7086), .ZN(n7085) );
  NAND2_X1 U8319 ( .A1(n9729), .A2(n12042), .ZN(n9978) );
  NAND2_X1 U8320 ( .A1(n8301), .A2(n8021), .ZN(n7401) );
  INV_X1 U8321 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U8322 ( .A1(n8299), .A2(n6981), .ZN(n6978) );
  NAND2_X1 U8323 ( .A1(n6983), .A2(n6980), .ZN(n8636) );
  AOI21_X1 U8324 ( .B1(n7375), .B2(n7377), .A(n6803), .ZN(n7372) );
  NAND2_X1 U8325 ( .A1(n8559), .A2(n7375), .ZN(n7373) );
  AOI21_X1 U8326 ( .B1(n8498), .B2(n8271), .A(n6972), .ZN(n6971) );
  INV_X1 U8327 ( .A(n8516), .ZN(n6972) );
  OR2_X1 U8328 ( .A1(n8257), .A2(n8256), .ZN(n8451) );
  AOI21_X1 U8329 ( .B1(n7380), .B2(n7382), .A(n6751), .ZN(n7378) );
  NAND2_X1 U8330 ( .A1(n8392), .A2(n8391), .ZN(n8394) );
  NAND2_X1 U8331 ( .A1(n8237), .A2(n8354), .ZN(n6942) );
  OR2_X1 U8332 ( .A1(n8237), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6941) );
  INV_X1 U8333 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6930) );
  OAI21_X1 U8334 ( .B1(n14377), .B2(n14378), .A(n6747), .ZN(n6893) );
  INV_X1 U8335 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14338) );
  XNOR2_X1 U8336 ( .A(n14343), .B(n14968), .ZN(n14376) );
  NOR2_X1 U8337 ( .A1(n14350), .A2(n14349), .ZN(n14375) );
  AND2_X1 U8338 ( .A1(n14414), .A2(n14444), .ZN(n7036) );
  NAND2_X1 U8339 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7040) );
  OR2_X1 U8340 ( .A1(n11295), .A2(n11303), .ZN(n7253) );
  AND2_X1 U8341 ( .A1(n7230), .A2(n8913), .ZN(n9794) );
  NOR2_X1 U8342 ( .A1(n12376), .A2(n7260), .ZN(n7259) );
  INV_X1 U8343 ( .A(n11876), .ZN(n7260) );
  OR2_X1 U8344 ( .A1(n8045), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U8345 ( .A1(n10596), .A2(n10595), .ZN(n7255) );
  OR2_X1 U8346 ( .A1(n8011), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U8347 ( .A1(n7695), .A2(n12431), .ZN(n8037) );
  INV_X1 U8348 ( .A(n8024), .ZN(n7695) );
  NAND2_X1 U8349 ( .A1(n7262), .A2(n6784), .ZN(n7261) );
  NAND2_X1 U8350 ( .A1(n11030), .A2(n7263), .ZN(n11137) );
  NOR2_X1 U8351 ( .A1(n7264), .A2(n6784), .ZN(n7263) );
  INV_X1 U8352 ( .A(n11029), .ZN(n7264) );
  INV_X1 U8353 ( .A(n8915), .ZN(n15106) );
  NAND2_X1 U8354 ( .A1(n7692), .A2(n7691), .ZN(n7933) );
  INV_X1 U8355 ( .A(n7947), .ZN(n7692) );
  OAI21_X1 U8356 ( .B1(n9506), .B2(n6850), .A(n9497), .ZN(n9498) );
  NOR2_X1 U8357 ( .A1(n9496), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n6850) );
  NOR2_X1 U8358 ( .A1(n9498), .A2(n15143), .ZN(n9522) );
  NOR2_X1 U8359 ( .A1(n9526), .A2(n9525), .ZN(n9542) );
  XNOR2_X1 U8360 ( .A(n9707), .B(n6995), .ZN(n9710) );
  XNOR2_X1 U8361 ( .A(n9702), .B(n9708), .ZN(n9544) );
  NOR2_X1 U8362 ( .A1(n9544), .A2(n9545), .ZN(n9703) );
  NAND2_X1 U8363 ( .A1(n10381), .A2(n10382), .ZN(n14974) );
  NAND2_X1 U8364 ( .A1(n10387), .A2(n10388), .ZN(n14980) );
  NAND2_X1 U8365 ( .A1(n14980), .A2(n14981), .ZN(n14979) );
  AND2_X1 U8366 ( .A1(n14979), .A2(n6959), .ZN(n10680) );
  NAND2_X1 U8367 ( .A1(n10390), .A2(n10389), .ZN(n6959) );
  AND2_X1 U8368 ( .A1(n6854), .A2(n6761), .ZN(n14992) );
  NAND2_X1 U8369 ( .A1(n10690), .A2(n10691), .ZN(n14994) );
  AOI21_X1 U8370 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10701), .A(n14990), .ZN(
        n10703) );
  XNOR2_X1 U8371 ( .A(n10692), .B(n10702), .ZN(n15022) );
  NAND2_X1 U8372 ( .A1(n6851), .A2(n7132), .ZN(n12721) );
  AND3_X1 U8373 ( .A1(n6851), .A2(n7132), .A3(n6815), .ZN(n12723) );
  NAND2_X1 U8374 ( .A1(n15029), .A2(n12777), .ZN(n15050) );
  AND2_X1 U8375 ( .A1(n15044), .A2(n12726), .ZN(n12727) );
  NAND2_X1 U8376 ( .A1(n15067), .A2(n12780), .ZN(n15086) );
  NAND2_X1 U8377 ( .A1(n15086), .A2(n15085), .ZN(n15084) );
  XNOR2_X1 U8378 ( .A(n12782), .B(n7970), .ZN(n14466) );
  AND2_X1 U8379 ( .A1(n7967), .A2(n7968), .ZN(n7955) );
  OAI21_X1 U8380 ( .B1(n14485), .B2(n14481), .A(n14483), .ZN(n14502) );
  NOR2_X1 U8381 ( .A1(n14502), .A2(n14501), .ZN(n14500) );
  XNOR2_X1 U8382 ( .A(n12763), .B(n12770), .ZN(n14517) );
  OR2_X1 U8383 ( .A1(n14505), .A2(n15481), .ZN(n7142) );
  NOR2_X1 U8384 ( .A1(n14500), .A2(n12762), .ZN(n12763) );
  NAND2_X1 U8385 ( .A1(n14512), .A2(n6991), .ZN(n6990) );
  OR2_X1 U8386 ( .A1(n14511), .A2(n13050), .ZN(n6991) );
  NAND2_X1 U8387 ( .A1(n6928), .A2(n12528), .ZN(n12462) );
  OR2_X1 U8388 ( .A1(n6997), .A2(n12529), .ZN(n6928) );
  OAI21_X1 U8389 ( .B1(n8063), .B2(n6998), .A(n6754), .ZN(n6997) );
  NAND2_X1 U8390 ( .A1(n8131), .A2(n12802), .ZN(n8132) );
  AND2_X1 U8391 ( .A1(n12528), .A2(n8133), .ZN(n12800) );
  OR2_X1 U8392 ( .A1(n8070), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8081) );
  AOI21_X1 U8393 ( .B1(n7106), .B2(n12498), .A(n7105), .ZN(n7104) );
  NOR2_X1 U8394 ( .A1(n13100), .A2(n11885), .ZN(n7105) );
  INV_X1 U8395 ( .A(n7109), .ZN(n7108) );
  OAI21_X1 U8396 ( .B1(n7111), .B2(n7952), .A(n8124), .ZN(n7109) );
  AND4_X1 U8397 ( .A1(n7937), .A2(n7936), .A3(n7935), .A4(n7934), .ZN(n12918)
         );
  OR2_X1 U8398 ( .A1(n12927), .A2(n7111), .ZN(n12916) );
  NOR2_X1 U8399 ( .A1(n12928), .A2(n12936), .ZN(n12927) );
  OR2_X1 U8400 ( .A1(n7960), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7947) );
  INV_X1 U8401 ( .A(n12517), .ZN(n12953) );
  AOI21_X1 U8402 ( .B1(n7097), .B2(n7099), .A(n7096), .ZN(n7095) );
  NOR2_X1 U8403 ( .A1(n13121), .A2(n12405), .ZN(n7096) );
  OR2_X1 U8404 ( .A1(n7975), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7977) );
  AND2_X1 U8405 ( .A1(n12608), .A2(n12964), .ZN(n12978) );
  NOR2_X1 U8406 ( .A1(n11149), .A2(n7565), .ZN(n12989) );
  NOR2_X1 U8407 ( .A1(n11150), .A2(n12599), .ZN(n11149) );
  NAND2_X1 U8408 ( .A1(n7116), .A2(n8110), .ZN(n8111) );
  OR2_X1 U8409 ( .A1(n7787), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U8410 ( .A1(n10503), .A2(n8104), .ZN(n10481) );
  NAND2_X1 U8411 ( .A1(n8097), .A2(n8103), .ZN(n10478) );
  INV_X1 U8412 ( .A(n15136), .ZN(n12990) );
  AND4_X1 U8413 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n10501)
         );
  INV_X1 U8414 ( .A(n12502), .ZN(n15114) );
  NAND2_X1 U8415 ( .A1(n15105), .A2(n15114), .ZN(n15104) );
  INV_X1 U8416 ( .A(n12769), .ZN(n12525) );
  AND4_X2 U8417 ( .A1(n7733), .A2(n7732), .A3(n7731), .A4(n7730), .ZN(n15135)
         );
  NAND2_X1 U8418 ( .A1(n12539), .A2(n12541), .ZN(n15139) );
  AND2_X1 U8419 ( .A1(n12472), .A2(n12471), .ZN(n12794) );
  NAND2_X1 U8420 ( .A1(n8023), .A2(n8022), .ZN(n11880) );
  OR2_X1 U8421 ( .A1(n7882), .A2(n8021), .ZN(n8022) );
  NAND2_X1 U8422 ( .A1(n10802), .A2(n12672), .ZN(n15136) );
  INV_X1 U8423 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7156) );
  NAND2_X1 U8424 ( .A1(n8182), .A2(n6684), .ZN(n9492) );
  AND2_X1 U8425 ( .A1(n7646), .A2(n7645), .ZN(n8019) );
  OR2_X1 U8426 ( .A1(n7940), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n7942) );
  INV_X1 U8427 ( .A(n7157), .ZN(n6912) );
  OR2_X1 U8428 ( .A1(n7779), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7781) );
  NOR2_X1 U8429 ( .A1(n7781), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7795) );
  XNOR2_X1 U8430 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7727) );
  NAND2_X1 U8431 ( .A1(n6915), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7726) );
  INV_X1 U8432 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6915) );
  AND2_X1 U8433 ( .A1(n7315), .A2(n10950), .ZN(n7314) );
  NAND2_X1 U8434 ( .A1(n7316), .A2(n7320), .ZN(n10942) );
  NAND2_X1 U8435 ( .A1(n10651), .A2(n7321), .ZN(n7316) );
  AND2_X1 U8436 ( .A1(n11075), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11173) );
  NOR2_X1 U8437 ( .A1(n11721), .A2(n6654), .ZN(n9647) );
  NAND2_X1 U8438 ( .A1(n10650), .A2(n7325), .ZN(n7324) );
  INV_X1 U8439 ( .A(n10652), .ZN(n7325) );
  AND2_X1 U8440 ( .A1(n13203), .A2(n13202), .ZN(n13205) );
  INV_X1 U8441 ( .A(n13286), .ZN(n13539) );
  NAND2_X1 U8442 ( .A1(n6656), .A2(n13349), .ZN(n11764) );
  NOR3_X1 U8444 ( .A1(n14771), .A2(n9464), .A3(n9065), .ZN(n14772) );
  NOR2_X1 U8445 ( .A1(n14788), .A2(n14787), .ZN(n14786) );
  NOR2_X1 U8446 ( .A1(n14804), .A2(n14803), .ZN(n14802) );
  NOR2_X1 U8447 ( .A1(n10317), .A2(n10316), .ZN(n10543) );
  AND2_X1 U8448 ( .A1(n11922), .A2(n11720), .ZN(n13372) );
  AND2_X1 U8449 ( .A1(n11657), .A2(n11656), .ZN(n13405) );
  NAND2_X1 U8450 ( .A1(n6935), .A2(n6671), .ZN(n6934) );
  NAND2_X1 U8451 ( .A1(n13475), .A2(n7066), .ZN(n13412) );
  NAND2_X1 U8452 ( .A1(n11942), .A2(n11941), .ZN(n13430) );
  AND2_X1 U8453 ( .A1(n13488), .A2(n13481), .ZN(n13475) );
  NAND2_X1 U8454 ( .A1(n13475), .A2(n13463), .ZN(n13457) );
  AOI21_X1 U8455 ( .B1(n7187), .B2(n7189), .A(n6737), .ZN(n7185) );
  NOR2_X1 U8456 ( .A1(n13611), .A2(n13523), .ZN(n13508) );
  NAND2_X1 U8457 ( .A1(n11908), .A2(n7273), .ZN(n6944) );
  NAND2_X1 U8458 ( .A1(n7061), .A2(n7060), .ZN(n13523) );
  NOR3_X1 U8459 ( .A1(n13627), .A2(n7063), .A3(n13616), .ZN(n7060) );
  AND2_X1 U8460 ( .A1(n7061), .A2(n7059), .ZN(n13548) );
  NOR2_X1 U8461 ( .A1(n7063), .A2(n13627), .ZN(n7059) );
  NAND2_X1 U8462 ( .A1(n7211), .A2(n11932), .ZN(n13537) );
  OR2_X1 U8463 ( .A1(n11934), .A2(n11933), .ZN(n7211) );
  OR2_X1 U8464 ( .A1(n13637), .A2(n11217), .ZN(n11215) );
  OR2_X1 U8465 ( .A1(n10767), .A2(n10766), .ZN(n10955) );
  NAND2_X1 U8466 ( .A1(n7200), .A2(n7202), .ZN(n11016) );
  INV_X1 U8467 ( .A(n7203), .ZN(n7202) );
  OAI21_X1 U8468 ( .B1(n10754), .B2(n7204), .A(n11014), .ZN(n7203) );
  NOR2_X1 U8469 ( .A1(n14558), .A2(n7071), .ZN(n7070) );
  NAND2_X1 U8470 ( .A1(n7075), .A2(n7074), .ZN(n7071) );
  NAND2_X1 U8471 ( .A1(n7290), .A2(n7293), .ZN(n11010) );
  NAND2_X1 U8472 ( .A1(n10368), .A2(n7073), .ZN(n14561) );
  NOR2_X1 U8473 ( .A1(n14558), .A2(n7072), .ZN(n7073) );
  INV_X1 U8474 ( .A(n7074), .ZN(n7072) );
  OR2_X1 U8475 ( .A1(n10357), .A2(n15532), .ZN(n10522) );
  INV_X1 U8476 ( .A(n7178), .ZN(n10747) );
  AOI21_X1 U8477 ( .B1(n10356), .B2(n7179), .A(n7182), .ZN(n7178) );
  INV_X1 U8478 ( .A(n7183), .ZN(n7179) );
  NAND2_X1 U8479 ( .A1(n10368), .A2(n14910), .ZN(n10534) );
  NAND2_X1 U8480 ( .A1(n10350), .A2(n10349), .ZN(n10512) );
  AOI21_X1 U8481 ( .B1(n10287), .B2(n7195), .A(n6735), .ZN(n7194) );
  OR2_X1 U8482 ( .A1(n10121), .A2(n10120), .ZN(n10213) );
  OR2_X1 U8483 ( .A1(n9856), .A2(n9855), .ZN(n10121) );
  NAND2_X1 U8484 ( .A1(n7196), .A2(n7199), .ZN(n10291) );
  NAND2_X1 U8485 ( .A1(n10172), .A2(n7197), .ZN(n7196) );
  NOR2_X1 U8486 ( .A1(n10459), .A2(n14874), .ZN(n10445) );
  NAND2_X1 U8487 ( .A1(n10092), .A2(n10091), .ZN(n10457) );
  INV_X1 U8488 ( .A(n11722), .ZN(n10227) );
  INV_X1 U8489 ( .A(n13470), .ZN(n13538) );
  NAND2_X1 U8490 ( .A1(n9061), .A2(n9460), .ZN(n13540) );
  AND2_X1 U8491 ( .A1(n13378), .A2(n13377), .ZN(n13566) );
  NAND2_X1 U8492 ( .A1(n11600), .A2(n11599), .ZN(n13573) );
  INV_X1 U8493 ( .A(n11392), .ZN(n14881) );
  NAND2_X1 U8494 ( .A1(n11764), .A2(n13653), .ZN(n14909) );
  INV_X1 U8495 ( .A(n14909), .ZN(n14917) );
  AND2_X1 U8496 ( .A1(n9441), .A2(n10010), .ZN(n9442) );
  INV_X1 U8497 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9441) );
  AND2_X1 U8498 ( .A1(n8988), .A2(n9038), .ZN(n9848) );
  OR2_X1 U8499 ( .A1(n8973), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U8500 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  OR2_X1 U8501 ( .A1(n12281), .A2(n12280), .ZN(n13706) );
  AND2_X1 U8502 ( .A1(n6716), .A2(n11827), .ZN(n7512) );
  AOI21_X1 U8503 ( .B1(n13696), .B2(n12312), .A(n12321), .ZN(n7489) );
  INV_X1 U8504 ( .A(n7489), .ZN(n7487) );
  NAND2_X1 U8505 ( .A1(n7482), .A2(n6695), .ZN(n13740) );
  AND2_X1 U8506 ( .A1(n13734), .A2(n12291), .ZN(n13765) );
  NAND2_X1 U8507 ( .A1(n7505), .A2(n7507), .ZN(n7504) );
  INV_X1 U8508 ( .A(n9804), .ZN(n7505) );
  AND2_X1 U8509 ( .A1(n9804), .A2(n9806), .ZN(n7508) );
  OR2_X1 U8510 ( .A1(n8460), .A2(n8459), .ZN(n8479) );
  AND2_X1 U8511 ( .A1(n13702), .A2(n11843), .ZN(n11845) );
  OR2_X1 U8512 ( .A1(n8533), .A2(n9030), .ZN(n7347) );
  NAND2_X1 U8513 ( .A1(n13736), .A2(n12304), .ZN(n13794) );
  AND2_X1 U8514 ( .A1(n12022), .A2(n14335), .ZN(n12201) );
  NAND2_X1 U8515 ( .A1(n6869), .A2(n6673), .ZN(n12208) );
  NOR2_X1 U8516 ( .A1(n12204), .A2(n6700), .ZN(n12247) );
  INV_X1 U8517 ( .A(n12178), .ZN(n8720) );
  INV_X1 U8518 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n13925) );
  OR3_X1 U8519 ( .A1(n8502), .A2(P1_IR_REG_10__SCAN_IN), .A3(n8501), .ZN(n8517) );
  NOR2_X1 U8520 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7466) );
  OR2_X1 U8521 ( .A1(n14032), .A2(n14042), .ZN(n6826) );
  NAND2_X1 U8522 ( .A1(n14113), .A2(n7093), .ZN(n14065) );
  NAND2_X1 U8523 ( .A1(n14113), .A2(n14091), .ZN(n14090) );
  NOR2_X1 U8524 ( .A1(n15519), .A2(n8687), .ZN(n8705) );
  OR2_X1 U8525 ( .A1(n14234), .A2(n13819), .ZN(n14104) );
  NAND2_X1 U8526 ( .A1(n14127), .A2(n14126), .ZN(n14125) );
  NOR2_X1 U8527 ( .A1(n14151), .A2(n14303), .ZN(n14136) );
  NAND2_X1 U8528 ( .A1(n7083), .A2(n7082), .ZN(n14151) );
  INV_X1 U8529 ( .A(n7083), .ZN(n14177) );
  INV_X1 U8530 ( .A(n7550), .ZN(n14174) );
  OAI21_X1 U8531 ( .B1(n11096), .B2(n7554), .A(n7551), .ZN(n7550) );
  NAND2_X1 U8532 ( .A1(n8621), .A2(n7558), .ZN(n7554) );
  AND2_X1 U8533 ( .A1(n6771), .A2(n7552), .ZN(n7551) );
  NOR2_X1 U8534 ( .A1(n7357), .A2(n7356), .ZN(n7355) );
  INV_X1 U8535 ( .A(n12108), .ZN(n7356) );
  NOR2_X1 U8536 ( .A1(n6663), .A2(n6699), .ZN(n7357) );
  OR2_X1 U8537 ( .A1(n11098), .A2(n14276), .ZN(n11157) );
  NOR2_X1 U8538 ( .A1(n11157), .A2(n13761), .ZN(n11287) );
  OR2_X1 U8539 ( .A1(n13815), .A2(n8575), .ZN(n12102) );
  NAND2_X1 U8540 ( .A1(n10576), .A2(n7088), .ZN(n10826) );
  NAND2_X1 U8541 ( .A1(n10576), .A2(n11135), .ZN(n10641) );
  NAND2_X1 U8542 ( .A1(n7531), .A2(n7530), .ZN(n10575) );
  AOI21_X1 U8543 ( .B1(n6660), .B2(n7533), .A(n6732), .ZN(n7530) );
  NAND2_X1 U8544 ( .A1(n7081), .A2(n7080), .ZN(n10420) );
  INV_X1 U8545 ( .A(n14663), .ZN(n7081) );
  NOR2_X1 U8546 ( .A1(n8479), .A2(n13925), .ZN(n8506) );
  NAND2_X1 U8547 ( .A1(n8477), .A2(n8476), .ZN(n14671) );
  NAND2_X1 U8548 ( .A1(n10024), .A2(n10068), .ZN(n14662) );
  NOR2_X1 U8549 ( .A1(n10052), .A2(n12064), .ZN(n10024) );
  NAND2_X1 U8550 ( .A1(n8784), .A2(n8783), .ZN(n10058) );
  NAND2_X1 U8551 ( .A1(n9947), .A2(n12211), .ZN(n9946) );
  INV_X1 U8552 ( .A(n6845), .ZN(n6844) );
  NAND2_X1 U8553 ( .A1(n12196), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6846) );
  OAI21_X1 U8554 ( .B1(n9036), .B2(n8369), .A(n8348), .ZN(n6845) );
  NAND2_X1 U8555 ( .A1(n9921), .A2(n9920), .ZN(n13990) );
  OR2_X1 U8556 ( .A1(n12214), .A2(n9990), .ZN(n9991) );
  XNOR2_X1 U8557 ( .A(n9350), .B(n12034), .ZN(n12214) );
  AND2_X1 U8558 ( .A1(n14015), .A2(n14014), .ZN(n14199) );
  AND2_X1 U8559 ( .A1(n14063), .A2(n14062), .ZN(n14215) );
  NAND2_X1 U8560 ( .A1(n7077), .A2(n14722), .ZN(n9981) );
  AND2_X1 U8561 ( .A1(n8860), .A2(n12023), .ZN(n14743) );
  OAI22_X1 U8562 ( .A1(n11680), .A2(n11681), .B1(n11615), .B2(n12464), .ZN(
        n11618) );
  XNOR2_X1 U8563 ( .A(n11680), .B(n11682), .ZN(n12266) );
  INV_X1 U8564 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8218) );
  NOR2_X1 U8565 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n6886) );
  XNOR2_X1 U8566 ( .A(n6961), .B(n11612), .ZN(n13682) );
  NAND2_X1 U8567 ( .A1(n7398), .A2(n7395), .ZN(n6961) );
  NAND2_X1 U8568 ( .A1(n8323), .A2(n8322), .ZN(n14328) );
  MUX2_X1 U8569 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8320), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n8323) );
  NOR2_X1 U8570 ( .A1(n8827), .A2(n8317), .ZN(n8828) );
  INV_X1 U8571 ( .A(n8829), .ZN(n8831) );
  AND2_X1 U8572 ( .A1(n8715), .A2(n8714), .ZN(n11651) );
  NAND2_X1 U8573 ( .A1(n6975), .A2(n8315), .ZN(n8715) );
  INV_X1 U8574 ( .A(n6976), .ZN(n6975) );
  INV_X1 U8575 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8826) );
  XNOR2_X1 U8576 ( .A(n6688), .B(n8336), .ZN(n11587) );
  OAI21_X1 U8577 ( .B1(n8683), .B2(n8305), .A(n8307), .ZN(n8698) );
  INV_X1 U8578 ( .A(n8681), .ZN(n8306) );
  NAND2_X1 U8579 ( .A1(n8842), .A2(n8841), .ZN(n8984) );
  NAND2_X1 U8580 ( .A1(n8825), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8840) );
  NAND2_X1 U8581 ( .A1(n7401), .A2(n8304), .ZN(n8669) );
  NAND2_X1 U8582 ( .A1(n6983), .A2(n6984), .ZN(n8623) );
  NAND2_X1 U8583 ( .A1(n7403), .A2(n7402), .ZN(n8611) );
  NAND2_X1 U8584 ( .A1(n8289), .A2(n15493), .ZN(n7402) );
  NOR2_X1 U8585 ( .A1(n8586), .A2(n7467), .ZN(n10880) );
  OR2_X1 U8586 ( .A1(n8499), .A2(n8498), .ZN(n6970) );
  NAND2_X1 U8587 ( .A1(n8467), .A2(n8466), .ZN(n8469) );
  XNOR2_X1 U8588 ( .A(n8439), .B(n8438), .ZN(n10116) );
  AND2_X1 U8589 ( .A1(n8426), .A2(n8425), .ZN(n9137) );
  AND2_X1 U8590 ( .A1(n7050), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14380) );
  XNOR2_X1 U8591 ( .A(n7051), .B(n14380), .ZN(n14381) );
  XNOR2_X1 U8592 ( .A(n7052), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n7051) );
  XNOR2_X1 U8593 ( .A(n6893), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14386) );
  NAND2_X1 U8594 ( .A1(n6889), .A2(n6696), .ZN(n6888) );
  OR2_X1 U8595 ( .A1(n15607), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6889) );
  NOR2_X1 U8596 ( .A1(n14346), .A2(n14345), .ZN(n14397) );
  INV_X1 U8597 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U8598 ( .A1(n14404), .A2(n14405), .ZN(n14406) );
  AOI21_X1 U8599 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n14355), .A(n14354), .ZN(
        n14371) );
  OAI21_X1 U8600 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15053), .A(n14358), .ZN(
        n14368) );
  NAND2_X1 U8601 ( .A1(n14421), .A2(n6899), .ZN(n6895) );
  AOI21_X1 U8602 ( .B1(n14422), .B2(n6897), .A(n6743), .ZN(n6896) );
  INV_X1 U8603 ( .A(n6902), .ZN(n6899) );
  AOI21_X1 U8604 ( .B1(n7240), .B2(n6669), .A(n6800), .ZN(n7237) );
  NAND2_X1 U8605 ( .A1(n11884), .A2(n6714), .ZN(n7236) );
  NAND2_X1 U8606 ( .A1(n8080), .A2(n8079), .ZN(n12822) );
  NAND2_X1 U8607 ( .A1(n7248), .A2(n7252), .ZN(n11308) );
  NAND2_X1 U8608 ( .A1(n11296), .A2(n7253), .ZN(n7248) );
  NAND2_X1 U8609 ( .A1(n12423), .A2(n11876), .ZN(n12375) );
  NAND2_X1 U8610 ( .A1(n7244), .A2(n11890), .ZN(n12382) );
  NAND2_X1 U8611 ( .A1(n7231), .A2(n7239), .ZN(n7244) );
  INV_X1 U8612 ( .A(n11891), .ZN(n7239) );
  NAND2_X1 U8613 ( .A1(n11861), .A2(n11860), .ZN(n12395) );
  INV_X1 U8614 ( .A(n12946), .ZN(n12405) );
  NAND2_X1 U8615 ( .A1(n12393), .A2(n11865), .ZN(n12403) );
  NAND2_X1 U8616 ( .A1(n8044), .A2(n8043), .ZN(n13021) );
  OR2_X1 U8617 ( .A1(n7882), .A2(n10897), .ZN(n8043) );
  NAND2_X1 U8618 ( .A1(n7255), .A2(n10605), .ZN(n10608) );
  NAND2_X1 U8619 ( .A1(n12425), .A2(n12424), .ZN(n12423) );
  NAND2_X1 U8620 ( .A1(n7261), .A2(n11137), .ZN(n11032) );
  AND4_X1 U8621 ( .A1(n7951), .A2(n7950), .A3(n7949), .A4(n7948), .ZN(n12930)
         );
  AND4_X1 U8622 ( .A1(n7807), .A2(n7806), .A3(n7805), .A4(n7804), .ZN(n12575)
         );
  NAND2_X1 U8623 ( .A1(n7233), .A2(n6729), .ZN(n7232) );
  NAND2_X1 U8624 ( .A1(n7247), .A2(n7245), .ZN(n11856) );
  AOI21_X1 U8625 ( .B1(n7249), .B2(n7251), .A(n7246), .ZN(n7245) );
  INV_X1 U8626 ( .A(n11309), .ZN(n7246) );
  INV_X1 U8627 ( .A(n9517), .ZN(n12693) );
  INV_X1 U8628 ( .A(n12353), .ZN(n12702) );
  INV_X1 U8629 ( .A(n12921), .ZN(n12706) );
  INV_X1 U8630 ( .A(n12930), .ZN(n12707) );
  NAND2_X1 U8631 ( .A1(n8138), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7114) );
  AND2_X1 U8632 ( .A1(n7853), .A2(n7852), .ZN(n7113) );
  INV_X1 U8633 ( .A(n10723), .ZN(n12714) );
  INV_X1 U8634 ( .A(n10501), .ZN(n12716) );
  INV_X1 U8635 ( .A(n15112), .ZN(n12719) );
  INV_X1 U8636 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14952) );
  XNOR2_X1 U8637 ( .A(n9518), .B(n6952), .ZN(n9520) );
  OAI21_X1 U8638 ( .B1(n7736), .B2(n7131), .A(n7129), .ZN(n7128) );
  NAND2_X1 U8639 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7131) );
  NOR2_X1 U8640 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7736) );
  AOI21_X1 U8641 ( .B1(n9697), .B2(n9696), .A(n6949), .ZN(n14954) );
  AND2_X1 U8642 ( .A1(n9695), .A2(n9708), .ZN(n6949) );
  NAND2_X1 U8643 ( .A1(n10373), .A2(n6694), .ZN(n10374) );
  OR2_X1 U8644 ( .A1(n6697), .A2(n10385), .ZN(n7127) );
  INV_X1 U8645 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14989) );
  XNOR2_X1 U8646 ( .A(n10703), .B(n10702), .ZN(n15011) );
  NOR2_X1 U8647 ( .A1(n15011), .A2(n15012), .ZN(n15010) );
  XNOR2_X1 U8648 ( .A(n12723), .B(n12775), .ZN(n15028) );
  NOR2_X1 U8649 ( .A1(n15028), .A2(n15498), .ZN(n15027) );
  NOR2_X1 U8650 ( .A1(n15036), .A2(n6953), .ZN(n15060) );
  AND2_X1 U8651 ( .A1(n12744), .A2(n12775), .ZN(n6953) );
  NAND2_X1 U8652 ( .A1(n15060), .A2(n15059), .ZN(n15058) );
  OR2_X1 U8653 ( .A1(n12726), .A2(n12749), .ZN(n7126) );
  NOR2_X1 U8654 ( .A1(n15074), .A2(n6948), .ZN(n15099) );
  AND2_X1 U8655 ( .A1(n12748), .A2(n12749), .ZN(n6948) );
  NAND2_X1 U8656 ( .A1(n15099), .A2(n15098), .ZN(n15097) );
  NAND2_X1 U8657 ( .A1(n6857), .A2(n6855), .ZN(n14492) );
  INV_X1 U8658 ( .A(n12733), .ZN(n6860) );
  NAND2_X1 U8659 ( .A1(n12805), .A2(n7570), .ZN(n8137) );
  XNOR2_X1 U8660 ( .A(n12462), .B(n12521), .ZN(n12336) );
  NAND2_X1 U8661 ( .A1(n8063), .A2(n12655), .ZN(n12831) );
  NAND2_X1 U8662 ( .A1(n8055), .A2(n8054), .ZN(n12845) );
  NAND2_X1 U8663 ( .A1(n12866), .A2(n12530), .ZN(n12855) );
  OAI21_X1 U8664 ( .B1(n12887), .B2(n12498), .A(n12499), .ZN(n12877) );
  NAND2_X1 U8665 ( .A1(n13039), .A2(n12638), .ZN(n12891) );
  OR2_X1 U8666 ( .A1(n12907), .A2(n12906), .ZN(n13039) );
  NAND2_X1 U8667 ( .A1(n7997), .A2(n7996), .ZN(n12905) );
  OAI21_X1 U8668 ( .B1(n11150), .B2(n7099), .A(n7098), .ZN(n12961) );
  NAND2_X1 U8669 ( .A1(n7011), .A2(n12596), .ZN(n11148) );
  INV_X1 U8670 ( .A(n11136), .ZN(n14535) );
  OR2_X1 U8671 ( .A1(n7882), .A2(n15521), .ZN(n7873) );
  AND3_X1 U8672 ( .A1(n7816), .A2(n7815), .A3(n7814), .ZN(n12534) );
  OR2_X1 U8673 ( .A1(n7882), .A2(n8996), .ZN(n7801) );
  NAND2_X1 U8674 ( .A1(n12848), .A2(n10397), .ZN(n15141) );
  NAND2_X1 U8675 ( .A1(n12690), .A2(n9938), .ZN(n15108) );
  OR2_X1 U8676 ( .A1(n9941), .A2(n9940), .ZN(n12998) );
  AND2_X2 U8677 ( .A1(n9936), .A2(n8196), .ZN(n15213) );
  INV_X1 U8678 ( .A(n12493), .ZN(n13076) );
  NOR2_X1 U8679 ( .A1(n12794), .A2(n12793), .ZN(n14531) );
  AND2_X1 U8680 ( .A1(n7678), .A2(n7677), .ZN(n12339) );
  OR2_X1 U8681 ( .A1(n7882), .A2(n13142), .ZN(n7677) );
  INV_X1 U8682 ( .A(n8136), .ZN(n13080) );
  OAI21_X1 U8683 ( .B1(n15172), .B2(n13006), .A(n13005), .ZN(n13077) );
  INV_X1 U8684 ( .A(n12822), .ZN(n8131) );
  AND2_X1 U8685 ( .A1(n8069), .A2(n8068), .ZN(n13087) );
  OR2_X1 U8686 ( .A1(n7882), .A2(n15444), .ZN(n8068) );
  INV_X1 U8687 ( .A(n12845), .ZN(n13091) );
  INV_X1 U8688 ( .A(n12651), .ZN(n13096) );
  INV_X1 U8689 ( .A(n11880), .ZN(n13100) );
  INV_X1 U8690 ( .A(n11877), .ZN(n13104) );
  INV_X1 U8691 ( .A(n12905), .ZN(n13108) );
  INV_X1 U8692 ( .A(n11869), .ZN(n13116) );
  NAND2_X1 U8693 ( .A1(n7896), .A2(n7895), .ZN(n13130) );
  NAND2_X1 U8694 ( .A1(n7862), .A2(n6728), .ZN(n11008) );
  INV_X1 U8695 ( .A(n8099), .ZN(n9943) );
  NAND2_X1 U8696 ( .A1(n15197), .A2(n15193), .ZN(n13131) );
  AND2_X1 U8697 ( .A1(n8158), .A2(n8157), .ZN(n13132) );
  NAND2_X1 U8698 ( .A1(n9492), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13133) );
  INV_X1 U8699 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n7700) );
  INV_X1 U8700 ( .A(n7704), .ZN(n13144) );
  XNOR2_X1 U8701 ( .A(n8088), .B(n8087), .ZN(n11320) );
  INV_X1 U8702 ( .A(SI_26_), .ZN(n15444) );
  XNOR2_X1 U8703 ( .A(n8154), .B(n8153), .ZN(n11043) );
  NAND2_X1 U8704 ( .A1(n8152), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U8705 ( .A1(n8151), .A2(n8152), .ZN(n10898) );
  NAND2_X1 U8706 ( .A1(n8018), .A2(n7646), .ZN(n8032) );
  INV_X1 U8707 ( .A(SI_23_), .ZN(n10475) );
  NOR2_X1 U8708 ( .A1(n9468), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13135) );
  NAND2_X1 U8709 ( .A1(n7167), .A2(n7164), .ZN(n8008) );
  NAND2_X1 U8710 ( .A1(n7167), .A2(n7642), .ZN(n8006) );
  NAND2_X1 U8711 ( .A1(n7596), .A2(n7666), .ZN(n10250) );
  XNOR2_X1 U8712 ( .A(n7592), .B(n7591), .ZN(n10049) );
  NAND2_X1 U8713 ( .A1(n7928), .A2(n7639), .ZN(n7916) );
  NAND2_X1 U8714 ( .A1(n7149), .A2(n7151), .ZN(n7939) );
  INV_X1 U8715 ( .A(SI_17_), .ZN(n15383) );
  INV_X1 U8716 ( .A(SI_16_), .ZN(n9418) );
  NAND2_X1 U8717 ( .A1(n7153), .A2(n7634), .ZN(n7954) );
  INV_X1 U8718 ( .A(SI_15_), .ZN(n9372) );
  INV_X1 U8719 ( .A(SI_13_), .ZN(n9237) );
  NAND2_X1 U8720 ( .A1(n7145), .A2(n7626), .ZN(n7889) );
  NAND2_X1 U8721 ( .A1(n7872), .A2(n7625), .ZN(n7145) );
  INV_X1 U8722 ( .A(SI_12_), .ZN(n9083) );
  INV_X1 U8723 ( .A(SI_11_), .ZN(n15521) );
  NAND2_X1 U8724 ( .A1(n6913), .A2(n7157), .ZN(n7838) );
  NAND2_X1 U8725 ( .A1(n6914), .A2(n7159), .ZN(n6913) );
  NAND2_X1 U8726 ( .A1(n7811), .A2(n7620), .ZN(n7831) );
  INV_X1 U8727 ( .A(n6927), .ZN(n7776) );
  NAND2_X1 U8728 ( .A1(n7168), .A2(n7612), .ZN(n7758) );
  NAND2_X1 U8729 ( .A1(n7610), .A2(n7609), .ZN(n7747) );
  OR2_X1 U8730 ( .A1(n9437), .A2(n9058), .ZN(n9060) );
  INV_X1 U8731 ( .A(n13573), .ZN(n13390) );
  NOR2_X1 U8732 ( .A1(n13146), .A2(n7327), .ZN(n7326) );
  INV_X1 U8733 ( .A(n12007), .ZN(n7327) );
  NAND2_X1 U8734 ( .A1(n13263), .A2(n12007), .ZN(n13147) );
  AND2_X1 U8735 ( .A1(n11630), .A2(n11603), .ZN(n13391) );
  AND2_X1 U8736 ( .A1(n11559), .A2(n11576), .ZN(n13461) );
  NAND2_X1 U8737 ( .A1(n7336), .A2(n7340), .ZN(n13172) );
  NAND2_X1 U8738 ( .A1(n13203), .A2(n7341), .ZN(n7336) );
  INV_X1 U8739 ( .A(n7342), .ZN(n7341) );
  NOR2_X1 U8740 ( .A1(n10207), .A2(n10206), .ZN(n10210) );
  OAI21_X1 U8741 ( .B1(n6837), .B2(n7311), .A(n7310), .ZN(n11199) );
  NAND2_X1 U8742 ( .A1(n11172), .A2(n11171), .ZN(n13632) );
  NOR2_X1 U8743 ( .A1(n9473), .A2(n11764), .ZN(n13268) );
  INV_X1 U8744 ( .A(n6839), .ZN(n6838) );
  NAND2_X1 U8745 ( .A1(n10651), .A2(n7324), .ZN(n10855) );
  NOR2_X1 U8746 ( .A1(n13217), .A2(n13540), .ZN(n13243) );
  AND2_X1 U8747 ( .A1(n11501), .A2(n11500), .ZN(n13541) );
  NOR2_X1 U8748 ( .A1(n13205), .A2(n11974), .ZN(n13256) );
  OAI21_X1 U8749 ( .B1(n7303), .B2(n7306), .A(n7302), .ZN(n9854) );
  AOI21_X1 U8750 ( .B1(n9674), .B2(n9675), .A(n6664), .ZN(n7302) );
  OAI21_X2 U8751 ( .B1(n9473), .B2(n10103), .A(n15592), .ZN(n13273) );
  NAND2_X1 U8752 ( .A1(n11072), .A2(n11071), .ZN(n11198) );
  NAND2_X1 U8753 ( .A1(n6837), .A2(n11069), .ZN(n11071) );
  INV_X1 U8754 ( .A(n13275), .ZN(n13249) );
  INV_X1 U8755 ( .A(n14857), .ZN(n11767) );
  NAND2_X1 U8756 ( .A1(n11752), .A2(n15591), .ZN(n11753) );
  INV_X1 U8757 ( .A(n11755), .ZN(n11752) );
  INV_X1 U8758 ( .A(n11930), .ZN(n13279) );
  INV_X1 U8759 ( .A(n11944), .ZN(n13423) );
  OR2_X1 U8760 ( .A1(n9466), .A2(n9573), .ZN(n9578) );
  OR2_X1 U8761 ( .A1(n9466), .A2(n9455), .ZN(n9458) );
  NOR2_X1 U8762 ( .A1(n14813), .A2(n14812), .ZN(n14810) );
  AOI21_X1 U8763 ( .B1(n9832), .B2(n9836), .A(n13314), .ZN(n14829) );
  INV_X1 U8764 ( .A(n11698), .ZN(n13558) );
  INV_X1 U8765 ( .A(n13359), .ZN(n13360) );
  NAND2_X1 U8766 ( .A1(n13428), .A2(n11918), .ZN(n13411) );
  NAND2_X1 U8767 ( .A1(n11575), .A2(n11574), .ZN(n13588) );
  NAND2_X1 U8768 ( .A1(n6938), .A2(n6666), .ZN(n13452) );
  NAND2_X1 U8769 ( .A1(n6939), .A2(n11914), .ZN(n13474) );
  OR2_X1 U8770 ( .A1(n13495), .A2(n11912), .ZN(n6939) );
  NAND2_X1 U8771 ( .A1(n7186), .A2(n11939), .ZN(n13468) );
  NAND2_X1 U8772 ( .A1(n11938), .A2(n6690), .ZN(n7186) );
  AND2_X1 U8773 ( .A1(n11525), .A2(n11524), .ZN(n13493) );
  NAND2_X1 U8774 ( .A1(n7210), .A2(n7212), .ZN(n13516) );
  INV_X1 U8775 ( .A(n13623), .ZN(n7063) );
  NAND2_X1 U8776 ( .A1(n11908), .A2(n11907), .ZN(n13533) );
  NAND2_X1 U8777 ( .A1(n7286), .A2(n7285), .ZN(n11276) );
  AND2_X1 U8778 ( .A1(n7286), .A2(n7287), .ZN(n11187) );
  NAND2_X1 U8779 ( .A1(n11184), .A2(n6698), .ZN(n7286) );
  NAND2_X1 U8780 ( .A1(n11225), .A2(n11168), .ZN(n11258) );
  NAND2_X1 U8781 ( .A1(n14552), .A2(n10754), .ZN(n11013) );
  NAND2_X1 U8782 ( .A1(n7292), .A2(n10776), .ZN(n14560) );
  NAND2_X1 U8783 ( .A1(n7300), .A2(n7299), .ZN(n7292) );
  NAND2_X1 U8784 ( .A1(n10353), .A2(n10352), .ZN(n11424) );
  NAND2_X1 U8785 ( .A1(n10290), .A2(n10262), .ZN(n10267) );
  NAND2_X1 U8786 ( .A1(n7272), .A2(n10261), .ZN(n10288) );
  NAND2_X1 U8787 ( .A1(n9556), .A2(n11767), .ZN(n15592) );
  NAND2_X1 U8788 ( .A1(n10172), .A2(n10171), .ZN(n10276) );
  OR2_X1 U8789 ( .A1(n15599), .A2(n10100), .ZN(n13496) );
  OR2_X1 U8790 ( .A1(n15599), .A2(n10103), .ZN(n13528) );
  OR2_X1 U8791 ( .A1(n15599), .A2(n11748), .ZN(n13550) );
  INV_X1 U8792 ( .A(n13550), .ZN(n15590) );
  NAND2_X1 U8793 ( .A1(n6947), .A2(n6727), .ZN(n13658) );
  OR2_X1 U8794 ( .A1(n13565), .A2(n14890), .ZN(n6947) );
  NOR2_X1 U8795 ( .A1(n13563), .A2(n6793), .ZN(n6946) );
  INV_X1 U8796 ( .A(n14851), .ZN(n14852) );
  OR2_X1 U8797 ( .A1(n9638), .A2(P2_U3088), .ZN(n14857) );
  NAND2_X1 U8798 ( .A1(n9055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U8799 ( .A1(n9055), .A2(n8896), .ZN(n11318) );
  NAND2_X1 U8800 ( .A1(n8900), .A2(n8899), .ZN(n11210) );
  XNOR2_X1 U8801 ( .A(n8883), .B(P2_IR_REG_24__SCAN_IN), .ZN(n10908) );
  OAI21_X1 U8802 ( .B1(n9047), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8883) );
  AND2_X1 U8803 ( .A1(n9560), .A2(P2_U3088), .ZN(n13676) );
  INV_X1 U8804 ( .A(n11757), .ZN(n11750) );
  INV_X1 U8805 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9761) );
  INV_X1 U8806 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9725) );
  INV_X1 U8807 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9218) );
  INV_X1 U8808 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9041) );
  INV_X1 U8809 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9021) );
  INV_X1 U8810 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8978) );
  INV_X1 U8811 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U8812 ( .A1(n8984), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8982) );
  INV_X1 U8813 ( .A(n7491), .ZN(n14580) );
  NAND2_X1 U8814 ( .A1(n6825), .A2(n6824), .ZN(n6823) );
  NAND2_X1 U8815 ( .A1(n7513), .A2(n11827), .ZN(n12268) );
  INV_X1 U8816 ( .A(n7499), .ZN(n7498) );
  AOI21_X1 U8817 ( .B1(n7499), .B2(n7497), .A(n6741), .ZN(n7496) );
  NAND2_X1 U8818 ( .A1(n13740), .A2(n11793), .ZN(n13755) );
  AND2_X1 U8819 ( .A1(n7509), .A2(n6675), .ZN(n10625) );
  NAND2_X1 U8820 ( .A1(n11119), .A2(n11118), .ZN(n14596) );
  INV_X1 U8821 ( .A(n12056), .ZN(n14732) );
  INV_X1 U8822 ( .A(n11787), .ZN(n7494) );
  AND2_X1 U8824 ( .A1(n10616), .A2(n14743), .ZN(n14602) );
  OAI21_X1 U8825 ( .B1(n14138), .B2(n6647), .A(n8668), .ZN(n13820) );
  NAND2_X1 U8826 ( .A1(n8609), .A2(n8608), .ZN(n13824) );
  OR2_X1 U8827 ( .A1(n6647), .A2(n9958), .ZN(n8360) );
  OR2_X1 U8828 ( .A1(n12179), .A2(n9005), .ZN(n8353) );
  OR2_X1 U8829 ( .A1(n6646), .A2(n9927), .ZN(n8352) );
  NOR2_X1 U8830 ( .A1(n7076), .A2(n14661), .ZN(n14192) );
  OR2_X1 U8831 ( .A1(n13981), .A2(n13980), .ZN(n14196) );
  NAND2_X1 U8832 ( .A1(n14004), .A2(n14003), .ZN(n14005) );
  NAND2_X1 U8833 ( .A1(n14069), .A2(n7545), .ZN(n14051) );
  AND2_X1 U8834 ( .A1(n14109), .A2(n8806), .ZN(n14084) );
  NAND2_X1 U8835 ( .A1(n8685), .A2(n8684), .ZN(n14110) );
  NAND2_X1 U8836 ( .A1(n14334), .A2(n7346), .ZN(n14234) );
  NAND2_X1 U8837 ( .A1(n7539), .A2(n8653), .ZN(n14134) );
  NAND2_X1 U8838 ( .A1(n7540), .A2(n14157), .ZN(n7539) );
  INV_X1 U8839 ( .A(n14150), .ZN(n7540) );
  NAND2_X1 U8840 ( .A1(n14161), .A2(n8800), .ZN(n14143) );
  OAI21_X1 U8841 ( .B1(n11096), .B2(n7557), .A(n7555), .ZN(n11286) );
  NAND2_X1 U8842 ( .A1(n11095), .A2(n8597), .ZN(n11156) );
  NAND2_X1 U8843 ( .A1(n11093), .A2(n8797), .ZN(n11160) );
  NAND2_X1 U8844 ( .A1(n10638), .A2(n8544), .ZN(n10825) );
  NAND2_X1 U8845 ( .A1(n8534), .A2(n6692), .ZN(n12092) );
  OR2_X1 U8846 ( .A1(n8533), .A2(n9364), .ZN(n7348) );
  NAND2_X1 U8847 ( .A1(n10302), .A2(n8793), .ZN(n10414) );
  OAI21_X1 U8848 ( .B1(n10308), .B2(n7533), .A(n6660), .ZN(n10417) );
  NAND2_X1 U8849 ( .A1(n10307), .A2(n8497), .ZN(n10419) );
  NAND2_X1 U8850 ( .A1(n10022), .A2(n8790), .ZN(n14655) );
  OAI21_X1 U8851 ( .B1(n9905), .B2(n12220), .A(n7520), .ZN(n14654) );
  NAND2_X1 U8852 ( .A1(n10017), .A2(n10019), .ZN(n10016) );
  NAND2_X1 U8853 ( .A1(n9905), .A2(n8450), .ZN(n10017) );
  OAI21_X1 U8854 ( .B1(n9972), .B2(n12216), .A(n7522), .ZN(n10051) );
  AOI21_X1 U8855 ( .B1(n7527), .B2(n9747), .A(n6685), .ZN(n7522) );
  NAND2_X1 U8856 ( .A1(n9745), .A2(n9747), .ZN(n9744) );
  NAND2_X1 U8857 ( .A1(n9972), .A2(n8404), .ZN(n9745) );
  NAND2_X1 U8858 ( .A1(n9736), .A2(n7077), .ZN(n9967) );
  NAND2_X1 U8859 ( .A1(n9924), .A2(n9923), .ZN(n14665) );
  INV_X1 U8860 ( .A(n9350), .ZN(n11962) );
  INV_X1 U8861 ( .A(n14156), .ZN(n14670) );
  INV_X1 U8862 ( .A(n14673), .ZN(n14165) );
  INV_X1 U8863 ( .A(n12202), .ZN(n14284) );
  INV_X1 U8864 ( .A(n11807), .ZN(n14314) );
  INV_X1 U8865 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U8866 ( .A1(n14321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8216) );
  XNOR2_X1 U8867 ( .A(n8752), .B(n8751), .ZN(n13686) );
  CLKBUF_X1 U8868 ( .A(n14328), .Z(n6843) );
  NAND2_X1 U8869 ( .A1(n8657), .A2(n8641), .ZN(n12262) );
  INV_X1 U8870 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9693) );
  INV_X1 U8871 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9767) );
  INV_X1 U8872 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9721) );
  INV_X1 U8873 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9364) );
  INV_X1 U8874 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9215) );
  INV_X1 U8875 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9196) );
  INV_X1 U8876 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9037) );
  INV_X1 U8877 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9023) );
  INV_X1 U8878 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9031) );
  OAI21_X1 U8879 ( .B1(n8420), .B2(n8419), .A(n8437), .ZN(n9847) );
  INV_X1 U8880 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9032) );
  INV_X1 U8881 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9033) );
  INV_X1 U8882 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9027) );
  AND2_X1 U8883 ( .A1(n8387), .A2(n8395), .ZN(n13869) );
  XNOR2_X1 U8884 ( .A(n14381), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n15616) );
  AND2_X1 U8885 ( .A1(n14384), .A2(n14385), .ZN(n14437) );
  AND2_X1 U8886 ( .A1(n7046), .A2(n7045), .ZN(n15614) );
  INV_X1 U8887 ( .A(n14438), .ZN(n7045) );
  OR2_X1 U8888 ( .A1(n14437), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n7046) );
  NOR2_X1 U8889 ( .A1(n15614), .A2(n15613), .ZN(n15612) );
  XNOR2_X1 U8890 ( .A(n6888), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n14441) );
  XNOR2_X1 U8891 ( .A(n14401), .B(n9103), .ZN(n15611) );
  XNOR2_X1 U8892 ( .A(n14406), .B(n14407), .ZN(n14442) );
  NAND2_X1 U8893 ( .A1(n7048), .A2(n14412), .ZN(n14446) );
  NAND2_X1 U8894 ( .A1(n14443), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7048) );
  OR2_X1 U8895 ( .A1(n14413), .A2(n14822), .ZN(n7037) );
  NAND2_X1 U8896 ( .A1(n6891), .A2(n14619), .ZN(n14626) );
  NAND2_X1 U8897 ( .A1(n6677), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6891) );
  INV_X1 U8898 ( .A(n14621), .ZN(n7042) );
  AOI21_X1 U8899 ( .B1(n14418), .B2(n14417), .A(n14629), .ZN(n14634) );
  INV_X1 U8900 ( .A(n14423), .ZN(n6901) );
  AND2_X1 U8901 ( .A1(n14427), .A2(n14428), .ZN(n14448) );
  NAND2_X1 U8902 ( .A1(n9888), .A2(n8921), .ZN(n10155) );
  INV_X1 U8903 ( .A(n6854), .ZN(n10699) );
  AOI21_X1 U8904 ( .B1(n12790), .B2(n15096), .A(n6987), .ZN(n12791) );
  NAND2_X1 U8905 ( .A1(n13161), .A2(n9656), .ZN(n9823) );
  NAND2_X1 U8906 ( .A1(n6836), .A2(n6834), .ZN(P2_U3233) );
  AOI21_X1 U8907 ( .B1(n13350), .B2(n13349), .A(n6835), .ZN(n6834) );
  NAND2_X1 U8908 ( .A1(n13351), .A2(n11748), .ZN(n6836) );
  OAI21_X1 U8909 ( .B1(n14823), .B2(n7674), .A(n13352), .ZN(n6835) );
  NAND2_X1 U8910 ( .A1(n7227), .A2(n7226), .ZN(P2_U3496) );
  NAND2_X1 U8911 ( .A1(n14923), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7226) );
  NAND2_X1 U8912 ( .A1(n13658), .A2(n14925), .ZN(n7227) );
  AND2_X1 U8913 ( .A1(n13701), .A2(n6802), .ZN(n6847) );
  OAI22_X1 U8914 ( .A1(n8868), .A2(n14273), .B1(n14764), .B2(n8861), .ZN(n8862) );
  OAI22_X1 U8915 ( .A1(n8868), .A2(n14318), .B1(n14755), .B2(n8867), .ZN(n8869) );
  NAND2_X1 U8916 ( .A1(n6829), .A2(n6828), .ZN(n14291) );
  OR2_X1 U8917 ( .A1(n14755), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U8918 ( .A1(n14290), .A2(n14755), .ZN(n6829) );
  XNOR2_X1 U8919 ( .A(n7044), .B(n6708), .ZN(SUB_1596_U4) );
  OAI21_X1 U8920 ( .B1(n14451), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6718), .ZN(
        n7044) );
  AND2_X1 U8921 ( .A1(n11914), .A2(n13467), .ZN(n6657) );
  AOI22_X1 U8922 ( .A1(n7242), .A2(n11891), .B1(n7241), .B2(n7243), .ZN(n7240)
         );
  INV_X1 U8923 ( .A(n9708), .ZN(n6995) );
  NOR2_X1 U8924 ( .A1(n7762), .A2(n7128), .ZN(n9523) );
  OR2_X1 U8925 ( .A1(n14157), .A2(n7364), .ZN(n6658) );
  AND2_X1 U8926 ( .A1(n11480), .A2(n7411), .ZN(n6659) );
  AND2_X1 U8927 ( .A1(n10418), .A2(n7532), .ZN(n6660) );
  INV_X1 U8928 ( .A(n14970), .ZN(n7138) );
  NAND2_X1 U8929 ( .A1(n7447), .A2(n12175), .ZN(n6661) );
  AND2_X1 U8930 ( .A1(n8213), .A2(n8214), .ZN(n6662) );
  XNOR2_X1 U8931 ( .A(n9448), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9456) );
  AND2_X1 U8932 ( .A1(n12102), .A2(n7556), .ZN(n6663) );
  NOR2_X1 U8933 ( .A1(n9845), .A2(n9846), .ZN(n6664) );
  AND2_X1 U8934 ( .A1(n7276), .A2(n11907), .ZN(n6665) );
  AND2_X1 U8935 ( .A1(n6940), .A2(n6722), .ZN(n6666) );
  AND2_X1 U8936 ( .A1(n6733), .A2(n7017), .ZN(n6667) );
  AOI21_X1 U8937 ( .B1(n7808), .B2(n7620), .A(n6750), .ZN(n7159) );
  AND2_X1 U8938 ( .A1(n6702), .A2(n11919), .ZN(n6668) );
  NOR2_X1 U8939 ( .A1(n12448), .A2(n7242), .ZN(n6669) );
  AND2_X1 U8940 ( .A1(n11589), .A2(n11588), .ZN(n13416) );
  INV_X1 U8941 ( .A(n13416), .ZN(n13584) );
  INV_X1 U8942 ( .A(n14032), .ZN(n14292) );
  NAND2_X1 U8943 ( .A1(n8326), .A2(n8325), .ZN(n14032) );
  INV_X1 U8944 ( .A(n12228), .ZN(n10639) );
  AND2_X1 U8945 ( .A1(n8796), .A2(n8543), .ZN(n12228) );
  AND2_X1 U8946 ( .A1(n6900), .A2(n6901), .ZN(n6670) );
  AND2_X1 U8947 ( .A1(n6748), .A2(n7288), .ZN(n6671) );
  OR2_X1 U8948 ( .A1(n6742), .A2(n6768), .ZN(n6672) );
  NAND2_X1 U8949 ( .A1(n14067), .A2(n14080), .ZN(n7545) );
  AND2_X1 U8950 ( .A1(n6868), .A2(n6740), .ZN(n6673) );
  AND2_X1 U8951 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n6674) );
  INV_X1 U8952 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U8953 ( .A1(n10618), .A2(n10617), .ZN(n6675) );
  AND2_X1 U8954 ( .A1(n12497), .A2(n12655), .ZN(n6676) );
  NAND2_X1 U8955 ( .A1(n7043), .A2(n7042), .ZN(n6677) );
  INV_X1 U8956 ( .A(n12192), .ZN(n7448) );
  AND2_X1 U8957 ( .A1(n11420), .A2(n6774), .ZN(n6678) );
  INV_X1 U8958 ( .A(n12174), .ZN(n7471) );
  NAND2_X1 U8959 ( .A1(n12071), .A2(n7453), .ZN(n7452) );
  AND2_X1 U8960 ( .A1(n7238), .A2(n11885), .ZN(n6679) );
  INV_X1 U8961 ( .A(n14157), .ZN(n7536) );
  AND2_X1 U8962 ( .A1(n8335), .A2(n8309), .ZN(n6680) );
  NAND2_X1 U8963 ( .A1(n8290), .A2(n15493), .ZN(n6681) );
  INV_X1 U8964 ( .A(n13818), .ZN(n14026) );
  NOR2_X1 U8965 ( .A1(n10136), .A2(n10135), .ZN(n10207) );
  INV_X1 U8966 ( .A(n11411), .ZN(n7056) );
  INV_X1 U8967 ( .A(n14491), .ZN(n6856) );
  AND2_X1 U8968 ( .A1(n6856), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6682) );
  INV_X1 U8969 ( .A(n9345), .ZN(n11836) );
  NAND2_X1 U8970 ( .A1(n9601), .A2(n9468), .ZN(n11572) );
  INV_X1 U8971 ( .A(n6645), .ZN(n7875) );
  INV_X1 U8972 ( .A(n9574), .ZN(n9858) );
  INV_X2 U8973 ( .A(n9858), .ZN(n11642) );
  OR2_X1 U8974 ( .A1(n12179), .A2(n9093), .ZN(n6683) );
  OR2_X1 U8975 ( .A1(n7666), .A2(n7266), .ZN(n6684) );
  AND2_X1 U8976 ( .A1(n10082), .A2(n10041), .ZN(n6685) );
  AOI21_X1 U8977 ( .B1(n10356), .B2(n7180), .A(n7176), .ZN(n7175) );
  OR2_X1 U8978 ( .A1(n14497), .A2(n12735), .ZN(n6686) );
  AND2_X1 U8979 ( .A1(n8273), .A2(n9083), .ZN(n6687) );
  NAND2_X1 U8980 ( .A1(n8700), .A2(n8309), .ZN(n6688) );
  NOR2_X1 U8981 ( .A1(n14169), .A2(n8633), .ZN(n7366) );
  NAND2_X1 U8982 ( .A1(n14113), .A2(n7090), .ZN(n6689) );
  NOR2_X1 U8983 ( .A1(n11940), .A2(n7190), .ZN(n6690) );
  AND2_X1 U8984 ( .A1(n7159), .A2(n7622), .ZN(n6691) );
  AND2_X1 U8985 ( .A1(n7349), .A2(n7348), .ZN(n6692) );
  OR2_X1 U8986 ( .A1(n11352), .A2(n11351), .ZN(n6693) );
  OR2_X1 U8987 ( .A1(n14956), .A2(n7127), .ZN(n6694) );
  NOR2_X1 U8988 ( .A1(n11789), .A2(n7481), .ZN(n6695) );
  OR2_X1 U8989 ( .A1(n14395), .A2(n14394), .ZN(n6696) );
  AND2_X1 U8990 ( .A1(n14955), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6697) );
  AND2_X1 U8991 ( .A1(n11222), .A2(n11183), .ZN(n6698) );
  OR2_X1 U8992 ( .A1(n8798), .A2(n7358), .ZN(n6699) );
  AND2_X1 U8993 ( .A1(n14284), .A2(n12203), .ZN(n6700) );
  NOR2_X1 U8994 ( .A1(n7334), .A2(n10206), .ZN(n6701) );
  AND2_X1 U8995 ( .A1(n13429), .A2(n11915), .ZN(n6702) );
  AND2_X1 U8996 ( .A1(n11462), .A2(n11461), .ZN(n6703) );
  NAND2_X1 U8997 ( .A1(n7637), .A2(n7173), .ZN(n7928) );
  OR2_X1 U8998 ( .A1(n8120), .A2(n8119), .ZN(n6704) );
  AND2_X1 U8999 ( .A1(n7579), .A2(n7762), .ZN(n7839) );
  AND2_X1 U9000 ( .A1(n14955), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6705) );
  OAI22_X1 U9001 ( .A1(n7799), .A2(n7618), .B1(P1_DATAO_REG_6__SCAN_IN), .B2(
        n9031), .ZN(n7809) );
  NAND2_X1 U9002 ( .A1(n11621), .A2(n11620), .ZN(n11698) );
  NAND2_X1 U9003 ( .A1(n6970), .A2(n8271), .ZN(n8515) );
  AND2_X1 U9004 ( .A1(n7822), .A2(n12567), .ZN(n6706) );
  INV_X1 U9005 ( .A(n11485), .ZN(n7033) );
  AND2_X1 U9006 ( .A1(n11492), .A2(n11491), .ZN(n13529) );
  INV_X1 U9007 ( .A(n13529), .ZN(n13616) );
  OR2_X1 U9008 ( .A1(n8324), .A2(n13861), .ZN(n6707) );
  XOR2_X1 U9009 ( .A(n14461), .B(n14460), .Z(n6708) );
  AND4_X1 U9010 ( .A1(n7587), .A2(n7586), .A3(n7585), .A4(n7968), .ZN(n6709)
         );
  AND2_X1 U9011 ( .A1(n12461), .A2(n12484), .ZN(n12521) );
  INV_X1 U9012 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14339) );
  AND2_X1 U9013 ( .A1(n11557), .A2(n11556), .ZN(n13463) );
  INV_X1 U9014 ( .A(n13463), .ZN(n13596) );
  NAND2_X1 U9015 ( .A1(n8389), .A2(n8388), .ZN(n6883) );
  NAND2_X1 U9016 ( .A1(n11653), .A2(n11652), .ZN(n13579) );
  INV_X1 U9017 ( .A(n13579), .ZN(n7065) );
  OR2_X1 U9018 ( .A1(n7797), .A2(n7796), .ZN(n14985) );
  AND2_X1 U9019 ( .A1(n12239), .A2(n7543), .ZN(n6710) );
  AND2_X1 U9020 ( .A1(n13761), .A2(n13824), .ZN(n6711) );
  OR2_X1 U9021 ( .A1(n14407), .A2(n14406), .ZN(n6712) );
  NAND2_X1 U9022 ( .A1(n8519), .A2(n8518), .ZN(n12082) );
  OR2_X1 U9023 ( .A1(n9591), .A2(n8369), .ZN(n6713) );
  AND2_X1 U9024 ( .A1(n7240), .A2(n7238), .ZN(n6714) );
  NAND2_X1 U9025 ( .A1(n13707), .A2(n13706), .ZN(n6715) );
  INV_X1 U9026 ( .A(n9675), .ZN(n7305) );
  NOR2_X1 U9027 ( .A1(n12278), .A2(n12281), .ZN(n6716) );
  AND2_X1 U9028 ( .A1(n7593), .A2(n7119), .ZN(n6717) );
  OR2_X1 U9029 ( .A1(n14453), .A2(n14452), .ZN(n6718) );
  INV_X1 U9030 ( .A(n13696), .ZN(n7490) );
  AND2_X1 U9031 ( .A1(n12124), .A2(n12125), .ZN(n14168) );
  OR2_X1 U9032 ( .A1(n13463), .A2(n13237), .ZN(n6719) );
  AND2_X1 U9033 ( .A1(n11431), .A2(n11430), .ZN(n6720) );
  AND2_X1 U9034 ( .A1(n11437), .A2(n11436), .ZN(n6721) );
  INV_X1 U9035 ( .A(n7558), .ZN(n7557) );
  NOR2_X1 U9036 ( .A1(n7576), .A2(n7559), .ZN(n7558) );
  INV_X1 U9037 ( .A(n13815), .ZN(n8817) );
  NAND2_X1 U9038 ( .A1(n8567), .A2(n8566), .ZN(n13815) );
  OR2_X1 U9039 ( .A1(n13481), .A2(n13451), .ZN(n6722) );
  INV_X1 U9040 ( .A(n12069), .ZN(n6881) );
  INV_X1 U9041 ( .A(n9950), .ZN(n12211) );
  AND2_X1 U9042 ( .A1(n8371), .A2(n8780), .ZN(n9950) );
  NAND2_X1 U9043 ( .A1(n13475), .A2(n7068), .ZN(n7069) );
  INV_X1 U9044 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n7052) );
  INV_X1 U9045 ( .A(n14094), .ZN(n14091) );
  NAND2_X1 U9046 ( .A1(n8702), .A2(n8701), .ZN(n14094) );
  OR2_X1 U9047 ( .A1(n12142), .A2(n12141), .ZN(n6723) );
  AND2_X1 U9048 ( .A1(n12423), .A2(n7259), .ZN(n6724) );
  AND2_X1 U9049 ( .A1(n7171), .A2(n7612), .ZN(n6725) );
  AND2_X1 U9050 ( .A1(n14584), .A2(n13827), .ZN(n6726) );
  AND2_X1 U9051 ( .A1(n12625), .A2(n12624), .ZN(n12936) );
  AND2_X1 U9052 ( .A1(n7228), .A2(n6946), .ZN(n6727) );
  INV_X1 U9053 ( .A(n12118), .ZN(n6876) );
  AND2_X1 U9054 ( .A1(n7861), .A2(n7002), .ZN(n6728) );
  AND2_X1 U9055 ( .A1(n7234), .A2(n7242), .ZN(n6729) );
  INV_X1 U9056 ( .A(n10788), .ZN(n12572) );
  AND2_X1 U9057 ( .A1(n7409), .A2(n7414), .ZN(n6730) );
  INV_X1 U9058 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9689) );
  INV_X1 U9059 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9056) );
  AND2_X1 U9060 ( .A1(n12866), .A2(n7006), .ZN(n6731) );
  NOR2_X1 U9061 ( .A1(n14607), .A2(n13830), .ZN(n6732) );
  OR2_X1 U9062 ( .A1(n11446), .A2(n11448), .ZN(n6733) );
  NOR2_X1 U9063 ( .A1(n12067), .A2(n13833), .ZN(n6734) );
  NOR2_X1 U9064 ( .A1(n11411), .A2(n11408), .ZN(n6735) );
  NOR2_X1 U9065 ( .A1(n14303), .A2(n13820), .ZN(n6736) );
  NOR2_X1 U9066 ( .A1(n13601), .A2(n13451), .ZN(n6737) );
  INV_X1 U9067 ( .A(n6937), .ZN(n6936) );
  NAND2_X1 U9068 ( .A1(n6666), .A2(n6719), .ZN(n6937) );
  NAND2_X1 U9069 ( .A1(n7668), .A2(n8153), .ZN(n6738) );
  INV_X1 U9070 ( .A(n7274), .ZN(n7273) );
  OAI21_X1 U9071 ( .B1(n6665), .B2(n7275), .A(n11910), .ZN(n7274) );
  NAND2_X1 U9072 ( .A1(n11783), .A2(n11782), .ZN(n6739) );
  OR2_X1 U9073 ( .A1(n7448), .A2(n12193), .ZN(n6740) );
  AND2_X1 U9074 ( .A1(n11122), .A2(n11121), .ZN(n6741) );
  AOI21_X1 U9075 ( .B1(n6914), .B2(n6691), .A(n6910), .ZN(n6907) );
  NAND2_X1 U9076 ( .A1(n7447), .A2(n12177), .ZN(n6742) );
  NAND2_X1 U9077 ( .A1(n12555), .A2(n12554), .ZN(n12501) );
  INV_X1 U9078 ( .A(n12501), .ZN(n8097) );
  NOR2_X1 U9079 ( .A1(n14423), .A2(n6903), .ZN(n6743) );
  AND2_X1 U9080 ( .A1(n12042), .A2(n12041), .ZN(n9731) );
  INV_X1 U9081 ( .A(n7091), .ZN(n7090) );
  NAND2_X1 U9082 ( .A1(n7092), .A2(n7093), .ZN(n7091) );
  NAND4_X1 U9083 ( .A1(n6958), .A2(n6709), .A3(n7579), .A4(n7581), .ZN(n6744)
         );
  OR2_X1 U9084 ( .A1(n11424), .A2(n11421), .ZN(n6745) );
  INV_X1 U9085 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6887) );
  AND2_X1 U9086 ( .A1(n8304), .A2(n8303), .ZN(n6746) );
  INV_X1 U9087 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8612) );
  INV_X1 U9088 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9030) );
  NAND2_X1 U9089 ( .A1(n14338), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6747) );
  OR2_X1 U9090 ( .A1(n13416), .A2(n13267), .ZN(n6748) );
  AND2_X1 U9091 ( .A1(n9037), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6749) );
  AND2_X1 U9092 ( .A1(n9041), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n6750) );
  NAND2_X1 U9093 ( .A1(n8436), .A2(n8254), .ZN(n6751) );
  AND2_X1 U9094 ( .A1(n6876), .A2(n12117), .ZN(n6752) );
  OR2_X1 U9095 ( .A1(n6912), .A2(n7621), .ZN(n6753) );
  OR2_X1 U9096 ( .A1(n6998), .A2(n6676), .ZN(n6754) );
  INV_X1 U9097 ( .A(n12500), .ZN(n7009) );
  NOR2_X1 U9098 ( .A1(n7429), .A2(n11447), .ZN(n6755) );
  AND2_X1 U9099 ( .A1(n12457), .A2(n12353), .ZN(n12665) );
  NOR2_X1 U9100 ( .A1(n13529), .A2(n13284), .ZN(n6756) );
  INV_X1 U9101 ( .A(n12237), .ZN(n14070) );
  AND2_X1 U9102 ( .A1(n8808), .A2(n8711), .ZN(n12237) );
  INV_X1 U9103 ( .A(n6900), .ZN(n6904) );
  INV_X1 U9104 ( .A(n12083), .ZN(n7458) );
  INV_X1 U9105 ( .A(n10777), .ZN(n7299) );
  INV_X1 U9106 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7054) );
  INV_X1 U9107 ( .A(n7231), .ZN(n12410) );
  NAND2_X1 U9108 ( .A1(n7233), .A2(n7234), .ZN(n7231) );
  INV_X1 U9109 ( .A(n7322), .ZN(n7321) );
  NAND2_X1 U9110 ( .A1(n7324), .A2(n7323), .ZN(n7322) );
  AND2_X1 U9111 ( .A1(n6904), .A2(n14423), .ZN(n6757) );
  INV_X1 U9112 ( .A(n11538), .ZN(n7422) );
  INV_X1 U9113 ( .A(n13505), .ZN(n13500) );
  OR2_X1 U9114 ( .A1(n11880), .A2(n12705), .ZN(n6758) );
  OR2_X1 U9115 ( .A1(n12399), .A2(n12946), .ZN(n6759) );
  INV_X1 U9116 ( .A(n11917), .ZN(n13429) );
  AND2_X1 U9117 ( .A1(n7240), .A2(n6679), .ZN(n6760) );
  OR2_X1 U9118 ( .A1(n10698), .A2(n10697), .ZN(n6761) );
  AND2_X1 U9119 ( .A1(n10624), .A2(n6675), .ZN(n6762) );
  OR2_X1 U9120 ( .A1(n14343), .A2(n14968), .ZN(n6763) );
  AND3_X1 U9121 ( .A1(n8765), .A2(n8211), .A3(n8773), .ZN(n6764) );
  AND2_X1 U9122 ( .A1(n12063), .A2(n12061), .ZN(n6765) );
  AND2_X1 U9123 ( .A1(n12063), .A2(n12057), .ZN(n6766) );
  AND2_X1 U9124 ( .A1(n6969), .A2(n8528), .ZN(n6767) );
  OAI21_X1 U9125 ( .B1(n13383), .B2(n13387), .A(n11947), .ZN(n11951) );
  AND2_X1 U9126 ( .A1(n7471), .A2(n12173), .ZN(n6768) );
  INV_X1 U9127 ( .A(n14067), .ZN(n14297) );
  NAND2_X1 U9128 ( .A1(n8338), .A2(n8337), .ZN(n14067) );
  AND2_X1 U9129 ( .A1(n6886), .A2(n8218), .ZN(n6769) );
  NAND2_X1 U9130 ( .A1(n13529), .A2(n13284), .ZN(n6770) );
  NAND2_X1 U9131 ( .A1(n11807), .A2(n13823), .ZN(n6771) );
  AND2_X1 U9132 ( .A1(n13995), .A2(n13989), .ZN(n6772) );
  INV_X1 U9133 ( .A(n11168), .ZN(n7224) );
  AND2_X1 U9134 ( .A1(n11916), .A2(n11915), .ZN(n6773) );
  INV_X1 U9135 ( .A(n7294), .ZN(n7293) );
  OAI21_X1 U9136 ( .B1(n10779), .B2(n7295), .A(n10780), .ZN(n7294) );
  AND2_X1 U9137 ( .A1(n11416), .A2(n11415), .ZN(n6774) );
  AND2_X1 U9138 ( .A1(n11862), .A2(n11860), .ZN(n6775) );
  INV_X1 U9139 ( .A(n11012), .ZN(n7204) );
  AND2_X1 U9140 ( .A1(n12222), .A2(n8790), .ZN(n6776) );
  INV_X1 U9141 ( .A(n7297), .ZN(n7296) );
  NOR2_X1 U9142 ( .A1(n10779), .A2(n7298), .ZN(n7297) );
  AND2_X1 U9143 ( .A1(n6668), .A2(n6657), .ZN(n6777) );
  AND2_X1 U9144 ( .A1(n7363), .A2(n14133), .ZN(n6778) );
  INV_X1 U9145 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7591) );
  INV_X1 U9146 ( .A(n6911), .ZN(n6910) );
  NAND2_X1 U9147 ( .A1(n6753), .A2(n7622), .ZN(n6911) );
  NAND2_X1 U9148 ( .A1(n12069), .A2(n6882), .ZN(n6779) );
  AND2_X1 U9149 ( .A1(n6861), .A2(n6860), .ZN(n6780) );
  AND2_X1 U9150 ( .A1(n7427), .A2(n7426), .ZN(n6781) );
  OR2_X1 U9151 ( .A1(n7422), .A2(n11540), .ZN(n6782) );
  INV_X1 U9152 ( .A(n7007), .ZN(n7006) );
  NAND2_X1 U9153 ( .A1(n7008), .A2(n12530), .ZN(n7007) );
  INV_X1 U9154 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8885) );
  OR2_X1 U9155 ( .A1(n7490), .A2(n7488), .ZN(n6783) );
  INV_X2 U9156 ( .A(n12066), .ZN(n12152) );
  INV_X1 U9157 ( .A(n8083), .ZN(n8142) );
  INV_X1 U9158 ( .A(n11689), .ZN(n10957) );
  NAND2_X1 U9159 ( .A1(n10758), .A2(n10757), .ZN(n11443) );
  INV_X1 U9160 ( .A(n11443), .ZN(n7075) );
  NOR2_X1 U9161 ( .A1(n11215), .A2(n13632), .ZN(n7061) );
  INV_X1 U9162 ( .A(n13536), .ZN(n7276) );
  XOR2_X1 U9163 ( .A(n11037), .B(n11895), .Z(n6784) );
  XNOR2_X1 U9164 ( .A(n7725), .B(n7724), .ZN(n9506) );
  INV_X1 U9165 ( .A(n9506), .ZN(n6952) );
  NAND2_X1 U9166 ( .A1(n10576), .A2(n7086), .ZN(n6785) );
  NAND2_X1 U9167 ( .A1(n12989), .A2(n12988), .ZN(n6786) );
  OR2_X1 U9168 ( .A1(n11215), .A2(n13632), .ZN(n6787) );
  NAND2_X1 U9169 ( .A1(n8717), .A2(n8716), .ZN(n14049) );
  INV_X1 U9170 ( .A(n14049), .ZN(n7092) );
  NAND2_X1 U9171 ( .A1(n6960), .A2(n11641), .ZN(n13564) );
  INV_X1 U9172 ( .A(n13564), .ZN(n7057) );
  AND2_X1 U9173 ( .A1(n7061), .A2(n7062), .ZN(n6788) );
  AND2_X1 U9174 ( .A1(n6681), .A2(n8287), .ZN(n6789) );
  AND2_X1 U9175 ( .A1(n13529), .A2(n13541), .ZN(n6790) );
  NOR2_X1 U9176 ( .A1(n12728), .A2(n15064), .ZN(n6791) );
  INV_X1 U9177 ( .A(n8891), .ZN(n9722) );
  AND2_X1 U9178 ( .A1(n11879), .A2(n11878), .ZN(n6792) );
  AND2_X1 U9179 ( .A1(n13564), .A2(n14917), .ZN(n6793) );
  AND2_X1 U9180 ( .A1(n10991), .A2(n12102), .ZN(n6794) );
  NOR2_X1 U9181 ( .A1(n8290), .A2(n15493), .ZN(n6795) );
  AND2_X1 U9182 ( .A1(n6944), .A2(n6945), .ZN(n6796) );
  NAND2_X1 U9183 ( .A1(n7624), .A2(n7623), .ZN(n6797) );
  AND2_X1 U9184 ( .A1(n10638), .A2(n7548), .ZN(n6798) );
  AND2_X1 U9185 ( .A1(n11119), .A2(n7499), .ZN(n6799) );
  NOR2_X1 U9186 ( .A1(n11894), .A2(n12702), .ZN(n6800) );
  INV_X1 U9187 ( .A(n6981), .ZN(n6980) );
  NAND2_X1 U9188 ( .A1(n6984), .A2(n6982), .ZN(n6981) );
  NAND2_X1 U9189 ( .A1(n8893), .A2(n10010), .ZN(n6801) );
  OR2_X1 U9190 ( .A1(n14292), .A2(n13792), .ZN(n6802) );
  AND2_X1 U9191 ( .A1(n8285), .A2(n9418), .ZN(n6803) );
  AND2_X1 U9192 ( .A1(n9339), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n6804) );
  NOR2_X1 U9193 ( .A1(n8311), .A2(SI_25_), .ZN(n6805) );
  OR2_X1 U9194 ( .A1(n8298), .A2(n8297), .ZN(n6806) );
  AND2_X1 U9195 ( .A1(n11184), .A2(n11183), .ZN(n6807) );
  NOR2_X1 U9196 ( .A1(n12927), .A2(n7564), .ZN(n6808) );
  INV_X1 U9197 ( .A(n12230), .ZN(n7556) );
  INV_X1 U9198 ( .A(n12579), .ZN(n7117) );
  AND2_X1 U9199 ( .A1(n10180), .A2(n10177), .ZN(n6809) );
  AND2_X1 U9200 ( .A1(n10368), .A2(n7074), .ZN(n6810) );
  INV_X1 U9201 ( .A(n13627), .ZN(n7062) );
  AND2_X1 U9202 ( .A1(n10654), .A2(n10653), .ZN(n6811) );
  OR2_X1 U9203 ( .A1(n7666), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n6812) );
  AND2_X1 U9204 ( .A1(n7301), .A2(n9674), .ZN(n6813) );
  NAND2_X1 U9205 ( .A1(n8643), .A2(n8642), .ZN(n14248) );
  INV_X1 U9206 ( .A(n14248), .ZN(n7082) );
  NOR2_X1 U9207 ( .A1(n15010), .A2(n10704), .ZN(n6814) );
  INV_X1 U9208 ( .A(n10135), .ZN(n7335) );
  NAND2_X1 U9209 ( .A1(n12722), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6815) );
  AND2_X1 U9210 ( .A1(n11613), .A2(n13142), .ZN(n6816) );
  INV_X1 U9211 ( .A(n7165), .ZN(n7164) );
  NAND2_X1 U9212 ( .A1(n7166), .A2(n7642), .ZN(n7165) );
  AND2_X1 U9213 ( .A1(n9693), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6817) );
  AND2_X1 U9214 ( .A1(n12726), .A2(n12749), .ZN(n6818) );
  AND2_X1 U9215 ( .A1(n7823), .A2(n7822), .ZN(n6819) );
  NAND2_X1 U9216 ( .A1(n9762), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n6820) );
  INV_X1 U9217 ( .A(n11185), .ZN(n7287) );
  INV_X1 U9218 ( .A(n14170), .ZN(n14082) );
  NAND2_X1 U9219 ( .A1(n8492), .A2(n8491), .ZN(n14744) );
  INV_X1 U9220 ( .A(n14744), .ZN(n7080) );
  AND3_X2 U9221 ( .A1(n9634), .A2(n14855), .A3(n9558), .ZN(n14925) );
  AND2_X1 U9222 ( .A1(n8815), .A2(n12183), .ZN(n14656) );
  INV_X1 U9223 ( .A(n14656), .ZN(n14144) );
  INV_X1 U9224 ( .A(n12216), .ZN(n9747) );
  NAND2_X1 U9225 ( .A1(n9705), .A2(n10385), .ZN(n10373) );
  AND2_X1 U9226 ( .A1(n7647), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6821) );
  OR2_X1 U9227 ( .A1(n14480), .A2(n6859), .ZN(n6822) );
  INV_X1 U9228 ( .A(SI_28_), .ZN(n7396) );
  INV_X1 U9229 ( .A(n11748), .ZN(n13349) );
  INV_X1 U9230 ( .A(n8858), .ZN(n10966) );
  INV_X1 U9231 ( .A(n9456), .ZN(n12267) );
  INV_X1 U9232 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n6859) );
  INV_X1 U9233 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7050) );
  AND2_X2 U9234 ( .A1(n9048), .A2(n9047), .ZN(n9581) );
  INV_X1 U9235 ( .A(n10559), .ZN(n6842) );
  XNOR2_X1 U9236 ( .A(n9649), .B(n9648), .ZN(n13181) );
  NAND2_X1 U9237 ( .A1(n10951), .A2(n10952), .ZN(n11070) );
  OAI21_X1 U9238 ( .B1(n13227), .B2(n13223), .A(n13224), .ZN(n13189) );
  AOI21_X1 U9239 ( .B1(n9652), .B2(n9651), .A(n13251), .ZN(n13163) );
  NAND2_X1 U9240 ( .A1(n13714), .A2(n11816), .ZN(n13716) );
  NAND2_X1 U9241 ( .A1(n8580), .A2(n8212), .ZN(n8825) );
  INV_X1 U9242 ( .A(n8838), .ZN(n8841) );
  OAI21_X2 U9243 ( .B1(n10186), .B2(n10185), .A(n10184), .ZN(n10190) );
  OAI21_X2 U9244 ( .B1(n11245), .B2(n11244), .A(n11243), .ZN(n11249) );
  INV_X1 U9245 ( .A(n9356), .ZN(n9354) );
  INV_X1 U9246 ( .A(n9352), .ZN(n6824) );
  INV_X1 U9247 ( .A(n9351), .ZN(n6825) );
  AOI21_X1 U9248 ( .B1(n7520), .B2(n12220), .A(n12222), .ZN(n7518) );
  NAND2_X1 U9249 ( .A1(n13997), .A2(n14752), .ZN(n7351) );
  NAND2_X1 U9250 ( .A1(n13782), .A2(n13783), .ZN(n13714) );
  NOR2_X2 U9251 ( .A1(n13812), .A2(n13811), .ZN(n13810) );
  INV_X1 U9252 ( .A(n7340), .ZN(n7339) );
  NAND2_X1 U9253 ( .A1(n13255), .A2(n7344), .ZN(n7343) );
  BUF_X4 U9254 ( .A(n8235), .Z(n9468) );
  NAND2_X1 U9255 ( .A1(n9344), .A2(n9343), .ZN(n9353) );
  OAI21_X2 U9256 ( .B1(n8805), .B2(n7369), .A(n7367), .ZN(n14057) );
  NAND2_X1 U9257 ( .A1(n8789), .A2(n12220), .ZN(n10022) );
  NAND2_X1 U9258 ( .A1(n9977), .A2(n8781), .ZN(n9748) );
  NAND2_X1 U9259 ( .A1(n14040), .A2(n8810), .ZN(n14024) );
  NAND2_X1 U9260 ( .A1(n7360), .A2(n7359), .ZN(n10413) );
  NAND2_X1 U9261 ( .A1(n10632), .A2(n12228), .ZN(n10636) );
  OAI21_X1 U9262 ( .B1(n14169), .B2(n7362), .A(n6778), .ZN(n8802) );
  OAI21_X2 U9263 ( .B1(n10991), .B2(n6699), .A(n7355), .ZN(n11284) );
  AND3_X2 U9264 ( .A1(n8212), .A2(n8580), .A3(n6885), .ZN(n8321) );
  NAND2_X1 U9265 ( .A1(n9949), .A2(n9950), .ZN(n9948) );
  AND2_X1 U9266 ( .A1(n13263), .A2(n6833), .ZN(n13276) );
  NAND2_X1 U9267 ( .A1(n13264), .A2(n13265), .ZN(n6833) );
  OR2_X2 U9268 ( .A1(n13264), .A2(n13265), .ZN(n13263) );
  MUX2_X1 U9269 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n8235), .Z(n8236) );
  NAND2_X1 U9270 ( .A1(n8346), .A2(n8239), .ZN(n8364) );
  NAND2_X1 U9271 ( .A1(n7328), .A2(n6838), .ZN(n10559) );
  OAI21_X1 U9272 ( .B1(n7332), .B2(n7335), .A(n7331), .ZN(n6839) );
  INV_X1 U9273 ( .A(n8344), .ZN(n7371) );
  NAND2_X1 U9274 ( .A1(n7379), .A2(n7378), .ZN(n8452) );
  NAND2_X1 U9275 ( .A1(n8342), .A2(n7371), .ZN(n8346) );
  NAND2_X1 U9276 ( .A1(n7309), .A2(n7307), .ZN(n11971) );
  OAI21_X1 U9277 ( .B1(SI_1_), .B2(n8236), .A(n8239), .ZN(n8344) );
  NAND2_X2 U9278 ( .A1(n10992), .A2(n12234), .ZN(n10991) );
  OR2_X1 U9279 ( .A1(n8866), .A2(n14753), .ZN(n8871) );
  OR2_X1 U9280 ( .A1(n8866), .A2(n14761), .ZN(n8864) );
  INV_X4 U9281 ( .A(n12295), .ZN(n12324) );
  NAND2_X1 U9282 ( .A1(n13716), .A2(n11820), .ZN(n13776) );
  NAND2_X2 U9283 ( .A1(n13794), .A2(n13795), .ZN(n13793) );
  NAND2_X1 U9284 ( .A1(n7502), .A2(n7507), .ZN(n7506) );
  NAND2_X1 U9285 ( .A1(n6772), .A2(n7351), .ZN(n7350) );
  NAND2_X1 U9286 ( .A1(n14653), .A2(n8486), .ZN(n10308) );
  NAND2_X1 U9287 ( .A1(n8467), .A2(n7386), .ZN(n7385) );
  OAI21_X1 U9288 ( .B1(n8405), .B2(n7382), .A(n8419), .ZN(n7381) );
  AND2_X2 U9289 ( .A1(n6842), .A2(n6841), .ZN(n10563) );
  NAND2_X1 U9290 ( .A1(n8804), .A2(n8803), .ZN(n14122) );
  NAND2_X1 U9291 ( .A1(n10819), .A2(n12097), .ZN(n10992) );
  NAND2_X1 U9292 ( .A1(n9730), .A2(n9731), .ZN(n9729) );
  NOR2_X1 U9293 ( .A1(n13987), .A2(n7350), .ZN(n8866) );
  XNOR2_X1 U9294 ( .A(n8814), .B(n12241), .ZN(n7354) );
  NAND2_X1 U9295 ( .A1(n7354), .A2(n14144), .ZN(n7353) );
  NAND2_X1 U9296 ( .A1(n6846), .A2(n6844), .ZN(n8356) );
  NAND2_X1 U9297 ( .A1(n13776), .A2(n13775), .ZN(n7513) );
  NAND2_X2 U9298 ( .A1(n10190), .A2(n10189), .ZN(n10434) );
  NAND2_X1 U9299 ( .A1(n6848), .A2(n6847), .ZN(P1_U3214) );
  NAND2_X1 U9300 ( .A1(n13697), .A2(n14585), .ZN(n6848) );
  INV_X1 U9301 ( .A(n7501), .ZN(n11128) );
  NAND2_X1 U9302 ( .A1(n11959), .A2(n11960), .ZN(n11958) );
  OAI21_X2 U9303 ( .B1(n9468), .B2(n9030), .A(n6849), .ZN(n8240) );
  NAND2_X1 U9304 ( .A1(n6643), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6849) );
  NAND2_X2 U9305 ( .A1(n8324), .A2(n9560), .ZN(n8369) );
  INV_X1 U9306 ( .A(n12728), .ZN(n6853) );
  NOR2_X1 U9307 ( .A1(n15065), .A2(n15066), .ZN(n15064) );
  INV_X1 U9308 ( .A(n12731), .ZN(n15082) );
  INV_X1 U9309 ( .A(n14463), .ZN(n6858) );
  INV_X1 U9310 ( .A(n6861), .ZN(n14462) );
  NAND3_X1 U9311 ( .A1(n12134), .A2(n12133), .A3(n6866), .ZN(n6865) );
  NAND2_X1 U9312 ( .A1(n7468), .A2(n6870), .ZN(n6869) );
  NAND3_X1 U9313 ( .A1(n6873), .A2(n6872), .A3(n12126), .ZN(n12129) );
  AND2_X1 U9314 ( .A1(n12110), .A2(n12109), .ZN(n6877) );
  NAND2_X1 U9315 ( .A1(n6879), .A2(n6878), .ZN(n7451) );
  NAND3_X1 U9316 ( .A1(n7443), .A2(n7440), .A3(n6779), .ZN(n6878) );
  AND3_X1 U9317 ( .A1(n8212), .A2(n8580), .A3(n6884), .ZN(n8217) );
  AND2_X1 U9318 ( .A1(n6662), .A2(n6886), .ZN(n6884) );
  NAND4_X1 U9319 ( .A1(n8212), .A2(n8580), .A3(n6662), .A4(n6769), .ZN(n14321)
         );
  NAND3_X1 U9320 ( .A1(n8212), .A2(n8580), .A3(n6662), .ZN(n8829) );
  INV_X1 U9321 ( .A(n6888), .ZN(n14399) );
  XNOR2_X1 U9322 ( .A(n14395), .B(n14394), .ZN(n15607) );
  OAI21_X1 U9323 ( .B1(n14376), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6763), .ZN(
        n6894) );
  NAND2_X1 U9324 ( .A1(n14422), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U9325 ( .A1(n6896), .A2(n6895), .ZN(n14427) );
  NOR2_X1 U9326 ( .A1(n6902), .A2(n6898), .ZN(n6897) );
  NAND2_X1 U9327 ( .A1(n14633), .A2(n6905), .ZN(n6900) );
  INV_X1 U9328 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6903) );
  NAND2_X1 U9329 ( .A1(n7809), .A2(n6911), .ZN(n6906) );
  INV_X1 U9330 ( .A(n7809), .ZN(n6914) );
  OAI21_X1 U9331 ( .B1(n8020), .B2(n6922), .A(n6920), .ZN(n7649) );
  INV_X1 U9332 ( .A(n7649), .ZN(n7648) );
  NAND2_X1 U9333 ( .A1(n7154), .A2(n6925), .ZN(n8053) );
  NAND2_X1 U9334 ( .A1(n7651), .A2(n6926), .ZN(n6925) );
  NAND2_X1 U9335 ( .A1(n8053), .A2(n7653), .ZN(n8065) );
  NAND3_X1 U9336 ( .A1(n6930), .A2(n6929), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7675) );
  AOI21_X1 U9337 ( .B1(n13495), .B2(n6777), .A(n6934), .ZN(n13400) );
  NAND3_X1 U9338 ( .A1(n11914), .A2(n11912), .A3(n13467), .ZN(n6940) );
  NAND2_X1 U9339 ( .A1(n6942), .A2(n6941), .ZN(n8238) );
  MUX2_X1 U9340 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n9560), .Z(n8681) );
  MUX2_X1 U9341 ( .A(n11211), .B(n11214), .S(n9560), .Z(n8310) );
  MUX2_X1 U9342 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n9560), .Z(n8750) );
  MUX2_X1 U9343 ( .A(n13692), .B(n14331), .S(n9560), .Z(n8730) );
  MUX2_X1 U9344 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n9560), .Z(n11614) );
  NAND2_X2 U9345 ( .A1(P1_U3086), .A2(n6643), .ZN(n14332) );
  NAND2_X1 U9346 ( .A1(n6944), .A2(n6943), .ZN(n13504) );
  NAND3_X1 U9347 ( .A1(n7725), .A2(n9504), .A3(n7130), .ZN(n6996) );
  AND2_X2 U9348 ( .A1(n6957), .A2(n6955), .ZN(n7593) );
  NAND3_X1 U9349 ( .A1(n6957), .A2(n6955), .A3(n7120), .ZN(n7003) );
  NAND3_X1 U9350 ( .A1(n6958), .A2(n7581), .A3(n7579), .ZN(n7588) );
  NAND3_X1 U9351 ( .A1(n11747), .A2(n11677), .A3(n6962), .ZN(n11676) );
  NAND2_X1 U9352 ( .A1(n8499), .A2(n6966), .ZN(n6965) );
  NAND2_X1 U9353 ( .A1(n6965), .A2(n6767), .ZN(n8277) );
  NAND2_X1 U9354 ( .A1(n8315), .A2(n6976), .ZN(n8732) );
  NAND2_X1 U9355 ( .A1(n8315), .A2(n8314), .ZN(n8713) );
  NAND2_X1 U9356 ( .A1(n8288), .A2(n6789), .ZN(n6983) );
  NAND2_X1 U9357 ( .A1(n8288), .A2(n8287), .ZN(n8289) );
  INV_X1 U9358 ( .A(n6996), .ZN(n7762) );
  NAND2_X1 U9359 ( .A1(n6996), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U9360 ( .A1(n8063), .A2(n6676), .ZN(n7000) );
  AND2_X1 U9361 ( .A1(n7000), .A2(n6999), .ZN(n12814) );
  OAI211_X2 U9362 ( .C1(n6706), .C2(n10788), .A(n12576), .B(n7001), .ZN(n10867) );
  NAND2_X1 U9363 ( .A1(n10793), .A2(n12572), .ZN(n10792) );
  NAND2_X1 U9364 ( .A1(n6706), .A2(n7823), .ZN(n10793) );
  NAND2_X1 U9365 ( .A1(n7011), .A2(n7010), .ZN(n7903) );
  NAND2_X1 U9366 ( .A1(n7012), .A2(n7013), .ZN(n8017) );
  NAND2_X1 U9367 ( .A1(n12907), .A2(n12638), .ZN(n7012) );
  NAND2_X1 U9368 ( .A1(n11440), .A2(n6667), .ZN(n7016) );
  INV_X1 U9369 ( .A(n6721), .ZN(n7019) );
  NAND2_X2 U9370 ( .A1(n8891), .A2(n8880), .ZN(n8892) );
  AOI21_X1 U9371 ( .B1(n7022), .B2(n7433), .A(n6678), .ZN(n7020) );
  NAND2_X1 U9372 ( .A1(n11414), .A2(n7022), .ZN(n7021) );
  NAND3_X1 U9373 ( .A1(n7029), .A2(n11520), .A3(n6782), .ZN(n7028) );
  NAND3_X1 U9374 ( .A1(n6656), .A2(n11757), .A3(n11748), .ZN(n11321) );
  OAI22_X1 U9375 ( .A1(n11395), .A2(n7030), .B1(n11394), .B2(n11393), .ZN(
        n11402) );
  NAND2_X1 U9376 ( .A1(n11402), .A2(n11403), .ZN(n11401) );
  NOR2_X1 U9377 ( .A1(n7031), .A2(n7032), .ZN(n7030) );
  INV_X1 U9378 ( .A(n11393), .ZN(n7031) );
  NAND3_X1 U9379 ( .A1(n11460), .A2(n11459), .A3(n6659), .ZN(n7034) );
  NAND2_X1 U9380 ( .A1(n7037), .A2(n14444), .ZN(n14616) );
  NAND2_X1 U9381 ( .A1(n7037), .A2(n7036), .ZN(n7035) );
  NOR2_X1 U9382 ( .A1(n14413), .A2(n7040), .ZN(n7038) );
  NOR2_X1 U9383 ( .A1(n14616), .A2(n14617), .ZN(n14615) );
  INV_X1 U9384 ( .A(n14617), .ZN(n7041) );
  INV_X1 U9385 ( .A(n7043), .ZN(n14620) );
  NAND3_X1 U9386 ( .A1(n7055), .A2(n9450), .A3(n7053), .ZN(n9061) );
  OR2_X2 U9387 ( .A1(n9055), .A2(n7428), .ZN(n9450) );
  INV_X1 U9388 ( .A(n7069), .ZN(n13443) );
  NAND2_X1 U9389 ( .A1(n10368), .A2(n7070), .ZN(n11019) );
  NOR2_X1 U9390 ( .A1(n14192), .A2(n14191), .ZN(n14281) );
  XNOR2_X1 U9391 ( .A(n13980), .B(n14284), .ZN(n7076) );
  NOR2_X2 U9392 ( .A1(n7077), .A2(n14722), .ZN(n9982) );
  NAND2_X1 U9393 ( .A1(n7079), .A2(n7078), .ZN(n7077) );
  OR2_X2 U9394 ( .A1(n14662), .A2(n14671), .ZN(n14663) );
  NAND2_X1 U9395 ( .A1(n10576), .A2(n7084), .ZN(n11098) );
  NAND2_X1 U9396 ( .A1(n7094), .A2(n7095), .ZN(n12945) );
  NAND2_X1 U9397 ( .A1(n11150), .A2(n7097), .ZN(n7094) );
  NAND2_X1 U9398 ( .A1(n12887), .A2(n7106), .ZN(n7103) );
  NAND2_X1 U9399 ( .A1(n7103), .A2(n7104), .ZN(n12862) );
  NAND2_X1 U9400 ( .A1(n12928), .A2(n7110), .ZN(n7107) );
  NAND2_X1 U9401 ( .A1(n7107), .A2(n7108), .ZN(n12897) );
  NAND3_X1 U9402 ( .A1(n7854), .A2(n7114), .A3(n7113), .ZN(n12710) );
  NAND2_X1 U9403 ( .A1(n12710), .A2(n11008), .ZN(n12586) );
  NAND3_X1 U9404 ( .A1(n10868), .A2(n12505), .A3(n7117), .ZN(n7116) );
  NAND3_X1 U9405 ( .A1(n7123), .A2(n7589), .A3(n7122), .ZN(n7121) );
  NAND2_X1 U9406 ( .A1(n15044), .A2(n6818), .ZN(n7125) );
  OAI211_X1 U9407 ( .C1(n15044), .C2(n12749), .A(n7126), .B(n7125), .ZN(n15065) );
  OR2_X1 U9408 ( .A1(n14956), .A2(n6697), .ZN(n9705) );
  AND2_X1 U9409 ( .A1(n7142), .A2(n6686), .ZN(n14522) );
  INV_X1 U9410 ( .A(n7142), .ZN(n14506) );
  NAND2_X1 U9411 ( .A1(n7872), .A2(n7146), .ZN(n7144) );
  NAND2_X1 U9412 ( .A1(n7966), .A2(n7633), .ZN(n7153) );
  NAND2_X1 U9413 ( .A1(n7966), .A2(n7150), .ZN(n7149) );
  OAI21_X1 U9414 ( .B1(n8042), .B2(n7156), .A(n7651), .ZN(n8051) );
  AOI21_X1 U9415 ( .B1(n7651), .B2(n7156), .A(n7155), .ZN(n7154) );
  INV_X1 U9416 ( .A(n8050), .ZN(n7155) );
  NAND2_X1 U9417 ( .A1(n7610), .A2(n7169), .ZN(n7168) );
  NAND2_X1 U9418 ( .A1(n7637), .A2(n7636), .ZN(n7926) );
  NAND2_X1 U9419 ( .A1(n7648), .A2(n10965), .ZN(n7651) );
  NAND2_X1 U9420 ( .A1(n8408), .A2(n8251), .ZN(n8420) );
  NAND2_X2 U9421 ( .A1(n12671), .A2(n12797), .ZN(n12816) );
  INV_X1 U9422 ( .A(n7175), .ZN(n14549) );
  NAND2_X1 U9423 ( .A1(n10356), .A2(n10355), .ZN(n10520) );
  NAND2_X1 U9424 ( .A1(n11938), .A2(n7187), .ZN(n7184) );
  NAND2_X1 U9425 ( .A1(n7184), .A2(n7185), .ZN(n13449) );
  NAND2_X1 U9426 ( .A1(n11938), .A2(n11937), .ZN(n13485) );
  INV_X1 U9427 ( .A(n11937), .ZN(n7190) );
  NAND2_X1 U9428 ( .A1(n10172), .A2(n7191), .ZN(n7192) );
  NAND2_X1 U9429 ( .A1(n7192), .A2(n7194), .ZN(n10354) );
  NAND2_X1 U9430 ( .A1(n7175), .A2(n7201), .ZN(n7200) );
  OR2_X1 U9431 ( .A1(n11934), .A2(n7208), .ZN(n7205) );
  NAND2_X1 U9432 ( .A1(n7205), .A2(n7206), .ZN(n13501) );
  INV_X1 U9433 ( .A(n11223), .ZN(n7225) );
  NAND2_X1 U9434 ( .A1(n7221), .A2(n7222), .ZN(n11260) );
  NAND2_X1 U9435 ( .A1(n11223), .A2(n11168), .ZN(n7221) );
  NAND3_X1 U9436 ( .A1(n11953), .A2(n11954), .A3(n7229), .ZN(n13562) );
  NAND2_X1 U9437 ( .A1(n9793), .A2(n7230), .ZN(n9898) );
  NAND2_X1 U9438 ( .A1(n8912), .A2(n15112), .ZN(n7230) );
  NAND2_X1 U9439 ( .A1(n12430), .A2(n11885), .ZN(n7233) );
  NAND2_X1 U9440 ( .A1(n12430), .A2(n6760), .ZN(n7235) );
  NAND2_X1 U9441 ( .A1(n7232), .A2(n7240), .ZN(n12447) );
  INV_X1 U9442 ( .A(n12383), .ZN(n7241) );
  NAND3_X1 U9443 ( .A1(n7236), .A2(n7235), .A3(n7237), .ZN(n12351) );
  NAND2_X1 U9444 ( .A1(n11296), .A2(n7249), .ZN(n7247) );
  NAND2_X1 U9445 ( .A1(n11861), .A2(n6775), .ZN(n12393) );
  NAND3_X1 U9446 ( .A1(n7261), .A2(n11137), .A3(n10742), .ZN(n11138) );
  NAND2_X1 U9447 ( .A1(n11030), .A2(n11029), .ZN(n7262) );
  NAND3_X1 U9448 ( .A1(n7579), .A2(n7581), .A3(n7762), .ZN(n7886) );
  NAND3_X1 U9449 ( .A1(n7270), .A2(n7269), .A3(n8180), .ZN(n7268) );
  NAND2_X2 U9450 ( .A1(n9061), .A2(n13691), .ZN(n9601) );
  NAND2_X1 U9451 ( .A1(n7279), .A2(n10092), .ZN(n7278) );
  NAND3_X1 U9452 ( .A1(n7278), .A2(n10160), .A3(n7277), .ZN(n10164) );
  INV_X1 U9453 ( .A(n10093), .ZN(n7281) );
  NAND2_X1 U9454 ( .A1(n10456), .A2(n10093), .ZN(n10161) );
  NAND2_X1 U9455 ( .A1(n10457), .A2(n11725), .ZN(n10456) );
  NAND2_X1 U9456 ( .A1(n10778), .A2(n7297), .ZN(n7290) );
  OAI21_X1 U9457 ( .B1(n10778), .B2(n7294), .A(n7291), .ZN(n11009) );
  NAND2_X1 U9458 ( .A1(n7306), .A2(n7305), .ZN(n7301) );
  INV_X1 U9459 ( .A(n9674), .ZN(n7303) );
  INV_X1 U9460 ( .A(n7306), .ZN(n9822) );
  NAND2_X1 U9461 ( .A1(n11070), .A2(n7310), .ZN(n7309) );
  XNOR2_X1 U9462 ( .A(n7312), .B(n11324), .ZN(n9648) );
  NAND2_X1 U9463 ( .A1(n10651), .A2(n7317), .ZN(n7313) );
  NAND2_X1 U9464 ( .A1(n7313), .A2(n7314), .ZN(n10951) );
  NAND2_X1 U9465 ( .A1(n10136), .A2(n7329), .ZN(n7328) );
  CLKBUF_X1 U9466 ( .A(n8324), .Z(n7346) );
  MUX2_X1 U9467 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14336), .S(n8324), .Z(n9995)
         );
  NAND2_X1 U9468 ( .A1(n10301), .A2(n8793), .ZN(n7360) );
  NAND2_X1 U9469 ( .A1(n10022), .A2(n6776), .ZN(n14658) );
  INV_X1 U9470 ( .A(n12222), .ZN(n7361) );
  NAND2_X1 U9471 ( .A1(n8800), .A2(n14168), .ZN(n7362) );
  INV_X1 U9472 ( .A(n7366), .ZN(n7365) );
  NAND2_X1 U9473 ( .A1(n7365), .A2(n12125), .ZN(n14158) );
  NOR2_X1 U9474 ( .A1(n8238), .A2(n15508), .ZN(n8342) );
  NAND2_X1 U9475 ( .A1(n8406), .A2(n7380), .ZN(n7379) );
  NAND2_X1 U9476 ( .A1(n8406), .A2(n8405), .ZN(n8408) );
  NAND2_X1 U9477 ( .A1(n8735), .A2(n7399), .ZN(n7398) );
  NAND2_X1 U9478 ( .A1(n8735), .A2(n8734), .ZN(n8752) );
  NAND2_X1 U9479 ( .A1(n8302), .A2(SI_22_), .ZN(n8304) );
  NAND2_X1 U9480 ( .A1(n8698), .A2(n6680), .ZN(n7405) );
  OR2_X1 U9481 ( .A1(n9466), .A2(n9465), .ZN(n7407) );
  NAND3_X1 U9482 ( .A1(n9456), .A2(n13683), .A3(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7406) );
  INV_X1 U9483 ( .A(n11463), .ZN(n7415) );
  NAND2_X1 U9484 ( .A1(n7420), .A2(n7416), .ZN(n11568) );
  NAND2_X1 U9485 ( .A1(n7418), .A2(n7417), .ZN(n7416) );
  NAND2_X1 U9486 ( .A1(n7419), .A2(n11553), .ZN(n7418) );
  NAND2_X1 U9487 ( .A1(n7421), .A2(n11552), .ZN(n7420) );
  NAND3_X1 U9488 ( .A1(n8891), .A2(n8890), .A3(n6781), .ZN(n7425) );
  NAND2_X1 U9489 ( .A1(n12135), .A2(n12137), .ZN(n7434) );
  OAI21_X1 U9490 ( .B1(n7435), .B2(n12037), .A(n9950), .ZN(n7439) );
  INV_X1 U9491 ( .A(n7436), .ZN(n7435) );
  OAI211_X1 U9492 ( .C1(n12033), .C2(n12152), .A(n7437), .B(n12214), .ZN(n7436) );
  NAND2_X1 U9493 ( .A1(n7078), .A2(n13838), .ZN(n12041) );
  NAND3_X1 U9494 ( .A1(n12031), .A2(n12152), .A3(n12030), .ZN(n7437) );
  NAND2_X1 U9495 ( .A1(n7439), .A2(n7438), .ZN(n12044) );
  NAND3_X1 U9496 ( .A1(n7442), .A2(n7441), .A3(n7446), .ZN(n7440) );
  NAND2_X1 U9497 ( .A1(n12062), .A2(n12061), .ZN(n7441) );
  NAND2_X1 U9498 ( .A1(n12058), .A2(n12057), .ZN(n7442) );
  NAND2_X1 U9499 ( .A1(n12062), .A2(n6765), .ZN(n7444) );
  NAND2_X1 U9500 ( .A1(n12058), .A2(n6766), .ZN(n7445) );
  NAND2_X4 U9501 ( .A1(n12188), .A2(n12028), .ZN(n12066) );
  AND2_X2 U9502 ( .A1(n12024), .A2(n7449), .ZN(n12188) );
  NAND3_X1 U9503 ( .A1(n8775), .A2(n14335), .A3(n12206), .ZN(n7449) );
  INV_X1 U9504 ( .A(n12070), .ZN(n7453) );
  NAND3_X1 U9505 ( .A1(n12080), .A2(n12081), .A3(n7457), .ZN(n7454) );
  NAND2_X1 U9506 ( .A1(n7454), .A2(n7455), .ZN(n12101) );
  AND2_X1 U9507 ( .A1(n12209), .A2(n12088), .ZN(n7459) );
  NAND2_X1 U9508 ( .A1(n7460), .A2(n7463), .ZN(n12155) );
  NAND3_X1 U9509 ( .A1(n12146), .A2(n7462), .A3(n7461), .ZN(n7460) );
  NAND2_X1 U9510 ( .A1(n8585), .A2(n7466), .ZN(n8624) );
  INV_X1 U9511 ( .A(n8600), .ZN(n7467) );
  NAND3_X1 U9512 ( .A1(n12172), .A2(n7469), .A3(n12171), .ZN(n7468) );
  NAND2_X1 U9513 ( .A1(n7472), .A2(n7474), .ZN(n12059) );
  NAND3_X1 U9514 ( .A1(n12051), .A2(n12050), .A3(n7473), .ZN(n7472) );
  INV_X1 U9515 ( .A(n12053), .ZN(n7475) );
  INV_X1 U9516 ( .A(n6827), .ZN(n7482) );
  NAND2_X1 U9517 ( .A1(n7477), .A2(n7476), .ZN(n11803) );
  NAND2_X1 U9518 ( .A1(n13810), .A2(n11793), .ZN(n7477) );
  NOR2_X1 U9519 ( .A1(n6827), .A2(n11789), .ZN(n13741) );
  OAI211_X1 U9520 ( .C1(n13793), .C2(n6783), .A(n7485), .B(n7483), .ZN(n12334)
         );
  OAI22_X1 U9521 ( .A1(n7487), .A2(n7484), .B1(n12329), .B2(n7489), .ZN(n7483)
         );
  NOR2_X1 U9522 ( .A1(n13696), .A2(n12329), .ZN(n7484) );
  NAND2_X1 U9523 ( .A1(n13793), .A2(n7486), .ZN(n7485) );
  NOR2_X1 U9524 ( .A1(n12329), .A2(n7487), .ZN(n7486) );
  INV_X1 U9525 ( .A(n12329), .ZN(n7488) );
  NAND2_X1 U9526 ( .A1(n11780), .A2(n11779), .ZN(n14581) );
  NOR2_X1 U9527 ( .A1(n14582), .A2(n7493), .ZN(n7492) );
  INV_X1 U9528 ( .A(n11779), .ZN(n7493) );
  INV_X1 U9529 ( .A(n7495), .ZN(n11788) );
  OAI21_X1 U9530 ( .B1(n10842), .B2(n7498), .A(n7496), .ZN(n7501) );
  NAND4_X1 U9531 ( .A1(n7506), .A2(n7503), .A3(n7504), .A4(n9868), .ZN(n9869)
         );
  NAND2_X1 U9532 ( .A1(n9805), .A2(n7508), .ZN(n9868) );
  INV_X1 U9533 ( .A(n9805), .ZN(n7502) );
  NAND3_X1 U9534 ( .A1(n7506), .A2(n9868), .A3(n7504), .ZN(n9808) );
  NAND2_X1 U9535 ( .A1(n10434), .A2(n10433), .ZN(n10435) );
  INV_X1 U9536 ( .A(n7509), .ZN(n10619) );
  NOR2_X1 U9537 ( .A1(n10436), .A2(n7511), .ZN(n7510) );
  INV_X1 U9538 ( .A(n10433), .ZN(n7511) );
  NAND2_X1 U9539 ( .A1(n7513), .A2(n7512), .ZN(n13707) );
  NAND2_X2 U9540 ( .A1(n12029), .A2(n9225), .ZN(n11834) );
  NAND2_X1 U9541 ( .A1(n12212), .A2(n7517), .ZN(n7516) );
  OAI21_X1 U9542 ( .B1(n9946), .B2(n9731), .A(n7515), .ZN(n9974) );
  NAND2_X1 U9543 ( .A1(n9727), .A2(n12212), .ZN(n9726) );
  NAND2_X1 U9544 ( .A1(n9946), .A2(n8372), .ZN(n9727) );
  NAND2_X1 U9545 ( .A1(n9905), .A2(n7520), .ZN(n7519) );
  NAND2_X1 U9546 ( .A1(n9972), .A2(n7526), .ZN(n7525) );
  NAND2_X2 U9547 ( .A1(n8695), .A2(n8694), .ZN(n14098) );
  NAND2_X1 U9548 ( .A1(n10308), .A2(n6660), .ZN(n7531) );
  NAND2_X1 U9549 ( .A1(n14150), .A2(n7537), .ZN(n7534) );
  OAI22_X2 U9550 ( .A1(n14071), .A2(n7542), .B1(n7541), .B2(n6710), .ZN(n14022) );
  INV_X1 U9551 ( .A(n6717), .ZN(n8152) );
  OAI211_X1 U9552 ( .C1(n13134), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9941)
         );
  NAND2_X1 U9553 ( .A1(n8100), .A2(n12502), .ZN(n15116) );
  INV_X1 U9554 ( .A(n8892), .ZN(n9443) );
  NAND2_X1 U9555 ( .A1(n9053), .A2(n8886), .ZN(n9047) );
  NAND2_X1 U9556 ( .A1(n13196), .A2(n12003), .ZN(n13264) );
  OR2_X1 U9557 ( .A1(n9050), .A2(n9049), .ZN(n9052) );
  NAND2_X1 U9558 ( .A1(n11322), .A2(n9569), .ZN(n11380) );
  INV_X2 U9559 ( .A(n9592), .ZN(n11683) );
  OR2_X1 U9560 ( .A1(n9271), .A2(n8169), .ZN(n8187) );
  OR2_X1 U9561 ( .A1(n9271), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U9562 ( .A1(n8180), .A2(n8179), .ZN(n8934) );
  OAI21_X1 U9563 ( .B1(n11571), .B2(n11570), .A(n11569), .ZN(n11584) );
  AOI21_X1 U9564 ( .B1(n13400), .B2(n11921), .A(n11920), .ZN(n13388) );
  INV_X1 U9565 ( .A(n11361), .ZN(n11364) );
  AOI21_X2 U9566 ( .B1(n13397), .B2(n11946), .A(n11945), .ZN(n13383) );
  AOI21_X1 U9567 ( .B1(n13180), .B2(n13247), .A(n13248), .ZN(n13251) );
  NOR2_X1 U9568 ( .A1(n11584), .A2(n11582), .ZN(n11585) );
  NAND2_X1 U9569 ( .A1(n8580), .A2(n8579), .ZN(n8583) );
  XNOR2_X1 U9570 ( .A(n8732), .B(n8316), .ZN(n13690) );
  AND2_X4 U9571 ( .A1(n7705), .A2(n13144), .ZN(n8083) );
  OR2_X1 U9572 ( .A1(n13990), .A2(n14114), .ZN(n14673) );
  NAND2_X1 U9573 ( .A1(n8313), .A2(SI_26_), .ZN(n8315) );
  OR2_X1 U9574 ( .A1(n12179), .A2(n9122), .ZN(n8358) );
  XNOR2_X1 U9575 ( .A(n8760), .B(n8813), .ZN(n13997) );
  INV_X1 U9576 ( .A(n8220), .ZN(n8222) );
  INV_X1 U9577 ( .A(n12568), .ZN(n10720) );
  AND2_X1 U9578 ( .A1(n12248), .A2(n12251), .ZN(n7560) );
  AND2_X2 U9579 ( .A1(n8865), .A2(n8859), .ZN(n14764) );
  OR2_X1 U9580 ( .A1(n12339), .A2(n13131), .ZN(n7561) );
  INV_X1 U9581 ( .A(n14497), .ZN(n12785) );
  AND2_X1 U9582 ( .A1(n7943), .A2(n7942), .ZN(n14497) );
  OR2_X1 U9583 ( .A1(n14000), .A2(n14009), .ZN(n7563) );
  INV_X1 U9584 ( .A(n11317), .ZN(n13685) );
  AND2_X1 U9585 ( .A1(n13116), .A2(n12918), .ZN(n7564) );
  AND2_X1 U9586 ( .A1(n13130), .A2(n11303), .ZN(n7565) );
  AND2_X1 U9587 ( .A1(n11995), .A2(n11332), .ZN(n7566) );
  INV_X1 U9588 ( .A(n13841), .ZN(n8777) );
  INV_X1 U9589 ( .A(n14332), .ZN(n14323) );
  INV_X1 U9590 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8459) );
  INV_X1 U9591 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13137) );
  OR2_X1 U9592 ( .A1(n12155), .A2(n12154), .ZN(n7567) );
  AND2_X1 U9593 ( .A1(n12155), .A2(n12154), .ZN(n7568) );
  INV_X1 U9594 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13678) );
  OR2_X1 U9595 ( .A1(n12339), .A2(n13073), .ZN(n7569) );
  AOI21_X1 U9596 ( .B1(n12823), .B2(n6645), .A(n8086), .ZN(n12802) );
  NAND2_X1 U9597 ( .A1(n11311), .A2(n12991), .ZN(n7571) );
  INV_X1 U9598 ( .A(SI_18_), .ZN(n15493) );
  AND3_X1 U9599 ( .A1(n11673), .A2(n11672), .A3(n11671), .ZN(n7572) );
  INV_X2 U9600 ( .A(n14556), .ZN(n13441) );
  CLKBUF_X2 U9601 ( .A(P2_U3947), .Z(n13301) );
  INV_X1 U9602 ( .A(n8580), .ZN(n8763) );
  NOR2_X1 U9603 ( .A1(n12268), .A2(n13723), .ZN(n7573) );
  AND3_X1 U9604 ( .A1(n14241), .A2(n14240), .A3(n14239), .ZN(n7574) );
  INV_X1 U9605 ( .A(n12220), .ZN(n10019) );
  NOR2_X1 U9606 ( .A1(n8113), .A2(n10982), .ZN(n7575) );
  NOR2_X2 U9607 ( .A1(n9225), .A2(n8982), .ZN(P1_U4016) );
  NAND2_X2 U9608 ( .A1(n13990), .A2(n14665), .ZN(n14668) );
  INV_X2 U9609 ( .A(n14668), .ZN(n14678) );
  INV_X1 U9610 ( .A(n6656), .ZN(n15591) );
  INV_X1 U9611 ( .A(n11950), .ZN(n11923) );
  NOR2_X1 U9612 ( .A1(n13761), .A2(n13824), .ZN(n7576) );
  OR2_X1 U9613 ( .A1(n11380), .A2(n11324), .ZN(n11325) );
  OAI21_X1 U9614 ( .B1(n11337), .B2(n11380), .A(n11336), .ZN(n11338) );
  NAND2_X1 U9615 ( .A1(n11716), .A2(n11346), .ZN(n11348) );
  INV_X1 U9616 ( .A(n11362), .ZN(n11363) );
  INV_X1 U9617 ( .A(n11375), .ZN(n11376) );
  NAND2_X1 U9618 ( .A1(n11377), .A2(n11376), .ZN(n11378) );
  NAND2_X1 U9619 ( .A1(n11407), .A2(n11406), .ZN(n11414) );
  AOI22_X1 U9620 ( .A1(n13553), .A2(n11692), .B1(n13285), .B2(n11693), .ZN(
        n11487) );
  OAI21_X1 U9621 ( .B1(n7568), .B2(n12156), .A(n7567), .ZN(n12159) );
  INV_X1 U9622 ( .A(n11502), .ZN(n11507) );
  OAI21_X1 U9623 ( .B1(n11519), .B2(n11518), .A(n11517), .ZN(n11520) );
  INV_X1 U9624 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9439) );
  INV_X1 U9625 ( .A(n14060), .ZN(n8809) );
  INV_X1 U9626 ( .A(n10373), .ZN(n10375) );
  AND2_X1 U9627 ( .A1(n10940), .A2(n10939), .ZN(n10941) );
  INV_X1 U9628 ( .A(n11775), .ZN(n11778) );
  INV_X1 U9629 ( .A(n11115), .ZN(n11116) );
  INV_X1 U9630 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8579) );
  INV_X1 U9631 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7582) );
  AND2_X1 U9632 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n11601), .ZN(n11602) );
  INV_X1 U9633 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9855) );
  INV_X1 U9634 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n11264) );
  INV_X1 U9635 ( .A(P2_B_REG_SCAN_IN), .ZN(n11948) );
  NAND2_X1 U9636 ( .A1(n11117), .A2(n11116), .ZN(n11118) );
  INV_X1 U9637 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8644) );
  AND2_X1 U9638 ( .A1(n9350), .A2(n14708), .ZN(n8778) );
  INV_X1 U9639 ( .A(n12241), .ZN(n8813) );
  INV_X1 U9640 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U9641 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7052), .ZN(n14337) );
  INV_X1 U9642 ( .A(n12396), .ZN(n11862) );
  INV_X1 U9643 ( .A(n10154), .ZN(n8924) );
  INV_X1 U9644 ( .A(n7998), .ZN(n7694) );
  OR2_X1 U9645 ( .A1(n8081), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8091) );
  INV_X1 U9646 ( .A(n15046), .ZN(n12725) );
  INV_X1 U9647 ( .A(n12672), .ZN(n12676) );
  AND2_X1 U9648 ( .A1(n12694), .A2(n12535), .ZN(n12672) );
  INV_X1 U9649 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7671) );
  OAI211_X1 U9650 ( .C1(n11670), .C2(n11669), .A(n11673), .B(n11667), .ZN(
        n11709) );
  AND2_X1 U9651 ( .A1(n11926), .A2(n11631), .ZN(n12016) );
  INV_X1 U9652 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10954) );
  NOR2_X1 U9653 ( .A1(n10213), .A2(n10212), .ZN(n10269) );
  NAND2_X1 U9654 ( .A1(n9605), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9454) );
  INV_X1 U9655 ( .A(n11951), .ZN(n13367) );
  OR2_X1 U9656 ( .A1(n11265), .A2(n11264), .ZN(n11494) );
  INV_X1 U9657 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10521) );
  OR2_X1 U9658 ( .A1(n9601), .A2(n9562), .ZN(n9563) );
  INV_X1 U9659 ( .A(n9572), .ZN(n9460) );
  NAND2_X1 U9660 ( .A1(n9689), .A2(n8885), .ZN(n9051) );
  INV_X1 U9661 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8535) );
  INV_X1 U9662 ( .A(n10430), .ZN(n10431) );
  INV_X1 U9663 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8662) );
  OR2_X1 U9664 ( .A1(n8645), .A2(n8644), .ZN(n8663) );
  OR2_X1 U9665 ( .A1(n8521), .A2(n11129), .ZN(n8536) );
  AND2_X1 U9666 ( .A1(n14200), .A2(n13818), .ZN(n8749) );
  INV_X1 U9667 ( .A(n14126), .ZN(n8803) );
  INV_X1 U9668 ( .A(n14168), .ZN(n8633) );
  OR2_X1 U9669 ( .A1(n8444), .A2(n10191), .ZN(n8460) );
  INV_X1 U9670 ( .A(n9962), .ZN(n12029) );
  NAND2_X1 U9671 ( .A1(n10413), .A2(n8794), .ZN(n10569) );
  INV_X1 U9672 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8827) );
  INV_X1 U9673 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8584) );
  INV_X1 U9674 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15445) );
  OR2_X1 U9675 ( .A1(n8037), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8045) );
  OR2_X1 U9676 ( .A1(n7933), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U9677 ( .A1(n7694), .A2(n7693), .ZN(n8011) );
  OR2_X1 U9678 ( .A1(n8950), .A2(n8949), .ZN(n12454) );
  AND2_X1 U9679 ( .A1(n8178), .A2(n8177), .ZN(n8179) );
  INV_X1 U9680 ( .A(n15017), .ZN(n10702) );
  INV_X1 U9681 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15462) );
  NAND2_X1 U9682 ( .A1(n12731), .A2(n12754), .ZN(n12732) );
  OR2_X1 U9683 ( .A1(n9503), .A2(n12693), .ZN(n15003) );
  INV_X1 U9684 ( .A(n8128), .ZN(n12863) );
  INV_X1 U9685 ( .A(n12906), .ZN(n8004) );
  INV_X1 U9686 ( .A(n11235), .ZN(n11230) );
  INV_X1 U9687 ( .A(n13132), .ZN(n9934) );
  AND2_X1 U9688 ( .A1(n8190), .A2(n12676), .ZN(n9937) );
  OR2_X1 U9689 ( .A1(n7882), .A2(n10047), .ZN(n7996) );
  INV_X1 U9690 ( .A(n7882), .ZN(n7972) );
  AND2_X1 U9691 ( .A1(n12596), .A2(n12597), .ZN(n12512) );
  AND2_X1 U9692 ( .A1(n7603), .A2(n8190), .ZN(n12868) );
  OR2_X1 U9693 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .ZN(
        n7699) );
  INV_X1 U9694 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U9695 ( .A1(n11173), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11265) );
  NAND2_X1 U9696 ( .A1(n9438), .A2(n11767), .ZN(n9473) );
  AND2_X1 U9697 ( .A1(n11628), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n11643) );
  AND2_X1 U9698 ( .A1(n11544), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n11558) );
  INV_X1 U9699 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9642) );
  INV_X1 U9700 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10120) );
  INV_X1 U9701 ( .A(n14843), .ZN(n14798) );
  INV_X1 U9702 ( .A(n13283), .ZN(n13190) );
  OR2_X1 U9703 ( .A1(n9569), .A2(n11750), .ZN(n9572) );
  NOR2_X1 U9704 ( .A1(n10522), .A2(n10521), .ZN(n10760) );
  INV_X1 U9705 ( .A(n11730), .ZN(n10277) );
  AND2_X1 U9706 ( .A1(n11764), .A2(n9460), .ZN(n10097) );
  INV_X1 U9707 ( .A(n11737), .ZN(n11186) );
  INV_X1 U9708 ( .A(n9472), .ZN(n9556) );
  NOR2_X1 U9709 ( .A1(n8536), .A2(n8535), .ZN(n8551) );
  AND2_X1 U9710 ( .A1(n13717), .A2(n13715), .ZN(n11816) );
  NAND2_X1 U9711 ( .A1(n10432), .A2(n10431), .ZN(n10433) );
  NAND2_X1 U9712 ( .A1(n11791), .A2(n11792), .ZN(n11793) );
  OAI21_X1 U9713 ( .B1(n8855), .B2(n8854), .A(n8853), .ZN(n9219) );
  NOR2_X1 U9714 ( .A1(n9389), .A2(P1_U3086), .ZN(n12257) );
  NOR2_X1 U9715 ( .A1(n8616), .A2(n8224), .ZN(n8629) );
  INV_X1 U9716 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9156) );
  INV_X1 U9717 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10191) );
  INV_X1 U9718 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14356) );
  INV_X1 U9719 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U9720 ( .A1(n12201), .A2(n9084), .ZN(n14170) );
  INV_X1 U9721 ( .A(n12052), .ZN(n10082) );
  NAND2_X1 U9722 ( .A1(n8776), .A2(n12324), .ZN(n14087) );
  INV_X1 U9723 ( .A(n14743), .ZN(n14731) );
  INV_X1 U9724 ( .A(n8982), .ZN(n9015) );
  OAI21_X1 U9725 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14362), .A(n14361), .ZN(
        n14420) );
  INV_X1 U9726 ( .A(n12454), .ZN(n12416) );
  AOI22_X1 U9727 ( .A1(n12351), .A2(n12352), .B1(n12802), .B2(n11896), .ZN(
        n11898) );
  INV_X1 U9728 ( .A(n12459), .ZN(n12436) );
  INV_X1 U9729 ( .A(n12446), .ZN(n12456) );
  OR2_X1 U9730 ( .A1(n10802), .A2(n12676), .ZN(n15134) );
  AND2_X1 U9731 ( .A1(n8076), .A2(n8075), .ZN(n12353) );
  AND4_X1 U9732 ( .A1(n8003), .A2(n8002), .A3(n8001), .A4(n8000), .ZN(n12921)
         );
  INV_X1 U9733 ( .A(n15043), .ZN(n15047) );
  XNOR2_X1 U9734 ( .A(n12735), .B(n14497), .ZN(n14505) );
  INV_X1 U9735 ( .A(n15134), .ZN(n12993) );
  NAND2_X1 U9736 ( .A1(n8171), .A2(n12492), .ZN(n12987) );
  INV_X1 U9737 ( .A(n15108), .ZN(n15140) );
  OAI21_X1 U9738 ( .B1(n9937), .B2(n9934), .A(n8195), .ZN(n8196) );
  AND2_X1 U9739 ( .A1(n12868), .A2(n15189), .ZN(n15172) );
  INV_X1 U9740 ( .A(n15182), .ZN(n15193) );
  INV_X1 U9741 ( .A(n15172), .ZN(n15187) );
  NOR2_X1 U9742 ( .A1(n9272), .A2(n13133), .ZN(n9277) );
  XNOR2_X1 U9743 ( .A(n7590), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12694) );
  INV_X1 U9744 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7968) );
  AND2_X1 U9745 ( .A1(n7860), .A2(n7883), .ZN(n12774) );
  INV_X1 U9746 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7763) );
  AND2_X1 U9747 ( .A1(n9060), .A2(n9059), .ZN(n9070) );
  AND4_X1 U9748 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(
        n11944) );
  INV_X1 U9749 ( .A(n11658), .ZN(n11551) );
  AND2_X1 U9750 ( .A1(n9076), .A2(n13691), .ZN(n14843) );
  INV_X1 U9751 ( .A(n14765), .ZN(n14841) );
  INV_X1 U9752 ( .A(n13496), .ZN(n14563) );
  INV_X1 U9753 ( .A(n13528), .ZN(n14557) );
  NOR2_X1 U9754 ( .A1(n10094), .A2(n10097), .ZN(n9633) );
  OR2_X1 U9755 ( .A1(n11327), .A2(n15591), .ZN(n13655) );
  INV_X1 U9756 ( .A(n13655), .ZN(n14915) );
  AND2_X1 U9757 ( .A1(n10094), .A2(n9557), .ZN(n9558) );
  XNOR2_X1 U9758 ( .A(n8903), .B(n8902), .ZN(n10851) );
  AND2_X1 U9759 ( .A1(n9192), .A2(n9191), .ZN(n14816) );
  AND2_X1 U9760 ( .A1(n8551), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8568) );
  INV_X1 U9761 ( .A(n9353), .ZN(n9357) );
  INV_X1 U9762 ( .A(n14598), .ZN(n14585) );
  AND2_X1 U9763 ( .A1(n8678), .A2(n8677), .ZN(n13724) );
  AND2_X1 U9764 ( .A1(n9092), .A2(n6843), .ZN(n13966) );
  AND2_X1 U9765 ( .A1(n9092), .A2(n9089), .ZN(n13963) );
  INV_X1 U9766 ( .A(n14167), .ZN(n14188) );
  INV_X1 U9767 ( .A(n14714), .ZN(n9961) );
  INV_X1 U9768 ( .A(n14752), .ZN(n14280) );
  NAND2_X1 U9769 ( .A1(n14087), .A2(n14221), .ZN(n14752) );
  NAND2_X1 U9770 ( .A1(n8852), .A2(n9017), .ZN(n9012) );
  INV_X1 U9771 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8545) );
  AND2_X1 U9772 ( .A1(n8489), .A2(n8475), .ZN(n9309) );
  AND2_X1 U9773 ( .A1(n9502), .A2(n9501), .ZN(n15095) );
  INV_X1 U9774 ( .A(n12451), .ZN(n12418) );
  NAND2_X1 U9775 ( .A1(n8947), .A2(n8946), .ZN(n12446) );
  AND2_X1 U9776 ( .A1(n12472), .A2(n8144), .ZN(n12487) );
  INV_X1 U9777 ( .A(n12650), .ZN(n12704) );
  OR2_X1 U9778 ( .A1(n8934), .A2(n13133), .ZN(n12720) );
  INV_X1 U9779 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14968) );
  INV_X1 U9780 ( .A(n15096), .ZN(n15077) );
  OR2_X1 U9781 ( .A1(n9503), .A2(n9499), .ZN(n15102) );
  INV_X1 U9782 ( .A(n15141), .ZN(n13002) );
  NAND2_X1 U9783 ( .A1(n15213), .A2(n15193), .ZN(n13073) );
  INV_X1 U9784 ( .A(n15213), .ZN(n15210) );
  INV_X1 U9785 ( .A(n15197), .ZN(n15195) );
  AND2_X2 U9786 ( .A1(n8184), .A2(n12690), .ZN(n15197) );
  INV_X1 U9787 ( .A(SI_29_), .ZN(n13142) );
  INV_X1 U9788 ( .A(SI_14_), .ZN(n15380) );
  INV_X1 U9789 ( .A(n15000), .ZN(n10701) );
  INV_X1 U9790 ( .A(n11424), .ZN(n14910) );
  INV_X1 U9791 ( .A(n14558), .ZN(n14573) );
  NAND2_X1 U9792 ( .A1(n9641), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13270) );
  INV_X1 U9793 ( .A(n13601), .ZN(n13481) );
  INV_X1 U9794 ( .A(n13273), .ZN(n13242) );
  INV_X1 U9795 ( .A(n13267), .ZN(n13281) );
  NAND2_X1 U9796 ( .A1(n11179), .A2(n11178), .ZN(n13286) );
  NAND2_X1 U9797 ( .A1(n14779), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14765) );
  NAND2_X1 U9798 ( .A1(n9076), .A2(n11766), .ZN(n14811) );
  INV_X1 U9799 ( .A(n13441), .ZN(n15599) );
  OR2_X1 U9800 ( .A1(n15599), .A2(n11321), .ZN(n15596) );
  AND2_X1 U9801 ( .A1(n10099), .A2(n15592), .ZN(n14556) );
  INV_X1 U9802 ( .A(n14943), .ZN(n14940) );
  AND3_X2 U9803 ( .A1(n9634), .A2(n14855), .A3(n9633), .ZN(n14943) );
  OR2_X1 U9804 ( .A1(n13625), .A2(n13624), .ZN(n13671) );
  AND4_X1 U9805 ( .A1(n14878), .A2(n14877), .A3(n14876), .A4(n14875), .ZN(
        n14930) );
  INV_X1 U9806 ( .A(n14925), .ZN(n14923) );
  NOR2_X1 U9807 ( .A1(n14857), .A2(n14850), .ZN(n14851) );
  INV_X1 U9808 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9691) );
  INV_X1 U9809 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9045) );
  INV_X2 U9810 ( .A(n13676), .ZN(n13693) );
  INV_X1 U9811 ( .A(n12082), .ZN(n11135) );
  OR3_X1 U9812 ( .A1(n9224), .A2(n9223), .A3(n9222), .ZN(n14598) );
  NAND4_X1 U9813 ( .A1(n8234), .A2(n8233), .A3(n8232), .A4(n8231), .ZN(n14042)
         );
  INV_X1 U9814 ( .A(n13724), .ZN(n13819) );
  CLKBUF_X1 U9815 ( .A(P1_U4016), .Z(n13847) );
  INV_X1 U9816 ( .A(n13966), .ZN(n14643) );
  INV_X1 U9817 ( .A(n13963), .ZN(n14645) );
  OR2_X1 U9818 ( .A1(n14678), .A2(n9925), .ZN(n14156) );
  OR2_X1 U9819 ( .A1(n14678), .A2(n9976), .ZN(n14167) );
  INV_X1 U9820 ( .A(n9995), .ZN(n9932) );
  INV_X1 U9821 ( .A(n14764), .ZN(n14761) );
  INV_X1 U9822 ( .A(n13985), .ZN(n14288) );
  INV_X1 U9823 ( .A(n14185), .ZN(n14310) );
  INV_X1 U9824 ( .A(n14755), .ZN(n14753) );
  AND2_X2 U9825 ( .A1(n8865), .A2(n9918), .ZN(n14755) );
  AND2_X2 U9826 ( .A1(n9924), .A2(n9012), .ZN(n14706) );
  INV_X1 U9827 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9762) );
  INV_X1 U9828 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9339) );
  INV_X1 U9829 ( .A(n12720), .ZN(P3_U3897) );
  NOR2_X1 U9830 ( .A1(n9060), .A2(P2_U3088), .ZN(P2_U3947) );
  NOR2_X1 U9831 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n7578) );
  AND4_X2 U9832 ( .A1(n7578), .A2(n7577), .A3(n7794), .A4(n7763), .ZN(n7579)
         );
  NOR2_X1 U9833 ( .A1(n7588), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U9834 ( .A1(n7955), .A2(n7582), .ZN(n7940) );
  NOR2_X1 U9835 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7587) );
  NOR2_X1 U9836 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7586) );
  NAND2_X1 U9837 ( .A1(n7666), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U9838 ( .A1(n6744), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7592) );
  NAND2_X1 U9839 ( .A1(n12694), .A2(n10049), .ZN(n7597) );
  INV_X1 U9840 ( .A(n7593), .ZN(n7594) );
  NAND2_X1 U9841 ( .A1(n7594), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7595) );
  MUX2_X1 U9842 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7595), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n7596) );
  AOI21_X1 U9843 ( .B1(n12525), .B2(n7597), .A(n12535), .ZN(n7600) );
  NAND2_X1 U9844 ( .A1(n10250), .A2(n10049), .ZN(n7598) );
  INV_X1 U9845 ( .A(n12694), .ZN(n8192) );
  AND2_X1 U9846 ( .A1(n7598), .A2(n8192), .ZN(n7599) );
  OR2_X1 U9847 ( .A1(n7600), .A2(n7599), .ZN(n8937) );
  NAND2_X1 U9848 ( .A1(n12769), .A2(n10049), .ZN(n12692) );
  NOR2_X1 U9849 ( .A1(n12692), .A2(n15193), .ZN(n7601) );
  NAND2_X1 U9850 ( .A1(n8937), .A2(n7601), .ZN(n7603) );
  AND2_X1 U9851 ( .A1(n12694), .A2(n8191), .ZN(n7602) );
  NAND2_X1 U9852 ( .A1(n12769), .A2(n7602), .ZN(n8190) );
  NAND2_X1 U9853 ( .A1(n12525), .A2(n10049), .ZN(n15137) );
  OR2_X1 U9854 ( .A1(n15137), .A2(n12694), .ZN(n15189) );
  INV_X1 U9855 ( .A(n7726), .ZN(n7604) );
  NAND2_X1 U9856 ( .A1(n7727), .A2(n7604), .ZN(n7606) );
  INV_X1 U9857 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U9858 ( .A1(n8959), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7605) );
  NAND2_X1 U9859 ( .A1(n7606), .A2(n7605), .ZN(n7735) );
  INV_X1 U9860 ( .A(n7735), .ZN(n7608) );
  INV_X1 U9861 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U9862 ( .A1(n9593), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U9863 ( .A1(n7608), .A2(n7607), .ZN(n7610) );
  NAND2_X1 U9864 ( .A1(n9030), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7609) );
  AND2_X1 U9865 ( .A1(n9027), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7611) );
  NAND2_X1 U9866 ( .A1(n8967), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7612) );
  NAND2_X1 U9867 ( .A1(n9033), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7614) );
  INV_X1 U9868 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8972) );
  NAND2_X1 U9869 ( .A1(n8972), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U9870 ( .A1(n7614), .A2(n7613), .ZN(n7757) );
  NAND2_X1 U9871 ( .A1(n9032), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U9872 ( .A1(n8978), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U9873 ( .A1(n7617), .A2(n7615), .ZN(n7775) );
  INV_X1 U9874 ( .A(n7775), .ZN(n7616) );
  NAND2_X1 U9875 ( .A1(n7777), .A2(n7617), .ZN(n7799) );
  INV_X1 U9876 ( .A(n7798), .ZN(n7618) );
  NAND2_X1 U9877 ( .A1(n9023), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7620) );
  NAND2_X1 U9878 ( .A1(n9021), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7619) );
  NAND2_X1 U9879 ( .A1(n7620), .A2(n7619), .ZN(n7808) );
  NOR2_X1 U9880 ( .A1(n9045), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7621) );
  NAND2_X1 U9881 ( .A1(n9045), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7622) );
  NAND2_X1 U9882 ( .A1(n9196), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7624) );
  INV_X1 U9883 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U9884 ( .A1(n9194), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7623) );
  NAND2_X1 U9885 ( .A1(n7856), .A2(n7624), .ZN(n7872) );
  NAND2_X1 U9886 ( .A1(n9218), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U9887 ( .A1(n9215), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7626) );
  XNOR2_X1 U9888 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n7888) );
  XNOR2_X1 U9889 ( .A(n7627), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U9890 ( .A1(n7892), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U9891 ( .A1(n7627), .A2(n9364), .ZN(n7628) );
  NAND2_X1 U9892 ( .A1(n7629), .A2(n7628), .ZN(n7905) );
  XNOR2_X1 U9893 ( .A(n9721), .B(P1_DATAO_REG_14__SCAN_IN), .ZN(n7904) );
  INV_X1 U9894 ( .A(n7904), .ZN(n7630) );
  NAND2_X1 U9895 ( .A1(n7905), .A2(n7630), .ZN(n7632) );
  NAND2_X1 U9896 ( .A1(n9721), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U9897 ( .A1(n7632), .A2(n7631), .ZN(n7966) );
  XNOR2_X1 U9898 ( .A(n9767), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n7965) );
  INV_X1 U9899 ( .A(n7965), .ZN(n7633) );
  NAND2_X1 U9900 ( .A1(n9767), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7634) );
  XNOR2_X1 U9901 ( .A(n9693), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n7953) );
  INV_X1 U9902 ( .A(n7953), .ZN(n7635) );
  NAND2_X1 U9903 ( .A1(n9761), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7636) );
  INV_X1 U9904 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U9905 ( .A1(n10014), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7639) );
  INV_X1 U9906 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U9907 ( .A1(n10012), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9908 ( .A1(n7639), .A2(n7638), .ZN(n7925) );
  XNOR2_X1 U9909 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n7915) );
  INV_X1 U9910 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10198) );
  NAND2_X1 U9911 ( .A1(n10198), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7640) );
  XNOR2_X1 U9912 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .ZN(n7994) );
  NAND2_X1 U9913 ( .A1(n12263), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7642) );
  INV_X1 U9914 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U9915 ( .A1(n10584), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7644) );
  INV_X1 U9916 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U9917 ( .A1(n10585), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7643) );
  NAND2_X1 U9918 ( .A1(n7644), .A2(n7643), .ZN(n8005) );
  INV_X1 U9919 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n15362) );
  NAND2_X1 U9920 ( .A1(n15362), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7646) );
  INV_X1 U9921 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15395) );
  NAND2_X1 U9922 ( .A1(n15395), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7645) );
  INV_X1 U9923 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7647) );
  XNOR2_X1 U9924 ( .A(n7647), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n8031) );
  INV_X1 U9925 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10965) );
  NAND2_X1 U9926 ( .A1(n7649), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7650) );
  INV_X1 U9927 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U9928 ( .A1(n11214), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7653) );
  INV_X1 U9929 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11211) );
  NAND2_X1 U9930 ( .A1(n11211), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7652) );
  AND2_X1 U9931 ( .A1(n7653), .A2(n7652), .ZN(n8050) );
  INV_X1 U9932 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15349) );
  NAND2_X1 U9933 ( .A1(n15349), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7655) );
  INV_X1 U9934 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11316) );
  NAND2_X1 U9935 ( .A1(n11316), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7654) );
  AND2_X1 U9936 ( .A1(n7655), .A2(n7654), .ZN(n8064) );
  NAND2_X1 U9937 ( .A1(n8065), .A2(n8064), .ZN(n8066) );
  INV_X1 U9938 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14331) );
  NAND2_X1 U9939 ( .A1(n14331), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7658) );
  INV_X1 U9940 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13692) );
  NAND2_X1 U9941 ( .A1(n13692), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U9942 ( .A1(n7658), .A2(n7656), .ZN(n8077) );
  INV_X1 U9943 ( .A(n8077), .ZN(n7657) );
  NAND2_X1 U9944 ( .A1(n8078), .A2(n7657), .ZN(n7659) );
  INV_X1 U9945 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13689) );
  NAND2_X1 U9946 ( .A1(n13689), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9947 ( .A1(n8088), .A2(n7660), .ZN(n7662) );
  INV_X1 U9948 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12265) );
  NAND2_X1 U9949 ( .A1(n12265), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U9950 ( .A1(n7662), .A2(n7661), .ZN(n7664) );
  XNOR2_X1 U9951 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n7663) );
  NAND2_X1 U9952 ( .A1(n7664), .A2(n7663), .ZN(n12345) );
  OR2_X1 U9953 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  NAND2_X1 U9954 ( .A1(n12345), .A2(n7665), .ZN(n13143) );
  INV_X1 U9955 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7667) );
  NAND3_X1 U9956 ( .A1(n7674), .A2(n7673), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7676) );
  OR2_X1 U9957 ( .A1(n13143), .A2(n8089), .ZN(n7678) );
  NAND2_X2 U9958 ( .A1(n9491), .A2(n9468), .ZN(n7882) );
  INV_X1 U9959 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n7740) );
  INV_X1 U9960 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U9961 ( .A1(n7740), .A2(n7679), .ZN(n7769) );
  INV_X1 U9962 ( .A(n7769), .ZN(n7680) );
  INV_X1 U9963 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U9964 ( .A1(n7680), .A2(n9713), .ZN(n7787) );
  INV_X1 U9965 ( .A(n7802), .ZN(n7682) );
  INV_X1 U9966 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U9967 ( .A1(n7682), .A2(n7681), .ZN(n7824) );
  OR2_X2 U9968 ( .A1(n7824), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7850) );
  INV_X1 U9969 ( .A(n7850), .ZN(n7684) );
  NOR2_X1 U9970 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_REG3_REG_9__SCAN_IN), 
        .ZN(n7683) );
  NAND2_X1 U9971 ( .A1(n7684), .A2(n7683), .ZN(n7863) );
  OR2_X2 U9972 ( .A1(n7876), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7897) );
  INV_X1 U9973 ( .A(n7897), .ZN(n7686) );
  INV_X1 U9974 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U9975 ( .A1(n7686), .A2(n7685), .ZN(n7909) );
  INV_X1 U9976 ( .A(n7909), .ZN(n7688) );
  INV_X1 U9977 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U9978 ( .A1(n7688), .A2(n7687), .ZN(n7975) );
  INV_X1 U9979 ( .A(n7977), .ZN(n7690) );
  INV_X1 U9980 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U9981 ( .A1(n7690), .A2(n7689), .ZN(n7960) );
  INV_X1 U9982 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7691) );
  INV_X1 U9983 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7693) );
  INV_X1 U9984 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12431) );
  INV_X1 U9985 ( .A(n8056), .ZN(n7696) );
  INV_X1 U9986 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n12384) );
  NAND2_X1 U9987 ( .A1(n7696), .A2(n12384), .ZN(n8070) );
  INV_X1 U9988 ( .A(n8091), .ZN(n7698) );
  INV_X1 U9989 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U9990 ( .A1(n7698), .A2(n7697), .ZN(n12337) );
  OR2_X1 U9991 ( .A1(n12337), .A2(n7875), .ZN(n12472) );
  INV_X1 U9992 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n7709) );
  NAND2_X1 U9993 ( .A1(n8083), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U9994 ( .A1(n8138), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7707) );
  OAI211_X1 U9995 ( .C1(n7709), .C2(n7919), .A(n7708), .B(n7707), .ZN(n7710)
         );
  INV_X1 U9996 ( .A(n7710), .ZN(n7711) );
  NAND2_X1 U9997 ( .A1(n12472), .A2(n7711), .ZN(n12700) );
  NAND2_X1 U9998 ( .A1(n12339), .A2(n12700), .ZN(n12461) );
  INV_X1 U9999 ( .A(n12339), .ZN(n7712) );
  INV_X1 U10000 ( .A(n12700), .ZN(n12803) );
  NAND2_X1 U10001 ( .A1(n7712), .A2(n12803), .ZN(n12484) );
  NAND2_X1 U10002 ( .A1(n8083), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7716) );
  INV_X2 U10003 ( .A(n7919), .ZN(n8058) );
  NAND2_X1 U10004 ( .A1(n8058), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U10005 ( .A1(n6644), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U10006 ( .A1(n8138), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7713) );
  INV_X1 U10007 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10008 ( .A1(n8354), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U10009 ( .A1(n7726), .A2(n7717), .ZN(n7718) );
  MUX2_X1 U10010 ( .A(n7718), .B(SI_0_), .S(n9468), .Z(n13145) );
  MUX2_X1 U10011 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13145), .S(n9491), .Z(n8099)
         );
  NOR2_X1 U10012 ( .A1(n15125), .A2(n9943), .ZN(n9791) );
  NAND2_X1 U10013 ( .A1(n8058), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U10014 ( .A1(n6645), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7722) );
  NAND2_X1 U10015 ( .A1(n7719), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7721) );
  NAND2_X1 U10016 ( .A1(n8083), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7720) );
  AND4_X2 U10017 ( .A1(n7723), .A2(n7722), .A3(n7721), .A4(n7720), .ZN(n15112)
         );
  INV_X1 U10018 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U10019 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n7724) );
  INV_X1 U10020 ( .A(SI_1_), .ZN(n8960) );
  OR2_X1 U10021 ( .A1(n7882), .A2(n8960), .ZN(n7729) );
  XNOR2_X1 U10022 ( .A(n7727), .B(n7726), .ZN(n8961) );
  OR2_X1 U10023 ( .A1(n8089), .A2(n8961), .ZN(n7728) );
  OAI211_X1 U10024 ( .C1(n9491), .C2(n9506), .A(n7729), .B(n7728), .ZN(n8911)
         );
  NAND2_X1 U10025 ( .A1(n9791), .A2(n12539), .ZN(n8908) );
  NAND2_X1 U10026 ( .A1(n15112), .A2(n8911), .ZN(n12541) );
  NAND2_X1 U10027 ( .A1(n8908), .A2(n12541), .ZN(n15105) );
  NAND2_X1 U10028 ( .A1(n8058), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U10029 ( .A1(n8138), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7732) );
  NAND2_X1 U10030 ( .A1(n6644), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U10031 ( .A1(n8083), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7730) );
  XNOR2_X1 U10032 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7734) );
  XNOR2_X1 U10033 ( .A(n7735), .B(n7734), .ZN(n9009) );
  OR2_X1 U10034 ( .A1(n8089), .A2(n9009), .ZN(n7738) );
  OR2_X1 U10035 ( .A1(n9491), .A2(n9523), .ZN(n7737) );
  NAND2_X1 U10036 ( .A1(n15135), .A2(n8915), .ZN(n12546) );
  INV_X1 U10037 ( .A(n15135), .ZN(n12718) );
  NAND2_X1 U10038 ( .A1(n12718), .A2(n15106), .ZN(n12545) );
  NAND2_X1 U10039 ( .A1(n12546), .A2(n12545), .ZN(n12502) );
  NAND2_X1 U10040 ( .A1(n15104), .A2(n12546), .ZN(n10500) );
  NAND2_X1 U10041 ( .A1(n8058), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U10042 ( .A1(n8083), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U10043 ( .A1(n6644), .A2(n7740), .ZN(n7743) );
  NAND2_X1 U10044 ( .A1(n12467), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7742) );
  OR2_X1 U10045 ( .A1(n7882), .A2(SI_3_), .ZN(n7751) );
  XNOR2_X1 U10046 ( .A(n9027), .B(P1_DATAO_REG_3__SCAN_IN), .ZN(n7746) );
  XNOR2_X1 U10047 ( .A(n7747), .B(n7746), .ZN(n8990) );
  OR2_X1 U10048 ( .A1(n8089), .A2(n8990), .ZN(n7750) );
  XNOR2_X1 U10049 ( .A(n7748), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9708) );
  OR2_X1 U10050 ( .A1(n9491), .A2(n9708), .ZN(n7749) );
  NAND2_X1 U10051 ( .A1(n15111), .A2(n15155), .ZN(n12549) );
  INV_X1 U10052 ( .A(n15111), .ZN(n12717) );
  INV_X1 U10053 ( .A(n15155), .ZN(n9892) );
  NAND2_X1 U10054 ( .A1(n12717), .A2(n9892), .ZN(n12550) );
  NAND2_X1 U10055 ( .A1(n10500), .A2(n12507), .ZN(n10499) );
  NAND2_X1 U10056 ( .A1(n10499), .A2(n12549), .ZN(n10244) );
  NAND2_X1 U10057 ( .A1(n8058), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U10058 ( .A1(n12467), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U10059 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7752) );
  NAND2_X1 U10060 ( .A1(n7769), .A2(n7752), .ZN(n10251) );
  NAND2_X1 U10061 ( .A1(n6644), .A2(n10251), .ZN(n7754) );
  NAND2_X1 U10062 ( .A1(n8083), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7753) );
  OR2_X1 U10063 ( .A1(n7882), .A2(SI_4_), .ZN(n7767) );
  NAND2_X1 U10064 ( .A1(n7758), .A2(n7757), .ZN(n7759) );
  AND2_X1 U10065 ( .A1(n7760), .A2(n7759), .ZN(n8962) );
  OR2_X1 U10066 ( .A1(n8089), .A2(n8962), .ZN(n7766) );
  INV_X1 U10067 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7761) );
  NAND2_X1 U10068 ( .A1(n7762), .A2(n7761), .ZN(n7779) );
  NAND2_X1 U10069 ( .A1(n7779), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7764) );
  XNOR2_X1 U10070 ( .A(n7764), .B(n7763), .ZN(n14955) );
  INV_X1 U10071 ( .A(n14955), .ZN(n9706) );
  OR2_X1 U10072 ( .A1(n9491), .A2(n9706), .ZN(n7765) );
  INV_X1 U10073 ( .A(n10252), .ZN(n15160) );
  NAND2_X1 U10074 ( .A1(n12716), .A2(n15160), .ZN(n12555) );
  NAND2_X1 U10075 ( .A1(n10501), .A2(n10252), .ZN(n12554) );
  NAND2_X1 U10076 ( .A1(n10244), .A2(n8097), .ZN(n7768) );
  NAND2_X1 U10077 ( .A1(n7768), .A2(n12554), .ZN(n10398) );
  NAND2_X1 U10078 ( .A1(n8083), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7774) );
  INV_X2 U10079 ( .A(n7919), .ZN(n8139) );
  NAND2_X1 U10080 ( .A1(n8139), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U10081 ( .A1(n7769), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U10082 ( .A1(n7787), .A2(n7770), .ZN(n10487) );
  NAND2_X1 U10083 ( .A1(n6645), .A2(n10487), .ZN(n7772) );
  NAND2_X1 U10084 ( .A1(n8138), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7771) );
  OR2_X1 U10085 ( .A1(n7882), .A2(SI_5_), .ZN(n7786) );
  NAND2_X1 U10086 ( .A1(n7776), .A2(n7775), .ZN(n7778) );
  AND2_X1 U10087 ( .A1(n7778), .A2(n7777), .ZN(n8998) );
  OR2_X1 U10088 ( .A1(n8089), .A2(n8998), .ZN(n7785) );
  NAND2_X1 U10089 ( .A1(n7781), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7780) );
  MUX2_X1 U10090 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7780), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n7783) );
  INV_X1 U10091 ( .A(n7795), .ZN(n7782) );
  NAND2_X1 U10092 ( .A1(n7783), .A2(n7782), .ZN(n10385) );
  INV_X1 U10093 ( .A(n10385), .ZN(n10380) );
  OR2_X1 U10094 ( .A1(n9491), .A2(n10380), .ZN(n7784) );
  NAND2_X1 U10095 ( .A1(n10405), .A2(n15165), .ZN(n12559) );
  INV_X1 U10096 ( .A(n10405), .ZN(n12715) );
  INV_X1 U10097 ( .A(n15165), .ZN(n8098) );
  NAND2_X1 U10098 ( .A1(n12715), .A2(n8098), .ZN(n12563) );
  NAND2_X1 U10099 ( .A1(n8083), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U10100 ( .A1(n8139), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U10101 ( .A1(n7787), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U10102 ( .A1(n7802), .A2(n7788), .ZN(n10409) );
  NAND2_X1 U10103 ( .A1(n6645), .A2(n10409), .ZN(n7790) );
  NAND2_X1 U10104 ( .A1(n12467), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7789) );
  AND4_X2 U10105 ( .A1(n7792), .A2(n7791), .A3(n7790), .A4(n7789), .ZN(n10723)
         );
  NOR2_X1 U10106 ( .A1(n7795), .A2(n13137), .ZN(n7793) );
  MUX2_X1 U10107 ( .A(n13137), .B(n7793), .S(P3_IR_REG_6__SCAN_IN), .Z(n7797)
         );
  NAND2_X1 U10108 ( .A1(n7795), .A2(n7794), .ZN(n7832) );
  INV_X1 U10109 ( .A(n7832), .ZN(n7796) );
  INV_X1 U10110 ( .A(SI_6_), .ZN(n8996) );
  XNOR2_X1 U10111 ( .A(n7799), .B(n7798), .ZN(n8997) );
  OR2_X1 U10112 ( .A1(n8089), .A2(n8997), .ZN(n7800) );
  OAI211_X1 U10113 ( .C1(n9491), .C2(n14985), .A(n7801), .B(n7800), .ZN(n10410) );
  NAND2_X1 U10114 ( .A1(n10723), .A2(n10410), .ZN(n12571) );
  INV_X1 U10115 ( .A(n10410), .ZN(n15171) );
  NAND2_X1 U10116 ( .A1(n8083), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10117 ( .A1(n8139), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U10118 ( .A1(n7802), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7803) );
  NAND2_X1 U10119 ( .A1(n7824), .A2(n7803), .ZN(n10729) );
  NAND2_X1 U10120 ( .A1(n6645), .A2(n10729), .ZN(n7805) );
  NAND2_X1 U10121 ( .A1(n12467), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7804) );
  OR2_X1 U10122 ( .A1(n7882), .A2(SI_7_), .ZN(n7816) );
  NAND2_X1 U10123 ( .A1(n7809), .A2(n7808), .ZN(n7810) );
  AND2_X1 U10124 ( .A1(n7811), .A2(n7810), .ZN(n8993) );
  OR2_X1 U10125 ( .A1(n8089), .A2(n8993), .ZN(n7815) );
  NAND2_X1 U10126 ( .A1(n7832), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7813) );
  INV_X1 U10127 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7812) );
  XNOR2_X1 U10128 ( .A(n7813), .B(n7812), .ZN(n10689) );
  INV_X1 U10129 ( .A(n10689), .ZN(n10698) );
  OR2_X1 U10130 ( .A1(n9491), .A2(n10698), .ZN(n7814) );
  NAND2_X1 U10131 ( .A1(n12575), .A2(n12534), .ZN(n12567) );
  INV_X1 U10132 ( .A(n12575), .ZN(n12713) );
  INV_X1 U10133 ( .A(n12534), .ZN(n15177) );
  NAND2_X1 U10134 ( .A1(n12713), .A2(n15177), .ZN(n7817) );
  NAND2_X1 U10135 ( .A1(n12567), .A2(n7817), .ZN(n12568) );
  AND2_X1 U10136 ( .A1(n10714), .A2(n10720), .ZN(n7818) );
  NAND2_X1 U10137 ( .A1(n10398), .A2(n7818), .ZN(n7823) );
  INV_X1 U10138 ( .A(n7819), .ZN(n7821) );
  AND2_X1 U10139 ( .A1(n12559), .A2(n12571), .ZN(n7820) );
  OR2_X1 U10140 ( .A1(n7821), .A2(n7820), .ZN(n10715) );
  OR2_X1 U10141 ( .A1(n12568), .A2(n10715), .ZN(n7822) );
  NAND2_X1 U10142 ( .A1(n8139), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U10143 ( .A1(n8138), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U10144 ( .A1(n7824), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U10145 ( .A1(n7850), .A2(n7825), .ZN(n10807) );
  NAND2_X1 U10146 ( .A1(n6645), .A2(n10807), .ZN(n7827) );
  NAND2_X1 U10147 ( .A1(n8083), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7826) );
  NAND4_X1 U10148 ( .A1(n7829), .A2(n7828), .A3(n7827), .A4(n7826), .ZN(n12712) );
  INV_X1 U10149 ( .A(SI_8_), .ZN(n8968) );
  OR2_X1 U10150 ( .A1(n7882), .A2(n8968), .ZN(n7836) );
  XNOR2_X1 U10151 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7830) );
  XNOR2_X1 U10152 ( .A(n7831), .B(n7830), .ZN(n8969) );
  OR2_X1 U10153 ( .A1(n8089), .A2(n8969), .ZN(n7835) );
  OAI21_X1 U10154 ( .B1(n7832), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7833) );
  XNOR2_X1 U10155 ( .A(n7833), .B(P3_IR_REG_8__SCAN_IN), .ZN(n15000) );
  OR2_X1 U10156 ( .A1(n9491), .A2(n10701), .ZN(n7834) );
  XNOR2_X1 U10157 ( .A(n12712), .B(n15183), .ZN(n10788) );
  INV_X1 U10158 ( .A(n12712), .ZN(n10611) );
  INV_X1 U10159 ( .A(n15183), .ZN(n10803) );
  NAND2_X1 U10160 ( .A1(n10611), .A2(n10803), .ZN(n12576) );
  XNOR2_X1 U10161 ( .A(n9045), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n7837) );
  XNOR2_X1 U10162 ( .A(n7838), .B(n7837), .ZN(n8979) );
  OR2_X1 U10163 ( .A1(n8089), .A2(n8979), .ZN(n7843) );
  OR2_X1 U10164 ( .A1(n7882), .A2(SI_9_), .ZN(n7842) );
  OR2_X1 U10165 ( .A1(n7839), .A2(n13137), .ZN(n7840) );
  XNOR2_X1 U10166 ( .A(n7840), .B(n7857), .ZN(n15017) );
  OR2_X1 U10167 ( .A1(n9491), .A2(n10702), .ZN(n7841) );
  NAND2_X1 U10168 ( .A1(n8083), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7847) );
  NAND2_X1 U10169 ( .A1(n8139), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7846) );
  XNOR2_X1 U10170 ( .A(n7850), .B(P3_REG3_REG_9__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U10171 ( .A1(n6645), .A2(n10874), .ZN(n7845) );
  NAND2_X1 U10172 ( .A1(n12467), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7844) );
  NAND4_X1 U10173 ( .A1(n7847), .A2(n7846), .A3(n7845), .A4(n7844), .ZN(n12711) );
  INV_X1 U10174 ( .A(n12711), .ZN(n10733) );
  OAI21_X1 U10175 ( .B1(n10867), .B2(n15194), .A(n10733), .ZN(n7849) );
  NAND2_X1 U10176 ( .A1(n10867), .A2(n15194), .ZN(n7848) );
  NAND2_X1 U10177 ( .A1(n7849), .A2(n7848), .ZN(n10923) );
  NAND2_X1 U10178 ( .A1(n8139), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7854) );
  OAI21_X1 U10179 ( .B1(n7850), .B2(P3_REG3_REG_9__SCAN_IN), .A(
        P3_REG3_REG_10__SCAN_IN), .ZN(n7851) );
  NAND2_X1 U10180 ( .A1(n7851), .A2(n7863), .ZN(n10925) );
  NAND2_X1 U10181 ( .A1(n6645), .A2(n10925), .ZN(n7853) );
  NAND2_X1 U10182 ( .A1(n8083), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7852) );
  NAND2_X1 U10183 ( .A1(n6907), .A2(n6797), .ZN(n7855) );
  AND2_X1 U10184 ( .A1(n7856), .A2(n7855), .ZN(n9024) );
  OR2_X1 U10185 ( .A1(n8089), .A2(n9024), .ZN(n7862) );
  NAND2_X1 U10186 ( .A1(n7839), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U10187 ( .A1(n7859), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7858) );
  MUX2_X1 U10188 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7858), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n7860) );
  OR2_X1 U10189 ( .A1(n9491), .A2(n12774), .ZN(n7861) );
  NAND2_X1 U10190 ( .A1(n11028), .A2(n10926), .ZN(n12585) );
  NAND2_X1 U10191 ( .A1(n12585), .A2(n12586), .ZN(n12505) );
  OR2_X2 U10192 ( .A1(n10923), .A2(n12505), .ZN(n11002) );
  NAND2_X1 U10193 ( .A1(n11002), .A2(n12586), .ZN(n10977) );
  NAND2_X1 U10194 ( .A1(n8083), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U10195 ( .A1(n8139), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U10196 ( .A1(n7863), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U10197 ( .A1(n7876), .A2(n7864), .ZN(n10978) );
  NAND2_X1 U10198 ( .A1(n6645), .A2(n10978), .ZN(n7867) );
  NAND2_X1 U10199 ( .A1(n8138), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7866) );
  NAND4_X1 U10200 ( .A1(n7869), .A2(n7868), .A3(n7867), .A4(n7866), .ZN(n12709) );
  NAND2_X1 U10201 ( .A1(n7883), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7870) );
  XNOR2_X1 U10202 ( .A(n7870), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12775) );
  INV_X1 U10203 ( .A(n12775), .ZN(n15031) );
  XNOR2_X1 U10204 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7871) );
  XNOR2_X1 U10205 ( .A(n7872), .B(n7871), .ZN(n9026) );
  OR2_X1 U10206 ( .A1(n9026), .A2(n8089), .ZN(n7874) );
  OAI211_X1 U10207 ( .C1(n9491), .C2(n15031), .A(n7874), .B(n7873), .ZN(n11037) );
  INV_X1 U10208 ( .A(n11037), .ZN(n14538) );
  XNOR2_X1 U10209 ( .A(n12709), .B(n14538), .ZN(n12511) );
  OR2_X2 U10210 ( .A1(n10977), .A2(n12511), .ZN(n10975) );
  INV_X1 U10211 ( .A(n12709), .ZN(n10742) );
  NAND2_X1 U10212 ( .A1(n10742), .A2(n11037), .ZN(n12593) );
  NAND2_X1 U10213 ( .A1(n10975), .A2(n12593), .ZN(n11087) );
  NAND2_X1 U10214 ( .A1(n8139), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U10215 ( .A1(n8083), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U10216 ( .A1(n7876), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U10217 ( .A1(n7897), .A2(n7877), .ZN(n11088) );
  NAND2_X1 U10218 ( .A1(n6645), .A2(n11088), .ZN(n7879) );
  NAND2_X1 U10219 ( .A1(n12467), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7878) );
  NAND4_X1 U10220 ( .A1(n7881), .A2(n7880), .A3(n7879), .A4(n7878), .ZN(n11235) );
  INV_X1 U10221 ( .A(n9491), .ZN(n7971) );
  OAI21_X1 U10222 ( .B1(n7883), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7885) );
  MUX2_X1 U10223 ( .A(n7885), .B(P3_IR_REG_31__SCAN_IN), .S(n7884), .Z(n7887)
         );
  NAND2_X1 U10224 ( .A1(n7887), .A2(n7886), .ZN(n15051) );
  AOI22_X1 U10225 ( .A1(n7972), .A2(n9083), .B1(n7971), .B2(n15051), .ZN(n7891) );
  XNOR2_X1 U10226 ( .A(n7889), .B(n7888), .ZN(n9082) );
  NAND2_X1 U10227 ( .A1(n9082), .A2(n12480), .ZN(n7890) );
  NAND2_X1 U10228 ( .A1(n11230), .A2(n11136), .ZN(n12596) );
  NAND2_X1 U10229 ( .A1(n11235), .A2(n14535), .ZN(n12597) );
  XNOR2_X1 U10230 ( .A(n7892), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U10231 ( .A1(n9236), .A2(n12480), .ZN(n7896) );
  NAND2_X1 U10232 ( .A1(n7886), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7893) );
  MUX2_X1 U10233 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7893), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n7894) );
  NAND2_X1 U10234 ( .A1(n7894), .A2(n7588), .ZN(n15071) );
  AOI22_X1 U10235 ( .A1(n7972), .A2(n9237), .B1(n7971), .B2(n15071), .ZN(n7895) );
  NAND2_X1 U10236 ( .A1(n8083), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10237 ( .A1(n8139), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U10238 ( .A1(n7897), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7898) );
  NAND2_X1 U10239 ( .A1(n7909), .A2(n7898), .ZN(n11239) );
  NAND2_X1 U10240 ( .A1(n6645), .A2(n11239), .ZN(n7900) );
  NAND2_X1 U10241 ( .A1(n8138), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7899) );
  NAND4_X1 U10242 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n12992) );
  OR2_X1 U10243 ( .A1(n13130), .A2(n12992), .ZN(n12603) );
  NAND2_X1 U10244 ( .A1(n13130), .A2(n12992), .ZN(n12602) );
  NAND2_X1 U10245 ( .A1(n7903), .A2(n12602), .ZN(n12986) );
  XNOR2_X1 U10246 ( .A(n7905), .B(n7904), .ZN(n9340) );
  NAND2_X1 U10247 ( .A1(n9340), .A2(n12480), .ZN(n7908) );
  NAND2_X1 U10248 ( .A1(n7588), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7906) );
  XNOR2_X1 U10249 ( .A(n7906), .B(P3_IR_REG_14__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U10250 ( .A1(n7972), .A2(SI_14_), .B1(n7971), .B2(n12751), .ZN(
        n7907) );
  NAND2_X1 U10251 ( .A1(n7908), .A2(n7907), .ZN(n13066) );
  NAND2_X1 U10252 ( .A1(n8083), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U10253 ( .A1(n8139), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10254 ( .A1(n7909), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7910) );
  NAND2_X1 U10255 ( .A1(n7975), .A2(n7910), .ZN(n12996) );
  NAND2_X1 U10256 ( .A1(n6645), .A2(n12996), .ZN(n7912) );
  NAND2_X1 U10257 ( .A1(n8138), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7911) );
  OR2_X1 U10258 ( .A1(n13066), .A2(n11297), .ZN(n12606) );
  NAND2_X1 U10259 ( .A1(n13066), .A2(n11297), .ZN(n12910) );
  NAND2_X1 U10260 ( .A1(n12606), .A2(n12910), .ZN(n12988) );
  OR2_X2 U10261 ( .A1(n12986), .A2(n12988), .ZN(n12911) );
  XNOR2_X1 U10262 ( .A(n7916), .B(n7915), .ZN(n9817) );
  NAND2_X1 U10263 ( .A1(n9817), .A2(n12480), .ZN(n7918) );
  INV_X1 U10264 ( .A(SI_19_), .ZN(n9816) );
  AOI22_X1 U10265 ( .A1(n7972), .A2(n9816), .B1(n7971), .B2(n12769), .ZN(n7917) );
  NAND2_X1 U10266 ( .A1(n8139), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U10267 ( .A1(n8083), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U10268 ( .A1(n7933), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10269 ( .A1(n7998), .A2(n7920), .ZN(n12922) );
  NAND2_X1 U10270 ( .A1(n6645), .A2(n12922), .ZN(n7922) );
  NAND2_X1 U10271 ( .A1(n8138), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n7921) );
  NAND4_X1 U10272 ( .A1(n7924), .A2(n7923), .A3(n7922), .A4(n7921), .ZN(n12899) );
  NAND2_X1 U10273 ( .A1(n13112), .A2(n12899), .ZN(n12634) );
  INV_X1 U10274 ( .A(n12634), .ZN(n7986) );
  NAND2_X1 U10275 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  NAND2_X1 U10276 ( .A1(n7928), .A2(n7927), .ZN(n9743) );
  OR2_X1 U10277 ( .A1(n9743), .A2(n8089), .ZN(n7931) );
  NAND2_X1 U10278 ( .A1(n7942), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7929) );
  XNOR2_X1 U10279 ( .A(n7929), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14511) );
  AOI22_X1 U10280 ( .A1(n7972), .A2(SI_18_), .B1(n7971), .B2(n14511), .ZN(
        n7930) );
  NAND2_X1 U10281 ( .A1(n7931), .A2(n7930), .ZN(n11869) );
  NAND2_X1 U10282 ( .A1(n8058), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U10283 ( .A1(n8083), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10284 ( .A1(n7947), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7932) );
  NAND2_X1 U10285 ( .A1(n7933), .A2(n7932), .ZN(n12940) );
  NAND2_X1 U10286 ( .A1(n6645), .A2(n12940), .ZN(n7935) );
  NAND2_X1 U10287 ( .A1(n12467), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7934) );
  INV_X1 U10288 ( .A(n12625), .ZN(n7985) );
  NAND2_X1 U10289 ( .A1(n11869), .A2(n12918), .ZN(n12624) );
  INV_X1 U10290 ( .A(n12936), .ZN(n7952) );
  XNOR2_X1 U10291 ( .A(n9761), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n7938) );
  XNOR2_X1 U10292 ( .A(n7939), .B(n7938), .ZN(n9554) );
  NAND2_X1 U10293 ( .A1(n9554), .A2(n12480), .ZN(n7945) );
  NAND2_X1 U10294 ( .A1(n7940), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7941) );
  MUX2_X1 U10295 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7941), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n7943) );
  AOI22_X1 U10296 ( .A1(n7972), .A2(SI_17_), .B1(n7971), .B2(n14497), .ZN(
        n7944) );
  NAND2_X1 U10297 ( .A1(n7945), .A2(n7944), .ZN(n13052) );
  NAND2_X1 U10298 ( .A1(n8058), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U10299 ( .A1(n8138), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10300 ( .A1(n7960), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7946) );
  NAND2_X1 U10301 ( .A1(n7947), .A2(n7946), .ZN(n12955) );
  NAND2_X1 U10302 ( .A1(n6645), .A2(n12955), .ZN(n7949) );
  NAND2_X1 U10303 ( .A1(n8083), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U10304 ( .A1(n13052), .A2(n12930), .ZN(n12937) );
  INV_X1 U10305 ( .A(n12937), .ZN(n12622) );
  NOR2_X1 U10306 ( .A1(n7952), .A2(n12622), .ZN(n7984) );
  OR2_X1 U10307 ( .A1(n13052), .A2(n12930), .ZN(n12626) );
  NAND2_X1 U10308 ( .A1(n12626), .A2(n12937), .ZN(n12517) );
  XNOR2_X1 U10309 ( .A(n7954), .B(n7953), .ZN(n9416) );
  NAND2_X1 U10310 ( .A1(n9416), .A2(n12480), .ZN(n7958) );
  OR2_X1 U10311 ( .A1(n7955), .A2(n13137), .ZN(n7956) );
  XNOR2_X1 U10312 ( .A(n7956), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14480) );
  AOI22_X1 U10313 ( .A1(n7972), .A2(SI_16_), .B1(n7971), .B2(n14480), .ZN(
        n7957) );
  NAND2_X1 U10314 ( .A1(n7958), .A2(n7957), .ZN(n12399) );
  NAND2_X1 U10315 ( .A1(n8083), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10316 ( .A1(n8139), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U10317 ( .A1(n7977), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U10318 ( .A1(n7960), .A2(n7959), .ZN(n12969) );
  NAND2_X1 U10319 ( .A1(n6645), .A2(n12969), .ZN(n7962) );
  NAND2_X1 U10320 ( .A1(n8138), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7961) );
  NAND4_X1 U10321 ( .A1(n7964), .A2(n7963), .A3(n7962), .A4(n7961), .ZN(n12946) );
  OR2_X1 U10322 ( .A1(n12399), .A2(n12405), .ZN(n12618) );
  INV_X1 U10323 ( .A(n12618), .ZN(n7983) );
  XNOR2_X1 U10324 ( .A(n7966), .B(n7965), .ZN(n9370) );
  NAND2_X1 U10325 ( .A1(n9370), .A2(n12480), .ZN(n7974) );
  OR2_X1 U10326 ( .A1(n7967), .A2(n13137), .ZN(n7969) );
  XNOR2_X1 U10327 ( .A(n7969), .B(n7968), .ZN(n14470) );
  INV_X1 U10328 ( .A(n14470), .ZN(n7970) );
  AOI22_X1 U10329 ( .A1(n7972), .A2(SI_15_), .B1(n7971), .B2(n7970), .ZN(n7973) );
  NAND2_X1 U10330 ( .A1(n7974), .A2(n7973), .ZN(n11311) );
  NAND2_X1 U10331 ( .A1(n8083), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7981) );
  NAND2_X1 U10332 ( .A1(n8058), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U10333 ( .A1(n7975), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U10334 ( .A1(n7977), .A2(n7976), .ZN(n12980) );
  NAND2_X1 U10335 ( .A1(n6645), .A2(n12980), .ZN(n7979) );
  NAND2_X1 U10336 ( .A1(n12467), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7978) );
  NAND4_X1 U10337 ( .A1(n7981), .A2(n7980), .A3(n7979), .A4(n7978), .ZN(n12991) );
  INV_X1 U10338 ( .A(n12991), .ZN(n11858) );
  NAND2_X1 U10339 ( .A1(n11311), .A2(n11858), .ZN(n12964) );
  NAND2_X1 U10340 ( .A1(n12399), .A2(n12405), .ZN(n12615) );
  AND2_X1 U10341 ( .A1(n12964), .A2(n12615), .ZN(n7982) );
  OR2_X1 U10342 ( .A1(n7983), .A2(n7982), .ZN(n12950) );
  OR2_X1 U10343 ( .A1(n12517), .A2(n12950), .ZN(n12934) );
  AND2_X1 U10344 ( .A1(n7984), .A2(n12934), .ZN(n12933) );
  OR2_X1 U10345 ( .A1(n7985), .A2(n12933), .ZN(n12913) );
  AND2_X1 U10346 ( .A1(n12910), .A2(n7988), .ZN(n7987) );
  NAND2_X1 U10347 ( .A1(n12911), .A2(n7987), .ZN(n7992) );
  INV_X1 U10348 ( .A(n7988), .ZN(n7990) );
  OR2_X1 U10349 ( .A1(n11311), .A2(n11858), .ZN(n12608) );
  AND2_X1 U10350 ( .A1(n12978), .A2(n12618), .ZN(n12949) );
  AND2_X1 U10351 ( .A1(n12949), .A2(n12953), .ZN(n12932) );
  AND2_X1 U10352 ( .A1(n12932), .A2(n12625), .ZN(n12912) );
  AND2_X1 U10353 ( .A1(n12912), .A2(n12634), .ZN(n7989) );
  OR2_X1 U10354 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  NAND2_X1 U10355 ( .A1(n7992), .A2(n7991), .ZN(n7993) );
  OR2_X1 U10356 ( .A1(n13112), .A2(n12899), .ZN(n12633) );
  NAND2_X1 U10357 ( .A1(n7993), .A2(n12633), .ZN(n12907) );
  XNOR2_X1 U10358 ( .A(n7995), .B(n7994), .ZN(n10046) );
  NAND2_X1 U10359 ( .A1(n10046), .A2(n12480), .ZN(n7997) );
  INV_X1 U10360 ( .A(SI_20_), .ZN(n10047) );
  NAND2_X1 U10361 ( .A1(n8058), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U10362 ( .A1(n8083), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U10363 ( .A1(n7998), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U10364 ( .A1(n8011), .A2(n7999), .ZN(n12901) );
  NAND2_X1 U10365 ( .A1(n6645), .A2(n12901), .ZN(n8001) );
  NAND2_X1 U10366 ( .A1(n8138), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8000) );
  OR2_X1 U10367 ( .A1(n12905), .A2(n12921), .ZN(n12638) );
  NAND2_X1 U10368 ( .A1(n12905), .A2(n12921), .ZN(n12637) );
  NAND2_X1 U10369 ( .A1(n12638), .A2(n12637), .ZN(n12906) );
  NAND2_X1 U10370 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  AND2_X1 U10371 ( .A1(n8008), .A2(n8007), .ZN(n10140) );
  NAND2_X1 U10372 ( .A1(n10140), .A2(n12480), .ZN(n8010) );
  INV_X1 U10373 ( .A(SI_21_), .ZN(n10141) );
  OR2_X1 U10374 ( .A1(n7882), .A2(n10141), .ZN(n8009) );
  NAND2_X1 U10375 ( .A1(n8010), .A2(n8009), .ZN(n11877) );
  NAND2_X1 U10376 ( .A1(n8139), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U10377 ( .A1(n12467), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U10378 ( .A1(n8011), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10379 ( .A1(n8024), .A2(n8012), .ZN(n12892) );
  NAND2_X1 U10380 ( .A1(n6645), .A2(n12892), .ZN(n8014) );
  NAND2_X1 U10381 ( .A1(n8083), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8013) );
  NAND4_X1 U10382 ( .A1(n8016), .A2(n8015), .A3(n8014), .A4(n8013), .ZN(n12898) );
  INV_X1 U10383 ( .A(n12898), .ZN(n11878) );
  NAND2_X1 U10384 ( .A1(n11877), .A2(n11878), .ZN(n12642) );
  NAND2_X1 U10385 ( .A1(n13104), .A2(n12898), .ZN(n12643) );
  NAND2_X1 U10386 ( .A1(n8017), .A2(n12643), .ZN(n12880) );
  OAI21_X1 U10387 ( .B1(n8020), .B2(n8019), .A(n8018), .ZN(n10243) );
  OR2_X1 U10388 ( .A1(n10243), .A2(n8089), .ZN(n8023) );
  INV_X1 U10389 ( .A(SI_22_), .ZN(n8021) );
  NAND2_X1 U10390 ( .A1(n8058), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10391 ( .A1(n8138), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10392 ( .A1(n8024), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8025) );
  NAND2_X1 U10393 ( .A1(n8037), .A2(n8025), .ZN(n12882) );
  NAND2_X1 U10394 ( .A1(n6645), .A2(n12882), .ZN(n8027) );
  NAND2_X1 U10395 ( .A1(n8083), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8026) );
  NAND4_X1 U10396 ( .A1(n8029), .A2(n8028), .A3(n8027), .A4(n8026), .ZN(n12705) );
  INV_X1 U10397 ( .A(n12705), .ZN(n11885) );
  NAND2_X1 U10398 ( .A1(n11880), .A2(n11885), .ZN(n12646) );
  NAND2_X1 U10399 ( .A1(n12880), .A2(n12646), .ZN(n8030) );
  NAND2_X1 U10400 ( .A1(n13100), .A2(n12705), .ZN(n12647) );
  NAND2_X1 U10401 ( .A1(n8030), .A2(n12647), .ZN(n12864) );
  XNOR2_X1 U10402 ( .A(n8032), .B(n8031), .ZN(n10473) );
  NAND2_X1 U10403 ( .A1(n10473), .A2(n12480), .ZN(n8034) );
  OR2_X1 U10404 ( .A1(n7882), .A2(n10475), .ZN(n8033) );
  NAND2_X1 U10405 ( .A1(n8139), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10406 ( .A1(n8138), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8035) );
  AND2_X1 U10407 ( .A1(n8036), .A2(n8035), .ZN(n8041) );
  NAND2_X1 U10408 ( .A1(n8037), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10409 ( .A1(n8045), .A2(n8038), .ZN(n12871) );
  NAND2_X1 U10410 ( .A1(n12871), .A2(n6645), .ZN(n8040) );
  NAND2_X1 U10411 ( .A1(n8083), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8039) );
  XNOR2_X1 U10412 ( .A(n12651), .B(n12650), .ZN(n8128) );
  OR2_X1 U10413 ( .A1(n12651), .A2(n12650), .ZN(n12530) );
  XNOR2_X1 U10414 ( .A(n8042), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n10895) );
  NAND2_X1 U10415 ( .A1(n10895), .A2(n12480), .ZN(n8044) );
  INV_X1 U10416 ( .A(SI_24_), .ZN(n10897) );
  INV_X1 U10417 ( .A(n12467), .ZN(n8095) );
  INV_X1 U10418 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10419 ( .A1(n8045), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10420 ( .A1(n8056), .A2(n8046), .ZN(n12856) );
  NAND2_X1 U10421 ( .A1(n12856), .A2(n6645), .ZN(n8048) );
  AOI22_X1 U10422 ( .A1(n8083), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n8058), .B2(
        P3_REG1_REG_24__SCAN_IN), .ZN(n8047) );
  OAI211_X1 U10423 ( .C1(n8095), .C2(n8049), .A(n8048), .B(n8047), .ZN(n12703)
         );
  OR2_X1 U10424 ( .A1(n13021), .A2(n12412), .ZN(n12531) );
  NAND2_X1 U10425 ( .A1(n13021), .A2(n12412), .ZN(n12532) );
  OR2_X1 U10426 ( .A1(n8051), .A2(n8050), .ZN(n8052) );
  AND2_X1 U10427 ( .A1(n8053), .A2(n8052), .ZN(n11040) );
  NAND2_X1 U10428 ( .A1(n11040), .A2(n12480), .ZN(n8055) );
  INV_X1 U10429 ( .A(SI_25_), .ZN(n11041) );
  OR2_X1 U10430 ( .A1(n7882), .A2(n11041), .ZN(n8054) );
  NAND2_X1 U10431 ( .A1(n8056), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10432 ( .A1(n8070), .A2(n8057), .ZN(n12844) );
  NAND2_X1 U10433 ( .A1(n12844), .A2(n6645), .ZN(n8061) );
  AOI22_X1 U10434 ( .A1(n8083), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n8058), .B2(
        P3_REG1_REG_25__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10435 ( .A1(n12467), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8059) );
  XNOR2_X1 U10436 ( .A(n12845), .B(n12656), .ZN(n12840) );
  INV_X1 U10437 ( .A(n12840), .ZN(n8062) );
  NAND2_X1 U10438 ( .A1(n12838), .A2(n8062), .ZN(n8063) );
  NAND2_X1 U10439 ( .A1(n12845), .A2(n12656), .ZN(n12655) );
  OR2_X1 U10440 ( .A1(n8065), .A2(n8064), .ZN(n8067) );
  AND2_X1 U10441 ( .A1(n8067), .A2(n8066), .ZN(n11058) );
  NAND2_X1 U10442 ( .A1(n11058), .A2(n12480), .ZN(n8069) );
  NAND2_X1 U10443 ( .A1(n8070), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10444 ( .A1(n8081), .A2(n8071), .ZN(n12833) );
  NAND2_X1 U10445 ( .A1(n12833), .A2(n6645), .ZN(n8076) );
  INV_X1 U10446 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13085) );
  NAND2_X1 U10447 ( .A1(n8058), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10448 ( .A1(n8083), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8072) );
  OAI211_X1 U10449 ( .C1(n13085), .C2(n8095), .A(n8073), .B(n8072), .ZN(n8074)
         );
  INV_X1 U10450 ( .A(n8074), .ZN(n8075) );
  NAND2_X1 U10451 ( .A1(n13087), .A2(n12702), .ZN(n12664) );
  XNOR2_X1 U10452 ( .A(n8078), .B(n8077), .ZN(n11111) );
  NAND2_X1 U10453 ( .A1(n11111), .A2(n12480), .ZN(n8080) );
  INV_X1 U10454 ( .A(SI_27_), .ZN(n11112) );
  OR2_X1 U10455 ( .A1(n7882), .A2(n11112), .ZN(n8079) );
  NAND2_X1 U10456 ( .A1(n8081), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8082) );
  NAND2_X1 U10457 ( .A1(n8091), .A2(n8082), .ZN(n12823) );
  INV_X1 U10458 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13082) );
  NAND2_X1 U10459 ( .A1(n8139), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8085) );
  NAND2_X1 U10460 ( .A1(n8083), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8084) );
  OAI211_X1 U10461 ( .C1(n13082), .C2(n8095), .A(n8085), .B(n8084), .ZN(n8086)
         );
  AOI22_X1 U10462 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13689), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n12265), .ZN(n8087) );
  NAND2_X1 U10463 ( .A1(n8091), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10464 ( .A1(n12337), .A2(n8092), .ZN(n12807) );
  INV_X1 U10465 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n15375) );
  NAND2_X1 U10466 ( .A1(n8139), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10467 ( .A1(n8083), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8093) );
  OAI211_X1 U10468 ( .C1(n8095), .C2(n15375), .A(n8094), .B(n8093), .ZN(n8096)
         );
  NAND2_X1 U10469 ( .A1(n8136), .A2(n12354), .ZN(n8133) );
  NAND2_X1 U10470 ( .A1(n8133), .A2(n12797), .ZN(n12529) );
  OR2_X1 U10471 ( .A1(n8136), .A2(n12354), .ZN(n12528) );
  NAND2_X1 U10472 ( .A1(n12716), .A2(n10252), .ZN(n8103) );
  OR2_X1 U10473 ( .A1(n12557), .A2(n10478), .ZN(n10480) );
  NAND2_X1 U10474 ( .A1(n10405), .A2(n8098), .ZN(n10402) );
  NAND2_X1 U10475 ( .A1(n15125), .A2(n8099), .ZN(n15126) );
  NAND2_X1 U10476 ( .A1(n15112), .A2(n15124), .ZN(n15113) );
  NAND2_X1 U10477 ( .A1(n15127), .A2(n15113), .ZN(n8100) );
  NAND2_X1 U10478 ( .A1(n15135), .A2(n15106), .ZN(n10502) );
  INV_X1 U10479 ( .A(n12507), .ZN(n8101) );
  AND2_X1 U10480 ( .A1(n10502), .A2(n8101), .ZN(n8102) );
  NAND2_X1 U10481 ( .A1(n12717), .A2(n15155), .ZN(n10245) );
  AND2_X1 U10482 ( .A1(n10245), .A2(n8103), .ZN(n10477) );
  INV_X1 U10483 ( .A(n12557), .ZN(n10483) );
  AND2_X1 U10484 ( .A1(n10477), .A2(n10483), .ZN(n8104) );
  NAND3_X1 U10485 ( .A1(n10403), .A2(n10481), .A3(n7009), .ZN(n10407) );
  NAND2_X1 U10486 ( .A1(n12714), .A2(n10410), .ZN(n8105) );
  NAND2_X1 U10487 ( .A1(n10407), .A2(n8105), .ZN(n10719) );
  AND2_X1 U10488 ( .A1(n12713), .A2(n12534), .ZN(n8106) );
  NAND2_X1 U10489 ( .A1(n12711), .A2(n15194), .ZN(n10917) );
  AND2_X1 U10490 ( .A1(n10788), .A2(n8110), .ZN(n8107) );
  NAND2_X1 U10491 ( .A1(n12710), .A2(n10926), .ZN(n8109) );
  AND2_X1 U10492 ( .A1(n8107), .A2(n8109), .ZN(n10980) );
  AND2_X1 U10493 ( .A1(n12709), .A2(n11037), .ZN(n8113) );
  INV_X1 U10494 ( .A(n8113), .ZN(n8108) );
  AND2_X1 U10495 ( .A1(n10980), .A2(n8108), .ZN(n8114) );
  INV_X1 U10496 ( .A(n8109), .ZN(n8112) );
  XNOR2_X1 U10497 ( .A(n12711), .B(n15194), .ZN(n12579) );
  NAND2_X1 U10498 ( .A1(n10611), .A2(n15183), .ZN(n10868) );
  OR2_X1 U10499 ( .A1(n8112), .A2(n8111), .ZN(n10982) );
  AOI21_X1 U10500 ( .B1(n10981), .B2(n8114), .A(n7575), .ZN(n8116) );
  NAND2_X1 U10501 ( .A1(n10742), .A2(n14538), .ZN(n8115) );
  NOR2_X1 U10502 ( .A1(n11235), .A2(n11136), .ZN(n8117) );
  INV_X1 U10503 ( .A(n12992), .ZN(n11303) );
  OR2_X1 U10504 ( .A1(n11311), .A2(n12991), .ZN(n8118) );
  AND2_X1 U10505 ( .A1(n12988), .A2(n8118), .ZN(n8121) );
  INV_X1 U10506 ( .A(n8118), .ZN(n8120) );
  INV_X1 U10507 ( .A(n11297), .ZN(n12708) );
  NAND2_X1 U10508 ( .A1(n13066), .A2(n12708), .ZN(n12973) );
  AND2_X1 U10509 ( .A1(n7571), .A2(n12973), .ZN(n8119) );
  INV_X1 U10510 ( .A(n12399), .ZN(n13121) );
  NAND2_X1 U10511 ( .A1(n12945), .A2(n12517), .ZN(n8123) );
  NAND2_X1 U10512 ( .A1(n13052), .A2(n12707), .ZN(n8122) );
  NAND2_X1 U10513 ( .A1(n8123), .A2(n8122), .ZN(n12928) );
  NAND2_X1 U10514 ( .A1(n12633), .A2(n12634), .ZN(n12917) );
  INV_X1 U10515 ( .A(n12899), .ZN(n12931) );
  OR2_X1 U10516 ( .A1(n13112), .A2(n12931), .ZN(n8124) );
  NAND2_X1 U10517 ( .A1(n12897), .A2(n12906), .ZN(n8126) );
  NAND2_X1 U10518 ( .A1(n12905), .A2(n12706), .ZN(n8125) );
  NAND2_X1 U10519 ( .A1(n8126), .A2(n8125), .ZN(n12887) );
  AND2_X1 U10520 ( .A1(n11877), .A2(n12898), .ZN(n12498) );
  INV_X1 U10521 ( .A(n12498), .ZN(n8127) );
  NAND2_X1 U10522 ( .A1(n13104), .A2(n11878), .ZN(n12499) );
  AOI22_X1 U10523 ( .A1(n12862), .A2(n8128), .B1(n12704), .B2(n12651), .ZN(
        n12851) );
  NAND2_X1 U10524 ( .A1(n13021), .A2(n12703), .ZN(n8129) );
  INV_X1 U10525 ( .A(n13021), .ZN(n12858) );
  AOI22_X1 U10526 ( .A1(n12851), .A2(n8129), .B1(n12858), .B2(n12412), .ZN(
        n12841) );
  NAND2_X1 U10527 ( .A1(n12841), .A2(n12840), .ZN(n12839) );
  OAI21_X1 U10528 ( .B1(n12656), .B2(n13091), .A(n12839), .ZN(n12828) );
  NAND2_X1 U10529 ( .A1(n13087), .A2(n12353), .ZN(n8130) );
  AOI22_X1 U10530 ( .A1(n12828), .A2(n8130), .B1(n12702), .B2(n12457), .ZN(
        n12817) );
  NAND2_X1 U10531 ( .A1(n12817), .A2(n12816), .ZN(n12815) );
  INV_X1 U10532 ( .A(n12802), .ZN(n12701) );
  NAND2_X1 U10533 ( .A1(n12815), .A2(n8132), .ZN(n12801) );
  INV_X1 U10534 ( .A(n12801), .ZN(n8135) );
  INV_X1 U10535 ( .A(n12800), .ZN(n8134) );
  XNOR2_X1 U10536 ( .A(n8137), .B(n12521), .ZN(n8147) );
  NAND2_X1 U10537 ( .A1(n12525), .A2(n12694), .ZN(n8171) );
  NAND2_X1 U10538 ( .A1(n12535), .A2(n8191), .ZN(n12492) );
  INV_X1 U10539 ( .A(n11319), .ZN(n9495) );
  NAND2_X1 U10540 ( .A1(n9495), .A2(n12693), .ZN(n9499) );
  NAND2_X1 U10541 ( .A1(n9491), .A2(n9499), .ZN(n10802) );
  INV_X1 U10542 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n15492) );
  NAND2_X1 U10543 ( .A1(n8138), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10544 ( .A1(n8139), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8140) );
  OAI211_X1 U10545 ( .C1(n8142), .C2(n15492), .A(n8141), .B(n8140), .ZN(n8143)
         );
  INV_X1 U10546 ( .A(n8143), .ZN(n8144) );
  AND2_X1 U10547 ( .A1(n9495), .A2(P3_B_REG_SCAN_IN), .ZN(n8145) );
  OR2_X1 U10548 ( .A1(n15136), .A2(n8145), .ZN(n12793) );
  OAI22_X1 U10549 ( .A1(n12354), .A2(n15134), .B1(n12487), .B2(n12793), .ZN(
        n8146) );
  AOI21_X2 U10550 ( .B1(n8147), .B2(n12987), .A(n8146), .ZN(n12343) );
  OAI21_X1 U10551 ( .B1(n15172), .B2(n12336), .A(n12343), .ZN(n8197) );
  NAND2_X1 U10552 ( .A1(n6717), .A2(n8153), .ZN(n8148) );
  NAND2_X1 U10553 ( .A1(n6684), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8150) );
  MUX2_X1 U10554 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8150), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8151) );
  XNOR2_X1 U10555 ( .A(n10898), .B(P3_B_REG_SCAN_IN), .ZN(n8155) );
  INV_X1 U10556 ( .A(n8180), .ZN(n11061) );
  NAND2_X1 U10557 ( .A1(n11061), .A2(n10898), .ZN(n8156) );
  NAND2_X1 U10558 ( .A1(n11061), .A2(n11043), .ZN(n8157) );
  NAND2_X1 U10559 ( .A1(n13134), .A2(n13132), .ZN(n8189) );
  INV_X1 U10560 ( .A(n8189), .ZN(n8170) );
  NOR2_X1 U10561 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .ZN(
        n8162) );
  NOR4_X1 U10562 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_D_REG_4__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8161) );
  NOR4_X1 U10563 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8160) );
  NOR4_X1 U10564 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8159) );
  NAND4_X1 U10565 ( .A1(n8162), .A2(n8161), .A3(n8160), .A4(n8159), .ZN(n8168)
         );
  NOR4_X1 U10566 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_26__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n8166) );
  NOR4_X1 U10567 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n8165) );
  NOR4_X1 U10568 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .A3(
        P3_D_REG_6__SCAN_IN), .A4(P3_D_REG_3__SCAN_IN), .ZN(n8164) );
  NOR4_X1 U10569 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_13__SCAN_IN), .ZN(n8163) );
  NAND4_X1 U10570 ( .A1(n8166), .A2(n8165), .A3(n8164), .A4(n8163), .ZN(n8167)
         );
  NOR2_X1 U10571 ( .A1(n8168), .A2(n8167), .ZN(n8169) );
  NAND2_X1 U10572 ( .A1(n8170), .A2(n8187), .ZN(n8945) );
  OR2_X1 U10573 ( .A1(n12676), .A2(n12692), .ZN(n9784) );
  NAND2_X1 U10574 ( .A1(n10250), .A2(n8191), .ZN(n12686) );
  OR2_X1 U10575 ( .A1(n8171), .A2(n12686), .ZN(n8932) );
  AND2_X1 U10576 ( .A1(n9784), .A2(n8932), .ZN(n8176) );
  INV_X1 U10577 ( .A(n8187), .ZN(n8172) );
  NOR2_X1 U10578 ( .A1(n13132), .A2(n8172), .ZN(n8174) );
  INV_X1 U10579 ( .A(n13134), .ZN(n8173) );
  NAND2_X1 U10580 ( .A1(n8174), .A2(n8173), .ZN(n8950) );
  INV_X1 U10581 ( .A(n8937), .ZN(n8175) );
  OAI22_X1 U10582 ( .A1(n8945), .A2(n8176), .B1(n8950), .B2(n8175), .ZN(n8184)
         );
  INV_X1 U10583 ( .A(n11043), .ZN(n8178) );
  INV_X1 U10584 ( .A(n10898), .ZN(n8177) );
  NAND2_X1 U10585 ( .A1(n6812), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8181) );
  MUX2_X1 U10586 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8181), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8182) );
  INV_X1 U10587 ( .A(n13133), .ZN(n8183) );
  MUX2_X1 U10588 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n8197), .S(n15197), .Z(
        n8185) );
  INV_X1 U10589 ( .A(n8185), .ZN(n8186) );
  NAND2_X1 U10590 ( .A1(n8186), .A2(n7561), .ZN(P3_U3456) );
  NAND2_X1 U10591 ( .A1(n12692), .A2(n12672), .ZN(n8933) );
  AND3_X1 U10592 ( .A1(n12690), .A2(n8187), .A3(n8933), .ZN(n8188) );
  OAI22_X1 U10593 ( .A1(n12525), .A2(n8192), .B1(n8191), .B2(n15182), .ZN(
        n8193) );
  AOI21_X1 U10594 ( .B1(n8193), .B2(n12692), .A(n12672), .ZN(n8194) );
  NAND2_X1 U10595 ( .A1(n13134), .A2(n8194), .ZN(n8195) );
  MUX2_X1 U10596 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n8197), .S(n15213), .Z(
        n8198) );
  INV_X1 U10597 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U10598 ( .A1(n8199), .A2(n7569), .ZN(P3_U3488) );
  AND3_X2 U10599 ( .A1(n8202), .A2(n8201), .A3(n8200), .ZN(n8422) );
  NOR2_X1 U10600 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .ZN(n8204) );
  NOR2_X2 U10601 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8500) );
  NOR2_X1 U10602 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .ZN(n8206) );
  NOR2_X1 U10603 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8205) );
  AND3_X4 U10604 ( .A1(n8422), .A2(n8208), .A3(n8207), .ZN(n8580) );
  XNOR2_X2 U10605 ( .A(n8216), .B(n8215), .ZN(n8220) );
  XNOR2_X2 U10606 ( .A(n8219), .B(n8218), .ZN(n8221) );
  NAND2_X1 U10607 ( .A1(n12178), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8234) );
  INV_X1 U10608 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14034) );
  OR2_X1 U10609 ( .A1(n6651), .A2(n14034), .ZN(n8233) );
  INV_X1 U10610 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n15519) );
  NAND2_X1 U10611 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8413) );
  NOR2_X1 U10612 ( .A1(n8413), .A2(n9156), .ZN(n8429) );
  NAND2_X1 U10613 ( .A1(n8429), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8444) );
  AND2_X1 U10614 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n8223) );
  NAND2_X1 U10615 ( .A1(n8506), .A2(n8223), .ZN(n8521) );
  NAND2_X1 U10616 ( .A1(n8568), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8590) );
  INV_X1 U10617 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U10618 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n8224) );
  NAND2_X1 U10619 ( .A1(n8629), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U10620 ( .A1(n8671), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U10621 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n8705), .ZN(n8704) );
  INV_X1 U10622 ( .A(n8704), .ZN(n8225) );
  NAND2_X1 U10623 ( .A1(n8225), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8722) );
  INV_X1 U10624 ( .A(n8722), .ZN(n8226) );
  NAND2_X1 U10625 ( .A1(n8226), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8724) );
  INV_X1 U10626 ( .A(n8724), .ZN(n8227) );
  NAND2_X1 U10627 ( .A1(n8227), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8741) );
  INV_X1 U10628 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10629 ( .A1(n8724), .A2(n8228), .ZN(n8229) );
  NAND2_X1 U10630 ( .A1(n8741), .A2(n8229), .ZN(n14033) );
  OR2_X1 U10631 ( .A1(n6647), .A2(n14033), .ZN(n8232) );
  INV_X1 U10632 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14207) );
  OR2_X1 U10633 ( .A1(n12179), .A2(n14207), .ZN(n8231) );
  NAND2_X1 U10634 ( .A1(n8236), .A2(SI_1_), .ZN(n8239) );
  NAND2_X1 U10635 ( .A1(n8240), .A2(SI_2_), .ZN(n8242) );
  OAI21_X1 U10636 ( .B1(n8240), .B2(SI_2_), .A(n8242), .ZN(n8365) );
  INV_X1 U10637 ( .A(n8365), .ZN(n8241) );
  NAND2_X1 U10638 ( .A1(n8364), .A2(n8241), .ZN(n8367) );
  NAND2_X1 U10639 ( .A1(n8367), .A2(n8242), .ZN(n8378) );
  MUX2_X1 U10640 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n9468), .Z(n8243) );
  NAND2_X1 U10641 ( .A1(n8243), .A2(SI_3_), .ZN(n8245) );
  OAI21_X1 U10642 ( .B1(n8243), .B2(SI_3_), .A(n8245), .ZN(n8244) );
  INV_X1 U10643 ( .A(n8244), .ZN(n8377) );
  NAND2_X1 U10644 ( .A1(n8378), .A2(n8377), .ZN(n8379) );
  NAND2_X1 U10645 ( .A1(n8379), .A2(n8245), .ZN(n8392) );
  MUX2_X1 U10646 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n9468), .Z(n8246) );
  NAND2_X1 U10647 ( .A1(n8246), .A2(SI_4_), .ZN(n8248) );
  OAI21_X1 U10648 ( .B1(n8246), .B2(SI_4_), .A(n8248), .ZN(n8247) );
  INV_X1 U10649 ( .A(n8247), .ZN(n8391) );
  MUX2_X1 U10650 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9468), .Z(n8249) );
  OAI21_X1 U10651 ( .B1(n8249), .B2(SI_5_), .A(n8251), .ZN(n8250) );
  INV_X1 U10652 ( .A(n8250), .ZN(n8405) );
  MUX2_X1 U10653 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6643), .Z(n8252) );
  NAND2_X1 U10654 ( .A1(n8252), .A2(SI_6_), .ZN(n8436) );
  OAI21_X1 U10655 ( .B1(SI_6_), .B2(n8252), .A(n8436), .ZN(n8253) );
  INV_X1 U10656 ( .A(n8253), .ZN(n8419) );
  MUX2_X1 U10657 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6643), .Z(n8255) );
  NAND2_X1 U10658 ( .A1(n8255), .A2(SI_7_), .ZN(n8254) );
  INV_X1 U10659 ( .A(n8254), .ZN(n8257) );
  OAI21_X1 U10660 ( .B1(n8255), .B2(SI_7_), .A(n8254), .ZN(n8438) );
  INV_X1 U10661 ( .A(n8438), .ZN(n8256) );
  MUX2_X1 U10662 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9468), .Z(n8258) );
  NAND2_X1 U10663 ( .A1(n8258), .A2(SI_8_), .ZN(n8261) );
  OAI21_X1 U10664 ( .B1(SI_8_), .B2(n8258), .A(n8261), .ZN(n8453) );
  INV_X1 U10665 ( .A(n8453), .ZN(n8259) );
  AND2_X1 U10666 ( .A1(n8451), .A2(n8259), .ZN(n8260) );
  NAND2_X1 U10667 ( .A1(n8452), .A2(n8260), .ZN(n8262) );
  MUX2_X1 U10668 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9468), .Z(n8263) );
  NAND2_X1 U10669 ( .A1(n8263), .A2(SI_9_), .ZN(n8265) );
  OAI21_X1 U10670 ( .B1(n8263), .B2(SI_9_), .A(n8265), .ZN(n8264) );
  INV_X1 U10671 ( .A(n8264), .ZN(n8466) );
  MUX2_X1 U10672 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9468), .Z(n8266) );
  NAND2_X1 U10673 ( .A1(n8266), .A2(SI_10_), .ZN(n8268) );
  OAI21_X1 U10674 ( .B1(SI_10_), .B2(n8266), .A(n8268), .ZN(n8487) );
  INV_X1 U10675 ( .A(n8487), .ZN(n8267) );
  MUX2_X1 U10676 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9468), .Z(n8269) );
  XNOR2_X1 U10677 ( .A(n8269), .B(SI_11_), .ZN(n8498) );
  INV_X1 U10678 ( .A(n8269), .ZN(n8270) );
  NAND2_X1 U10679 ( .A1(n8270), .A2(n15521), .ZN(n8271) );
  MUX2_X1 U10680 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n9468), .Z(n8272) );
  XNOR2_X1 U10681 ( .A(n8272), .B(n9083), .ZN(n8516) );
  INV_X1 U10682 ( .A(n8272), .ZN(n8273) );
  MUX2_X1 U10683 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n9468), .Z(n8274) );
  XNOR2_X1 U10684 ( .A(n8274), .B(n9237), .ZN(n8528) );
  INV_X1 U10685 ( .A(n8274), .ZN(n8275) );
  NAND2_X1 U10686 ( .A1(n8275), .A2(n9237), .ZN(n8276) );
  MUX2_X1 U10687 ( .A(n9721), .B(n9725), .S(n9468), .Z(n8561) );
  MUX2_X1 U10688 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n9468), .Z(n8563) );
  NAND2_X1 U10689 ( .A1(n8563), .A2(SI_15_), .ZN(n8282) );
  OAI21_X1 U10690 ( .B1(n15380), .B2(n8561), .A(n8282), .ZN(n8278) );
  INV_X1 U10691 ( .A(n8278), .ZN(n8279) );
  INV_X1 U10692 ( .A(n8561), .ZN(n8280) );
  NOR2_X1 U10693 ( .A1(n8280), .A2(SI_14_), .ZN(n8283) );
  INV_X1 U10694 ( .A(n8563), .ZN(n8281) );
  AOI22_X1 U10695 ( .A1(n8283), .A2(n8282), .B1(n9372), .B2(n8281), .ZN(n8284)
         );
  MUX2_X1 U10696 ( .A(n9693), .B(n9691), .S(n9468), .Z(n8285) );
  XNOR2_X1 U10697 ( .A(n8285), .B(SI_16_), .ZN(n8577) );
  MUX2_X1 U10698 ( .A(n9762), .B(n9761), .S(n9468), .Z(n8286) );
  XNOR2_X1 U10699 ( .A(n8286), .B(SI_17_), .ZN(n8598) );
  NAND2_X1 U10700 ( .A1(n8286), .A2(n15383), .ZN(n8287) );
  MUX2_X1 U10701 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9468), .Z(n8610) );
  INV_X1 U10702 ( .A(n8610), .ZN(n8290) );
  MUX2_X1 U10703 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6643), .Z(n8291) );
  XNOR2_X1 U10704 ( .A(n8291), .B(SI_19_), .ZN(n8622) );
  INV_X1 U10705 ( .A(n8291), .ZN(n8292) );
  NAND2_X1 U10706 ( .A1(n8292), .A2(n9816), .ZN(n8635) );
  MUX2_X1 U10707 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9468), .Z(n8293) );
  NAND2_X1 U10708 ( .A1(n8293), .A2(SI_21_), .ZN(n8300) );
  OAI21_X1 U10709 ( .B1(SI_21_), .B2(n8293), .A(n8300), .ZN(n8654) );
  MUX2_X1 U10710 ( .A(n10648), .B(n12263), .S(n9468), .Z(n8639) );
  NOR2_X1 U10711 ( .A1(n8296), .A2(SI_20_), .ZN(n8294) );
  NOR2_X1 U10712 ( .A1(n8654), .A2(n8294), .ZN(n8295) );
  AND2_X1 U10713 ( .A1(n8635), .A2(n8295), .ZN(n8299) );
  INV_X1 U10714 ( .A(n8295), .ZN(n8298) );
  NAND2_X1 U10715 ( .A1(n8296), .A2(SI_20_), .ZN(n8297) );
  NAND2_X1 U10716 ( .A1(n8658), .A2(n8300), .ZN(n8302) );
  INV_X1 U10717 ( .A(n8302), .ZN(n8301) );
  MUX2_X1 U10718 ( .A(n15362), .B(n15395), .S(n9468), .Z(n10810) );
  NOR2_X1 U10719 ( .A1(n8306), .A2(n10475), .ZN(n8305) );
  NAND2_X1 U10720 ( .A1(n8306), .A2(n10475), .ZN(n8307) );
  MUX2_X1 U10721 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9468), .Z(n8308) );
  NAND2_X1 U10722 ( .A1(n8308), .A2(SI_24_), .ZN(n8309) );
  OAI21_X1 U10723 ( .B1(SI_24_), .B2(n8308), .A(n8309), .ZN(n8697) );
  XNOR2_X1 U10724 ( .A(n8310), .B(SI_25_), .ZN(n8335) );
  INV_X1 U10725 ( .A(n8310), .ZN(n8311) );
  NAND2_X1 U10726 ( .A1(n8312), .A2(n15444), .ZN(n8314) );
  MUX2_X1 U10727 ( .A(n15349), .B(n11316), .S(n6643), .Z(n8712) );
  INV_X1 U10728 ( .A(n8730), .ZN(n8733) );
  XNOR2_X1 U10729 ( .A(n8733), .B(SI_27_), .ZN(n8316) );
  INV_X1 U10730 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8317) );
  OR2_X2 U10731 ( .A1(n8321), .A2(n8317), .ZN(n8319) );
  XNOR2_X2 U10732 ( .A(n8319), .B(n8318), .ZN(n8816) );
  NAND2_X1 U10733 ( .A1(n8829), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8320) );
  INV_X1 U10734 ( .A(n8321), .ZN(n8322) );
  NAND2_X2 U10735 ( .A1(n8816), .A2(n14328), .ZN(n8324) );
  NAND2_X1 U10736 ( .A1(n13690), .A2(n12195), .ZN(n8326) );
  NAND2_X2 U10737 ( .A1(n8324), .A2(n6643), .ZN(n8533) );
  INV_X4 U10738 ( .A(n8533), .ZN(n12196) );
  NAND2_X1 U10739 ( .A1(n12196), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U10740 ( .A1(n12178), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8334) );
  INV_X1 U10741 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8327) );
  OR2_X1 U10742 ( .A1(n6651), .A2(n8327), .ZN(n8333) );
  INV_X1 U10743 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10744 ( .A1(n8704), .A2(n8328), .ZN(n8329) );
  NAND2_X1 U10745 ( .A1(n8722), .A2(n8329), .ZN(n14064) );
  OR2_X1 U10746 ( .A1(n6647), .A2(n14064), .ZN(n8332) );
  INV_X1 U10747 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8330) );
  OR2_X1 U10748 ( .A1(n12179), .A2(n8330), .ZN(n8331) );
  NAND4_X1 U10749 ( .A1(n8334), .A2(n8333), .A3(n8332), .A4(n8331), .ZN(n14080) );
  INV_X1 U10750 ( .A(n14080), .ZN(n13799) );
  INV_X1 U10751 ( .A(n8335), .ZN(n8336) );
  NAND2_X1 U10752 ( .A1(n11587), .A2(n12195), .ZN(n8338) );
  NAND2_X1 U10753 ( .A1(n12196), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8337) );
  INV_X1 U10754 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9086) );
  OR2_X1 U10755 ( .A1(n8819), .A2(n9086), .ZN(n8341) );
  INV_X1 U10756 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9999) );
  INV_X1 U10757 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U10758 ( .A1(n12178), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8339) );
  INV_X1 U10759 ( .A(n8342), .ZN(n8343) );
  NAND2_X1 U10760 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  AND2_X1 U10761 ( .A1(n8346), .A2(n8345), .ZN(n9559) );
  INV_X1 U10762 ( .A(n9559), .ZN(n9036) );
  NAND2_X1 U10763 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8347) );
  XNOR2_X1 U10764 ( .A(n8347), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U10765 ( .A1(n8381), .A2(n9130), .ZN(n8348) );
  INV_X1 U10766 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9005) );
  INV_X1 U10767 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9927) );
  INV_X1 U10768 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8349) );
  OR2_X1 U10769 ( .A1(n6651), .A2(n8349), .ZN(n8351) );
  NAND2_X1 U10770 ( .A1(n12178), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8350) );
  NOR2_X1 U10771 ( .A1(n9468), .A2(n15508), .ZN(n8355) );
  XNOR2_X1 U10772 ( .A(n8355), .B(n8354), .ZN(n14336) );
  AND2_X1 U10773 ( .A1(n13841), .A2(n9995), .ZN(n9990) );
  INV_X1 U10774 ( .A(n8356), .ZN(n14708) );
  NAND2_X1 U10775 ( .A1(n11962), .A2(n14708), .ZN(n8357) );
  NAND2_X1 U10776 ( .A1(n9991), .A2(n8357), .ZN(n9947) );
  NAND2_X1 U10777 ( .A1(n12178), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8361) );
  INV_X1 U10778 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9958) );
  INV_X1 U10779 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9129) );
  OR2_X1 U10780 ( .A1(n6650), .A2(n9129), .ZN(n8359) );
  INV_X1 U10781 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9122) );
  INV_X1 U10782 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13844) );
  INV_X1 U10783 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10784 ( .A1(n13844), .A2(n8362), .ZN(n8382) );
  NAND2_X1 U10785 ( .A1(n8382), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8363) );
  INV_X1 U10786 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8383) );
  XNOR2_X1 U10787 ( .A(n8363), .B(n8383), .ZN(n13861) );
  INV_X1 U10788 ( .A(n8364), .ZN(n8366) );
  NAND2_X1 U10789 ( .A1(n8366), .A2(n8365), .ZN(n8368) );
  NAND2_X1 U10790 ( .A1(n8368), .A2(n8367), .ZN(n9591) );
  INV_X1 U10791 ( .A(n12039), .ZN(n8371) );
  INV_X1 U10792 ( .A(n12038), .ZN(n8780) );
  INV_X1 U10793 ( .A(n13839), .ZN(n9732) );
  NAND2_X1 U10794 ( .A1(n9732), .A2(n14714), .ZN(n8372) );
  NAND2_X1 U10795 ( .A1(n12178), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8376) );
  OR2_X1 U10796 ( .A1(n6647), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8375) );
  INV_X1 U10797 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9125) );
  OR2_X1 U10798 ( .A1(n12179), .A2(n9125), .ZN(n8374) );
  INV_X1 U10799 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9966) );
  OR2_X1 U10800 ( .A1(n6650), .A2(n9966), .ZN(n8373) );
  NAND4_X1 U10801 ( .A1(n8376), .A2(n8375), .A3(n8374), .A4(n8373), .ZN(n13838) );
  OR2_X1 U10802 ( .A1(n8378), .A2(n8377), .ZN(n8380) );
  AND2_X1 U10803 ( .A1(n8380), .A2(n8379), .ZN(n9600) );
  NAND2_X1 U10804 ( .A1(n9600), .A2(n12195), .ZN(n8389) );
  INV_X1 U10805 ( .A(n8382), .ZN(n8384) );
  NAND2_X1 U10806 ( .A1(n8384), .A2(n8383), .ZN(n8386) );
  NAND2_X1 U10807 ( .A1(n8386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8385) );
  MUX2_X1 U10808 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8385), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8387) );
  OR2_X1 U10809 ( .A1(n8386), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8395) );
  AOI22_X1 U10810 ( .A1(n12196), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n8626), 
        .B2(n13869), .ZN(n8388) );
  NAND2_X1 U10811 ( .A1(n6649), .A2(n7078), .ZN(n8390) );
  OR2_X1 U10812 ( .A1(n8392), .A2(n8391), .ZN(n8393) );
  AND2_X1 U10813 ( .A1(n8394), .A2(n8393), .ZN(n9658) );
  NAND2_X1 U10814 ( .A1(n9658), .A2(n12195), .ZN(n8398) );
  NAND2_X1 U10815 ( .A1(n8395), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8396) );
  XNOR2_X1 U10816 ( .A(n8396), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9133) );
  AOI22_X1 U10817 ( .A1(n12196), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8626), 
        .B2(n9133), .ZN(n8397) );
  NAND2_X1 U10818 ( .A1(n8398), .A2(n8397), .ZN(n14722) );
  NAND2_X1 U10819 ( .A1(n12178), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8403) );
  INV_X1 U10820 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n8399) );
  OR2_X1 U10821 ( .A1(n12179), .A2(n8399), .ZN(n8402) );
  OAI21_X1 U10822 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n8413), .ZN(n9984) );
  OR2_X1 U10823 ( .A1(n6647), .A2(n9984), .ZN(n8401) );
  INV_X1 U10824 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9134) );
  OR2_X1 U10825 ( .A1(n6650), .A2(n9134), .ZN(n8400) );
  XNOR2_X1 U10826 ( .A(n14722), .B(n13837), .ZN(n12213) );
  INV_X1 U10827 ( .A(n12213), .ZN(n9973) );
  NAND2_X1 U10828 ( .A1(n9974), .A2(n9973), .ZN(n9972) );
  OR2_X1 U10829 ( .A1(n14722), .A2(n13837), .ZN(n8404) );
  OR2_X1 U10830 ( .A1(n8406), .A2(n8405), .ZN(n8407) );
  NAND2_X1 U10831 ( .A1(n8408), .A2(n8407), .ZN(n9665) );
  OR2_X1 U10832 ( .A1(n9665), .A2(n8369), .ZN(n8411) );
  OR2_X1 U10833 ( .A1(n8422), .A2(n8317), .ZN(n8409) );
  XNOR2_X1 U10834 ( .A(n8409), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9136) );
  AOI22_X1 U10835 ( .A1(n12196), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8626), 
        .B2(n9136), .ZN(n8410) );
  NAND2_X1 U10836 ( .A1(n12178), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8418) );
  INV_X1 U10837 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8412) );
  OR2_X1 U10838 ( .A1(n12179), .A2(n8412), .ZN(n8417) );
  AND2_X1 U10839 ( .A1(n8413), .A2(n9156), .ZN(n8414) );
  OR2_X1 U10840 ( .A1(n8414), .A2(n8429), .ZN(n10083) );
  OR2_X1 U10841 ( .A1(n6647), .A2(n10083), .ZN(n8416) );
  INV_X1 U10842 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9135) );
  OR2_X1 U10843 ( .A1(n6651), .A2(n9135), .ZN(n8415) );
  NAND4_X1 U10844 ( .A1(n8418), .A2(n8417), .A3(n8416), .A4(n8415), .ZN(n13836) );
  XNOR2_X1 U10845 ( .A(n12052), .B(n13836), .ZN(n12216) );
  INV_X1 U10846 ( .A(n13836), .ZN(n10041) );
  OR2_X1 U10847 ( .A1(n9847), .A2(n8369), .ZN(n8428) );
  INV_X1 U10848 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U10849 ( .A1(n8422), .A2(n8421), .ZN(n8423) );
  NOR2_X1 U10850 ( .A1(n8423), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8456) );
  INV_X1 U10851 ( .A(n8456), .ZN(n8426) );
  NAND2_X1 U10852 ( .A1(n8423), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8424) );
  MUX2_X1 U10853 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8424), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n8425) );
  AOI22_X1 U10854 ( .A1(n12196), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8626), 
        .B2(n9137), .ZN(n8427) );
  NAND2_X1 U10855 ( .A1(n12178), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8434) );
  INV_X1 U10856 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10061) );
  OR2_X1 U10857 ( .A1(n6651), .A2(n10061), .ZN(n8433) );
  OR2_X1 U10858 ( .A1(n8429), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U10859 ( .A1(n8444), .A2(n8430), .ZN(n10054) );
  OR2_X1 U10860 ( .A1(n6647), .A2(n10054), .ZN(n8432) );
  INV_X1 U10861 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9198) );
  OR2_X1 U10862 ( .A1(n12179), .A2(n9198), .ZN(n8431) );
  NAND4_X1 U10863 ( .A1(n8434), .A2(n8433), .A3(n8432), .A4(n8431), .ZN(n13835) );
  INV_X1 U10864 ( .A(n13835), .ZN(n9910) );
  OR2_X1 U10865 ( .A1(n12056), .A2(n13835), .ZN(n8435) );
  NAND2_X1 U10866 ( .A1(n8437), .A2(n8436), .ZN(n8439) );
  NAND2_X1 U10867 ( .A1(n10116), .A2(n12195), .ZN(n8442) );
  OR2_X1 U10868 ( .A1(n8456), .A2(n8317), .ZN(n8440) );
  XNOR2_X1 U10869 ( .A(n8440), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13910) );
  AOI22_X1 U10870 ( .A1(n12196), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8626), 
        .B2(n13910), .ZN(n8441) );
  NAND2_X1 U10871 ( .A1(n8442), .A2(n8441), .ZN(n12064) );
  NAND2_X1 U10872 ( .A1(n8718), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8449) );
  INV_X1 U10873 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8443) );
  OR2_X1 U10874 ( .A1(n8720), .A2(n8443), .ZN(n8448) );
  NAND2_X1 U10875 ( .A1(n8444), .A2(n10191), .ZN(n8445) );
  NAND2_X1 U10876 ( .A1(n8460), .A2(n8445), .ZN(n10192) );
  OR2_X1 U10877 ( .A1(n6647), .A2(n10192), .ZN(n8447) );
  INV_X1 U10878 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9205) );
  OR2_X1 U10879 ( .A1(n6650), .A2(n9205), .ZN(n8446) );
  NAND4_X1 U10880 ( .A1(n8449), .A2(n8448), .A3(n8447), .A4(n8446), .ZN(n13834) );
  XNOR2_X1 U10881 ( .A(n12064), .B(n13834), .ZN(n12219) );
  INV_X1 U10882 ( .A(n12219), .ZN(n9908) );
  OR2_X1 U10883 ( .A1(n12064), .A2(n13834), .ZN(n8450) );
  AND2_X1 U10884 ( .A1(n8452), .A2(n8451), .ZN(n8454) );
  NAND2_X1 U10885 ( .A1(n10201), .A2(n12195), .ZN(n8458) );
  INV_X1 U10886 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10887 ( .A1(n8456), .A2(n8455), .ZN(n8502) );
  NAND2_X1 U10888 ( .A1(n8502), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8471) );
  XNOR2_X1 U10889 ( .A(n8471), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9207) );
  AOI22_X1 U10890 ( .A1(n12196), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8626), 
        .B2(n9207), .ZN(n8457) );
  NAND2_X1 U10891 ( .A1(n12178), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8465) );
  INV_X1 U10892 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9307) );
  OR2_X1 U10893 ( .A1(n6651), .A2(n9307), .ZN(n8464) );
  NAND2_X1 U10894 ( .A1(n8460), .A2(n8459), .ZN(n8461) );
  NAND2_X1 U10895 ( .A1(n8479), .A2(n8461), .ZN(n10439) );
  OR2_X1 U10896 ( .A1(n6647), .A2(n10439), .ZN(n8463) );
  INV_X1 U10897 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9197) );
  OR2_X1 U10898 ( .A1(n12179), .A2(n9197), .ZN(n8462) );
  NAND4_X1 U10899 ( .A1(n8465), .A2(n8464), .A3(n8463), .A4(n8462), .ZN(n13833) );
  XNOR2_X1 U10900 ( .A(n12067), .B(n13833), .ZN(n12220) );
  OR2_X1 U10901 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  NAND2_X1 U10902 ( .A1(n8469), .A2(n8468), .ZN(n10263) );
  OR2_X1 U10903 ( .A1(n10263), .A2(n8369), .ZN(n8477) );
  INV_X1 U10904 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10905 ( .A1(n8471), .A2(n8470), .ZN(n8472) );
  NAND2_X1 U10906 ( .A1(n8472), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8474) );
  INV_X1 U10907 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10908 ( .A1(n8474), .A2(n8473), .ZN(n8489) );
  OR2_X1 U10909 ( .A1(n8474), .A2(n8473), .ZN(n8475) );
  AOI22_X1 U10910 ( .A1(n12196), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8626), 
        .B2(n9309), .ZN(n8476) );
  NAND2_X1 U10911 ( .A1(n12178), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8485) );
  INV_X1 U10912 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n8478) );
  OR2_X1 U10913 ( .A1(n12179), .A2(n8478), .ZN(n8484) );
  INV_X1 U10914 ( .A(n8506), .ZN(n8481) );
  NAND2_X1 U10915 ( .A1(n8479), .A2(n13925), .ZN(n8480) );
  NAND2_X1 U10916 ( .A1(n8481), .A2(n8480), .ZN(n14666) );
  OR2_X1 U10917 ( .A1(n6647), .A2(n14666), .ZN(n8483) );
  INV_X1 U10918 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n14667) );
  OR2_X1 U10919 ( .A1(n6650), .A2(n14667), .ZN(n8482) );
  NAND4_X1 U10920 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n13832) );
  XNOR2_X1 U10921 ( .A(n14671), .B(n13832), .ZN(n12222) );
  OR2_X1 U10922 ( .A1(n14671), .A2(n13832), .ZN(n8486) );
  XNOR2_X1 U10923 ( .A(n8488), .B(n8487), .ZN(n10351) );
  NAND2_X1 U10924 ( .A1(n10351), .A2(n12195), .ZN(n8492) );
  NAND2_X1 U10925 ( .A1(n8489), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8490) );
  XNOR2_X1 U10926 ( .A(n8490), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9404) );
  AOI22_X1 U10927 ( .A1(n12196), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9404), 
        .B2(n8626), .ZN(n8491) );
  NAND2_X1 U10928 ( .A1(n8718), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8496) );
  OR2_X1 U10929 ( .A1(n8720), .A2(n14754), .ZN(n8495) );
  XNOR2_X1 U10930 ( .A(n8506), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n10845) );
  OR2_X1 U10931 ( .A1(n6647), .A2(n10845), .ZN(n8494) );
  INV_X1 U10932 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10309) );
  OR2_X1 U10933 ( .A1(n6651), .A2(n10309), .ZN(n8493) );
  NAND4_X1 U10934 ( .A1(n8496), .A2(n8495), .A3(n8494), .A4(n8493), .ZN(n13831) );
  INV_X1 U10935 ( .A(n13831), .ZN(n14595) );
  XNOR2_X1 U10936 ( .A(n14744), .B(n14595), .ZN(n12224) );
  OR2_X1 U10937 ( .A1(n14744), .A2(n13831), .ZN(n8497) );
  XNOR2_X1 U10938 ( .A(n8499), .B(n8498), .ZN(n10515) );
  NAND2_X1 U10939 ( .A1(n10515), .A2(n12195), .ZN(n8505) );
  INV_X1 U10940 ( .A(n8500), .ZN(n8501) );
  NAND2_X1 U10941 ( .A1(n8517), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8503) );
  XNOR2_X1 U10942 ( .A(n8503), .B(P1_IR_REG_11__SCAN_IN), .ZN(n13945) );
  AOI22_X1 U10943 ( .A1(n12196), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8626), 
        .B2(n13945), .ZN(n8504) );
  NAND2_X1 U10944 ( .A1(n12178), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U10945 ( .A1(n8506), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8508) );
  INV_X1 U10946 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U10947 ( .A1(n8508), .A2(n8507), .ZN(n8509) );
  NAND2_X1 U10948 ( .A1(n8509), .A2(n8521), .ZN(n14605) );
  OR2_X1 U10949 ( .A1(n6647), .A2(n14605), .ZN(n8513) );
  INV_X1 U10950 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9399) );
  OR2_X1 U10951 ( .A1(n6650), .A2(n9399), .ZN(n8512) );
  INV_X1 U10952 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8510) );
  OR2_X1 U10953 ( .A1(n12179), .A2(n8510), .ZN(n8511) );
  NAND4_X1 U10954 ( .A1(n8514), .A2(n8513), .A3(n8512), .A4(n8511), .ZN(n13830) );
  XNOR2_X1 U10955 ( .A(n14607), .B(n13830), .ZN(n12225) );
  INV_X1 U10956 ( .A(n12225), .ZN(n10418) );
  XNOR2_X1 U10957 ( .A(n8515), .B(n8516), .ZN(n10749) );
  NAND2_X1 U10958 ( .A1(n10749), .A2(n12195), .ZN(n8519) );
  OAI21_X1 U10959 ( .B1(n8517), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8531) );
  XNOR2_X1 U10960 ( .A(n8531), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9406) );
  AOI22_X1 U10961 ( .A1(n12196), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8626), 
        .B2(n9406), .ZN(n8518) );
  NAND2_X1 U10962 ( .A1(n8718), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8526) );
  INV_X1 U10963 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8520) );
  OR2_X1 U10964 ( .A1(n8720), .A2(n8520), .ZN(n8525) );
  NAND2_X1 U10965 ( .A1(n8521), .A2(n11129), .ZN(n8522) );
  NAND2_X1 U10966 ( .A1(n8536), .A2(n8522), .ZN(n10578) );
  OR2_X1 U10967 ( .A1(n6647), .A2(n10578), .ZN(n8524) );
  INV_X1 U10968 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9397) );
  OR2_X1 U10969 ( .A1(n6650), .A2(n9397), .ZN(n8523) );
  NAND4_X1 U10970 ( .A1(n8526), .A2(n8525), .A3(n8524), .A4(n8523), .ZN(n13829) );
  XNOR2_X1 U10971 ( .A(n12082), .B(n13829), .ZN(n12226) );
  INV_X1 U10972 ( .A(n12226), .ZN(n10574) );
  NAND2_X1 U10973 ( .A1(n10575), .A2(n10574), .ZN(n10573) );
  OR2_X1 U10974 ( .A1(n12082), .A2(n13829), .ZN(n8527) );
  XNOR2_X1 U10975 ( .A(n8529), .B(n8528), .ZN(n10755) );
  NAND2_X1 U10976 ( .A1(n10755), .A2(n12195), .ZN(n8534) );
  INV_X1 U10977 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U10978 ( .A1(n8531), .A2(n8530), .ZN(n8532) );
  NAND2_X1 U10979 ( .A1(n8532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8546) );
  XNOR2_X1 U10980 ( .A(n8546), .B(n8545), .ZN(n9778) );
  INV_X1 U10981 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15496) );
  OR2_X1 U10982 ( .A1(n8720), .A2(n15496), .ZN(n8542) );
  INV_X1 U10983 ( .A(n8551), .ZN(n8538) );
  NAND2_X1 U10984 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  NAND2_X1 U10985 ( .A1(n8538), .A2(n8537), .ZN(n11251) );
  OR2_X1 U10986 ( .A1(n6647), .A2(n11251), .ZN(n8541) );
  INV_X1 U10987 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9482) );
  OR2_X1 U10988 ( .A1(n6651), .A2(n9482), .ZN(n8540) );
  INV_X1 U10989 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9772) );
  OR2_X1 U10990 ( .A1(n12179), .A2(n9772), .ZN(n8539) );
  NAND4_X1 U10991 ( .A1(n8542), .A2(n8541), .A3(n8540), .A4(n8539), .ZN(n13828) );
  INV_X1 U10992 ( .A(n13828), .ZN(n12090) );
  OR2_X1 U10993 ( .A1(n12092), .A2(n12090), .ZN(n8796) );
  NAND2_X1 U10994 ( .A1(n12092), .A2(n12090), .ZN(n8543) );
  OR2_X1 U10995 ( .A1(n12092), .A2(n13828), .ZN(n8544) );
  XNOR2_X1 U10996 ( .A(n8559), .B(SI_14_), .ZN(n8562) );
  XNOR2_X1 U10997 ( .A(n8562), .B(n8561), .ZN(n10932) );
  NAND2_X1 U10998 ( .A1(n10932), .A2(n12195), .ZN(n8550) );
  NAND2_X1 U10999 ( .A1(n8546), .A2(n8545), .ZN(n8547) );
  NAND2_X1 U11000 ( .A1(n8547), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8548) );
  XNOR2_X1 U11001 ( .A(n8548), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U11002 ( .A1(n9768), .A2(n8626), .B1(n12196), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8549) );
  INV_X1 U11003 ( .A(n6647), .ZN(n8604) );
  NOR2_X1 U11004 ( .A1(n8551), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8552) );
  OR2_X1 U11005 ( .A1(n8568), .A2(n8552), .ZN(n14591) );
  INV_X1 U11006 ( .A(n14591), .ZN(n10828) );
  NAND2_X1 U11007 ( .A1(n8604), .A2(n10828), .ZN(n8557) );
  INV_X1 U11008 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8553) );
  OR2_X1 U11009 ( .A1(n8720), .A2(n8553), .ZN(n8556) );
  INV_X1 U11010 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10664) );
  OR2_X1 U11011 ( .A1(n6650), .A2(n10664), .ZN(n8555) );
  INV_X1 U11012 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10668) );
  OR2_X1 U11013 ( .A1(n12179), .A2(n10668), .ZN(n8554) );
  NAND4_X1 U11014 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(n13827) );
  INV_X1 U11015 ( .A(n13827), .ZN(n8558) );
  OR2_X1 U11016 ( .A1(n14584), .A2(n8558), .ZN(n12097) );
  NAND2_X1 U11017 ( .A1(n14584), .A2(n8558), .ZN(n12089) );
  AND2_X1 U11018 ( .A1(n8559), .A2(n15380), .ZN(n8560) );
  XNOR2_X1 U11019 ( .A(n8563), .B(SI_15_), .ZN(n8564) );
  NAND2_X1 U11020 ( .A1(n11062), .A2(n12195), .ZN(n8567) );
  NAND2_X1 U11021 ( .A1(n8763), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8565) );
  XNOR2_X1 U11022 ( .A(n8565), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U11023 ( .A1(n12196), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8626), 
        .B2(n10670), .ZN(n8566) );
  OR2_X1 U11024 ( .A1(n8568), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8569) );
  AND2_X1 U11025 ( .A1(n8590), .A2(n8569), .ZN(n13805) );
  NAND2_X1 U11026 ( .A1(n8604), .A2(n13805), .ZN(n8574) );
  INV_X1 U11027 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11109) );
  OR2_X1 U11028 ( .A1(n12179), .A2(n11109), .ZN(n8573) );
  INV_X1 U11029 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15452) );
  OR2_X1 U11030 ( .A1(n8720), .A2(n15452), .ZN(n8572) );
  INV_X1 U11031 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8570) );
  OR2_X1 U11032 ( .A1(n6650), .A2(n8570), .ZN(n8571) );
  NAND4_X1 U11033 ( .A1(n8574), .A2(n8573), .A3(n8572), .A4(n8571), .ZN(n13826) );
  INV_X1 U11034 ( .A(n13826), .ZN(n8575) );
  NAND2_X1 U11035 ( .A1(n13815), .A2(n8575), .ZN(n12103) );
  OR2_X1 U11036 ( .A1(n13815), .A2(n13826), .ZN(n8576) );
  XNOR2_X1 U11037 ( .A(n8578), .B(n8577), .ZN(n11169) );
  NAND2_X1 U11038 ( .A1(n11169), .A2(n12195), .ZN(n8588) );
  NAND2_X1 U11039 ( .A1(n8583), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8581) );
  MUX2_X1 U11040 ( .A(n8581), .B(P1_IR_REG_31__SCAN_IN), .S(n8584), .Z(n8582)
         );
  INV_X1 U11041 ( .A(n8582), .ZN(n8586) );
  AOI22_X1 U11042 ( .A1(n12196), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8626), 
        .B2(n10880), .ZN(n8587) );
  NAND2_X1 U11043 ( .A1(n8590), .A2(n8589), .ZN(n8591) );
  NAND2_X1 U11044 ( .A1(n8616), .A2(n8591), .ZN(n13746) );
  INV_X1 U11045 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8592) );
  OR2_X1 U11046 ( .A1(n8720), .A2(n8592), .ZN(n8594) );
  INV_X1 U11047 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n15418) );
  OR2_X1 U11048 ( .A1(n12179), .A2(n15418), .ZN(n8593) );
  AND2_X1 U11049 ( .A1(n8594), .A2(n8593), .ZN(n8596) );
  INV_X1 U11050 ( .A(n6651), .ZN(n8755) );
  NAND2_X1 U11051 ( .A1(n8755), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8595) );
  OAI211_X1 U11052 ( .C1(n13746), .C2(n6647), .A(n8596), .B(n8595), .ZN(n13825) );
  INV_X1 U11053 ( .A(n13825), .ZN(n12104) );
  XNOR2_X1 U11054 ( .A(n14276), .B(n12104), .ZN(n12230) );
  OR2_X1 U11055 ( .A1(n14276), .A2(n13825), .ZN(n8597) );
  XNOR2_X1 U11056 ( .A(n8599), .B(n8598), .ZN(n11261) );
  NAND2_X1 U11057 ( .A1(n11261), .A2(n12195), .ZN(n8603) );
  NAND2_X1 U11058 ( .A1(n8600), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8601) );
  XNOR2_X1 U11059 ( .A(n8601), .B(n8612), .ZN(n11051) );
  INV_X1 U11060 ( .A(n11051), .ZN(n10883) );
  AOI22_X1 U11061 ( .A1(n12196), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8626), 
        .B2(n10883), .ZN(n8602) );
  XNOR2_X1 U11062 ( .A(n8616), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n13756) );
  NAND2_X1 U11063 ( .A1(n13756), .A2(n8604), .ZN(n8609) );
  INV_X1 U11064 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11048) );
  NAND2_X1 U11065 ( .A1(n12178), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8606) );
  INV_X1 U11066 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14271) );
  OR2_X1 U11067 ( .A1(n12179), .A2(n14271), .ZN(n8605) );
  OAI211_X1 U11068 ( .C1(n11048), .C2(n6651), .A(n8606), .B(n8605), .ZN(n8607)
         );
  INV_X1 U11069 ( .A(n8607), .ZN(n8608) );
  XNOR2_X1 U11070 ( .A(n8611), .B(n8610), .ZN(n11481) );
  NAND2_X1 U11071 ( .A1(n11481), .A2(n12195), .ZN(n8615) );
  NAND2_X1 U11072 ( .A1(n8624), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8613) );
  XNOR2_X1 U11073 ( .A(n8613), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13959) );
  AOI22_X1 U11074 ( .A1(n12196), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8626), 
        .B2(n13959), .ZN(n8614) );
  INV_X1 U11075 ( .A(n8616), .ZN(n8617) );
  AOI21_X1 U11076 ( .B1(n8617), .B2(P1_REG3_REG_17__SCAN_IN), .A(
        P1_REG3_REG_18__SCAN_IN), .ZN(n8618) );
  OR2_X1 U11077 ( .A1(n8618), .A2(n8629), .ZN(n13786) );
  AOI22_X1 U11078 ( .A1(n12178), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n8718), 
        .B2(P1_REG1_REG_18__SCAN_IN), .ZN(n8620) );
  INV_X1 U11079 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n11288) );
  OR2_X1 U11080 ( .A1(n6650), .A2(n11288), .ZN(n8619) );
  OAI211_X1 U11081 ( .C1(n13786), .C2(n6647), .A(n8620), .B(n8619), .ZN(n13823) );
  OR2_X1 U11082 ( .A1(n11807), .A2(n13823), .ZN(n8621) );
  XNOR2_X1 U11083 ( .A(n8623), .B(n8622), .ZN(n11489) );
  NAND2_X1 U11084 ( .A1(n11489), .A2(n12195), .ZN(n8628) );
  XNOR2_X2 U11085 ( .A(n8625), .B(P1_IR_REG_19__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U11086 ( .A1(n12196), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14114), 
        .B2(n8626), .ZN(n8627) );
  OR2_X1 U11087 ( .A1(n8629), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U11088 ( .A1(n8645), .A2(n8630), .ZN(n14179) );
  AOI22_X1 U11089 ( .A1(n12178), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n8718), 
        .B2(P1_REG1_REG_19__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U11090 ( .A1(n8755), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8631) );
  OAI211_X1 U11091 ( .C1(n14179), .C2(n6647), .A(n8632), .B(n8631), .ZN(n13822) );
  INV_X1 U11092 ( .A(n13822), .ZN(n14261) );
  OR2_X1 U11093 ( .A1(n14185), .A2(n14261), .ZN(n12124) );
  NAND2_X1 U11094 ( .A1(n14185), .A2(n14261), .ZN(n12125) );
  OR2_X1 U11095 ( .A1(n14185), .A2(n13822), .ZN(n8634) );
  NAND2_X1 U11096 ( .A1(n8636), .A2(n8635), .ZN(n8637) );
  NAND2_X1 U11097 ( .A1(n8637), .A2(n10047), .ZN(n8638) );
  NAND2_X1 U11098 ( .A1(n8655), .A2(n8638), .ZN(n8640) );
  NAND2_X1 U11099 ( .A1(n8640), .A2(n8639), .ZN(n8641) );
  NAND2_X1 U11100 ( .A1(n12196), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11101 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND2_X1 U11102 ( .A1(n8663), .A2(n8646), .ZN(n14153) );
  OR2_X1 U11103 ( .A1(n14153), .A2(n6647), .ZN(n8652) );
  INV_X1 U11104 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U11105 ( .A1(n8718), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U11106 ( .A1(n12178), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8647) );
  OAI211_X1 U11107 ( .C1(n8649), .C2(n6650), .A(n8648), .B(n8647), .ZN(n8650)
         );
  INV_X1 U11108 ( .A(n8650), .ZN(n8651) );
  NAND2_X1 U11109 ( .A1(n8652), .A2(n8651), .ZN(n13821) );
  XNOR2_X1 U11110 ( .A(n14248), .B(n14253), .ZN(n14157) );
  NAND2_X1 U11111 ( .A1(n14248), .A2(n13821), .ZN(n8653) );
  AND2_X1 U11112 ( .A1(n8655), .A2(n8654), .ZN(n8656) );
  NAND2_X1 U11113 ( .A1(n8657), .A2(n8656), .ZN(n8659) );
  NAND2_X1 U11114 ( .A1(n8659), .A2(n8658), .ZN(n11523) );
  OR2_X1 U11115 ( .A1(n11523), .A2(n8369), .ZN(n8661) );
  NAND2_X1 U11116 ( .A1(n12196), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8660) );
  AND2_X1 U11117 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  OR2_X1 U11118 ( .A1(n8671), .A2(n8664), .ZN(n14138) );
  INV_X1 U11119 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U11120 ( .A1(n8718), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U11121 ( .A1(n12178), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8665) );
  OAI211_X1 U11122 ( .C1(n14139), .C2(n6651), .A(n8666), .B(n8665), .ZN(n8667)
         );
  INV_X1 U11123 ( .A(n8667), .ZN(n8668) );
  INV_X1 U11124 ( .A(n13820), .ZN(n14159) );
  XNOR2_X1 U11125 ( .A(n14303), .B(n14159), .ZN(n14142) );
  OR2_X1 U11126 ( .A1(n8669), .A2(n9468), .ZN(n8670) );
  XNOR2_X1 U11127 ( .A(n8670), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14334) );
  OR2_X1 U11128 ( .A1(n8671), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U11129 ( .A1(n8672), .A2(n8687), .ZN(n11850) );
  OR2_X1 U11130 ( .A1(n11850), .A2(n6647), .ZN(n8678) );
  INV_X1 U11131 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11132 ( .A1(n8718), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U11133 ( .A1(n8755), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8673) );
  OAI211_X1 U11134 ( .C1(n8720), .C2(n8675), .A(n8674), .B(n8673), .ZN(n8676)
         );
  INV_X1 U11135 ( .A(n8676), .ZN(n8677) );
  NAND2_X1 U11136 ( .A1(n14234), .A2(n13819), .ZN(n8679) );
  NAND2_X1 U11137 ( .A1(n14104), .A2(n8679), .ZN(n14126) );
  NAND2_X1 U11138 ( .A1(n14234), .A2(n13724), .ZN(n8680) );
  NAND2_X1 U11139 ( .A1(n14125), .A2(n8680), .ZN(n14100) );
  INV_X1 U11140 ( .A(n14100), .ZN(n8695) );
  XNOR2_X1 U11141 ( .A(n8681), .B(SI_23_), .ZN(n8682) );
  XNOR2_X1 U11142 ( .A(n8683), .B(n8682), .ZN(n11555) );
  NAND2_X1 U11143 ( .A1(n11555), .A2(n12195), .ZN(n8685) );
  NAND2_X1 U11144 ( .A1(n12196), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U11145 ( .A1(n8718), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8693) );
  INV_X1 U11146 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8686) );
  OR2_X1 U11147 ( .A1(n8720), .A2(n8686), .ZN(n8692) );
  INV_X1 U11148 ( .A(n8687), .ZN(n8689) );
  INV_X1 U11149 ( .A(n8705), .ZN(n8688) );
  OAI21_X1 U11150 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8689), .A(n8688), .ZN(
        n14101) );
  OR2_X1 U11151 ( .A1(n6647), .A2(n14101), .ZN(n8691) );
  INV_X1 U11152 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14102) );
  OR2_X1 U11153 ( .A1(n6650), .A2(n14102), .ZN(n8690) );
  NAND4_X1 U11154 ( .A1(n8693), .A2(n8692), .A3(n8691), .A4(n8690), .ZN(n14081) );
  XNOR2_X1 U11155 ( .A(n14110), .B(n14081), .ZN(n14106) );
  INV_X1 U11156 ( .A(n14106), .ZN(n8694) );
  NAND2_X1 U11157 ( .A1(n14110), .A2(n14081), .ZN(n8696) );
  NAND2_X1 U11158 ( .A1(n8698), .A2(n8697), .ZN(n8699) );
  NAND2_X1 U11159 ( .A1(n8700), .A2(n8699), .ZN(n11573) );
  NAND2_X1 U11160 ( .A1(n12196), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U11161 ( .A1(n8718), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8709) );
  INV_X1 U11162 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8703) );
  OR2_X1 U11163 ( .A1(n8720), .A2(n8703), .ZN(n8708) );
  OAI21_X1 U11164 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8705), .A(n8704), .ZN(
        n14088) );
  OR2_X1 U11165 ( .A1(n6647), .A2(n14088), .ZN(n8707) );
  INV_X1 U11166 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14089) );
  OR2_X1 U11167 ( .A1(n6651), .A2(n14089), .ZN(n8706) );
  NAND4_X1 U11168 ( .A1(n8709), .A2(n8708), .A3(n8707), .A4(n8706), .ZN(n14061) );
  XNOR2_X1 U11169 ( .A(n14094), .B(n14061), .ZN(n14083) );
  INV_X1 U11170 ( .A(n14061), .ZN(n12149) );
  NAND2_X1 U11171 ( .A1(n14091), .A2(n12149), .ZN(n8710) );
  NAND2_X1 U11172 ( .A1(n14067), .A2(n13799), .ZN(n8808) );
  OR2_X1 U11173 ( .A1(n14067), .A2(n13799), .ZN(n8711) );
  NAND2_X1 U11174 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  NAND2_X1 U11175 ( .A1(n11651), .A2(n12195), .ZN(n8717) );
  NAND2_X1 U11176 ( .A1(n12196), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U11177 ( .A1(n8718), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8728) );
  INV_X1 U11178 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8719) );
  OR2_X1 U11179 ( .A1(n8720), .A2(n8719), .ZN(n8727) );
  INV_X1 U11180 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U11181 ( .A1(n8722), .A2(n8721), .ZN(n8723) );
  NAND2_X1 U11182 ( .A1(n8724), .A2(n8723), .ZN(n14044) );
  OR2_X1 U11183 ( .A1(n6647), .A2(n14044), .ZN(n8726) );
  INV_X1 U11184 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14045) );
  OR2_X1 U11185 ( .A1(n6650), .A2(n14045), .ZN(n8725) );
  NAND4_X1 U11186 ( .A1(n8728), .A2(n8727), .A3(n8726), .A4(n8725), .ZN(n14060) );
  XNOR2_X1 U11187 ( .A(n14049), .B(n8809), .ZN(n12239) );
  INV_X1 U11188 ( .A(n14042), .ZN(n8729) );
  NAND2_X1 U11189 ( .A1(n14032), .A2(n8729), .ZN(n8811) );
  OAI21_X1 U11190 ( .B1(n14032), .B2(n8729), .A(n8811), .ZN(n14021) );
  NAND2_X1 U11191 ( .A1(n8730), .A2(n11112), .ZN(n8731) );
  NAND2_X1 U11192 ( .A1(n8733), .A2(SI_27_), .ZN(n8734) );
  XNOR2_X1 U11193 ( .A(n8750), .B(SI_28_), .ZN(n8751) );
  NAND2_X1 U11194 ( .A1(n13686), .A2(n12195), .ZN(n8737) );
  NAND2_X1 U11195 ( .A1(n12196), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U11196 ( .A1(n12178), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8747) );
  INV_X1 U11197 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8738) );
  OR2_X1 U11198 ( .A1(n12179), .A2(n8738), .ZN(n8746) );
  INV_X1 U11199 ( .A(n8741), .ZN(n8739) );
  NAND2_X1 U11200 ( .A1(n8739), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13988) );
  INV_X1 U11201 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U11202 ( .A1(n8741), .A2(n8740), .ZN(n8742) );
  NAND2_X1 U11203 ( .A1(n13988), .A2(n8742), .ZN(n14012) );
  OR2_X1 U11204 ( .A1(n6647), .A2(n14012), .ZN(n8745) );
  INV_X1 U11205 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8743) );
  OR2_X1 U11206 ( .A1(n6650), .A2(n8743), .ZN(n8744) );
  NAND4_X1 U11207 ( .A1(n8747), .A2(n8746), .A3(n8745), .A4(n8744), .ZN(n13818) );
  NAND2_X1 U11208 ( .A1(n14200), .A2(n14026), .ZN(n8812) );
  OR2_X1 U11209 ( .A1(n14200), .A2(n14026), .ZN(n8748) );
  NAND2_X1 U11210 ( .A1(n8812), .A2(n8748), .ZN(n12240) );
  INV_X1 U11211 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14326) );
  INV_X1 U11212 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13684) );
  MUX2_X1 U11213 ( .A(n14326), .B(n13684), .S(n9468), .Z(n11613) );
  XNOR2_X1 U11214 ( .A(n11613), .B(SI_29_), .ZN(n11612) );
  NAND2_X1 U11215 ( .A1(n13682), .A2(n12195), .ZN(n8754) );
  NAND2_X1 U11216 ( .A1(n12196), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11217 ( .A1(n12178), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U11218 ( .A1(n8755), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8758) );
  INV_X1 U11219 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8861) );
  OR2_X1 U11220 ( .A1(n12179), .A2(n8861), .ZN(n8757) );
  OR2_X1 U11221 ( .A1(n6647), .A2(n13988), .ZN(n8756) );
  NAND4_X1 U11222 ( .A1(n8759), .A2(n8758), .A3(n8757), .A4(n8756), .ZN(n14002) );
  XNOR2_X1 U11223 ( .A(n13992), .B(n14002), .ZN(n12241) );
  INV_X1 U11224 ( .A(n8761), .ZN(n8762) );
  NOR2_X2 U11225 ( .A1(n8768), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n8766) );
  INV_X1 U11226 ( .A(n8766), .ZN(n8770) );
  NAND2_X1 U11227 ( .A1(n8770), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11228 ( .A1(n8766), .A2(n8765), .ZN(n8772) );
  NAND2_X1 U11229 ( .A1(n8768), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8769) );
  MUX2_X1 U11230 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8769), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8771) );
  NOR2_X2 U11231 ( .A1(n12206), .A2(n12205), .ZN(n9962) );
  OR2_X1 U11232 ( .A1(n12029), .A2(n12027), .ZN(n9975) );
  AND2_X1 U11233 ( .A1(n9975), .A2(n8775), .ZN(n8776) );
  AND2_X2 U11234 ( .A1(n12027), .A2(n12029), .ZN(n12295) );
  AND2_X1 U11235 ( .A1(n12025), .A2(n10649), .ZN(n12200) );
  NAND2_X1 U11236 ( .A1(n12200), .A2(n14114), .ZN(n14221) );
  NAND2_X1 U11237 ( .A1(n9948), .A2(n8780), .ZN(n9730) );
  NAND2_X1 U11238 ( .A1(n9978), .A2(n12213), .ZN(n9977) );
  INV_X1 U11239 ( .A(n13837), .ZN(n12046) );
  NAND2_X1 U11240 ( .A1(n14722), .A2(n12046), .ZN(n8781) );
  NAND2_X1 U11241 ( .A1(n10082), .A2(n13836), .ZN(n8782) );
  NAND2_X1 U11242 ( .A1(n9748), .A2(n8782), .ZN(n8784) );
  NAND2_X1 U11243 ( .A1(n12052), .A2(n10041), .ZN(n8783) );
  INV_X1 U11244 ( .A(n12218), .ZN(n10057) );
  NAND2_X1 U11245 ( .A1(n10058), .A2(n10057), .ZN(n8786) );
  NAND2_X1 U11246 ( .A1(n12056), .A2(n9910), .ZN(n8785) );
  NAND2_X1 U11247 ( .A1(n8786), .A2(n8785), .ZN(n9907) );
  NAND2_X1 U11248 ( .A1(n9907), .A2(n12219), .ZN(n8788) );
  INV_X1 U11249 ( .A(n13834), .ZN(n10040) );
  NAND2_X1 U11250 ( .A1(n12064), .A2(n10040), .ZN(n8787) );
  NAND2_X1 U11251 ( .A1(n8788), .A2(n8787), .ZN(n10018) );
  INV_X1 U11252 ( .A(n10018), .ZN(n8789) );
  INV_X1 U11253 ( .A(n13833), .ZN(n9909) );
  OR2_X1 U11254 ( .A1(n12067), .A2(n9909), .ZN(n8790) );
  INV_X1 U11255 ( .A(n13832), .ZN(n8791) );
  NAND2_X1 U11256 ( .A1(n14671), .A2(n8791), .ZN(n8792) );
  NAND2_X1 U11257 ( .A1(n14658), .A2(n8792), .ZN(n10301) );
  OR2_X1 U11258 ( .A1(n14744), .A2(n14595), .ZN(n8793) );
  INV_X1 U11259 ( .A(n13830), .ZN(n10844) );
  OR2_X1 U11260 ( .A1(n14607), .A2(n10844), .ZN(n8794) );
  NAND2_X1 U11261 ( .A1(n10569), .A2(n12226), .ZN(n10568) );
  INV_X1 U11262 ( .A(n13829), .ZN(n14592) );
  OR2_X1 U11263 ( .A1(n12082), .A2(n14592), .ZN(n8795) );
  NAND2_X1 U11264 ( .A1(n10568), .A2(n8795), .ZN(n10632) );
  NAND2_X1 U11265 ( .A1(n10636), .A2(n8796), .ZN(n10820) );
  NAND2_X1 U11266 ( .A1(n10820), .A2(n12209), .ZN(n10819) );
  NAND2_X1 U11267 ( .A1(n14276), .A2(n12104), .ZN(n8797) );
  NAND2_X1 U11268 ( .A1(n13761), .A2(n13745), .ZN(n12107) );
  INV_X1 U11269 ( .A(n12107), .ZN(n8798) );
  OR2_X1 U11270 ( .A1(n13761), .A2(n13745), .ZN(n12108) );
  INV_X1 U11271 ( .A(n13823), .ZN(n14171) );
  OR2_X1 U11272 ( .A1(n11807), .A2(n14171), .ZN(n12120) );
  NAND2_X1 U11273 ( .A1(n11807), .A2(n14171), .ZN(n12119) );
  NAND2_X1 U11274 ( .A1(n12120), .A2(n12119), .ZN(n12118) );
  NAND2_X1 U11275 ( .A1(n11284), .A2(n6876), .ZN(n8799) );
  NAND2_X1 U11276 ( .A1(n8799), .A2(n12120), .ZN(n14169) );
  OR2_X1 U11277 ( .A1(n14248), .A2(n14253), .ZN(n8800) );
  OR2_X1 U11278 ( .A1(n14303), .A2(n14159), .ZN(n8801) );
  NAND2_X1 U11279 ( .A1(n8802), .A2(n8801), .ZN(n14120) );
  INV_X1 U11280 ( .A(n14120), .ZN(n8804) );
  NAND2_X1 U11281 ( .A1(n14122), .A2(n14104), .ZN(n8805) );
  INV_X1 U11282 ( .A(n14081), .ZN(n13770) );
  NAND2_X1 U11283 ( .A1(n14110), .A2(n13770), .ZN(n8806) );
  NAND2_X1 U11284 ( .A1(n14091), .A2(n14061), .ZN(n14055) );
  AND2_X1 U11285 ( .A1(n12237), .A2(n14055), .ZN(n8807) );
  NAND2_X1 U11286 ( .A1(n14057), .A2(n8808), .ZN(n14041) );
  INV_X1 U11287 ( .A(n12239), .ZN(n14050) );
  NAND2_X1 U11288 ( .A1(n14041), .A2(n14050), .ZN(n14040) );
  NAND2_X1 U11289 ( .A1(n14049), .A2(n8809), .ZN(n8810) );
  INV_X1 U11290 ( .A(n14021), .ZN(n14025) );
  NAND2_X1 U11291 ( .A1(n14024), .A2(n14025), .ZN(n14023) );
  NAND2_X1 U11292 ( .A1(n14023), .A2(n8811), .ZN(n14000) );
  NAND2_X1 U11293 ( .A1(n14000), .A2(n14009), .ZN(n14001) );
  NAND2_X1 U11294 ( .A1(n14001), .A2(n8812), .ZN(n8814) );
  NAND2_X1 U11295 ( .A1(n14114), .A2(n14335), .ZN(n8815) );
  INV_X1 U11296 ( .A(n12206), .ZN(n12022) );
  NAND2_X1 U11297 ( .A1(n12022), .A2(n12205), .ZN(n12183) );
  INV_X1 U11298 ( .A(n8816), .ZN(n9084) );
  INV_X1 U11299 ( .A(n12067), .ZN(n10068) );
  NOR2_X2 U11300 ( .A1(n12034), .A2(n9995), .ZN(n9994) );
  NAND2_X1 U11301 ( .A1(n9994), .A2(n14714), .ZN(n9957) );
  AND2_X1 U11302 ( .A1(n9982), .A2(n10082), .ZN(n10053) );
  NAND2_X1 U11303 ( .A1(n14732), .A2(n10053), .ZN(n10052) );
  NOR2_X2 U11304 ( .A1(n14607), .A2(n10420), .ZN(n10576) );
  NAND2_X1 U11305 ( .A1(n11287), .A2(n14314), .ZN(n14175) );
  OR2_X2 U11306 ( .A1(n14030), .A2(n14200), .ZN(n14014) );
  AND2_X2 U11307 ( .A1(n12025), .A2(n12206), .ZN(n12023) );
  AND2_X4 U11308 ( .A1(n12023), .A2(n10649), .ZN(n14176) );
  AOI21_X1 U11309 ( .B1(n13992), .B2(n14014), .A(n14661), .ZN(n8818) );
  OR2_X2 U11310 ( .A1(n14014), .A2(n13992), .ZN(n13978) );
  NAND2_X1 U11311 ( .A1(n8818), .A2(n13978), .ZN(n13995) );
  INV_X1 U11312 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n13982) );
  INV_X1 U11313 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8820) );
  OR2_X1 U11314 ( .A1(n12179), .A2(n8820), .ZN(n8822) );
  NAND2_X1 U11315 ( .A1(n12178), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8821) );
  OAI211_X1 U11316 ( .C1(n6651), .C2(n13982), .A(n8822), .B(n8821), .ZN(n13817) );
  NAND2_X1 U11317 ( .A1(n12201), .A2(n8816), .ZN(n14260) );
  INV_X1 U11318 ( .A(P1_B_REG_SCAN_IN), .ZN(n8823) );
  NOR2_X1 U11319 ( .A1(n6843), .A2(n8823), .ZN(n8824) );
  NOR2_X1 U11320 ( .A1(n14260), .A2(n8824), .ZN(n13974) );
  NAND2_X1 U11321 ( .A1(n13817), .A2(n13974), .ZN(n13989) );
  NAND2_X1 U11322 ( .A1(n8838), .A2(n8826), .ZN(n8834) );
  NAND2_X1 U11323 ( .A1(n8834), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8835) );
  MUX2_X1 U11324 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8835), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8836) );
  MUX2_X1 U11325 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8840), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8842) );
  NAND2_X1 U11326 ( .A1(n8775), .A2(n10649), .ZN(n8860) );
  NAND2_X1 U11327 ( .A1(n8860), .A2(n12201), .ZN(n9233) );
  NAND3_X1 U11328 ( .A1(n9225), .A2(n8984), .A3(n9233), .ZN(n9389) );
  NOR4_X1 U11329 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n8846) );
  NOR4_X1 U11330 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8845) );
  NOR4_X1 U11331 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8844) );
  NOR4_X1 U11332 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n8843) );
  NAND4_X1 U11333 ( .A1(n8846), .A2(n8845), .A3(n8844), .A4(n8843), .ZN(n8855)
         );
  NOR2_X1 U11334 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n8850) );
  NOR4_X1 U11335 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8849) );
  NOR4_X1 U11336 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n8848) );
  NOR4_X1 U11337 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n8847) );
  NAND4_X1 U11338 ( .A1(n8850), .A2(n8849), .A3(n8848), .A4(n8847), .ZN(n8854)
         );
  NAND2_X1 U11339 ( .A1(n11212), .A2(P1_B_REG_SCAN_IN), .ZN(n8851) );
  MUX2_X1 U11340 ( .A(n8851), .B(P1_B_REG_SCAN_IN), .S(n8858), .Z(n8852) );
  INV_X1 U11341 ( .A(n9012), .ZN(n8853) );
  NAND2_X1 U11342 ( .A1(n11968), .A2(n11212), .ZN(n8856) );
  OAI21_X1 U11343 ( .B1(n9012), .B2(P1_D_REG_1__SCAN_IN), .A(n8856), .ZN(n9917) );
  NAND2_X1 U11344 ( .A1(n14176), .A2(n14114), .ZN(n9922) );
  AND2_X1 U11345 ( .A1(n9917), .A2(n9922), .ZN(n8857) );
  AND2_X1 U11346 ( .A1(n9921), .A2(n8857), .ZN(n8865) );
  OAI22_X1 U11347 ( .A1(n9012), .A2(P1_D_REG_0__SCAN_IN), .B1(n9017), .B2(
        n8858), .ZN(n9918) );
  INV_X1 U11348 ( .A(n9918), .ZN(n8859) );
  INV_X1 U11349 ( .A(n13992), .ZN(n8868) );
  NAND2_X1 U11350 ( .A1(n14764), .A2(n14743), .ZN(n14273) );
  INV_X1 U11351 ( .A(n8862), .ZN(n8863) );
  NAND2_X1 U11352 ( .A1(n8864), .A2(n8863), .ZN(P1_U3557) );
  NAND2_X1 U11353 ( .A1(n14755), .A2(n14743), .ZN(n14318) );
  INV_X1 U11354 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8867) );
  INV_X1 U11355 ( .A(n8869), .ZN(n8870) );
  NAND2_X1 U11356 ( .A1(n8871), .A2(n8870), .ZN(P1_U3525) );
  INV_X1 U11357 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8873) );
  INV_X1 U11358 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8872) );
  INV_X1 U11359 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8956) );
  AND2_X2 U11360 ( .A1(n8876), .A2(n8965), .ZN(n9043) );
  NOR2_X1 U11361 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), 
        .ZN(n8878) );
  INV_X1 U11362 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8880) );
  NOR2_X1 U11363 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n8882) );
  NAND4_X1 U11364 ( .A1(n8882), .A2(n8881), .A3(n9757), .A4(n9444), .ZN(n8888)
         );
  NOR2_X2 U11365 ( .A1(n8892), .A2(n8888), .ZN(n9050) );
  AND2_X2 U11366 ( .A1(n9050), .A2(n8885), .ZN(n9053) );
  NAND4_X1 U11367 ( .A1(n8886), .A2(n8885), .A3(n8902), .A4(n8884), .ZN(n8887)
         );
  NOR3_X1 U11368 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .A3(P2_IR_REG_26__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U11369 ( .A1(n8893), .A2(n8894), .ZN(n8897) );
  NAND2_X1 U11370 ( .A1(n8899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U11371 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8895), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8896) );
  NAND2_X1 U11372 ( .A1(n8897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8898) );
  MUX2_X1 U11373 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8898), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8900) );
  NOR2_X1 U11374 ( .A1(n11318), .A2(n11210), .ZN(n8901) );
  NAND2_X1 U11375 ( .A1(n10908), .A2(n8901), .ZN(n9437) );
  NAND2_X1 U11376 ( .A1(n9047), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8903) );
  INV_X1 U11377 ( .A(n10851), .ZN(n9058) );
  INV_X1 U11378 ( .A(n12686), .ZN(n8904) );
  OAI21_X1 U11379 ( .B1(n12769), .B2(n12535), .A(n10049), .ZN(n8905) );
  AND2_X4 U11380 ( .A1(n8906), .A2(n8905), .ZN(n11886) );
  INV_X2 U11381 ( .A(n11886), .ZN(n11895) );
  XNOR2_X1 U11382 ( .A(n10410), .B(n11895), .ZN(n10592) );
  XNOR2_X1 U11383 ( .A(n10723), .B(n10592), .ZN(n8931) );
  NAND2_X1 U11384 ( .A1(n15126), .A2(n11886), .ZN(n8907) );
  NAND2_X1 U11385 ( .A1(n8908), .A2(n8907), .ZN(n8914) );
  NAND2_X1 U11386 ( .A1(n8911), .A2(n11886), .ZN(n8909) );
  OR2_X1 U11387 ( .A1(n15112), .A2(n8909), .ZN(n8913) );
  INV_X1 U11388 ( .A(n11886), .ZN(n8910) );
  XNOR2_X1 U11389 ( .A(n8911), .B(n8910), .ZN(n8912) );
  NAND2_X1 U11390 ( .A1(n8914), .A2(n9794), .ZN(n9793) );
  XNOR2_X1 U11391 ( .A(n8915), .B(n11886), .ZN(n8916) );
  XNOR2_X1 U11392 ( .A(n8916), .B(n15135), .ZN(n9899) );
  NAND2_X1 U11393 ( .A1(n9898), .A2(n9899), .ZN(n9889) );
  XNOR2_X1 U11394 ( .A(n15155), .B(n11886), .ZN(n8919) );
  XNOR2_X1 U11395 ( .A(n8919), .B(n15111), .ZN(n9890) );
  INV_X1 U11396 ( .A(n8916), .ZN(n8917) );
  NAND2_X1 U11397 ( .A1(n8917), .A2(n15135), .ZN(n9891) );
  AND2_X1 U11398 ( .A1(n9890), .A2(n9891), .ZN(n8918) );
  INV_X1 U11399 ( .A(n8919), .ZN(n8920) );
  OR2_X1 U11400 ( .A1(n15111), .A2(n8920), .ZN(n8921) );
  XNOR2_X1 U11401 ( .A(n10252), .B(n11895), .ZN(n8922) );
  NAND2_X1 U11402 ( .A1(n8922), .A2(n10501), .ZN(n8925) );
  OR2_X1 U11403 ( .A1(n10501), .A2(n8922), .ZN(n8923) );
  NAND2_X1 U11404 ( .A1(n8925), .A2(n8923), .ZN(n10154) );
  XNOR2_X1 U11405 ( .A(n15165), .B(n11886), .ZN(n8926) );
  XNOR2_X1 U11406 ( .A(n8926), .B(n10405), .ZN(n10342) );
  NAND2_X1 U11407 ( .A1(n10341), .A2(n10342), .ZN(n10596) );
  INV_X1 U11408 ( .A(n8926), .ZN(n8927) );
  NAND2_X1 U11409 ( .A1(n8927), .A2(n10405), .ZN(n10594) );
  NAND2_X1 U11410 ( .A1(n10596), .A2(n10594), .ZN(n8930) );
  NAND2_X1 U11411 ( .A1(n8937), .A2(n15182), .ZN(n8928) );
  OAI22_X1 U11412 ( .A1(n8945), .A2(n8928), .B1(n8950), .B2(n8932), .ZN(n8929)
         );
  NOR2_X1 U11413 ( .A1(n8930), .A2(n8931), .ZN(n10586) );
  AOI211_X1 U11414 ( .C1(n8931), .C2(n8930), .A(n12459), .B(n10586), .ZN(n8954) );
  INV_X1 U11415 ( .A(n8932), .ZN(n8936) );
  NAND3_X1 U11416 ( .A1(n8934), .A2(n9492), .A3(n8933), .ZN(n8935) );
  AOI21_X1 U11417 ( .B1(n8950), .B2(n8936), .A(n8935), .ZN(n8939) );
  NAND2_X1 U11418 ( .A1(n8945), .A2(n8937), .ZN(n8938) );
  NAND2_X1 U11419 ( .A1(n8939), .A2(n8938), .ZN(n8940) );
  NAND2_X1 U11420 ( .A1(n8940), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8943) );
  INV_X1 U11421 ( .A(n9784), .ZN(n8941) );
  NAND3_X1 U11422 ( .A1(n8950), .A2(n8941), .A3(n12690), .ZN(n8942) );
  INV_X1 U11423 ( .A(n10409), .ZN(n8944) );
  NOR2_X1 U11424 ( .A1(n12418), .A2(n8944), .ZN(n8953) );
  NAND2_X1 U11425 ( .A1(n8945), .A2(n15137), .ZN(n8947) );
  AND2_X1 U11426 ( .A1(n12690), .A2(n15193), .ZN(n8946) );
  NAND2_X1 U11427 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14987) );
  OAI21_X1 U11428 ( .B1(n12446), .B2(n15171), .A(n14987), .ZN(n8952) );
  INV_X1 U11429 ( .A(n12692), .ZN(n8948) );
  NAND2_X1 U11430 ( .A1(n12690), .A2(n8948), .ZN(n8949) );
  NOR2_X1 U11431 ( .A1(n12454), .A2(n15134), .ZN(n11899) );
  INV_X1 U11432 ( .A(n11899), .ZN(n12442) );
  NAND2_X1 U11433 ( .A1(n12416), .A2(n12990), .ZN(n12368) );
  OAI22_X1 U11434 ( .A1(n10405), .A2(n12442), .B1(n12575), .B2(n12368), .ZN(
        n8951) );
  OR4_X1 U11435 ( .A1(n8954), .A2(n8953), .A3(n8952), .A4(n8951), .ZN(P3_U3179) );
  OR2_X1 U11436 ( .A1(n8955), .A2(n9689), .ZN(n8957) );
  XNOR2_X1 U11437 ( .A(n8957), .B(n8956), .ZN(n14780) );
  NAND2_X2 U11438 ( .A1(n6643), .A2(P2_U3088), .ZN(n11317) );
  OAI222_X1 U11439 ( .A1(P2_U3088), .A2(n14780), .B1(n11317), .B2(n9591), .C1(
        n9593), .C2(n13693), .ZN(P2_U3325) );
  NAND2_X1 U11440 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8958) );
  XNOR2_X1 U11441 ( .A(n8958), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9561) );
  OAI222_X1 U11442 ( .A1(P2_U3088), .A2(n9562), .B1(n11317), .B2(n9036), .C1(
        n8959), .C2(n13693), .ZN(P2_U3326) );
  INV_X2 U11443 ( .A(n13135), .ZN(n11060) );
  OAI222_X1 U11444 ( .A1(n11060), .A2(n8961), .B1(n12350), .B2(n8960), .C1(
        P3_U3151), .C2(n9506), .ZN(P3_U3294) );
  INV_X1 U11445 ( .A(SI_4_), .ZN(n8964) );
  INV_X1 U11446 ( .A(n8962), .ZN(n8963) );
  OAI222_X1 U11447 ( .A1(P3_U3151), .A2(n14955), .B1(n12350), .B2(n8964), .C1(
        n11060), .C2(n8963), .ZN(P3_U3291) );
  OR2_X1 U11448 ( .A1(n8965), .A2(n9689), .ZN(n8966) );
  XNOR2_X1 U11449 ( .A(n8966), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9602) );
  INV_X1 U11450 ( .A(n9602), .ZN(n9114) );
  INV_X1 U11451 ( .A(n9600), .ZN(n9028) );
  OAI222_X1 U11452 ( .A1(P2_U3088), .A2(n9114), .B1(n11317), .B2(n9028), .C1(
        n8967), .C2(n13693), .ZN(P2_U3324) );
  OAI222_X1 U11453 ( .A1(n11060), .A2(n8969), .B1(n12350), .B2(n8968), .C1(
        P3_U3151), .C2(n10701), .ZN(P3_U3287) );
  INV_X1 U11454 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U11455 ( .A1(n8965), .A2(n8970), .ZN(n8973) );
  NAND2_X1 U11456 ( .A1(n8973), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8971) );
  XNOR2_X1 U11457 ( .A(n8971), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9659) );
  INV_X1 U11458 ( .A(n9659), .ZN(n9265) );
  INV_X1 U11459 ( .A(n9658), .ZN(n9034) );
  OAI222_X1 U11460 ( .A1(P2_U3088), .A2(n9265), .B1(n11317), .B2(n9034), .C1(
        n8972), .C2(n13693), .ZN(P2_U3323) );
  NAND2_X1 U11461 ( .A1(n8975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8974) );
  MUX2_X1 U11462 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8974), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8977) );
  INV_X1 U11463 ( .A(n8975), .ZN(n8976) );
  INV_X1 U11464 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n15472) );
  NAND2_X1 U11465 ( .A1(n8976), .A2(n15472), .ZN(n8987) );
  NAND2_X1 U11466 ( .A1(n8977), .A2(n8987), .ZN(n9172) );
  OAI222_X1 U11467 ( .A1(P2_U3088), .A2(n9172), .B1(n11317), .B2(n9665), .C1(
        n8978), .C2(n13693), .ZN(P2_U3322) );
  INV_X1 U11468 ( .A(SI_9_), .ZN(n8981) );
  INV_X1 U11469 ( .A(n8979), .ZN(n8980) );
  OAI222_X1 U11470 ( .A1(P3_U3151), .A2(n15017), .B1(n12350), .B2(n8981), .C1(
        n11060), .C2(n8980), .ZN(P3_U3286) );
  INV_X1 U11471 ( .A(n9924), .ZN(n9223) );
  INV_X1 U11472 ( .A(n8984), .ZN(n8983) );
  NAND2_X1 U11473 ( .A1(n8983), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12260) );
  NAND2_X1 U11474 ( .A1(n9223), .A2(n12260), .ZN(n9003) );
  NAND2_X1 U11475 ( .A1(n12201), .A2(n8984), .ZN(n8985) );
  AND2_X1 U11476 ( .A1(n9003), .A2(n9001), .ZN(n13929) );
  NOR2_X1 U11477 ( .A1(n13929), .A2(P1_U4016), .ZN(P1_U3085) );
  NAND2_X1 U11478 ( .A1(n8987), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8986) );
  MUX2_X1 U11479 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8986), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n8988) );
  INV_X1 U11480 ( .A(n9848), .ZN(n14794) );
  INV_X1 U11481 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n8989) );
  OAI222_X1 U11482 ( .A1(P2_U3088), .A2(n14794), .B1(n11317), .B2(n9847), .C1(
        n8989), .C2(n13693), .ZN(P2_U3321) );
  INV_X1 U11483 ( .A(SI_3_), .ZN(n8992) );
  INV_X1 U11484 ( .A(n8990), .ZN(n8991) );
  OAI222_X1 U11485 ( .A1(P3_U3151), .A2(n6995), .B1(n12350), .B2(n8992), .C1(
        n11060), .C2(n8991), .ZN(P3_U3292) );
  INV_X1 U11486 ( .A(SI_7_), .ZN(n8995) );
  INV_X1 U11487 ( .A(n8993), .ZN(n8994) );
  OAI222_X1 U11488 ( .A1(P3_U3151), .A2(n10689), .B1(n12350), .B2(n8995), .C1(
        n11060), .C2(n8994), .ZN(P3_U3288) );
  OAI222_X1 U11489 ( .A1(n11060), .A2(n8997), .B1(n12350), .B2(n8996), .C1(
        P3_U3151), .C2(n14985), .ZN(P3_U3289) );
  INV_X1 U11490 ( .A(SI_5_), .ZN(n9000) );
  INV_X1 U11491 ( .A(n8998), .ZN(n8999) );
  OAI222_X1 U11492 ( .A1(P3_U3151), .A2(n10385), .B1(n12350), .B2(n9000), .C1(
        n11060), .C2(n8999), .ZN(P3_U3290) );
  INV_X1 U11493 ( .A(n13929), .ZN(n14651) );
  INV_X1 U11494 ( .A(n9001), .ZN(n9002) );
  AND2_X1 U11495 ( .A1(n9003), .A2(n9002), .ZN(n9092) );
  INV_X1 U11496 ( .A(n6843), .ZN(n12256) );
  NAND2_X1 U11497 ( .A1(n12256), .A2(n8349), .ZN(n9004) );
  NAND2_X1 U11498 ( .A1(n9084), .A2(n9004), .ZN(n13845) );
  AOI21_X1 U11499 ( .B1(n6843), .B2(n9005), .A(n13845), .ZN(n9006) );
  XNOR2_X1 U11500 ( .A(n9006), .B(n13844), .ZN(n9007) );
  AOI22_X1 U11501 ( .A1(n9092), .A2(n9007), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9008) );
  OAI21_X1 U11502 ( .B1(n14651), .B2(n7050), .A(n9008), .ZN(P1_U3243) );
  INV_X1 U11503 ( .A(n9523), .ZN(n9543) );
  INV_X1 U11504 ( .A(n9009), .ZN(n9011) );
  INV_X1 U11505 ( .A(SI_2_), .ZN(n9010) );
  OAI222_X1 U11506 ( .A1(n9543), .A2(P3_U3151), .B1(n11060), .B2(n9011), .C1(
        n9010), .C2(n12350), .ZN(P3_U3293) );
  NAND3_X1 U11507 ( .A1(n11968), .A2(n9015), .A3(n11212), .ZN(n9013) );
  OAI21_X1 U11508 ( .B1(n14706), .B2(P1_D_REG_1__SCAN_IN), .A(n9013), .ZN(
        n9014) );
  INV_X1 U11509 ( .A(n9014), .ZN(P1_U3446) );
  NAND2_X1 U11510 ( .A1(n10966), .A2(n9015), .ZN(n9016) );
  OAI22_X1 U11511 ( .A1(n14706), .A2(P1_D_REG_0__SCAN_IN), .B1(n9017), .B2(
        n9016), .ZN(n9018) );
  INV_X1 U11512 ( .A(n9018), .ZN(P1_U3445) );
  INV_X1 U11513 ( .A(n10116), .ZN(n9022) );
  NAND2_X1 U11514 ( .A1(n9038), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9019) );
  XNOR2_X1 U11515 ( .A(n9019), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10117) );
  INV_X1 U11516 ( .A(n10117), .ZN(n9020) );
  OAI222_X1 U11517 ( .A1(n13693), .A2(n9021), .B1(n11317), .B2(n9022), .C1(
        P2_U3088), .C2(n9020), .ZN(P2_U3320) );
  INV_X1 U11518 ( .A(n13910), .ZN(n13899) );
  OAI222_X1 U11519 ( .A1(n14332), .A2(n9023), .B1(n14330), .B2(n9022), .C1(
        P1_U3086), .C2(n13899), .ZN(P1_U3348) );
  INV_X1 U11520 ( .A(n12774), .ZN(n12722) );
  INV_X1 U11521 ( .A(SI_10_), .ZN(n15378) );
  INV_X1 U11522 ( .A(n9024), .ZN(n9025) );
  OAI222_X1 U11523 ( .A1(P3_U3151), .A2(n12722), .B1(n12350), .B2(n15378), 
        .C1(n11060), .C2(n9025), .ZN(P3_U3285) );
  OAI222_X1 U11524 ( .A1(n12350), .A2(n15521), .B1(n11060), .B2(n9026), .C1(
        n15031), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U11525 ( .A(n13869), .ZN(n9029) );
  OAI222_X1 U11526 ( .A1(P1_U3086), .A2(n9029), .B1(n14330), .B2(n9028), .C1(
        n9027), .C2(n14332), .ZN(P1_U3352) );
  OAI222_X1 U11527 ( .A1(P1_U3086), .A2(n13861), .B1(n14330), .B2(n9591), .C1(
        n9030), .C2(n14332), .ZN(P1_U3353) );
  INV_X1 U11528 ( .A(n9137), .ZN(n9204) );
  OAI222_X1 U11529 ( .A1(P1_U3086), .A2(n9204), .B1(n14330), .B2(n9847), .C1(
        n9031), .C2(n14332), .ZN(P1_U3349) );
  INV_X1 U11530 ( .A(n9136), .ZN(n9159) );
  OAI222_X1 U11531 ( .A1(P1_U3086), .A2(n9159), .B1(n14330), .B2(n9665), .C1(
        n9032), .C2(n14332), .ZN(P1_U3350) );
  INV_X1 U11532 ( .A(n9133), .ZN(n13892) );
  OAI222_X1 U11533 ( .A1(P1_U3086), .A2(n13892), .B1(n14330), .B2(n9034), .C1(
        n9033), .C2(n14332), .ZN(P1_U3351) );
  INV_X1 U11534 ( .A(n9130), .ZN(n9102) );
  INV_X1 U11535 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9035) );
  OAI222_X1 U11536 ( .A1(P1_U3086), .A2(n9102), .B1(n14330), .B2(n9036), .C1(
        n9035), .C2(n14332), .ZN(P1_U3354) );
  INV_X1 U11537 ( .A(n10201), .ZN(n9040) );
  INV_X1 U11538 ( .A(n9207), .ZN(n9308) );
  OAI222_X1 U11539 ( .A1(n14332), .A2(n9037), .B1(n14330), .B2(n9040), .C1(
        P1_U3086), .C2(n9308), .ZN(P1_U3347) );
  OAI21_X1 U11540 ( .B1(n9038), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9039) );
  XNOR2_X1 U11541 ( .A(n9039), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10202) );
  INV_X1 U11542 ( .A(n10202), .ZN(n9178) );
  OAI222_X1 U11543 ( .A1(n13693), .A2(n9041), .B1(n11317), .B2(n9040), .C1(
        P2_U3088), .C2(n9178), .ZN(P2_U3319) );
  INV_X1 U11544 ( .A(n9309), .ZN(n13926) );
  INV_X1 U11545 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9042) );
  OAI222_X1 U11546 ( .A1(P1_U3086), .A2(n13926), .B1(n14330), .B2(n10263), 
        .C1(n9042), .C2(n14332), .ZN(P1_U3346) );
  OR2_X1 U11547 ( .A1(n9043), .A2(n9689), .ZN(n9044) );
  XNOR2_X1 U11548 ( .A(n9044), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10264) );
  INV_X1 U11549 ( .A(n10264), .ZN(n9319) );
  OAI222_X1 U11550 ( .A1(P2_U3088), .A2(n9319), .B1(n11317), .B2(n10263), .C1(
        n9045), .C2(n13693), .ZN(P2_U3318) );
  NAND2_X1 U11551 ( .A1(n9052), .A2(n9051), .ZN(n9054) );
  NOR2_X4 U11552 ( .A1(n9054), .A2(n9053), .ZN(n11757) );
  OAI21_X1 U11553 ( .B1(n9572), .B2(n9058), .A(n9601), .ZN(n9059) );
  INV_X1 U11554 ( .A(n9070), .ZN(n9064) );
  AND2_X1 U11555 ( .A1(n9064), .A2(n9061), .ZN(n14779) );
  INV_X1 U11556 ( .A(n9061), .ZN(n9062) );
  NAND2_X1 U11557 ( .A1(n9062), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13687) );
  INV_X1 U11558 ( .A(n13687), .ZN(n9063) );
  AND2_X1 U11559 ( .A1(n9064), .A2(n9063), .ZN(n9076) );
  INV_X1 U11560 ( .A(n13691), .ZN(n11766) );
  INV_X1 U11561 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10147) );
  MUX2_X1 U11562 ( .A(n10147), .B(P2_REG2_REG_1__SCAN_IN), .S(n9561), .Z(
        n14771) );
  INV_X1 U11563 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9464) );
  INV_X1 U11564 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9065) );
  AOI21_X1 U11565 ( .B1(n9561), .B2(P2_REG2_REG_1__SCAN_IN), .A(n14772), .ZN(
        n14788) );
  INV_X1 U11566 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10236) );
  MUX2_X1 U11567 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10236), .S(n14780), .Z(
        n14787) );
  NOR2_X1 U11568 ( .A1(n14780), .A2(n10236), .ZN(n9067) );
  INV_X1 U11569 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9606) );
  MUX2_X1 U11570 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9606), .S(n9602), .Z(n9066)
         );
  OAI21_X1 U11571 ( .B1(n14786), .B2(n9067), .A(n9066), .ZN(n9104) );
  INV_X1 U11572 ( .A(n9104), .ZN(n9069) );
  NOR3_X1 U11573 ( .A1(n14786), .A2(n9067), .A3(n9066), .ZN(n9068) );
  NOR3_X1 U11574 ( .A1(n14811), .A2(n9069), .A3(n9068), .ZN(n9072) );
  AND2_X1 U11575 ( .A1(n9070), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14835) );
  INV_X1 U11576 ( .A(n14835), .ZN(n14823) );
  INV_X1 U11577 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14388) );
  INV_X1 U11578 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n13165) );
  OAI22_X1 U11579 ( .A1(n14823), .A2(n14388), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13165), .ZN(n9071) );
  NOR2_X1 U11580 ( .A1(n9072), .A2(n9071), .ZN(n9081) );
  INV_X1 U11581 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9073) );
  MUX2_X1 U11582 ( .A(n9073), .B(P2_REG1_REG_1__SCAN_IN), .S(n9561), .Z(n14769) );
  NAND2_X1 U11583 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14768) );
  NOR2_X1 U11584 ( .A1(n14769), .A2(n14768), .ZN(n14767) );
  AOI21_X1 U11585 ( .B1(n9561), .B2(P2_REG1_REG_1__SCAN_IN), .A(n14767), .ZN(
        n14784) );
  INV_X1 U11586 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n14926) );
  MUX2_X1 U11587 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n14926), .S(n14780), .Z(
        n14783) );
  NOR2_X1 U11588 ( .A1(n14784), .A2(n14783), .ZN(n14782) );
  INV_X1 U11589 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9637) );
  MUX2_X1 U11590 ( .A(n9637), .B(P2_REG1_REG_3__SCAN_IN), .S(n9602), .Z(n9075)
         );
  NOR2_X1 U11591 ( .A1(n14780), .A2(n14926), .ZN(n9078) );
  INV_X1 U11592 ( .A(n9078), .ZN(n9074) );
  NAND2_X1 U11593 ( .A1(n9075), .A2(n9074), .ZN(n9079) );
  MUX2_X1 U11594 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9637), .S(n9602), .Z(n9077)
         );
  OAI21_X1 U11595 ( .B1(n14782), .B2(n9078), .A(n9077), .ZN(n9113) );
  OAI211_X1 U11596 ( .C1(n14782), .C2(n9079), .A(n14843), .B(n9113), .ZN(n9080) );
  OAI211_X1 U11597 ( .C1(n14765), .C2(n9114), .A(n9081), .B(n9080), .ZN(
        P2_U3217) );
  OAI222_X1 U11598 ( .A1(P3_U3151), .A2(n15051), .B1(n12350), .B2(n9083), .C1(
        n11060), .C2(n9082), .ZN(P3_U3283) );
  INV_X1 U11599 ( .A(n9092), .ZN(n9085) );
  OR2_X1 U11600 ( .A1(n9085), .A2(n9084), .ZN(n14647) );
  AND2_X1 U11601 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9087) );
  INV_X1 U11602 ( .A(n9087), .ZN(n13843) );
  MUX2_X1 U11603 ( .A(n9086), .B(P1_REG2_REG_1__SCAN_IN), .S(n9130), .Z(n9091)
         );
  MUX2_X1 U11604 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9086), .S(n9130), .Z(n9088)
         );
  NAND2_X1 U11605 ( .A1(n9088), .A2(n9087), .ZN(n13855) );
  INV_X1 U11606 ( .A(n13855), .ZN(n9090) );
  NOR2_X1 U11607 ( .A1(n8816), .A2(n6843), .ZN(n9089) );
  AOI211_X1 U11608 ( .C1(n13843), .C2(n9091), .A(n9090), .B(n14645), .ZN(n9099) );
  MUX2_X1 U11609 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9093), .S(n9130), .Z(n9095)
         );
  AND2_X1 U11610 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9094) );
  NAND2_X1 U11611 ( .A1(n9095), .A2(n9094), .ZN(n13851) );
  MUX2_X1 U11612 ( .A(n9093), .B(P1_REG1_REG_1__SCAN_IN), .S(n9130), .Z(n9096)
         );
  OAI21_X1 U11613 ( .B1(n9005), .B2(n13844), .A(n9096), .ZN(n9097) );
  AND3_X1 U11614 ( .A1(n13966), .A2(n13851), .A3(n9097), .ZN(n9098) );
  NOR2_X1 U11615 ( .A1(n9099), .A2(n9098), .ZN(n9101) );
  AOI22_X1 U11616 ( .A1(n13929), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9100) );
  OAI211_X1 U11617 ( .C1(n9102), .C2(n14647), .A(n9101), .B(n9100), .ZN(
        P1_U3244) );
  INV_X1 U11618 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11619 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10129) );
  OAI21_X1 U11620 ( .B1(n14823), .B2(n9103), .A(n10129), .ZN(n9112) );
  INV_X1 U11621 ( .A(n9172), .ZN(n9666) );
  OAI21_X1 U11622 ( .B1(n9606), .B2(n9114), .A(n9104), .ZN(n9259) );
  INV_X1 U11623 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9619) );
  MUX2_X1 U11624 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9619), .S(n9659), .Z(n9258)
         );
  NAND2_X1 U11625 ( .A1(n9259), .A2(n9258), .ZN(n9257) );
  NAND2_X1 U11626 ( .A1(n9659), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9161) );
  INV_X1 U11627 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9105) );
  MUX2_X1 U11628 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9105), .S(n9172), .Z(n9160)
         );
  AOI21_X1 U11629 ( .B1(n9257), .B2(n9161), .A(n9160), .ZN(n9163) );
  AOI21_X1 U11630 ( .B1(n9666), .B2(P2_REG2_REG_5__SCAN_IN), .A(n9163), .ZN(
        n14804) );
  INV_X1 U11631 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9106) );
  MUX2_X1 U11632 ( .A(n9106), .B(P2_REG2_REG_6__SCAN_IN), .S(n9848), .Z(n14803) );
  NOR2_X1 U11633 ( .A1(n14794), .A2(n9106), .ZN(n9108) );
  INV_X1 U11634 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10176) );
  MUX2_X1 U11635 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10176), .S(n10117), .Z(
        n9107) );
  OAI21_X1 U11636 ( .B1(n14802), .B2(n9108), .A(n9107), .ZN(n9176) );
  INV_X1 U11637 ( .A(n9176), .ZN(n9110) );
  NOR3_X1 U11638 ( .A1(n14802), .A2(n9108), .A3(n9107), .ZN(n9109) );
  NOR3_X1 U11639 ( .A1(n9110), .A2(n9109), .A3(n14811), .ZN(n9111) );
  AOI211_X1 U11640 ( .C1(n14841), .C2(n10117), .A(n9112), .B(n9111), .ZN(n9121) );
  OAI21_X1 U11641 ( .B1(n9637), .B2(n9114), .A(n9113), .ZN(n9256) );
  INV_X1 U11642 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15327) );
  MUX2_X1 U11643 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15327), .S(n9659), .Z(n9255) );
  NAND2_X1 U11644 ( .A1(n9256), .A2(n9255), .ZN(n9254) );
  NAND2_X1 U11645 ( .A1(n9659), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9167) );
  INV_X1 U11646 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14929) );
  MUX2_X1 U11647 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n14929), .S(n9172), .Z(n9166) );
  AOI21_X1 U11648 ( .B1(n9254), .B2(n9167), .A(n9166), .ZN(n9165) );
  AOI21_X1 U11649 ( .B1(n9666), .B2(P2_REG1_REG_5__SCAN_IN), .A(n9165), .ZN(
        n14800) );
  INV_X1 U11650 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14931) );
  MUX2_X1 U11651 ( .A(n14931), .B(P2_REG1_REG_6__SCAN_IN), .S(n9848), .Z(
        n14799) );
  NOR2_X1 U11652 ( .A1(n14800), .A2(n14799), .ZN(n14797) );
  NOR2_X1 U11653 ( .A1(n14794), .A2(n14931), .ZN(n9118) );
  INV_X1 U11654 ( .A(n9118), .ZN(n9116) );
  INV_X1 U11655 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n14933) );
  MUX2_X1 U11656 ( .A(n14933), .B(P2_REG1_REG_7__SCAN_IN), .S(n10117), .Z(
        n9115) );
  NAND2_X1 U11657 ( .A1(n9116), .A2(n9115), .ZN(n9119) );
  MUX2_X1 U11658 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n14933), .S(n10117), .Z(
        n9117) );
  OAI21_X1 U11659 ( .B1(n14797), .B2(n9118), .A(n9117), .ZN(n9182) );
  OAI211_X1 U11660 ( .C1(n14797), .C2(n9119), .A(n9182), .B(n14843), .ZN(n9120) );
  NAND2_X1 U11661 ( .A1(n9121), .A2(n9120), .ZN(P2_U3221) );
  MUX2_X1 U11662 ( .A(n9122), .B(P1_REG1_REG_2__SCAN_IN), .S(n13861), .Z(n9124) );
  NAND2_X1 U11663 ( .A1(n9130), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n13850) );
  NAND2_X1 U11664 ( .A1(n13851), .A2(n13850), .ZN(n9123) );
  AND2_X1 U11665 ( .A1(n9124), .A2(n9123), .ZN(n13849) );
  NOR2_X1 U11666 ( .A1(n13861), .A2(n9122), .ZN(n13868) );
  MUX2_X1 U11667 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9125), .S(n13869), .Z(n9126) );
  OAI21_X1 U11668 ( .B1(n13849), .B2(n13868), .A(n9126), .ZN(n13883) );
  NAND2_X1 U11669 ( .A1(n13869), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13882) );
  MUX2_X1 U11670 ( .A(n8399), .B(P1_REG1_REG_4__SCAN_IN), .S(n9133), .Z(n13881) );
  AOI21_X1 U11671 ( .B1(n13883), .B2(n13882), .A(n13881), .ZN(n13885) );
  AOI21_X1 U11672 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9133), .A(n13885), .ZN(
        n9147) );
  MUX2_X1 U11673 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n8412), .S(n9136), .Z(n9148)
         );
  NAND2_X1 U11674 ( .A1(n9147), .A2(n9148), .ZN(n9146) );
  OAI21_X1 U11675 ( .B1(n9136), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9146), .ZN(
        n9128) );
  MUX2_X1 U11676 ( .A(n9198), .B(P1_REG1_REG_6__SCAN_IN), .S(n9137), .Z(n9127)
         );
  NOR2_X1 U11677 ( .A1(n9128), .A2(n9127), .ZN(n13908) );
  AOI211_X1 U11678 ( .C1(n9128), .C2(n9127), .A(n13908), .B(n14643), .ZN(n9142) );
  MUX2_X1 U11679 ( .A(n9129), .B(P1_REG2_REG_2__SCAN_IN), .S(n13861), .Z(n9132) );
  NAND2_X1 U11680 ( .A1(n9130), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n13854) );
  NAND2_X1 U11681 ( .A1(n13855), .A2(n13854), .ZN(n9131) );
  AND2_X1 U11682 ( .A1(n9132), .A2(n9131), .ZN(n13875) );
  NOR2_X1 U11683 ( .A1(n13861), .A2(n9129), .ZN(n13874) );
  MUX2_X1 U11684 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9966), .S(n13869), .Z(
        n13876) );
  OAI21_X1 U11685 ( .B1(n13875), .B2(n13874), .A(n13876), .ZN(n13888) );
  NAND2_X1 U11686 ( .A1(n13869), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13887) );
  MUX2_X1 U11687 ( .A(n9134), .B(P1_REG2_REG_4__SCAN_IN), .S(n9133), .Z(n13886) );
  AOI21_X1 U11688 ( .B1(n13888), .B2(n13887), .A(n13886), .ZN(n13890) );
  NOR2_X1 U11689 ( .A1(n13892), .A2(n9134), .ZN(n9151) );
  MUX2_X1 U11690 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9135), .S(n9136), .Z(n9150)
         );
  OAI21_X1 U11691 ( .B1(n13890), .B2(n9151), .A(n9150), .ZN(n9149) );
  NAND2_X1 U11692 ( .A1(n9136), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9139) );
  MUX2_X1 U11693 ( .A(n10061), .B(P1_REG2_REG_6__SCAN_IN), .S(n9137), .Z(n9138) );
  AOI21_X1 U11694 ( .B1(n9149), .B2(n9139), .A(n9138), .ZN(n13915) );
  AND3_X1 U11695 ( .A1(n9149), .A2(n9139), .A3(n9138), .ZN(n9140) );
  NOR3_X1 U11696 ( .A1(n14645), .A2(n13915), .A3(n9140), .ZN(n9141) );
  NOR2_X1 U11697 ( .A1(n9142), .A2(n9141), .ZN(n9145) );
  INV_X1 U11698 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9143) );
  NOR2_X1 U11699 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9143), .ZN(n10043) );
  AOI21_X1 U11700 ( .B1(n13929), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10043), .ZN(
        n9144) );
  OAI211_X1 U11701 ( .C1(n9204), .C2(n14647), .A(n9145), .B(n9144), .ZN(
        P1_U3249) );
  OAI21_X1 U11702 ( .B1(n9148), .B2(n9147), .A(n9146), .ZN(n9155) );
  INV_X1 U11703 ( .A(n9149), .ZN(n9153) );
  NOR3_X1 U11704 ( .A1(n13890), .A2(n9151), .A3(n9150), .ZN(n9152) );
  NOR3_X1 U11705 ( .A1(n14645), .A2(n9153), .A3(n9152), .ZN(n9154) );
  AOI21_X1 U11706 ( .B1(n13966), .B2(n9155), .A(n9154), .ZN(n9158) );
  NOR2_X1 U11707 ( .A1(n9156), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9879) );
  AOI21_X1 U11708 ( .B1(n13929), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9879), .ZN(
        n9157) );
  OAI211_X1 U11709 ( .C1(n9159), .C2(n14647), .A(n9158), .B(n9157), .ZN(
        P1_U3248) );
  NOR2_X1 U11710 ( .A1(n9642), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9686) );
  AND3_X1 U11711 ( .A1(n9257), .A2(n9161), .A3(n9160), .ZN(n9162) );
  NOR3_X1 U11712 ( .A1(n14811), .A2(n9163), .A3(n9162), .ZN(n9164) );
  AOI211_X1 U11713 ( .C1(n14835), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n9686), .B(
        n9164), .ZN(n9171) );
  INV_X1 U11714 ( .A(n9165), .ZN(n9169) );
  NAND3_X1 U11715 ( .A1(n9254), .A2(n9167), .A3(n9166), .ZN(n9168) );
  NAND3_X1 U11716 ( .A1(n14843), .A2(n9169), .A3(n9168), .ZN(n9170) );
  OAI211_X1 U11717 ( .C1(n14765), .C2(n9172), .A(n9171), .B(n9170), .ZN(
        P2_U3219) );
  NAND2_X1 U11718 ( .A1(n10117), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9175) );
  INV_X1 U11719 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9173) );
  MUX2_X1 U11720 ( .A(n9173), .B(P2_REG2_REG_8__SCAN_IN), .S(n10202), .Z(n9174) );
  AOI21_X1 U11721 ( .B1(n9176), .B2(n9175), .A(n9174), .ZN(n9238) );
  NAND3_X1 U11722 ( .A1(n9176), .A2(n9175), .A3(n9174), .ZN(n9177) );
  INV_X1 U11723 ( .A(n14811), .ZN(n14837) );
  NAND2_X1 U11724 ( .A1(n9177), .A2(n14837), .ZN(n9187) );
  NOR2_X1 U11725 ( .A1(n10120), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10220) );
  NOR2_X1 U11726 ( .A1(n14765), .A2(n9178), .ZN(n9179) );
  AOI211_X1 U11727 ( .C1(n14835), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10220), .B(
        n9179), .ZN(n9186) );
  NAND2_X1 U11728 ( .A1(n10117), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9181) );
  INV_X1 U11729 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14935) );
  MUX2_X1 U11730 ( .A(n14935), .B(P2_REG1_REG_8__SCAN_IN), .S(n10202), .Z(
        n9180) );
  AOI21_X1 U11731 ( .B1(n9182), .B2(n9181), .A(n9180), .ZN(n9239) );
  INV_X1 U11732 ( .A(n9239), .ZN(n9184) );
  NAND3_X1 U11733 ( .A1(n9182), .A2(n9181), .A3(n9180), .ZN(n9183) );
  NAND3_X1 U11734 ( .A1(n9184), .A2(n14843), .A3(n9183), .ZN(n9185) );
  OAI211_X1 U11735 ( .C1(n9238), .C2(n9187), .A(n9186), .B(n9185), .ZN(
        P2_U3222) );
  INV_X1 U11736 ( .A(n10351), .ZN(n9195) );
  NAND2_X1 U11737 ( .A1(n9043), .A2(n9188), .ZN(n9189) );
  NOR2_X1 U11738 ( .A1(n9189), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n9335) );
  INV_X1 U11739 ( .A(n9335), .ZN(n9192) );
  NAND2_X1 U11740 ( .A1(n9189), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9190) );
  MUX2_X1 U11741 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9190), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n9191) );
  INV_X1 U11742 ( .A(n14816), .ZN(n9193) );
  OAI222_X1 U11743 ( .A1(n13693), .A2(n9194), .B1(n11317), .B2(n9195), .C1(
        P2_U3088), .C2(n9193), .ZN(P2_U3317) );
  INV_X1 U11744 ( .A(n9404), .ZN(n9398) );
  OAI222_X1 U11745 ( .A1(n14332), .A2(n9196), .B1(n14330), .B2(n9195), .C1(
        P1_U3086), .C2(n9398), .ZN(P1_U3345) );
  MUX2_X1 U11746 ( .A(n9197), .B(P1_REG1_REG_8__SCAN_IN), .S(n9207), .Z(n9201)
         );
  INV_X1 U11747 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n13903) );
  NOR2_X1 U11748 ( .A1(n9204), .A2(n9198), .ZN(n13902) );
  MUX2_X1 U11749 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n13903), .S(n13910), .Z(
        n9199) );
  OAI21_X1 U11750 ( .B1(n13908), .B2(n13902), .A(n9199), .ZN(n13906) );
  OAI21_X1 U11751 ( .B1(n13903), .B2(n13899), .A(n13906), .ZN(n9200) );
  NOR2_X1 U11752 ( .A1(n9200), .A2(n9201), .ZN(n13922) );
  AOI21_X1 U11753 ( .B1(n9201), .B2(n9200), .A(n13922), .ZN(n9214) );
  NOR2_X1 U11754 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8459), .ZN(n9203) );
  NOR2_X1 U11755 ( .A1(n14647), .A2(n9308), .ZN(n9202) );
  AOI211_X1 U11756 ( .C1(n13929), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9203), .B(
        n9202), .ZN(n9213) );
  NOR2_X1 U11757 ( .A1(n9204), .A2(n10061), .ZN(n13909) );
  MUX2_X1 U11758 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9205), .S(n13910), .Z(n9206) );
  OAI21_X1 U11759 ( .B1(n13915), .B2(n13909), .A(n9206), .ZN(n13913) );
  NAND2_X1 U11760 ( .A1(n13910), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9209) );
  MUX2_X1 U11761 ( .A(n9307), .B(P1_REG2_REG_8__SCAN_IN), .S(n9207), .Z(n9208)
         );
  AOI21_X1 U11762 ( .B1(n13913), .B2(n9209), .A(n9208), .ZN(n13932) );
  INV_X1 U11763 ( .A(n13932), .ZN(n9211) );
  NAND3_X1 U11764 ( .A1(n13913), .A2(n9209), .A3(n9208), .ZN(n9210) );
  NAND3_X1 U11765 ( .A1(n9211), .A2(n13963), .A3(n9210), .ZN(n9212) );
  OAI211_X1 U11766 ( .C1(n9214), .C2(n14643), .A(n9213), .B(n9212), .ZN(
        P1_U3251) );
  INV_X1 U11767 ( .A(n10515), .ZN(n9217) );
  INV_X1 U11768 ( .A(n13945), .ZN(n9405) );
  OAI222_X1 U11769 ( .A1(n14332), .A2(n9215), .B1(n14330), .B2(n9217), .C1(
        P1_U3086), .C2(n9405), .ZN(P1_U3344) );
  OR2_X1 U11770 ( .A1(n9335), .A2(n9689), .ZN(n9216) );
  XNOR2_X1 U11771 ( .A(n9216), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10516) );
  INV_X1 U11772 ( .A(n10516), .ZN(n9831) );
  OAI222_X1 U11773 ( .A1(n13693), .A2(n9218), .B1(n11317), .B2(n9217), .C1(
        P2_U3088), .C2(n9831), .ZN(P2_U3316) );
  NOR2_X1 U11774 ( .A1(n9918), .A2(n9917), .ZN(n9232) );
  NAND2_X1 U11775 ( .A1(n9232), .A2(n9219), .ZN(n9224) );
  AND2_X1 U11776 ( .A1(n9224), .A2(n9922), .ZN(n9390) );
  INV_X1 U11777 ( .A(n9390), .ZN(n9220) );
  AND2_X1 U11778 ( .A1(n9220), .A2(n9924), .ZN(n10616) );
  INV_X1 U11779 ( .A(n14602), .ZN(n13792) );
  INV_X1 U11780 ( .A(n12201), .ZN(n9221) );
  NAND2_X1 U11781 ( .A1(n14731), .A2(n9221), .ZN(n9222) );
  NAND2_X1 U11782 ( .A1(n13841), .A2(n11811), .ZN(n9227) );
  INV_X1 U11783 ( .A(n9225), .ZN(n9228) );
  AOI22_X1 U11784 ( .A1(n9345), .A2(n9995), .B1(n9228), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9226) );
  AND2_X1 U11785 ( .A1(n9227), .A2(n9226), .ZN(n9231) );
  NAND2_X1 U11786 ( .A1(n13841), .A2(n9345), .ZN(n9230) );
  AOI22_X1 U11787 ( .A1(n9346), .A2(n9995), .B1(n9228), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U11788 ( .A1(n9230), .A2(n9229), .ZN(n9342) );
  NAND2_X1 U11789 ( .A1(n9231), .A2(n9342), .ZN(n9343) );
  OAI21_X1 U11790 ( .B1(n9231), .B2(n9342), .A(n9343), .ZN(n13842) );
  NAND2_X1 U11791 ( .A1(n9232), .A2(n9921), .ZN(n13808) );
  NOR2_X1 U11792 ( .A1(n13808), .A2(n14260), .ZN(n13797) );
  AOI22_X1 U11793 ( .A1(n14585), .A2(n13842), .B1(n13797), .B2(n9350), .ZN(
        n9235) );
  NAND2_X1 U11794 ( .A1(n10616), .A2(n9233), .ZN(n11964) );
  NAND2_X1 U11795 ( .A1(n11964), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9234) );
  OAI211_X1 U11796 ( .C1(n13792), .C2(n9932), .A(n9235), .B(n9234), .ZN(
        P1_U3232) );
  OAI222_X1 U11797 ( .A1(P3_U3151), .A2(n15071), .B1(n12350), .B2(n9237), .C1(
        n11060), .C2(n9236), .ZN(P3_U3282) );
  AOI21_X1 U11798 ( .B1(n10202), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9238), .ZN(
        n9244) );
  INV_X1 U11799 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9242) );
  NOR3_X1 U11800 ( .A1(n9244), .A2(n9242), .A3(n14811), .ZN(n9241) );
  AOI21_X1 U11801 ( .B1(n10202), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9239), .ZN(
        n9249) );
  INV_X1 U11802 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n14937) );
  NOR3_X1 U11803 ( .A1(n9249), .A2(n14937), .A3(n14798), .ZN(n9240) );
  NOR3_X1 U11804 ( .A1(n9241), .A2(n14841), .A3(n9240), .ZN(n9253) );
  NAND2_X1 U11805 ( .A1(n9319), .A2(n9242), .ZN(n9324) );
  MUX2_X1 U11806 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9242), .S(n10264), .Z(n9243) );
  NAND2_X1 U11807 ( .A1(n9244), .A2(n9243), .ZN(n9325) );
  OAI21_X1 U11808 ( .B1(n9244), .B2(n9324), .A(n9325), .ZN(n9247) );
  INV_X1 U11809 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9245) );
  NAND2_X1 U11810 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10335) );
  OAI21_X1 U11811 ( .B1(n14823), .B2(n9245), .A(n10335), .ZN(n9246) );
  AOI21_X1 U11812 ( .B1(n9247), .B2(n14837), .A(n9246), .ZN(n9252) );
  NOR3_X1 U11813 ( .A1(n9249), .A2(n10264), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n9250) );
  MUX2_X1 U11814 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14937), .S(n10264), .Z(
        n9248) );
  AND2_X1 U11815 ( .A1(n9249), .A2(n9248), .ZN(n9318) );
  OAI21_X1 U11816 ( .B1(n9250), .B2(n9318), .A(n14843), .ZN(n9251) );
  OAI211_X1 U11817 ( .C1(n9253), .C2(n9319), .A(n9252), .B(n9251), .ZN(
        P2_U3223) );
  OAI211_X1 U11818 ( .C1(n9256), .C2(n9255), .A(n14843), .B(n9254), .ZN(n9261)
         );
  OAI211_X1 U11819 ( .C1(n9259), .C2(n9258), .A(n14837), .B(n9257), .ZN(n9260)
         );
  NAND2_X1 U11820 ( .A1(n9261), .A2(n9260), .ZN(n9263) );
  NAND2_X1 U11821 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n9825) );
  INV_X1 U11822 ( .A(n9825), .ZN(n9262) );
  AOI211_X1 U11823 ( .C1(n14835), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n9263), .B(
        n9262), .ZN(n9264) );
  OAI21_X1 U11824 ( .B1(n9265), .B2(n14765), .A(n9264), .ZN(P2_U3218) );
  AOI22_X1 U11825 ( .A1(n14837), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n14843), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n9268) );
  OAI21_X1 U11826 ( .B1(n14798), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14765), .ZN(
        n9266) );
  AOI21_X1 U11827 ( .B1(n14837), .B2(n9464), .A(n9266), .ZN(n9267) );
  MUX2_X1 U11828 ( .A(n9268), .B(n9267), .S(P2_IR_REG_0__SCAN_IN), .Z(n9270)
         );
  AOI22_X1 U11829 ( .A1(n14835), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9269) );
  NAND2_X1 U11830 ( .A1(n9270), .A2(n9269), .ZN(P2_U3214) );
  INV_X1 U11831 ( .A(n9271), .ZN(n9272) );
  CLKBUF_X1 U11832 ( .A(n9277), .Z(n9298) );
  INV_X1 U11833 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9273) );
  NOR2_X1 U11834 ( .A1(n9298), .A2(n9273), .ZN(P3_U3256) );
  INV_X1 U11835 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9274) );
  NOR2_X1 U11836 ( .A1(n9298), .A2(n9274), .ZN(P3_U3257) );
  INV_X1 U11837 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9275) );
  NOR2_X1 U11838 ( .A1(n9298), .A2(n9275), .ZN(P3_U3261) );
  INV_X1 U11839 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9276) );
  NOR2_X1 U11840 ( .A1(n9298), .A2(n9276), .ZN(P3_U3259) );
  INV_X1 U11841 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n15393) );
  NOR2_X1 U11842 ( .A1(n9298), .A2(n15393), .ZN(P3_U3263) );
  INV_X1 U11843 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9278) );
  NOR2_X1 U11844 ( .A1(n9298), .A2(n9278), .ZN(P3_U3244) );
  INV_X1 U11845 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9279) );
  NOR2_X1 U11846 ( .A1(n9277), .A2(n9279), .ZN(P3_U3262) );
  INV_X1 U11847 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9280) );
  NOR2_X1 U11848 ( .A1(n9298), .A2(n9280), .ZN(P3_U3246) );
  INV_X1 U11849 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n15382) );
  NOR2_X1 U11850 ( .A1(n9277), .A2(n15382), .ZN(P3_U3234) );
  INV_X1 U11851 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9281) );
  NOR2_X1 U11852 ( .A1(n9277), .A2(n9281), .ZN(P3_U3235) );
  INV_X1 U11853 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n15482) );
  NOR2_X1 U11854 ( .A1(n9277), .A2(n15482), .ZN(P3_U3236) );
  INV_X1 U11855 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9282) );
  NOR2_X1 U11856 ( .A1(n9277), .A2(n9282), .ZN(P3_U3237) );
  INV_X1 U11857 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9283) );
  NOR2_X1 U11858 ( .A1(n9277), .A2(n9283), .ZN(P3_U3238) );
  INV_X1 U11859 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9284) );
  NOR2_X1 U11860 ( .A1(n9277), .A2(n9284), .ZN(P3_U3239) );
  INV_X1 U11861 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9285) );
  NOR2_X1 U11862 ( .A1(n9298), .A2(n9285), .ZN(P3_U3253) );
  INV_X1 U11863 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n15339) );
  NOR2_X1 U11864 ( .A1(n9277), .A2(n15339), .ZN(P3_U3258) );
  INV_X1 U11865 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9286) );
  NOR2_X1 U11866 ( .A1(n9298), .A2(n9286), .ZN(P3_U3255) );
  INV_X1 U11867 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9287) );
  NOR2_X1 U11868 ( .A1(n9298), .A2(n9287), .ZN(P3_U3252) );
  INV_X1 U11869 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9288) );
  NOR2_X1 U11870 ( .A1(n9277), .A2(n9288), .ZN(P3_U3240) );
  INV_X1 U11871 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9289) );
  NOR2_X1 U11872 ( .A1(n9277), .A2(n9289), .ZN(P3_U3241) );
  INV_X1 U11873 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9290) );
  NOR2_X1 U11874 ( .A1(n9277), .A2(n9290), .ZN(P3_U3242) );
  INV_X1 U11875 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9291) );
  NOR2_X1 U11876 ( .A1(n9298), .A2(n9291), .ZN(P3_U3260) );
  INV_X1 U11877 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9292) );
  NOR2_X1 U11878 ( .A1(n9298), .A2(n9292), .ZN(P3_U3249) );
  INV_X1 U11879 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9293) );
  NOR2_X1 U11880 ( .A1(n9298), .A2(n9293), .ZN(P3_U3245) );
  INV_X1 U11881 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n15483) );
  NOR2_X1 U11882 ( .A1(n9298), .A2(n15483), .ZN(P3_U3251) );
  INV_X1 U11883 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9294) );
  NOR2_X1 U11884 ( .A1(n9298), .A2(n9294), .ZN(P3_U3247) );
  INV_X1 U11885 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9295) );
  NOR2_X1 U11886 ( .A1(n9298), .A2(n9295), .ZN(P3_U3248) );
  INV_X1 U11887 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9296) );
  NOR2_X1 U11888 ( .A1(n9298), .A2(n9296), .ZN(P3_U3254) );
  INV_X1 U11889 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9297) );
  NOR2_X1 U11890 ( .A1(n9298), .A2(n9297), .ZN(P3_U3250) );
  INV_X1 U11891 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n15495) );
  NOR2_X1 U11892 ( .A1(n9298), .A2(n15495), .ZN(P3_U3243) );
  INV_X1 U11893 ( .A(n12023), .ZN(n9926) );
  NOR2_X1 U11894 ( .A1(n14752), .A2(n14144), .ZN(n9300) );
  NAND2_X1 U11895 ( .A1(n13841), .A2(n9932), .ZN(n12030) );
  NAND2_X1 U11896 ( .A1(n12032), .A2(n12030), .ZN(n12210) );
  INV_X1 U11897 ( .A(n12210), .ZN(n9299) );
  OAI222_X1 U11898 ( .A1(n9932), .A2(n9926), .B1(n9300), .B2(n9299), .C1(
        n14260), .C2(n11962), .ZN(n9302) );
  NAND2_X1 U11899 ( .A1(n9302), .A2(n14764), .ZN(n9301) );
  OAI21_X1 U11900 ( .B1(n14764), .B2(n9005), .A(n9301), .ZN(P1_U3528) );
  INV_X1 U11901 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U11902 ( .A1(n9302), .A2(n14755), .ZN(n9303) );
  OAI21_X1 U11903 ( .B1(n14755), .B2(n9304), .A(n9303), .ZN(P1_U3459) );
  AND2_X1 U11904 ( .A1(n9308), .A2(n9197), .ZN(n13920) );
  MUX2_X1 U11905 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n8478), .S(n9309), .Z(n13921) );
  OAI21_X1 U11906 ( .B1(n13922), .B2(n13920), .A(n13921), .ZN(n13919) );
  OAI21_X1 U11907 ( .B1(n9309), .B2(P1_REG1_REG_9__SCAN_IN), .A(n13919), .ZN(
        n9306) );
  INV_X1 U11908 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14762) );
  MUX2_X1 U11909 ( .A(n14762), .B(P1_REG1_REG_10__SCAN_IN), .S(n9404), .Z(
        n9305) );
  NOR2_X1 U11910 ( .A1(n9306), .A2(n9305), .ZN(n9403) );
  AOI211_X1 U11911 ( .C1(n9306), .C2(n9305), .A(n14643), .B(n9403), .ZN(n9317)
         );
  NOR2_X1 U11912 ( .A1(n9308), .A2(n9307), .ZN(n13931) );
  MUX2_X1 U11913 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n14667), .S(n9309), .Z(
        n13930) );
  OAI21_X1 U11914 ( .B1(n13932), .B2(n13931), .A(n13930), .ZN(n13934) );
  NAND2_X1 U11915 ( .A1(n9309), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9311) );
  MUX2_X1 U11916 ( .A(n10309), .B(P1_REG2_REG_10__SCAN_IN), .S(n9404), .Z(
        n9310) );
  AOI21_X1 U11917 ( .B1(n13934), .B2(n9311), .A(n9310), .ZN(n13950) );
  INV_X1 U11918 ( .A(n13950), .ZN(n9313) );
  NAND3_X1 U11919 ( .A1(n13934), .A2(n9311), .A3(n9310), .ZN(n9312) );
  NAND3_X1 U11920 ( .A1(n9313), .A2(n13963), .A3(n9312), .ZN(n9315) );
  AOI22_X1 U11921 ( .A1(n13929), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(
        P1_REG3_REG_10__SCAN_IN), .B2(P1_U3086), .ZN(n9314) );
  OAI211_X1 U11922 ( .C1(n14647), .C2(n9398), .A(n9315), .B(n9314), .ZN(n9316)
         );
  OR2_X1 U11923 ( .A1(n9317), .A2(n9316), .ZN(P1_U3253) );
  AOI21_X1 U11924 ( .B1(n14937), .B2(n9319), .A(n9318), .ZN(n14819) );
  INV_X1 U11925 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9320) );
  MUX2_X1 U11926 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9320), .S(n14816), .Z(
        n14818) );
  NAND2_X1 U11927 ( .A1(n14819), .A2(n14818), .ZN(n14817) );
  NAND2_X1 U11928 ( .A1(n14816), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9322) );
  INV_X1 U11929 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14941) );
  MUX2_X1 U11930 ( .A(n14941), .B(P2_REG1_REG_11__SCAN_IN), .S(n10516), .Z(
        n9321) );
  AOI21_X1 U11931 ( .B1(n14817), .B2(n9322), .A(n9321), .ZN(n9835) );
  NAND3_X1 U11932 ( .A1(n14817), .A2(n9322), .A3(n9321), .ZN(n9323) );
  NAND2_X1 U11933 ( .A1(n9323), .A2(n14843), .ZN(n9333) );
  NAND2_X1 U11934 ( .A1(n9325), .A2(n9324), .ZN(n14813) );
  INV_X1 U11935 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9326) );
  MUX2_X1 U11936 ( .A(n9326), .B(P2_REG2_REG_10__SCAN_IN), .S(n14816), .Z(
        n14812) );
  AOI21_X1 U11937 ( .B1(n14816), .B2(P2_REG2_REG_10__SCAN_IN), .A(n14810), 
        .ZN(n9328) );
  INV_X1 U11938 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9830) );
  MUX2_X1 U11939 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9830), .S(n10516), .Z(
        n9327) );
  NAND2_X1 U11940 ( .A1(n9328), .A2(n9327), .ZN(n13312) );
  OAI21_X1 U11941 ( .B1(n9328), .B2(n9327), .A(n13312), .ZN(n9329) );
  NAND2_X1 U11942 ( .A1(n9329), .A2(n14837), .ZN(n9332) );
  INV_X1 U11943 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14414) );
  NAND2_X1 U11944 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10658)
         );
  OAI21_X1 U11945 ( .B1(n14823), .B2(n14414), .A(n10658), .ZN(n9330) );
  AOI21_X1 U11946 ( .B1(n10516), .B2(n14841), .A(n9330), .ZN(n9331) );
  OAI211_X1 U11947 ( .C1(n9835), .C2(n9333), .A(n9332), .B(n9331), .ZN(
        P2_U3225) );
  INV_X1 U11948 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9337) );
  INV_X1 U11949 ( .A(n10749), .ZN(n9338) );
  NAND2_X1 U11950 ( .A1(n9335), .A2(n9334), .ZN(n9365) );
  NAND2_X1 U11951 ( .A1(n9365), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9336) );
  XNOR2_X1 U11952 ( .A(n9336), .B(P2_IR_REG_12__SCAN_IN), .ZN(n13309) );
  INV_X1 U11953 ( .A(n13309), .ZN(n9836) );
  OAI222_X1 U11954 ( .A1(n13693), .A2(n9337), .B1(n11317), .B2(n9338), .C1(
        n9836), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U11955 ( .A(n9406), .ZN(n9481) );
  OAI222_X1 U11956 ( .A1(n14332), .A2(n9339), .B1(n14330), .B2(n9338), .C1(
        n9481), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U11957 ( .A(n12751), .ZN(n15091) );
  INV_X1 U11958 ( .A(n9340), .ZN(n9341) );
  OAI222_X1 U11959 ( .A1(P3_U3151), .A2(n15091), .B1(n12350), .B2(n15380), 
        .C1(n11060), .C2(n9341), .ZN(P3_U3281) );
  OR2_X1 U11960 ( .A1(n9342), .A2(n12295), .ZN(n9344) );
  NAND2_X1 U11961 ( .A1(n9350), .A2(n9345), .ZN(n9348) );
  NAND2_X1 U11962 ( .A1(n9346), .A2(n8356), .ZN(n9347) );
  NAND2_X1 U11963 ( .A1(n9348), .A2(n9347), .ZN(n9349) );
  XNOR2_X1 U11964 ( .A(n9349), .B(n12295), .ZN(n9352) );
  NAND2_X1 U11965 ( .A1(n9352), .A2(n9351), .ZN(n9373) );
  INV_X1 U11966 ( .A(n9374), .ZN(n9355) );
  AOI21_X1 U11967 ( .B1(n9357), .B2(n9356), .A(n9355), .ZN(n9361) );
  NOR2_X1 U11968 ( .A1(n13808), .A2(n14170), .ZN(n13789) );
  INV_X1 U11969 ( .A(n13789), .ZN(n14594) );
  INV_X1 U11970 ( .A(n13797), .ZN(n14593) );
  OAI22_X1 U11971 ( .A1(n8777), .A2(n14594), .B1(n14593), .B2(n9732), .ZN(
        n9359) );
  NOR2_X1 U11972 ( .A1(n13792), .A2(n14708), .ZN(n9358) );
  AOI211_X1 U11973 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n11964), .A(n9359), .B(
        n9358), .ZN(n9360) );
  OAI21_X1 U11974 ( .B1(n9361), .B2(n14598), .A(n9360), .ZN(P1_U3222) );
  INV_X1 U11975 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U11976 ( .A1(n11235), .A2(P3_U3897), .ZN(n9362) );
  OAI21_X1 U11977 ( .B1(P3_U3897), .B2(n9363), .A(n9362), .ZN(P3_U3503) );
  INV_X1 U11978 ( .A(n10755), .ZN(n9369) );
  OAI222_X1 U11979 ( .A1(n14332), .A2(n9364), .B1(n14330), .B2(n9369), .C1(
        n9778), .C2(P1_U3086), .ZN(P1_U3342) );
  OAI21_X1 U11980 ( .B1(n9365), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9367) );
  INV_X1 U11981 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9366) );
  XNOR2_X1 U11982 ( .A(n9367), .B(n9366), .ZN(n10756) );
  INV_X1 U11983 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9368) );
  OAI222_X1 U11984 ( .A1(P2_U3088), .A2(n10756), .B1(n11317), .B2(n9369), .C1(
        n9368), .C2(n13693), .ZN(P2_U3314) );
  INV_X1 U11985 ( .A(n9370), .ZN(n9371) );
  OAI222_X1 U11986 ( .A1(P3_U3151), .A2(n14470), .B1(n12350), .B2(n9372), .C1(
        n11060), .C2(n9371), .ZN(P3_U3280) );
  NAND2_X1 U11987 ( .A1(n9374), .A2(n9373), .ZN(n11959) );
  NAND2_X1 U11988 ( .A1(n13839), .A2(n9345), .ZN(n9376) );
  INV_X2 U11989 ( .A(n11834), .ZN(n12326) );
  NAND2_X1 U11990 ( .A1(n9961), .A2(n9346), .ZN(n9375) );
  NAND2_X1 U11991 ( .A1(n9376), .A2(n9375), .ZN(n9377) );
  XNOR2_X1 U11992 ( .A(n9377), .B(n12324), .ZN(n9378) );
  AOI22_X1 U11993 ( .A1(n13839), .A2(n11811), .B1(n6648), .B2(n9961), .ZN(
        n9379) );
  XNOR2_X1 U11994 ( .A(n9378), .B(n9379), .ZN(n11960) );
  INV_X1 U11995 ( .A(n9378), .ZN(n9380) );
  NAND2_X1 U11996 ( .A1(n9380), .A2(n9379), .ZN(n9381) );
  NAND2_X1 U11997 ( .A1(n13838), .A2(n6648), .ZN(n9383) );
  NAND2_X1 U11998 ( .A1(n6883), .A2(n12326), .ZN(n9382) );
  NAND2_X1 U11999 ( .A1(n9383), .A2(n9382), .ZN(n9384) );
  XNOR2_X1 U12000 ( .A(n9384), .B(n12295), .ZN(n9801) );
  NAND2_X1 U12001 ( .A1(n13838), .A2(n12322), .ZN(n9386) );
  NAND2_X1 U12002 ( .A1(n6883), .A2(n6648), .ZN(n9385) );
  NAND2_X1 U12003 ( .A1(n9386), .A2(n9385), .ZN(n9802) );
  XNOR2_X1 U12004 ( .A(n9801), .B(n9802), .ZN(n9387) );
  OAI211_X1 U12005 ( .C1(n9388), .C2(n9387), .A(n9805), .B(n14585), .ZN(n9395)
         );
  OAI21_X2 U12006 ( .B1(n9390), .B2(n9389), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n14606) );
  INV_X1 U12007 ( .A(n14606), .ZN(n13806) );
  INV_X1 U12008 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9393) );
  NAND2_X1 U12009 ( .A1(n13797), .A2(n13837), .ZN(n9391) );
  NAND2_X1 U12010 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13865) );
  OAI211_X1 U12011 ( .C1(n14594), .C2(n9732), .A(n9391), .B(n13865), .ZN(n9392) );
  AOI21_X1 U12012 ( .B1(n13806), .B2(n9393), .A(n9392), .ZN(n9394) );
  OAI211_X1 U12013 ( .C1(n7078), .C2(n13792), .A(n9395), .B(n9394), .ZN(
        P1_U3218) );
  INV_X1 U12014 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n15347) );
  NAND2_X1 U12015 ( .A1(n12991), .A2(P3_U3897), .ZN(n9396) );
  OAI21_X1 U12016 ( .B1(P3_U3897), .B2(n15347), .A(n9396), .ZN(P3_U3506) );
  MUX2_X1 U12017 ( .A(n9397), .B(P1_REG2_REG_12__SCAN_IN), .S(n9406), .Z(n9402) );
  NOR2_X1 U12018 ( .A1(n9398), .A2(n10309), .ZN(n13944) );
  MUX2_X1 U12019 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n9399), .S(n13945), .Z(
        n9400) );
  OAI21_X1 U12020 ( .B1(n13950), .B2(n13944), .A(n9400), .ZN(n13948) );
  OAI21_X1 U12021 ( .B1(n9399), .B2(n9405), .A(n13948), .ZN(n9401) );
  NOR2_X1 U12022 ( .A1(n9401), .A2(n9402), .ZN(n9480) );
  AOI21_X1 U12023 ( .B1(n9402), .B2(n9401), .A(n9480), .ZN(n9415) );
  AOI21_X1 U12024 ( .B1(n9404), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9403), .ZN(
        n13939) );
  MUX2_X1 U12025 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n8510), .S(n13945), .Z(
        n13940) );
  NAND2_X1 U12026 ( .A1(n13939), .A2(n13940), .ZN(n13938) );
  NAND2_X1 U12027 ( .A1(n9405), .A2(n8510), .ZN(n9409) );
  OR2_X1 U12028 ( .A1(n9406), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U12029 ( .A1(n9406), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9407) );
  NAND2_X1 U12030 ( .A1(n9477), .A2(n9407), .ZN(n9408) );
  AOI21_X1 U12031 ( .B1(n13938), .B2(n9409), .A(n9408), .ZN(n9479) );
  AND3_X1 U12032 ( .A1(n13938), .A2(n9409), .A3(n9408), .ZN(n9410) );
  OAI21_X1 U12033 ( .B1(n9479), .B2(n9410), .A(n13966), .ZN(n9414) );
  NOR2_X1 U12034 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11129), .ZN(n9412) );
  NOR2_X1 U12035 ( .A1(n14647), .A2(n9481), .ZN(n9411) );
  AOI211_X1 U12036 ( .C1(n13929), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9412), .B(
        n9411), .ZN(n9413) );
  OAI211_X1 U12037 ( .C1(n9415), .C2(n14645), .A(n9414), .B(n9413), .ZN(
        P1_U3255) );
  INV_X1 U12038 ( .A(n9416), .ZN(n9417) );
  INV_X1 U12039 ( .A(n14480), .ZN(n12772) );
  OAI222_X1 U12040 ( .A1(n12350), .A2(n9418), .B1(n11060), .B2(n9417), .C1(
        n12772), .C2(P3_U3151), .ZN(P3_U3279) );
  XNOR2_X1 U12041 ( .A(n10908), .B(n11948), .ZN(n9419) );
  NAND2_X1 U12042 ( .A1(n9419), .A2(n11210), .ZN(n9420) );
  INV_X1 U12043 ( .A(n11318), .ZN(n9421) );
  INV_X1 U12044 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14854) );
  NAND2_X1 U12045 ( .A1(n14850), .A2(n14854), .ZN(n9423) );
  OR2_X1 U12046 ( .A1(n9421), .A2(n10908), .ZN(n9422) );
  NAND2_X1 U12047 ( .A1(n9423), .A2(n9422), .ZN(n10094) );
  INV_X1 U12048 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14856) );
  NAND2_X1 U12049 ( .A1(n14850), .A2(n14856), .ZN(n9425) );
  NAND2_X1 U12050 ( .A1(n11318), .A2(n11210), .ZN(n9424) );
  NAND2_X1 U12051 ( .A1(n9425), .A2(n9424), .ZN(n10096) );
  NOR2_X1 U12052 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .ZN(
        n9429) );
  NOR4_X1 U12053 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n9428) );
  NOR4_X1 U12054 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9427) );
  NOR4_X1 U12055 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9426) );
  AND4_X1 U12056 ( .A1(n9429), .A2(n9428), .A3(n9427), .A4(n9426), .ZN(n9435)
         );
  NOR4_X1 U12057 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n9433) );
  NOR4_X1 U12058 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n9432) );
  NOR4_X1 U12059 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9431) );
  NOR4_X1 U12060 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9430) );
  AND4_X1 U12061 ( .A1(n9433), .A2(n9432), .A3(n9431), .A4(n9430), .ZN(n9434)
         );
  NAND2_X1 U12062 ( .A1(n9435), .A2(n9434), .ZN(n9436) );
  AND2_X1 U12063 ( .A1(n14850), .A2(n9436), .ZN(n10095) );
  OR3_X1 U12064 ( .A1(n10094), .A2(n10096), .A3(n10095), .ZN(n9461) );
  INV_X1 U12065 ( .A(n9461), .ZN(n9438) );
  NAND2_X1 U12066 ( .A1(n9437), .A2(n10851), .ZN(n9638) );
  NAND2_X1 U12067 ( .A1(n9439), .A2(n9757), .ZN(n9440) );
  NOR2_X1 U12068 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(n9440), .ZN(n10010) );
  NAND2_X1 U12069 ( .A1(n9443), .A2(n9442), .ZN(n9446) );
  NAND2_X1 U12070 ( .A1(n9446), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9447) );
  INV_X1 U12071 ( .A(n13268), .ZN(n13217) );
  INV_X1 U12072 ( .A(n13243), .ZN(n13258) );
  NAND2_X1 U12073 ( .A1(n9450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9449) );
  OR2_X2 U12074 ( .A1(n9450), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n13677) );
  NAND2_X2 U12075 ( .A1(n9451), .A2(n13677), .ZN(n13683) );
  AND2_X2 U12076 ( .A1(n12267), .A2(n9452), .ZN(n9574) );
  NAND2_X1 U12077 ( .A1(n9574), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9453) );
  AND2_X1 U12078 ( .A1(n9454), .A2(n9453), .ZN(n9459) );
  INV_X1 U12079 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U12080 ( .A1(n10957), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9457) );
  NAND3_X2 U12081 ( .A1(n9459), .A2(n9458), .A3(n9457), .ZN(n11323) );
  NAND2_X1 U12082 ( .A1(n11748), .A2(n9569), .ZN(n11327) );
  OR2_X1 U12083 ( .A1(n13655), .A2(n11757), .ZN(n9472) );
  AOI21_X1 U12084 ( .B1(n9461), .B2(n9472), .A(n10097), .ZN(n9640) );
  NAND2_X1 U12085 ( .A1(n9640), .A2(n11767), .ZN(n13245) );
  INV_X1 U12086 ( .A(n9473), .ZN(n9463) );
  AND2_X1 U12087 ( .A1(n14909), .A2(n9572), .ZN(n9462) );
  NAND2_X1 U12088 ( .A1(n6656), .A2(n13653), .ZN(n9657) );
  NAND2_X1 U12089 ( .A1(n9605), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9467) );
  INV_X1 U12090 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9465) );
  CLKBUF_X1 U12091 ( .A(n11331), .Z(n13302) );
  INV_X1 U12092 ( .A(n13302), .ZN(n9579) );
  NAND2_X1 U12093 ( .A1(n9468), .A2(SI_0_), .ZN(n9469) );
  XNOR2_X1 U12094 ( .A(n9469), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13694) );
  NAND2_X1 U12095 ( .A1(n11331), .A2(n13654), .ZN(n11721) );
  INV_X1 U12096 ( .A(n11721), .ZN(n9567) );
  NOR4_X1 U12097 ( .A1(n13275), .A2(n10936), .A3(n9579), .A4(n9567), .ZN(n9470) );
  AOI21_X1 U12098 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n13245), .A(n9470), .ZN(
        n9476) );
  INV_X1 U12099 ( .A(n13653), .ZN(n9471) );
  OR2_X1 U12100 ( .A1(n6656), .A2(n9471), .ZN(n10103) );
  OAI21_X1 U12101 ( .B1(n9647), .B2(n13275), .A(n13242), .ZN(n9474) );
  NAND2_X1 U12102 ( .A1(n9474), .A2(n13654), .ZN(n9475) );
  OAI211_X1 U12103 ( .C1(n13258), .C2(n11337), .A(n9476), .B(n9475), .ZN(
        P2_U3204) );
  INV_X1 U12104 ( .A(n9477), .ZN(n9478) );
  NOR2_X1 U12105 ( .A1(n9479), .A2(n9478), .ZN(n9770) );
  XNOR2_X1 U12106 ( .A(n9778), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9769) );
  XNOR2_X1 U12107 ( .A(n9770), .B(n9769), .ZN(n9489) );
  NAND2_X1 U12108 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11250)
         );
  AOI21_X1 U12109 ( .B1(n9397), .B2(n9481), .A(n9480), .ZN(n9484) );
  MUX2_X1 U12110 ( .A(n9482), .B(P1_REG2_REG_13__SCAN_IN), .S(n9778), .Z(n9483) );
  NAND2_X1 U12111 ( .A1(n9484), .A2(n9483), .ZN(n9777) );
  OAI211_X1 U12112 ( .C1(n9484), .C2(n9483), .A(n13963), .B(n9777), .ZN(n9485)
         );
  NAND2_X1 U12113 ( .A1(n11250), .A2(n9485), .ZN(n9487) );
  NOR2_X1 U12114 ( .A1(n14647), .A2(n9778), .ZN(n9486) );
  AOI211_X1 U12115 ( .C1(n13929), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n9487), .B(
        n9486), .ZN(n9488) );
  OAI21_X1 U12116 ( .B1(n9489), .B2(n14643), .A(n9488), .ZN(P1_U3256) );
  INV_X1 U12117 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9496) );
  INV_X1 U12118 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9885) );
  MUX2_X1 U12119 ( .A(n9496), .B(n9885), .S(n9517), .Z(n14946) );
  AND2_X1 U12120 ( .A1(n14946), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14949) );
  MUX2_X1 U12121 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n9517), .Z(n9518) );
  XOR2_X1 U12122 ( .A(n14949), .B(n9520), .Z(n9516) );
  NAND2_X1 U12123 ( .A1(n9492), .A2(n12672), .ZN(n9490) );
  NAND2_X1 U12124 ( .A1(n9491), .A2(n9490), .ZN(n9501) );
  INV_X1 U12125 ( .A(n9492), .ZN(n9493) );
  NAND2_X1 U12126 ( .A1(n9493), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12697) );
  INV_X1 U12127 ( .A(n12697), .ZN(n9494) );
  NOR2_X1 U12128 ( .A1(n12690), .A2(n9494), .ZN(n9500) );
  OR2_X1 U12129 ( .A1(n9501), .A2(n9500), .ZN(n9503) );
  MUX2_X1 U12130 ( .A(n9503), .B(n12720), .S(n9495), .Z(n15092) );
  INV_X1 U12131 ( .A(n15092), .ZN(n14999) );
  INV_X1 U12132 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15143) );
  NOR3_X1 U12133 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n9496), .ZN(n9521) );
  INV_X1 U12134 ( .A(n9521), .ZN(n9497) );
  AOI21_X1 U12135 ( .B1(n15143), .B2(n9498), .A(n9522), .ZN(n9513) );
  INV_X1 U12136 ( .A(n9500), .ZN(n9502) );
  AOI22_X1 U12137 ( .A1(n15095), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9512) );
  INV_X1 U12138 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9504) );
  AND2_X1 U12139 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9504), .ZN(n9505) );
  OR3_X1 U12140 ( .A1(n9885), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n9528) );
  OAI21_X1 U12141 ( .B1(n9506), .B2(n9505), .A(n9528), .ZN(n9508) );
  INV_X1 U12142 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9507) );
  OR2_X1 U12143 ( .A1(n9508), .A2(n9507), .ZN(n9529) );
  NAND2_X1 U12144 ( .A1(n9508), .A2(n9507), .ZN(n9509) );
  NAND2_X1 U12145 ( .A1(n9529), .A2(n9509), .ZN(n9510) );
  NAND2_X1 U12146 ( .A1(n15087), .A2(n9510), .ZN(n9511) );
  OAI211_X1 U12147 ( .C1(n9513), .C2(n15102), .A(n9512), .B(n9511), .ZN(n9514)
         );
  AOI21_X1 U12148 ( .B1(n6952), .B2(n14999), .A(n9514), .ZN(n9515) );
  OAI21_X1 U12149 ( .B1(n15077), .B2(n9516), .A(n9515), .ZN(P3_U3183) );
  MUX2_X1 U12150 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n9517), .Z(n9539) );
  XOR2_X1 U12151 ( .A(n9523), .B(n9539), .Z(n9540) );
  INV_X1 U12152 ( .A(n9518), .ZN(n9519) );
  XOR2_X1 U12153 ( .A(n9540), .B(n9541), .Z(n9538) );
  NOR2_X1 U12154 ( .A1(n9522), .A2(n9521), .ZN(n9526) );
  INV_X1 U12155 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9524) );
  MUX2_X1 U12156 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n9524), .S(n9523), .Z(n9525)
         );
  AOI21_X1 U12157 ( .B1(n9526), .B2(n9525), .A(n9542), .ZN(n9535) );
  AOI22_X1 U12158 ( .A1(n15095), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n9534) );
  INV_X1 U12159 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9527) );
  MUX2_X1 U12160 ( .A(n9527), .B(P3_REG1_REG_2__SCAN_IN), .S(n9523), .Z(n9531)
         );
  NAND2_X1 U12161 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  NAND2_X1 U12162 ( .A1(n9531), .A2(n9530), .ZN(n9546) );
  OAI21_X1 U12163 ( .B1(n9531), .B2(n9530), .A(n9546), .ZN(n9532) );
  NAND2_X1 U12164 ( .A1(n15087), .A2(n9532), .ZN(n9533) );
  OAI211_X1 U12165 ( .C1(n9535), .C2(n15102), .A(n9534), .B(n9533), .ZN(n9536)
         );
  AOI21_X1 U12166 ( .B1(n9523), .B2(n14999), .A(n9536), .ZN(n9537) );
  OAI21_X1 U12167 ( .B1(n9538), .B2(n15077), .A(n9537), .ZN(P3_U3184) );
  MUX2_X1 U12168 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12758), .Z(n9694) );
  XNOR2_X1 U12169 ( .A(n9694), .B(n9708), .ZN(n9696) );
  XOR2_X1 U12170 ( .A(n9696), .B(n9697), .Z(n9553) );
  INV_X1 U12171 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9545) );
  AOI21_X1 U12172 ( .B1(n9545), .B2(n9544), .A(n9703), .ZN(n9550) );
  AOI22_X1 U12173 ( .A1(n15095), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n9549) );
  OAI21_X1 U12174 ( .B1(n9523), .B2(n9527), .A(n9546), .ZN(n9707) );
  XOR2_X1 U12175 ( .A(P3_REG1_REG_3__SCAN_IN), .B(n9710), .Z(n9547) );
  NAND2_X1 U12176 ( .A1(n15087), .A2(n9547), .ZN(n9548) );
  OAI211_X1 U12177 ( .C1(n9550), .C2(n15102), .A(n9549), .B(n9548), .ZN(n9551)
         );
  AOI21_X1 U12178 ( .B1(n9708), .B2(n14999), .A(n9551), .ZN(n9552) );
  OAI21_X1 U12179 ( .B1(n9553), .B2(n15077), .A(n9552), .ZN(P3_U3185) );
  INV_X1 U12180 ( .A(n9554), .ZN(n9555) );
  OAI222_X1 U12181 ( .A1(n12350), .A2(n15383), .B1(n11060), .B2(n9555), .C1(
        n12785), .C2(P3_U3151), .ZN(P3_U3278) );
  NOR2_X1 U12182 ( .A1(n10095), .A2(n9556), .ZN(n9634) );
  AND2_X1 U12183 ( .A1(n10096), .A2(n11767), .ZN(n14855) );
  INV_X1 U12184 ( .A(n10097), .ZN(n9557) );
  NAND2_X1 U12185 ( .A1(n11619), .A2(n9559), .ZN(n9565) );
  INV_X1 U12186 ( .A(n9561), .ZN(n9562) );
  INV_X1 U12187 ( .A(n9570), .ZN(n9566) );
  NAND2_X1 U12188 ( .A1(n9566), .A2(n11721), .ZN(n9590) );
  NAND2_X1 U12189 ( .A1(n9570), .A2(n9567), .ZN(n9568) );
  AND2_X1 U12190 ( .A1(n9590), .A2(n9568), .ZN(n10143) );
  NAND2_X1 U12191 ( .A1(n15591), .A2(n11757), .ZN(n11756) );
  NAND2_X1 U12192 ( .A1(n11748), .A2(n9581), .ZN(n11690) );
  INV_X1 U12193 ( .A(n13654), .ZN(n11332) );
  NOR2_X1 U12194 ( .A1(n13302), .A2(n11332), .ZN(n9571) );
  OAI21_X1 U12195 ( .B1(n9571), .B2(n9570), .A(n10226), .ZN(n9585) );
  NOR2_X2 U12196 ( .A1(n9572), .A2(n9061), .ZN(n13470) );
  INV_X1 U12197 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U12198 ( .A1(n9605), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U12199 ( .A1(n9574), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9576) );
  OR2_X1 U12200 ( .A1(n11689), .A2(n10236), .ZN(n9575) );
  INV_X1 U12201 ( .A(n11346), .ZN(n9598) );
  OAI22_X1 U12202 ( .A1(n9579), .A2(n13538), .B1(n9598), .B2(n13540), .ZN(
        n9584) );
  NOR2_X1 U12203 ( .A1(n10143), .A2(n13647), .ZN(n9583) );
  AOI211_X1 U12204 ( .C1(n13521), .C2(n9585), .A(n9584), .B(n9583), .ZN(n10151) );
  NAND2_X1 U12205 ( .A1(n11324), .A2(n11332), .ZN(n10232) );
  INV_X1 U12206 ( .A(n10232), .ZN(n9586) );
  AOI211_X1 U12207 ( .C1(n13654), .C2(n13179), .A(n13459), .B(n9586), .ZN(
        n10145) );
  AOI21_X1 U12208 ( .B1(n14917), .B2(n13179), .A(n10145), .ZN(n9587) );
  OAI211_X1 U12209 ( .C1(n10143), .C2(n13655), .A(n10151), .B(n9587), .ZN(
        n13646) );
  NAND2_X1 U12210 ( .A1(n13646), .A2(n14925), .ZN(n9588) );
  OAI21_X1 U12211 ( .B1(n14925), .B2(n9455), .A(n9588), .ZN(P2_U3433) );
  INV_X1 U12212 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12213 ( .A1(n11337), .A2(n11324), .ZN(n9589) );
  NAND2_X1 U12214 ( .A1(n9590), .A2(n9589), .ZN(n10224) );
  NOR2_X1 U12215 ( .A1(n9591), .A2(n11572), .ZN(n9595) );
  OAI22_X1 U12216 ( .A1(n9592), .A2(n9593), .B1(n9601), .B2(n14780), .ZN(n9594) );
  OR2_X1 U12217 ( .A1(n9595), .A2(n9594), .ZN(n9596) );
  NAND2_X1 U12218 ( .A1(n9598), .A2(n13246), .ZN(n9616) );
  INV_X1 U12219 ( .A(n9596), .ZN(n9646) );
  NAND2_X1 U12220 ( .A1(n11346), .A2(n9646), .ZN(n9597) );
  NAND2_X1 U12221 ( .A1(n10224), .A2(n10227), .ZN(n10223) );
  NAND2_X1 U12222 ( .A1(n9598), .A2(n9646), .ZN(n9599) );
  NAND2_X1 U12223 ( .A1(n10223), .A2(n9599), .ZN(n9611) );
  NAND2_X1 U12224 ( .A1(n9600), .A2(n6652), .ZN(n9604) );
  AOI22_X1 U12225 ( .A1(n11683), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n11490), 
        .B2(n9602), .ZN(n9603) );
  NAND2_X1 U12226 ( .A1(n11686), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U12227 ( .A1(n11658), .A2(n13165), .ZN(n9609) );
  NAND2_X1 U12228 ( .A1(n9574), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9608) );
  OR2_X1 U12229 ( .A1(n11689), .A2(n9606), .ZN(n9607) );
  NAND4_X1 U12230 ( .A1(n9610), .A2(n9609), .A3(n9608), .A4(n9607), .ZN(n13300) );
  XNOR2_X1 U12231 ( .A(n11354), .B(n13300), .ZN(n11723) );
  NAND2_X1 U12232 ( .A1(n9611), .A2(n11723), .ZN(n10092) );
  OR2_X1 U12233 ( .A1(n9611), .A2(n11723), .ZN(n9612) );
  NAND2_X1 U12234 ( .A1(n10092), .A2(n9612), .ZN(n10496) );
  NOR2_X1 U12235 ( .A1(n10232), .A2(n13246), .ZN(n10234) );
  NAND2_X1 U12236 ( .A1(n10234), .A2(n11354), .ZN(n10458) );
  OAI211_X1 U12237 ( .C1(n10234), .C2(n11354), .A(n10458), .B(n10936), .ZN(
        n10492) );
  OAI21_X1 U12238 ( .B1(n11354), .B2(n14909), .A(n10492), .ZN(n9630) );
  INV_X1 U12239 ( .A(n13647), .ZN(n14873) );
  NAND2_X1 U12240 ( .A1(n10496), .A2(n14873), .ZN(n9629) );
  NAND2_X1 U12241 ( .A1(n11337), .A2(n13179), .ZN(n10225) );
  NAND2_X1 U12242 ( .A1(n10226), .A2(n10225), .ZN(n9613) );
  NAND2_X1 U12243 ( .A1(n9613), .A2(n11722), .ZN(n10228) );
  NAND2_X1 U12244 ( .A1(n10228), .A2(n9616), .ZN(n9615) );
  INV_X1 U12245 ( .A(n11723), .ZN(n9614) );
  NAND2_X1 U12246 ( .A1(n9615), .A2(n9614), .ZN(n10464) );
  NAND3_X1 U12247 ( .A1(n10228), .A2(n11723), .A3(n9616), .ZN(n9617) );
  NAND2_X1 U12248 ( .A1(n10464), .A2(n9617), .ZN(n9627) );
  NAND2_X1 U12249 ( .A1(n9574), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12250 ( .A1(n11686), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U12251 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9643) );
  OAI21_X1 U12252 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9643), .ZN(n9618) );
  INV_X1 U12253 ( .A(n9618), .ZN(n10461) );
  NAND2_X1 U12254 ( .A1(n11658), .A2(n10461), .ZN(n9621) );
  OR2_X1 U12255 ( .A1(n11689), .A2(n9619), .ZN(n9620) );
  NAND2_X1 U12256 ( .A1(n13650), .A2(n13299), .ZN(n9625) );
  NAND2_X1 U12257 ( .A1(n11346), .A2(n13470), .ZN(n9624) );
  NAND2_X1 U12258 ( .A1(n9625), .A2(n9624), .ZN(n9626) );
  AOI21_X1 U12259 ( .B1(n9627), .B2(n13521), .A(n9626), .ZN(n9628) );
  NAND2_X1 U12260 ( .A1(n9629), .A2(n9628), .ZN(n10493) );
  AOI211_X1 U12261 ( .C1(n14915), .C2(n10496), .A(n9630), .B(n10493), .ZN(
        n9635) );
  OR2_X1 U12262 ( .A1(n9635), .A2(n14923), .ZN(n9631) );
  OAI21_X1 U12263 ( .B1(n14925), .B2(n9632), .A(n9631), .ZN(P2_U3439) );
  OR2_X1 U12264 ( .A1(n9635), .A2(n14940), .ZN(n9636) );
  OAI21_X1 U12265 ( .B1(n14943), .B2(n9637), .A(n9636), .ZN(P2_U3502) );
  INV_X1 U12266 ( .A(n9638), .ZN(n9639) );
  NAND2_X1 U12267 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  NOR2_X1 U12268 ( .A1(n9643), .A2(n9642), .ZN(n9677) );
  AND2_X1 U12269 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  NOR2_X1 U12270 ( .A1(n9677), .A2(n9644), .ZN(n9669) );
  INV_X1 U12271 ( .A(n9669), .ZN(n10104) );
  XNOR2_X1 U12272 ( .A(n9850), .B(n9646), .ZN(n9652) );
  NAND2_X1 U12273 ( .A1(n11346), .A2(n9657), .ZN(n9651) );
  NAND2_X1 U12274 ( .A1(n11323), .A2(n9657), .ZN(n9649) );
  NOR2_X1 U12275 ( .A1(n9647), .A2(n7566), .ZN(n13182) );
  NAND2_X1 U12276 ( .A1(n13181), .A2(n13182), .ZN(n13180) );
  INV_X1 U12277 ( .A(n9648), .ZN(n9650) );
  NAND2_X1 U12278 ( .A1(n9650), .A2(n9649), .ZN(n13247) );
  XNOR2_X1 U12279 ( .A(n9652), .B(n9651), .ZN(n13248) );
  XNOR2_X1 U12280 ( .A(n12012), .B(n11354), .ZN(n9654) );
  NAND2_X1 U12281 ( .A1(n13300), .A2(n9657), .ZN(n9653) );
  NOR2_X1 U12282 ( .A1(n9654), .A2(n9653), .ZN(n9655) );
  AOI21_X1 U12283 ( .B1(n9654), .B2(n9653), .A(n9655), .ZN(n13162) );
  NAND2_X1 U12284 ( .A1(n13163), .A2(n13162), .ZN(n13161) );
  INV_X1 U12285 ( .A(n9655), .ZN(n9656) );
  NAND2_X1 U12286 ( .A1(n13299), .A2(n9657), .ZN(n9662) );
  NAND2_X1 U12287 ( .A1(n9658), .A2(n6652), .ZN(n9661) );
  AOI22_X1 U12288 ( .A1(n11683), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n11490), 
        .B2(n9659), .ZN(n9660) );
  NAND2_X1 U12289 ( .A1(n9661), .A2(n9660), .ZN(n11370) );
  XNOR2_X1 U12290 ( .A(n12012), .B(n11370), .ZN(n9664) );
  XOR2_X1 U12291 ( .A(n9662), .B(n9664), .Z(n9824) );
  INV_X1 U12292 ( .A(n9662), .ZN(n9663) );
  NOR2_X1 U12293 ( .A1(n9664), .A2(n9663), .ZN(n9675) );
  OR2_X1 U12294 ( .A1(n9665), .A2(n11572), .ZN(n9668) );
  AOI22_X1 U12295 ( .A1(n11683), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n11490), 
        .B2(n9666), .ZN(n9667) );
  XNOR2_X1 U12296 ( .A(n14874), .B(n12012), .ZN(n9845) );
  NAND2_X1 U12297 ( .A1(n11686), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U12298 ( .A1(n11642), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U12299 ( .A1(n11658), .A2(n9669), .ZN(n9671) );
  OR2_X1 U12300 ( .A1(n11605), .A2(n9105), .ZN(n9670) );
  NAND4_X1 U12301 ( .A1(n9673), .A2(n9672), .A3(n9671), .A4(n9670), .ZN(n13298) );
  NAND2_X1 U12302 ( .A1(n13298), .A2(n10208), .ZN(n9844) );
  XNOR2_X1 U12303 ( .A(n9845), .B(n9844), .ZN(n9674) );
  NOR3_X1 U12304 ( .A1(n9822), .A2(n9675), .A3(n9674), .ZN(n9676) );
  OAI21_X1 U12305 ( .B1(n6813), .B2(n9676), .A(n13249), .ZN(n9688) );
  NAND2_X1 U12306 ( .A1(n11686), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9682) );
  NAND2_X1 U12307 ( .A1(n11642), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9681) );
  NAND2_X1 U12308 ( .A1(n9677), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9856) );
  OR2_X1 U12309 ( .A1(n9677), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9678) );
  AND2_X1 U12310 ( .A1(n9856), .A2(n9678), .ZN(n10446) );
  NAND2_X1 U12311 ( .A1(n11658), .A2(n10446), .ZN(n9680) );
  OR2_X1 U12312 ( .A1(n11605), .A2(n9106), .ZN(n9679) );
  NAND4_X1 U12313 ( .A1(n9682), .A2(n9681), .A3(n9680), .A4(n9679), .ZN(n13297) );
  NAND2_X1 U12314 ( .A1(n13650), .A2(n13297), .ZN(n9684) );
  NAND2_X1 U12315 ( .A1(n13299), .A2(n13470), .ZN(n9683) );
  NAND2_X1 U12316 ( .A1(n9684), .A2(n9683), .ZN(n10111) );
  INV_X1 U12317 ( .A(n14874), .ZN(n10162) );
  NOR2_X1 U12318 ( .A1(n13242), .A2(n10162), .ZN(n9685) );
  AOI211_X1 U12319 ( .C1(n13268), .C2(n10111), .A(n9686), .B(n9685), .ZN(n9687) );
  OAI211_X1 U12320 ( .C1(n13270), .C2(n10104), .A(n9688), .B(n9687), .ZN(
        P2_U3199) );
  NOR2_X1 U12321 ( .A1(n8892), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n9758) );
  OR2_X1 U12322 ( .A1(n9758), .A2(n9689), .ZN(n9690) );
  XNOR2_X1 U12323 ( .A(n9690), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11170) );
  INV_X1 U12324 ( .A(n11170), .ZN(n13327) );
  INV_X1 U12325 ( .A(n11169), .ZN(n9692) );
  OAI222_X1 U12326 ( .A1(P2_U3088), .A2(n13327), .B1(n11317), .B2(n9692), .C1(
        n9691), .C2(n13693), .ZN(P2_U3311) );
  INV_X1 U12327 ( .A(n10880), .ZN(n10887) );
  OAI222_X1 U12328 ( .A1(n14332), .A2(n9693), .B1(n14330), .B2(n9692), .C1(
        n10887), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12329 ( .A(n9694), .ZN(n9695) );
  MUX2_X1 U12330 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12758), .Z(n9698) );
  XNOR2_X1 U12331 ( .A(n9698), .B(n14955), .ZN(n14953) );
  OAI22_X1 U12332 ( .A1(n14954), .A2(n14953), .B1(n9698), .B2(n14955), .ZN(
        n9700) );
  MUX2_X1 U12333 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12758), .Z(n10386) );
  XNOR2_X1 U12334 ( .A(n10386), .B(n10380), .ZN(n9699) );
  NAND2_X1 U12335 ( .A1(n9700), .A2(n9699), .ZN(n10387) );
  OAI21_X1 U12336 ( .B1(n9700), .B2(n9699), .A(n10387), .ZN(n9701) );
  NAND2_X1 U12337 ( .A1(n9701), .A2(n15096), .ZN(n9720) );
  INV_X1 U12338 ( .A(n15102), .ZN(n14520) );
  INV_X1 U12339 ( .A(n9702), .ZN(n9704) );
  INV_X1 U12340 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U12341 ( .A1(n9706), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n10254), .B2(
        n14955), .ZN(n14957) );
  INV_X1 U12342 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10486) );
  XNOR2_X1 U12343 ( .A(n10374), .B(n10486), .ZN(n9718) );
  INV_X1 U12344 ( .A(n15095), .ZN(n15054) );
  INV_X1 U12345 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9716) );
  INV_X1 U12346 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15201) );
  AOI22_X1 U12347 ( .A1(n9706), .A2(n15201), .B1(P3_REG1_REG_4__SCAN_IN), .B2(
        n14955), .ZN(n14960) );
  INV_X1 U12348 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n9709) );
  XNOR2_X1 U12349 ( .A(n10379), .B(n10385), .ZN(n9711) );
  NAND2_X1 U12350 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n9711), .ZN(n10381) );
  OAI21_X1 U12351 ( .B1(n9711), .B2(P3_REG1_REG_5__SCAN_IN), .A(n10381), .ZN(
        n9712) );
  NAND2_X1 U12352 ( .A1(n15087), .A2(n9712), .ZN(n9715) );
  NOR2_X1 U12353 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9713), .ZN(n10345) );
  INV_X1 U12354 ( .A(n10345), .ZN(n9714) );
  OAI211_X1 U12355 ( .C1(n15054), .C2(n9716), .A(n9715), .B(n9714), .ZN(n9717)
         );
  AOI21_X1 U12356 ( .B1(n14520), .B2(n9718), .A(n9717), .ZN(n9719) );
  OAI211_X1 U12357 ( .C1(n15092), .C2(n10385), .A(n9720), .B(n9719), .ZN(
        P3_U3187) );
  INV_X1 U12358 ( .A(n10932), .ZN(n9724) );
  INV_X1 U12359 ( .A(n9768), .ZN(n10669) );
  OAI222_X1 U12360 ( .A1(n14332), .A2(n9721), .B1(n14330), .B2(n9724), .C1(
        n10669), .C2(P1_U3086), .ZN(P1_U3341) );
  NAND2_X1 U12361 ( .A1(n9722), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9723) );
  XNOR2_X1 U12362 ( .A(n9723), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10933) );
  INV_X1 U12363 ( .A(n10933), .ZN(n10321) );
  OAI222_X1 U12364 ( .A1(n13693), .A2(n9725), .B1(n11317), .B2(n9724), .C1(
        n10321), .C2(P2_U3088), .ZN(P2_U3313) );
  OAI21_X1 U12365 ( .B1(n9727), .B2(n12212), .A(n9726), .ZN(n9728) );
  INV_X1 U12366 ( .A(n9728), .ZN(n9971) );
  OAI21_X1 U12367 ( .B1(n9731), .B2(n9730), .A(n9729), .ZN(n9735) );
  OAI22_X1 U12368 ( .A1(n12046), .A2(n14260), .B1(n9732), .B2(n14170), .ZN(
        n9734) );
  NOR2_X1 U12369 ( .A1(n9971), .A2(n14087), .ZN(n9733) );
  AOI211_X1 U12370 ( .C1(n14144), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9965)
         );
  AOI21_X1 U12371 ( .B1(n9957), .B2(n6883), .A(n14661), .ZN(n9736) );
  OAI211_X1 U12372 ( .C1(n9971), .C2(n14221), .A(n9965), .B(n9967), .ZN(n9741)
         );
  OAI22_X1 U12373 ( .A1(n14273), .A2(n7078), .B1(n14764), .B2(n9125), .ZN(
        n9737) );
  AOI21_X1 U12374 ( .B1(n9741), .B2(n14764), .A(n9737), .ZN(n9738) );
  INV_X1 U12375 ( .A(n9738), .ZN(P1_U3531) );
  INV_X1 U12376 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9739) );
  OAI22_X1 U12377 ( .A1(n14318), .A2(n7078), .B1(n14755), .B2(n9739), .ZN(
        n9740) );
  AOI21_X1 U12378 ( .B1(n9741), .B2(n14755), .A(n9740), .ZN(n9742) );
  INV_X1 U12379 ( .A(n9742), .ZN(P1_U3468) );
  INV_X1 U12380 ( .A(n14511), .ZN(n12770) );
  OAI222_X1 U12381 ( .A1(P3_U3151), .A2(n12770), .B1(n12350), .B2(n15493), 
        .C1(n11060), .C2(n9743), .ZN(P3_U3277) );
  OAI21_X1 U12382 ( .B1(n9745), .B2(n9747), .A(n9744), .ZN(n10087) );
  INV_X1 U12383 ( .A(n9982), .ZN(n9746) );
  AOI211_X1 U12384 ( .C1(n12052), .C2(n9746), .A(n14661), .B(n10053), .ZN(
        n10086) );
  XNOR2_X1 U12385 ( .A(n9748), .B(n9747), .ZN(n9750) );
  OAI22_X1 U12386 ( .A1(n12046), .A2(n14170), .B1(n9910), .B2(n14260), .ZN(
        n9880) );
  INV_X1 U12387 ( .A(n9880), .ZN(n9749) );
  OAI21_X1 U12388 ( .B1(n9750), .B2(n14656), .A(n9749), .ZN(n10081) );
  AOI211_X1 U12389 ( .C1(n14752), .C2(n10087), .A(n10086), .B(n10081), .ZN(
        n9756) );
  OAI22_X1 U12390 ( .A1(n14273), .A2(n10082), .B1(n14764), .B2(n8412), .ZN(
        n9751) );
  INV_X1 U12391 ( .A(n9751), .ZN(n9752) );
  OAI21_X1 U12392 ( .B1(n9756), .B2(n14761), .A(n9752), .ZN(P1_U3533) );
  INV_X1 U12393 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9753) );
  OAI22_X1 U12394 ( .A1(n14318), .A2(n10082), .B1(n14755), .B2(n9753), .ZN(
        n9754) );
  INV_X1 U12395 ( .A(n9754), .ZN(n9755) );
  OAI21_X1 U12396 ( .B1(n9756), .B2(n14753), .A(n9755), .ZN(P1_U3474) );
  NAND2_X1 U12397 ( .A1(n9758), .A2(n9757), .ZN(n9759) );
  NAND2_X1 U12398 ( .A1(n9759), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9760) );
  XNOR2_X1 U12399 ( .A(n9760), .B(n9439), .ZN(n13328) );
  INV_X1 U12400 ( .A(n11261), .ZN(n9763) );
  OAI222_X1 U12401 ( .A1(P2_U3088), .A2(n13328), .B1(n11317), .B2(n9763), .C1(
        n9761), .C2(n13693), .ZN(P2_U3310) );
  OAI222_X1 U12402 ( .A1(P1_U3086), .A2(n11051), .B1(n14330), .B2(n9763), .C1(
        n9762), .C2(n14332), .ZN(P1_U3338) );
  NAND2_X1 U12403 ( .A1(n8892), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9764) );
  XNOR2_X1 U12404 ( .A(n9764), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11063) );
  INV_X1 U12405 ( .A(n11063), .ZN(n10327) );
  INV_X1 U12406 ( .A(n11062), .ZN(n9766) );
  INV_X1 U12407 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9765) );
  OAI222_X1 U12408 ( .A1(P2_U3088), .A2(n10327), .B1(n11317), .B2(n9766), .C1(
        n9765), .C2(n13693), .ZN(P2_U3312) );
  INV_X1 U12409 ( .A(n10670), .ZN(n14646) );
  OAI222_X1 U12410 ( .A1(n14332), .A2(n9767), .B1(n14330), .B2(n9766), .C1(
        n14646), .C2(P1_U3086), .ZN(P1_U3340) );
  AOI22_X1 U12411 ( .A1(n9768), .A2(n10668), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10669), .ZN(n9774) );
  NAND2_X1 U12412 ( .A1(n9770), .A2(n9769), .ZN(n9771) );
  OAI21_X1 U12413 ( .B1(n9778), .B2(n9772), .A(n9771), .ZN(n9773) );
  NOR2_X1 U12414 ( .A1(n9774), .A2(n9773), .ZN(n10667) );
  AOI21_X1 U12415 ( .B1(n9774), .B2(n9773), .A(n10667), .ZN(n9783) );
  NAND2_X1 U12416 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14589)
         );
  NAND2_X1 U12417 ( .A1(n13929), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n9775) );
  OAI211_X1 U12418 ( .C1(n14647), .C2(n10669), .A(n14589), .B(n9775), .ZN(
        n9776) );
  INV_X1 U12419 ( .A(n9776), .ZN(n9782) );
  OAI21_X1 U12420 ( .B1(n9482), .B2(n9778), .A(n9777), .ZN(n9780) );
  XNOR2_X1 U12421 ( .A(n10669), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n9779) );
  NAND2_X1 U12422 ( .A1(n9779), .A2(n9780), .ZN(n10663) );
  OAI211_X1 U12423 ( .C1(n9780), .C2(n9779), .A(n13963), .B(n10663), .ZN(n9781) );
  OAI211_X1 U12424 ( .C1(n9783), .C2(n14643), .A(n9782), .B(n9781), .ZN(
        P1_U3257) );
  NAND2_X1 U12425 ( .A1(n15125), .A2(n9943), .ZN(n12536) );
  INV_X1 U12426 ( .A(n12536), .ZN(n12542) );
  NOR2_X1 U12427 ( .A1(n9791), .A2(n12542), .ZN(n12506) );
  NAND2_X1 U12428 ( .A1(n9784), .A2(n15182), .ZN(n9785) );
  OR2_X1 U12429 ( .A1(n12506), .A2(n9785), .ZN(n9787) );
  OR2_X1 U12430 ( .A1(n15112), .A2(n15136), .ZN(n9786) );
  NAND2_X1 U12431 ( .A1(n9787), .A2(n9786), .ZN(n9939) );
  INV_X1 U12432 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9788) );
  OAI22_X1 U12433 ( .A1(n13131), .A2(n9943), .B1(n15197), .B2(n9788), .ZN(
        n9789) );
  AOI21_X1 U12434 ( .B1(n9939), .B2(n15197), .A(n9789), .ZN(n9790) );
  INV_X1 U12435 ( .A(n9790), .ZN(P3_U3390) );
  NOR2_X1 U12436 ( .A1(n12451), .A2(P3_U3151), .ZN(n9904) );
  INV_X1 U12437 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n9799) );
  INV_X1 U12438 ( .A(n9791), .ZN(n15138) );
  NAND3_X1 U12439 ( .A1(n15138), .A2(n15139), .A3(n11895), .ZN(n9792) );
  OAI211_X1 U12440 ( .C1(n9794), .C2(n15126), .A(n9793), .B(n9792), .ZN(n9795)
         );
  NAND2_X1 U12441 ( .A1(n9795), .A2(n12436), .ZN(n9798) );
  OAI22_X1 U12442 ( .A1(n15135), .A2(n12368), .B1(n15124), .B2(n12446), .ZN(
        n9796) );
  AOI21_X1 U12443 ( .B1(n11899), .B2(n15125), .A(n9796), .ZN(n9797) );
  OAI211_X1 U12444 ( .C1(n9904), .C2(n9799), .A(n9798), .B(n9797), .ZN(
        P3_U3162) );
  AOI22_X1 U12445 ( .A1(n14722), .A2(n12326), .B1(n12323), .B2(n13837), .ZN(
        n9800) );
  XOR2_X1 U12446 ( .A(n12324), .B(n9800), .Z(n9809) );
  INV_X1 U12447 ( .A(n9801), .ZN(n9803) );
  NAND2_X1 U12448 ( .A1(n9803), .A2(n9802), .ZN(n9804) );
  AOI22_X1 U12449 ( .A1(n14722), .A2(n12323), .B1(n12322), .B2(n13837), .ZN(
        n9806) );
  INV_X1 U12450 ( .A(n9869), .ZN(n9807) );
  AOI21_X1 U12451 ( .B1(n9809), .B2(n9808), .A(n9807), .ZN(n9815) );
  NAND2_X1 U12452 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13891) );
  INV_X1 U12453 ( .A(n13808), .ZN(n14587) );
  NAND2_X1 U12454 ( .A1(n13838), .A2(n14082), .ZN(n9811) );
  NAND2_X1 U12455 ( .A1(n13836), .A2(n14079), .ZN(n9810) );
  NAND2_X1 U12456 ( .A1(n9811), .A2(n9810), .ZN(n14721) );
  NAND2_X1 U12457 ( .A1(n14587), .A2(n14721), .ZN(n9812) );
  OAI211_X1 U12458 ( .C1(n14606), .C2(n9984), .A(n13891), .B(n9812), .ZN(n9813) );
  AOI21_X1 U12459 ( .B1(n14602), .B2(n14722), .A(n9813), .ZN(n9814) );
  OAI21_X1 U12460 ( .B1(n9815), .B2(n14598), .A(n9814), .ZN(P1_U3230) );
  OAI222_X1 U12461 ( .A1(n11060), .A2(n9817), .B1(n12350), .B2(n9816), .C1(
        P3_U3151), .C2(n12769), .ZN(P3_U3276) );
  INV_X1 U12462 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9942) );
  INV_X1 U12463 ( .A(n12368), .ZN(n12440) );
  NAND2_X1 U12464 ( .A1(P3_U3151), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n14944) );
  OAI21_X1 U12465 ( .B1(n12446), .B2(n9943), .A(n14944), .ZN(n9819) );
  NOR2_X1 U12466 ( .A1(n12506), .A2(n12459), .ZN(n9818) );
  AOI211_X1 U12467 ( .C1(n12440), .C2(n12719), .A(n9819), .B(n9818), .ZN(n9820) );
  OAI21_X1 U12468 ( .B1(n12418), .B2(n9942), .A(n9820), .ZN(P3_U3172) );
  NAND2_X1 U12469 ( .A1(n12720), .A2(P3_DATAO_REG_25__SCAN_IN), .ZN(n9821) );
  OAI21_X1 U12470 ( .B1(n12656), .B2(n12720), .A(n9821), .ZN(P3_U3516) );
  AOI21_X1 U12471 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9829) );
  INV_X1 U12472 ( .A(n13270), .ZN(n13219) );
  INV_X1 U12473 ( .A(n11370), .ZN(n14866) );
  OAI21_X1 U12474 ( .B1(n13242), .B2(n14866), .A(n9825), .ZN(n9827) );
  INV_X1 U12475 ( .A(n13300), .ZN(n11358) );
  NOR2_X2 U12476 ( .A1(n13217), .A2(n13538), .ZN(n13244) );
  INV_X1 U12477 ( .A(n13244), .ZN(n13257) );
  OAI22_X1 U12478 ( .A1(n11358), .A2(n13257), .B1(n13258), .B2(n11384), .ZN(
        n9826) );
  AOI211_X1 U12479 ( .C1(n10461), .C2(n13219), .A(n9827), .B(n9826), .ZN(n9828) );
  OAI21_X1 U12480 ( .B1(n9829), .B2(n13275), .A(n9828), .ZN(P2_U3202) );
  INV_X1 U12481 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9833) );
  INV_X1 U12482 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9832) );
  NAND2_X1 U12483 ( .A1(n9831), .A2(n9830), .ZN(n13310) );
  MUX2_X1 U12484 ( .A(n9832), .B(P2_REG2_REG_12__SCAN_IN), .S(n13309), .Z(
        n13311) );
  AOI21_X1 U12485 ( .B1(n13312), .B2(n13310), .A(n13311), .ZN(n13314) );
  MUX2_X1 U12486 ( .A(n9833), .B(P2_REG2_REG_13__SCAN_IN), .S(n10756), .Z(
        n14828) );
  NAND2_X1 U12487 ( .A1(n14829), .A2(n14828), .ZN(n14827) );
  OAI21_X1 U12488 ( .B1(n9833), .B2(n10756), .A(n14827), .ZN(n10315) );
  XOR2_X1 U12489 ( .A(n10315), .B(n10321), .Z(n9834) );
  NOR2_X1 U12490 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9834), .ZN(n10316) );
  AOI21_X1 U12491 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9834), .A(n10316), .ZN(
        n9843) );
  INV_X1 U12492 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14570) );
  INV_X1 U12493 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14576) );
  AOI21_X1 U12494 ( .B1(n10516), .B2(P2_REG1_REG_11__SCAN_IN), .A(n9835), .ZN(
        n13304) );
  MUX2_X1 U12495 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14576), .S(n13309), .Z(
        n13303) );
  AND2_X1 U12496 ( .A1(n13304), .A2(n13303), .ZN(n13305) );
  AOI21_X1 U12497 ( .B1(n14576), .B2(n9836), .A(n13305), .ZN(n14826) );
  MUX2_X1 U12498 ( .A(n14570), .B(P2_REG1_REG_13__SCAN_IN), .S(n10756), .Z(
        n14825) );
  NAND2_X1 U12499 ( .A1(n14826), .A2(n14825), .ZN(n14824) );
  OAI21_X1 U12500 ( .B1(n14570), .B2(n10756), .A(n14824), .ZN(n9838) );
  XNOR2_X1 U12501 ( .A(n10321), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U12502 ( .A1(n9837), .A2(n9838), .ZN(n10319) );
  OAI211_X1 U12503 ( .C1(n9838), .C2(n9837), .A(n14843), .B(n10319), .ZN(n9840) );
  AND2_X1 U12504 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n10962) );
  AOI21_X1 U12505 ( .B1(n14835), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n10962), 
        .ZN(n9839) );
  OAI211_X1 U12506 ( .C1(n14765), .C2(n10321), .A(n9840), .B(n9839), .ZN(n9841) );
  INV_X1 U12507 ( .A(n9841), .ZN(n9842) );
  OAI21_X1 U12508 ( .B1(n9843), .B2(n14811), .A(n9842), .ZN(P2_U3228) );
  INV_X1 U12509 ( .A(n9844), .ZN(n9846) );
  AOI22_X1 U12510 ( .A1(n11683), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n11490), 
        .B2(n9848), .ZN(n9849) );
  XNOR2_X1 U12511 ( .A(n11392), .B(n12012), .ZN(n9852) );
  AND2_X1 U12512 ( .A1(n13297), .A2(n10208), .ZN(n9851) );
  NAND2_X1 U12513 ( .A1(n9852), .A2(n9851), .ZN(n10130) );
  OAI21_X1 U12514 ( .B1(n9852), .B2(n9851), .A(n10130), .ZN(n9853) );
  AOI211_X1 U12515 ( .C1(n9854), .C2(n9853), .A(n13275), .B(n10132), .ZN(n9867) );
  INV_X1 U12516 ( .A(n10446), .ZN(n9865) );
  NAND2_X1 U12517 ( .A1(n11686), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U12518 ( .A1(n9856), .A2(n9855), .ZN(n9857) );
  AND2_X1 U12519 ( .A1(n10121), .A2(n9857), .ZN(n10178) );
  NAND2_X1 U12520 ( .A1(n11658), .A2(n10178), .ZN(n9861) );
  NAND2_X1 U12521 ( .A1(n11642), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9860) );
  OR2_X1 U12522 ( .A1(n11605), .A2(n10176), .ZN(n9859) );
  NAND4_X1 U12523 ( .A1(n9862), .A2(n9861), .A3(n9860), .A4(n9859), .ZN(n13296) );
  AOI22_X1 U12524 ( .A1(n13244), .A2(n13298), .B1(n13243), .B2(n13296), .ZN(
        n9864) );
  AOI22_X1 U12525 ( .A1(n13273), .A2(n11392), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9863) );
  OAI211_X1 U12526 ( .C1(n9865), .C2(n13270), .A(n9864), .B(n9863), .ZN(n9866)
         );
  OR2_X1 U12527 ( .A1(n9867), .A2(n9866), .ZN(P2_U3211) );
  NAND2_X1 U12528 ( .A1(n9869), .A2(n9868), .ZN(n10035) );
  NAND2_X1 U12529 ( .A1(n12052), .A2(n12326), .ZN(n9871) );
  NAND2_X1 U12530 ( .A1(n13836), .A2(n12323), .ZN(n9870) );
  NAND2_X1 U12531 ( .A1(n9871), .A2(n9870), .ZN(n9872) );
  XNOR2_X1 U12532 ( .A(n9872), .B(n12324), .ZN(n9876) );
  NAND2_X1 U12533 ( .A1(n12052), .A2(n12323), .ZN(n9874) );
  NAND2_X1 U12534 ( .A1(n13836), .A2(n12322), .ZN(n9873) );
  NAND2_X1 U12535 ( .A1(n9874), .A2(n9873), .ZN(n9875) );
  NOR2_X1 U12536 ( .A1(n9876), .A2(n9875), .ZN(n10034) );
  INV_X1 U12537 ( .A(n10034), .ZN(n9877) );
  NAND2_X1 U12538 ( .A1(n9876), .A2(n9875), .ZN(n10033) );
  NAND2_X1 U12539 ( .A1(n9877), .A2(n10033), .ZN(n9878) );
  XNOR2_X1 U12540 ( .A(n10035), .B(n9878), .ZN(n9884) );
  AOI21_X1 U12541 ( .B1(n9880), .B2(n14587), .A(n9879), .ZN(n9881) );
  OAI21_X1 U12542 ( .B1(n14606), .B2(n10083), .A(n9881), .ZN(n9882) );
  AOI21_X1 U12543 ( .B1(n14602), .B2(n12052), .A(n9882), .ZN(n9883) );
  OAI21_X1 U12544 ( .B1(n9884), .B2(n14598), .A(n9883), .ZN(P1_U3227) );
  OAI22_X1 U12545 ( .A1(n13073), .A2(n9943), .B1(n15213), .B2(n9885), .ZN(
        n9886) );
  AOI21_X1 U12546 ( .B1(n9939), .B2(n15213), .A(n9886), .ZN(n9887) );
  INV_X1 U12547 ( .A(n9887), .ZN(P3_U3459) );
  NAND2_X1 U12548 ( .A1(n9888), .A2(n12436), .ZN(n9897) );
  AOI21_X1 U12549 ( .B1(n9889), .B2(n9891), .A(n9890), .ZN(n9896) );
  OAI22_X1 U12550 ( .A1(n9892), .A2(n12446), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n7740), .ZN(n9894) );
  OAI22_X1 U12551 ( .A1(n15135), .A2(n12442), .B1(n10501), .B2(n12368), .ZN(
        n9893) );
  AOI211_X1 U12552 ( .C1(n7740), .C2(n12451), .A(n9894), .B(n9893), .ZN(n9895)
         );
  OAI21_X1 U12553 ( .B1(n9897), .B2(n9896), .A(n9895), .ZN(P3_U3158) );
  INV_X1 U12554 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15107) );
  OAI21_X1 U12555 ( .B1(n9899), .B2(n9898), .A(n9889), .ZN(n9900) );
  NAND2_X1 U12556 ( .A1(n9900), .A2(n12436), .ZN(n9903) );
  OAI22_X1 U12557 ( .A1(n15111), .A2(n12368), .B1(n12446), .B2(n15106), .ZN(
        n9901) );
  AOI21_X1 U12558 ( .B1(n11899), .B2(n12719), .A(n9901), .ZN(n9902) );
  OAI211_X1 U12559 ( .C1(n9904), .C2(n15107), .A(n9903), .B(n9902), .ZN(
        P3_U3177) );
  OAI21_X1 U12560 ( .B1(n9906), .B2(n9908), .A(n9905), .ZN(n10077) );
  AOI211_X1 U12561 ( .C1(n12064), .C2(n10052), .A(n14661), .B(n10024), .ZN(
        n10076) );
  XNOR2_X1 U12562 ( .A(n9907), .B(n9908), .ZN(n9912) );
  OAI22_X1 U12563 ( .A1(n9910), .A2(n14170), .B1(n9909), .B2(n14260), .ZN(
        n10194) );
  INV_X1 U12564 ( .A(n10194), .ZN(n9911) );
  OAI21_X1 U12565 ( .B1(n9912), .B2(n14656), .A(n9911), .ZN(n10073) );
  AOI211_X1 U12566 ( .C1(n14752), .C2(n10077), .A(n10076), .B(n10073), .ZN(
        n9916) );
  INV_X1 U12567 ( .A(n14273), .ZN(n14245) );
  AOI22_X1 U12568 ( .A1(n12064), .A2(n14245), .B1(n14761), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n9913) );
  OAI21_X1 U12569 ( .B1(n9916), .B2(n14761), .A(n9913), .ZN(P1_U3535) );
  INV_X1 U12570 ( .A(n12064), .ZN(n10197) );
  OAI22_X1 U12571 ( .A1(n10197), .A2(n14318), .B1(n14755), .B2(n8443), .ZN(
        n9914) );
  INV_X1 U12572 ( .A(n9914), .ZN(n9915) );
  OAI21_X1 U12573 ( .B1(n9916), .B2(n14753), .A(n9915), .ZN(P1_U3480) );
  INV_X1 U12574 ( .A(n9917), .ZN(n9919) );
  AND2_X1 U12575 ( .A1(n9919), .A2(n9918), .ZN(n9920) );
  INV_X1 U12576 ( .A(n9922), .ZN(n9923) );
  NAND2_X1 U12577 ( .A1(n12023), .A2(n12205), .ZN(n9925) );
  AOI21_X1 U12578 ( .B1(n14176), .B2(n14165), .A(n14670), .ZN(n9933) );
  NAND3_X1 U12579 ( .A1(n12210), .A2(n9926), .A3(n9975), .ZN(n9928) );
  OAI22_X1 U12580 ( .A1(n14678), .A2(n9928), .B1(n9927), .B2(n14665), .ZN(
        n9930) );
  NAND2_X1 U12581 ( .A1(n14668), .A2(n14079), .ZN(n14183) );
  NOR2_X1 U12582 ( .A1(n14183), .A2(n11962), .ZN(n9929) );
  AOI211_X1 U12583 ( .C1(n14678), .C2(P1_REG2_REG_0__SCAN_IN), .A(n9930), .B(
        n9929), .ZN(n9931) );
  OAI21_X1 U12584 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(P1_U3293) );
  NAND2_X1 U12585 ( .A1(n9934), .A2(n9937), .ZN(n9935) );
  NOR2_X1 U12586 ( .A1(n15137), .A2(n15182), .ZN(n9938) );
  MUX2_X1 U12587 ( .A(n9939), .B(P3_REG2_REG_0__SCAN_IN), .S(n15146), .Z(n9945) );
  NAND2_X1 U12588 ( .A1(n15137), .A2(n15193), .ZN(n9940) );
  OAI22_X1 U12589 ( .A1(n12998), .A2(n9943), .B1(n15108), .B2(n9942), .ZN(
        n9944) );
  OR2_X1 U12590 ( .A1(n9945), .A2(n9944), .ZN(P3_U3233) );
  OAI21_X1 U12591 ( .B1(n9947), .B2(n12211), .A(n9946), .ZN(n14717) );
  INV_X1 U12592 ( .A(n14087), .ZN(n14660) );
  NAND2_X1 U12593 ( .A1(n14717), .A2(n14660), .ZN(n9956) );
  OAI21_X1 U12594 ( .B1(n9950), .B2(n9949), .A(n9948), .ZN(n9954) );
  NAND2_X1 U12595 ( .A1(n9350), .A2(n14082), .ZN(n9952) );
  NAND2_X1 U12596 ( .A1(n13838), .A2(n14079), .ZN(n9951) );
  NAND2_X1 U12597 ( .A1(n9952), .A2(n9951), .ZN(n9953) );
  AOI21_X1 U12598 ( .B1(n9954), .B2(n14144), .A(n9953), .ZN(n9955) );
  AND2_X1 U12599 ( .A1(n9956), .A2(n9955), .ZN(n14719) );
  OAI211_X1 U12600 ( .C1(n9994), .C2(n14714), .A(n9957), .B(n14176), .ZN(
        n14713) );
  OAI22_X1 U12601 ( .A1(n14673), .A2(n14713), .B1(n9958), .B2(n14665), .ZN(
        n9960) );
  NOR2_X1 U12602 ( .A1(n14668), .A2(n9129), .ZN(n9959) );
  AOI211_X1 U12603 ( .C1(n14670), .C2(n9961), .A(n9960), .B(n9959), .ZN(n9964)
         );
  NAND2_X1 U12604 ( .A1(n9962), .A2(n14114), .ZN(n12199) );
  OR2_X1 U12605 ( .A1(n14678), .A2(n12199), .ZN(n14097) );
  INV_X1 U12606 ( .A(n14097), .ZN(n14675) );
  NAND2_X1 U12607 ( .A1(n14717), .A2(n14675), .ZN(n9963) );
  OAI211_X1 U12608 ( .C1(n14678), .C2(n14719), .A(n9964), .B(n9963), .ZN(
        P1_U3291) );
  MUX2_X1 U12609 ( .A(n9966), .B(n9965), .S(n14668), .Z(n9970) );
  OAI22_X1 U12610 ( .A1(n14673), .A2(n9967), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n14665), .ZN(n9968) );
  AOI21_X1 U12611 ( .B1(n14670), .B2(n6883), .A(n9968), .ZN(n9969) );
  OAI211_X1 U12612 ( .C1(n9971), .C2(n14097), .A(n9970), .B(n9969), .ZN(
        P1_U3290) );
  OAI21_X1 U12613 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(n14727) );
  INV_X1 U12614 ( .A(n14727), .ZN(n9989) );
  NAND2_X1 U12615 ( .A1(n12324), .A2(n9975), .ZN(n9976) );
  OAI21_X1 U12616 ( .B1(n9978), .B2(n12213), .A(n9977), .ZN(n9979) );
  NAND2_X1 U12617 ( .A1(n9979), .A2(n14144), .ZN(n14725) );
  INV_X1 U12618 ( .A(n14725), .ZN(n9980) );
  OAI21_X1 U12619 ( .B1(n9980), .B2(n14721), .A(n14668), .ZN(n9988) );
  NAND2_X1 U12620 ( .A1(n9981), .A2(n14176), .ZN(n9983) );
  OR2_X1 U12621 ( .A1(n9983), .A2(n9982), .ZN(n14723) );
  NOR2_X1 U12622 ( .A1(n14723), .A2(n14673), .ZN(n9986) );
  OAI22_X1 U12623 ( .A1(n14668), .A2(n9134), .B1(n9984), .B2(n14665), .ZN(
        n9985) );
  AOI211_X1 U12624 ( .C1(n14670), .C2(n14722), .A(n9986), .B(n9985), .ZN(n9987) );
  OAI211_X1 U12625 ( .C1(n9989), .C2(n14167), .A(n9988), .B(n9987), .ZN(
        P1_U3289) );
  INV_X1 U12626 ( .A(n12214), .ZN(n9993) );
  INV_X1 U12627 ( .A(n9990), .ZN(n9992) );
  OAI21_X1 U12628 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(n14711) );
  INV_X1 U12629 ( .A(n14711), .ZN(n10009) );
  INV_X1 U12630 ( .A(n9994), .ZN(n9997) );
  NAND2_X1 U12631 ( .A1(n12034), .A2(n9995), .ZN(n9996) );
  NAND2_X1 U12632 ( .A1(n9997), .A2(n9996), .ZN(n10002) );
  INV_X1 U12633 ( .A(n10002), .ZN(n9998) );
  NAND2_X1 U12634 ( .A1(n9998), .A2(n14176), .ZN(n14707) );
  OAI22_X1 U12635 ( .A1(n14673), .A2(n14707), .B1(n9999), .B2(n14665), .ZN(
        n10001) );
  NOR2_X1 U12636 ( .A1(n14668), .A2(n9086), .ZN(n10000) );
  AOI211_X1 U12637 ( .C1(n14670), .C2(n12034), .A(n10001), .B(n10000), .ZN(
        n10008) );
  XNOR2_X1 U12638 ( .A(n10002), .B(n11962), .ZN(n10003) );
  MUX2_X1 U12639 ( .A(n10003), .B(n12214), .S(n13841), .Z(n10006) );
  NAND2_X1 U12640 ( .A1(n14711), .A2(n14660), .ZN(n10005) );
  AOI22_X1 U12641 ( .A1(n14082), .A2(n13841), .B1(n13839), .B2(n14079), .ZN(
        n10004) );
  OAI211_X1 U12642 ( .C1(n10006), .C2(n14656), .A(n10005), .B(n10004), .ZN(
        n14709) );
  NAND2_X1 U12643 ( .A1(n14709), .A2(n14668), .ZN(n10007) );
  OAI211_X1 U12644 ( .C1(n10009), .C2(n14097), .A(n10008), .B(n10007), .ZN(
        P1_U3292) );
  NAND2_X1 U12645 ( .A1(n6801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10011) );
  XNOR2_X1 U12646 ( .A(n10011), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13340) );
  INV_X1 U12647 ( .A(n13340), .ZN(n10013) );
  INV_X1 U12648 ( .A(n11481), .ZN(n10015) );
  OAI222_X1 U12649 ( .A1(P2_U3088), .A2(n10013), .B1(n11317), .B2(n10015), 
        .C1(n10012), .C2(n13693), .ZN(P2_U3309) );
  INV_X1 U12650 ( .A(n13959), .ZN(n11057) );
  OAI222_X1 U12651 ( .A1(P1_U3086), .A2(n11057), .B1(n14330), .B2(n10015), 
        .C1(n10014), .C2(n14332), .ZN(P1_U3337) );
  OAI21_X1 U12652 ( .B1(n10017), .B2(n10019), .A(n10016), .ZN(n10070) );
  INV_X1 U12653 ( .A(n10070), .ZN(n10028) );
  AOI21_X1 U12654 ( .B1(n10018), .B2(n10019), .A(n14656), .ZN(n10023) );
  NAND2_X1 U12655 ( .A1(n13834), .A2(n14082), .ZN(n10021) );
  NAND2_X1 U12656 ( .A1(n13832), .A2(n14079), .ZN(n10020) );
  NAND2_X1 U12657 ( .A1(n10021), .A2(n10020), .ZN(n10437) );
  AOI21_X1 U12658 ( .B1(n10023), .B2(n10022), .A(n10437), .ZN(n10072) );
  INV_X1 U12659 ( .A(n10024), .ZN(n10026) );
  INV_X1 U12660 ( .A(n14662), .ZN(n10025) );
  AOI21_X1 U12661 ( .B1(n12067), .B2(n10026), .A(n10025), .ZN(n10064) );
  AOI22_X1 U12662 ( .A1(n10064), .A2(n14176), .B1(n14743), .B2(n12067), .ZN(
        n10027) );
  OAI211_X1 U12663 ( .C1(n10028), .C2(n14280), .A(n10072), .B(n10027), .ZN(
        n10030) );
  NAND2_X1 U12664 ( .A1(n10030), .A2(n14764), .ZN(n10029) );
  OAI21_X1 U12665 ( .B1(n14764), .B2(n9197), .A(n10029), .ZN(P1_U3536) );
  INV_X1 U12666 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10032) );
  NAND2_X1 U12667 ( .A1(n10030), .A2(n14755), .ZN(n10031) );
  OAI21_X1 U12668 ( .B1(n14755), .B2(n10032), .A(n10031), .ZN(P1_U3483) );
  OAI21_X2 U12669 ( .B1(n10035), .B2(n10034), .A(n10033), .ZN(n10039) );
  AND2_X1 U12670 ( .A1(n13835), .A2(n12322), .ZN(n10036) );
  AOI21_X1 U12671 ( .B1(n12056), .B2(n12323), .A(n10036), .ZN(n10186) );
  AOI22_X1 U12672 ( .A1(n12056), .A2(n12326), .B1(n12323), .B2(n13835), .ZN(
        n10037) );
  XNOR2_X1 U12673 ( .A(n10037), .B(n12324), .ZN(n10185) );
  XOR2_X1 U12674 ( .A(n10186), .B(n10185), .Z(n10038) );
  NAND2_X1 U12675 ( .A1(n10039), .A2(n10038), .ZN(n10184) );
  OAI211_X1 U12676 ( .C1(n10039), .C2(n10038), .A(n10184), .B(n14585), .ZN(
        n10045) );
  OAI22_X1 U12677 ( .A1(n10041), .A2(n14170), .B1(n10040), .B2(n14260), .ZN(
        n10059) );
  NOR2_X1 U12678 ( .A1(n14606), .A2(n10054), .ZN(n10042) );
  AOI211_X1 U12679 ( .C1(n14587), .C2(n10059), .A(n10043), .B(n10042), .ZN(
        n10044) );
  OAI211_X1 U12680 ( .C1(n14732), .C2(n13792), .A(n10045), .B(n10044), .ZN(
        P1_U3239) );
  INV_X1 U12681 ( .A(n10046), .ZN(n10048) );
  OAI222_X1 U12682 ( .A1(P3_U3151), .A2(n10049), .B1(n11060), .B2(n10048), 
        .C1(n10047), .C2(n12350), .ZN(P3_U3275) );
  OAI21_X1 U12683 ( .B1(n10051), .B2(n12218), .A(n10050), .ZN(n14734) );
  OAI211_X1 U12684 ( .C1(n14732), .C2(n10053), .A(n14176), .B(n10052), .ZN(
        n14729) );
  NOR2_X1 U12685 ( .A1(n14729), .A2(n14673), .ZN(n10056) );
  OAI22_X1 U12686 ( .A1(n14732), .A2(n14156), .B1(n10054), .B2(n14665), .ZN(
        n10055) );
  AOI211_X1 U12687 ( .C1(n14734), .C2(n14188), .A(n10056), .B(n10055), .ZN(
        n10063) );
  XNOR2_X1 U12688 ( .A(n10058), .B(n10057), .ZN(n10060) );
  AOI21_X1 U12689 ( .B1(n10060), .B2(n14144), .A(n10059), .ZN(n14730) );
  MUX2_X1 U12690 ( .A(n10061), .B(n14730), .S(n14668), .Z(n10062) );
  NAND2_X1 U12691 ( .A1(n10063), .A2(n10062), .ZN(P1_U3287) );
  NAND3_X1 U12692 ( .A1(n10064), .A2(n14176), .A3(n14165), .ZN(n10067) );
  INV_X1 U12693 ( .A(n10439), .ZN(n10065) );
  INV_X1 U12694 ( .A(n14665), .ZN(n14180) );
  AOI22_X1 U12695 ( .A1(n14678), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n10065), 
        .B2(n14180), .ZN(n10066) );
  OAI211_X1 U12696 ( .C1(n10068), .C2(n14156), .A(n10067), .B(n10066), .ZN(
        n10069) );
  AOI21_X1 U12697 ( .B1(n10070), .B2(n14188), .A(n10069), .ZN(n10071) );
  OAI21_X1 U12698 ( .B1(n14678), .B2(n10072), .A(n10071), .ZN(P1_U3285) );
  INV_X1 U12699 ( .A(n10073), .ZN(n10080) );
  NOR2_X1 U12700 ( .A1(n10197), .A2(n14156), .ZN(n10075) );
  OAI22_X1 U12701 ( .A1(n14668), .A2(n9205), .B1(n10192), .B2(n14665), .ZN(
        n10074) );
  AOI211_X1 U12702 ( .C1(n10076), .C2(n14165), .A(n10075), .B(n10074), .ZN(
        n10079) );
  NAND2_X1 U12703 ( .A1(n10077), .A2(n14188), .ZN(n10078) );
  OAI211_X1 U12704 ( .C1(n10080), .C2(n14678), .A(n10079), .B(n10078), .ZN(
        P1_U3286) );
  INV_X1 U12705 ( .A(n10081), .ZN(n10090) );
  NOR2_X1 U12706 ( .A1(n14156), .A2(n10082), .ZN(n10085) );
  OAI22_X1 U12707 ( .A1(n14668), .A2(n9135), .B1(n10083), .B2(n14665), .ZN(
        n10084) );
  AOI211_X1 U12708 ( .C1(n10086), .C2(n14165), .A(n10085), .B(n10084), .ZN(
        n10089) );
  NAND2_X1 U12709 ( .A1(n10087), .A2(n14188), .ZN(n10088) );
  OAI211_X1 U12710 ( .C1(n10090), .C2(n14678), .A(n10089), .B(n10088), .ZN(
        P1_U3288) );
  NAND2_X1 U12711 ( .A1(n11358), .A2(n11354), .ZN(n10091) );
  INV_X1 U12712 ( .A(n13299), .ZN(n11367) );
  XNOR2_X1 U12713 ( .A(n11370), .B(n11367), .ZN(n11725) );
  OR2_X1 U12714 ( .A1(n11370), .A2(n13299), .ZN(n10093) );
  XNOR2_X1 U12715 ( .A(n14874), .B(n11384), .ZN(n11726) );
  XNOR2_X1 U12716 ( .A(n10161), .B(n11726), .ZN(n14872) );
  INV_X1 U12717 ( .A(n14872), .ZN(n10115) );
  AND2_X1 U12718 ( .A1(n10094), .A2(n11767), .ZN(n14853) );
  NOR3_X1 U12719 ( .A1(n10097), .A2(n10096), .A3(n10095), .ZN(n10098) );
  NAND2_X1 U12720 ( .A1(n14853), .A2(n10098), .ZN(n10099) );
  AND2_X1 U12721 ( .A1(n13647), .A2(n11321), .ZN(n10100) );
  OR2_X1 U12722 ( .A1(n10458), .A2(n11370), .ZN(n10459) );
  NAND2_X1 U12723 ( .A1(n10459), .A2(n14874), .ZN(n10101) );
  NAND2_X1 U12724 ( .A1(n10101), .A2(n10936), .ZN(n10102) );
  OR2_X1 U12725 ( .A1(n10102), .A2(n10445), .ZN(n14875) );
  INV_X1 U12726 ( .A(n14875), .ZN(n10106) );
  OAI22_X1 U12727 ( .A1(n13528), .A2(n10162), .B1(n15592), .B2(n10104), .ZN(
        n10105) );
  AOI21_X1 U12728 ( .B1(n15590), .B2(n10106), .A(n10105), .ZN(n10114) );
  INV_X1 U12729 ( .A(n11354), .ZN(n13164) );
  NAND2_X1 U12730 ( .A1(n13164), .A2(n11358), .ZN(n10463) );
  NAND2_X1 U12731 ( .A1(n10464), .A2(n10463), .ZN(n10108) );
  INV_X1 U12732 ( .A(n11725), .ZN(n10107) );
  NAND2_X1 U12733 ( .A1(n10108), .A2(n10107), .ZN(n10466) );
  NAND2_X1 U12734 ( .A1(n11370), .A2(n11367), .ZN(n10109) );
  NAND2_X1 U12735 ( .A1(n10466), .A2(n10109), .ZN(n10168) );
  INV_X1 U12736 ( .A(n11726), .ZN(n10110) );
  XNOR2_X1 U12737 ( .A(n10168), .B(n10110), .ZN(n10112) );
  AOI21_X1 U12738 ( .B1(n10112), .B2(n13521), .A(n10111), .ZN(n14877) );
  MUX2_X1 U12739 ( .A(n9105), .B(n14877), .S(n13441), .Z(n10113) );
  OAI211_X1 U12740 ( .C1(n10115), .C2(n13496), .A(n10114), .B(n10113), .ZN(
        P2_U3260) );
  NAND2_X1 U12741 ( .A1(n10116), .A2(n6652), .ZN(n10119) );
  AOI22_X1 U12742 ( .A1(n11683), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11490), 
        .B2(n10117), .ZN(n10118) );
  NAND2_X1 U12743 ( .A1(n11686), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n10127) );
  NAND2_X1 U12744 ( .A1(n11642), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U12745 ( .A1(n10121), .A2(n10120), .ZN(n10122) );
  NAND2_X1 U12746 ( .A1(n10213), .A2(n10122), .ZN(n10295) );
  INV_X1 U12747 ( .A(n10295), .ZN(n10123) );
  NAND2_X1 U12748 ( .A1(n11658), .A2(n10123), .ZN(n10125) );
  OR2_X1 U12749 ( .A1(n11605), .A2(n9173), .ZN(n10124) );
  NAND4_X1 U12750 ( .A1(n10127), .A2(n10126), .A3(n10125), .A4(n10124), .ZN(
        n13295) );
  AOI22_X1 U12751 ( .A1(n13650), .A2(n13295), .B1(n13297), .B2(n13470), .ZN(
        n10173) );
  NAND2_X1 U12752 ( .A1(n13219), .A2(n10178), .ZN(n10128) );
  OAI211_X1 U12753 ( .C1(n13217), .C2(n10173), .A(n10129), .B(n10128), .ZN(
        n10138) );
  INV_X1 U12754 ( .A(n10130), .ZN(n10131) );
  XNOR2_X1 U12755 ( .A(n14887), .B(n12012), .ZN(n10134) );
  AND2_X1 U12756 ( .A1(n13296), .A2(n10208), .ZN(n10133) );
  NAND2_X1 U12757 ( .A1(n10134), .A2(n10133), .ZN(n10205) );
  OAI21_X1 U12758 ( .B1(n10134), .B2(n10133), .A(n10205), .ZN(n10135) );
  AOI211_X1 U12759 ( .C1(n10136), .C2(n10135), .A(n13275), .B(n10207), .ZN(
        n10137) );
  AOI211_X1 U12760 ( .C1(n14887), .C2(n13273), .A(n10138), .B(n10137), .ZN(
        n10139) );
  INV_X1 U12761 ( .A(n10139), .ZN(P2_U3185) );
  INV_X1 U12762 ( .A(n10140), .ZN(n10142) );
  OAI222_X1 U12763 ( .A1(n11060), .A2(n10142), .B1(n12350), .B2(n10141), .C1(
        P3_U3151), .C2(n10250), .ZN(P3_U3274) );
  INV_X1 U12764 ( .A(n15596), .ZN(n10497) );
  INV_X1 U12765 ( .A(n10143), .ZN(n10144) );
  AOI22_X1 U12766 ( .A1(n15590), .A2(n10145), .B1(n10497), .B2(n10144), .ZN(
        n10150) );
  INV_X1 U12767 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10146) );
  OAI22_X1 U12768 ( .A1(n13441), .A2(n10147), .B1(n10146), .B2(n15592), .ZN(
        n10148) );
  AOI21_X1 U12769 ( .B1(n14557), .B2(n13179), .A(n10148), .ZN(n10149) );
  OAI211_X1 U12770 ( .C1(n10151), .C2(n14556), .A(n10150), .B(n10149), .ZN(
        P2_U3264) );
  INV_X1 U12771 ( .A(n10152), .ZN(n10153) );
  AOI21_X1 U12772 ( .B1(n10155), .B2(n10154), .A(n10153), .ZN(n10159) );
  NAND2_X1 U12773 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n14966) );
  OAI21_X1 U12774 ( .B1(n15160), .B2(n12446), .A(n14966), .ZN(n10157) );
  OAI22_X1 U12775 ( .A1(n15111), .A2(n12442), .B1(n10405), .B2(n12368), .ZN(
        n10156) );
  AOI211_X1 U12776 ( .C1(n10251), .C2(n12451), .A(n10157), .B(n10156), .ZN(
        n10158) );
  OAI21_X1 U12777 ( .B1(n10159), .B2(n12459), .A(n10158), .ZN(P3_U3170) );
  NAND2_X1 U12778 ( .A1(n14874), .A2(n13298), .ZN(n10160) );
  NAND2_X1 U12779 ( .A1(n10162), .A2(n11384), .ZN(n10163) );
  NAND2_X1 U12780 ( .A1(n10164), .A2(n10163), .ZN(n10443) );
  INV_X1 U12781 ( .A(n11727), .ZN(n10165) );
  NAND2_X1 U12782 ( .A1(n10443), .A2(n10165), .ZN(n10167) );
  OR2_X1 U12783 ( .A1(n11392), .A2(n13297), .ZN(n10166) );
  NAND2_X1 U12784 ( .A1(n10167), .A2(n10166), .ZN(n10260) );
  XNOR2_X1 U12785 ( .A(n14887), .B(n13296), .ZN(n11728) );
  XNOR2_X1 U12786 ( .A(n10260), .B(n11728), .ZN(n14891) );
  OAI21_X1 U12787 ( .B1(n10168), .B2(n11384), .A(n14874), .ZN(n10170) );
  NAND2_X1 U12788 ( .A1(n10168), .A2(n11384), .ZN(n10169) );
  NAND2_X1 U12789 ( .A1(n10170), .A2(n10169), .ZN(n10448) );
  NAND2_X1 U12790 ( .A1(n10448), .A2(n11727), .ZN(n10172) );
  INV_X1 U12791 ( .A(n13297), .ZN(n11389) );
  NAND2_X1 U12792 ( .A1(n11392), .A2(n11389), .ZN(n10171) );
  XNOR2_X1 U12793 ( .A(n10276), .B(n11728), .ZN(n10175) );
  INV_X1 U12794 ( .A(n10173), .ZN(n10174) );
  AOI21_X1 U12795 ( .B1(n10175), .B2(n13521), .A(n10174), .ZN(n14888) );
  MUX2_X1 U12796 ( .A(n10176), .B(n14888), .S(n13441), .Z(n10183) );
  INV_X1 U12797 ( .A(n10177), .ZN(n10444) );
  INV_X1 U12798 ( .A(n14887), .ZN(n10180) );
  AOI211_X1 U12799 ( .C1(n14887), .C2(n10444), .A(n13459), .B(n6809), .ZN(
        n14886) );
  INV_X1 U12800 ( .A(n10178), .ZN(n10179) );
  OAI22_X1 U12801 ( .A1(n10180), .A2(n13528), .B1(n15592), .B2(n10179), .ZN(
        n10181) );
  AOI21_X1 U12802 ( .B1(n14886), .B2(n15590), .A(n10181), .ZN(n10182) );
  OAI211_X1 U12803 ( .C1(n13496), .C2(n14891), .A(n10183), .B(n10182), .ZN(
        P2_U3258) );
  AND2_X1 U12804 ( .A1(n13834), .A2(n12322), .ZN(n10187) );
  AOI21_X1 U12805 ( .B1(n12064), .B2(n12323), .A(n10187), .ZN(n10430) );
  AOI22_X1 U12806 ( .A1(n12064), .A2(n12326), .B1(n12323), .B2(n13834), .ZN(
        n10188) );
  XNOR2_X1 U12807 ( .A(n10188), .B(n12324), .ZN(n10429) );
  XOR2_X1 U12808 ( .A(n10430), .B(n10429), .Z(n10189) );
  OAI211_X1 U12809 ( .C1(n10190), .C2(n10189), .A(n10434), .B(n14585), .ZN(
        n10196) );
  NOR2_X1 U12810 ( .A1(n10191), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13901) );
  NOR2_X1 U12811 ( .A1(n14606), .A2(n10192), .ZN(n10193) );
  AOI211_X1 U12812 ( .C1(n14587), .C2(n10194), .A(n13901), .B(n10193), .ZN(
        n10195) );
  OAI211_X1 U12813 ( .C1(n10197), .C2(n13792), .A(n10196), .B(n10195), .ZN(
        P1_U3213) );
  INV_X1 U12814 ( .A(n11489), .ZN(n10199) );
  OAI222_X1 U12815 ( .A1(n13693), .A2(n10198), .B1(n11317), .B2(n10199), .C1(
        n13349), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U12816 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10200) );
  OAI222_X1 U12817 ( .A1(n14332), .A2(n10200), .B1(n14330), .B2(n10199), .C1(
        P1_U3086), .C2(n8775), .ZN(P1_U3336) );
  NAND2_X1 U12818 ( .A1(n10201), .A2(n6652), .ZN(n10204) );
  AOI22_X1 U12819 ( .A1(n11683), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11490), 
        .B2(n10202), .ZN(n10203) );
  XNOR2_X1 U12820 ( .A(n12012), .B(n11411), .ZN(n10328) );
  NAND2_X1 U12821 ( .A1(n13295), .A2(n10208), .ZN(n10329) );
  XNOR2_X1 U12822 ( .A(n10328), .B(n10329), .ZN(n10209) );
  OAI21_X1 U12823 ( .B1(n10210), .B2(n10209), .A(n10333), .ZN(n10211) );
  NAND2_X1 U12824 ( .A1(n10211), .A2(n13249), .ZN(n10222) );
  NAND2_X1 U12825 ( .A1(n11686), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U12826 ( .A1(n11642), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10217) );
  AND2_X1 U12827 ( .A1(n10213), .A2(n10212), .ZN(n10214) );
  NOR2_X1 U12828 ( .A1(n10269), .A2(n10214), .ZN(n10281) );
  NAND2_X1 U12829 ( .A1(n11658), .A2(n10281), .ZN(n10216) );
  OR2_X1 U12830 ( .A1(n11605), .A2(n9242), .ZN(n10215) );
  NAND4_X1 U12831 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n13294) );
  INV_X1 U12832 ( .A(n13294), .ZN(n11419) );
  OAI22_X1 U12833 ( .A1(n13258), .A2(n11419), .B1(n13270), .B2(n10295), .ZN(
        n10219) );
  AOI211_X1 U12834 ( .C1(n13244), .C2(n13296), .A(n10220), .B(n10219), .ZN(
        n10221) );
  OAI211_X1 U12835 ( .C1(n7056), .C2(n13242), .A(n10222), .B(n10221), .ZN(
        P2_U3193) );
  OAI21_X1 U12836 ( .B1(n10224), .B2(n10227), .A(n10223), .ZN(n14864) );
  OAI22_X1 U12837 ( .A1(n11337), .A2(n13538), .B1(n11358), .B2(n13540), .ZN(
        n10231) );
  NAND3_X1 U12838 ( .A1(n10227), .A2(n10226), .A3(n10225), .ZN(n10229) );
  INV_X1 U12839 ( .A(n13521), .ZN(n14548) );
  AOI21_X1 U12840 ( .B1(n10229), .B2(n10228), .A(n14548), .ZN(n10230) );
  AOI211_X1 U12841 ( .C1(n14873), .C2(n14864), .A(n10231), .B(n10230), .ZN(
        n14861) );
  NAND2_X1 U12842 ( .A1(n10232), .A2(n13246), .ZN(n10233) );
  NAND2_X1 U12843 ( .A1(n10233), .A2(n10936), .ZN(n10235) );
  OR2_X1 U12844 ( .A1(n10235), .A2(n10234), .ZN(n14860) );
  NOR2_X1 U12845 ( .A1(n13550), .A2(n14860), .ZN(n10239) );
  INV_X1 U12846 ( .A(n15592), .ZN(n14555) );
  AOI22_X1 U12847 ( .A1(n14556), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14555), .ZN(n10237) );
  OAI21_X1 U12848 ( .B1(n13528), .B2(n9646), .A(n10237), .ZN(n10238) );
  AOI211_X1 U12849 ( .C1(n10497), .C2(n14864), .A(n10239), .B(n10238), .ZN(
        n10240) );
  OAI21_X1 U12850 ( .B1(n14556), .B2(n14861), .A(n10240), .ZN(P2_U3263) );
  NAND2_X1 U12851 ( .A1(n12720), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10241) );
  OAI21_X1 U12852 ( .B1(n12354), .B2(n12720), .A(n10241), .ZN(P3_U3519) );
  OAI22_X1 U12853 ( .A1(n12694), .A2(P3_U3151), .B1(SI_22_), .B2(n12350), .ZN(
        n10242) );
  AOI21_X1 U12854 ( .B1(n10243), .B2(n13135), .A(n10242), .ZN(P3_U3273) );
  XNOR2_X1 U12855 ( .A(n10244), .B(n12501), .ZN(n15161) );
  NAND2_X1 U12856 ( .A1(n10503), .A2(n10245), .ZN(n10246) );
  XNOR2_X1 U12857 ( .A(n10246), .B(n8097), .ZN(n10248) );
  OAI22_X1 U12858 ( .A1(n15111), .A2(n15134), .B1(n10405), .B2(n15136), .ZN(
        n10247) );
  AOI21_X1 U12859 ( .B1(n10248), .B2(n12987), .A(n10247), .ZN(n10249) );
  OAI21_X1 U12860 ( .B1(n12868), .B2(n15161), .A(n10249), .ZN(n15163) );
  INV_X1 U12861 ( .A(n15163), .ZN(n10258) );
  INV_X1 U12862 ( .A(n15161), .ZN(n10256) );
  NOR2_X1 U12863 ( .A1(n15137), .A2(n10250), .ZN(n15122) );
  NAND2_X1 U12864 ( .A1(n15144), .A2(n15122), .ZN(n12848) );
  INV_X1 U12865 ( .A(n12848), .ZN(n12874) );
  AOI22_X1 U12866 ( .A1(n14528), .A2(n10252), .B1(n15140), .B2(n10251), .ZN(
        n10253) );
  OAI21_X1 U12867 ( .B1(n10254), .B2(n15144), .A(n10253), .ZN(n10255) );
  AOI21_X1 U12868 ( .B1(n10256), .B2(n12874), .A(n10255), .ZN(n10257) );
  OAI21_X1 U12869 ( .B1(n10258), .B2(n15146), .A(n10257), .ZN(P3_U3229) );
  INV_X1 U12870 ( .A(n11728), .ZN(n10259) );
  OR2_X1 U12871 ( .A1(n14887), .A2(n13296), .ZN(n10261) );
  INV_X1 U12872 ( .A(n13295), .ZN(n11408) );
  XNOR2_X1 U12873 ( .A(n11411), .B(n11408), .ZN(n11732) );
  INV_X1 U12874 ( .A(n11732), .ZN(n10287) );
  NAND2_X1 U12875 ( .A1(n11411), .A2(n13295), .ZN(n10262) );
  OR2_X1 U12876 ( .A1(n10263), .A2(n11572), .ZN(n10266) );
  AOI22_X1 U12877 ( .A1(n11683), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n11490), 
        .B2(n10264), .ZN(n10265) );
  XNOR2_X1 U12878 ( .A(n11417), .B(n13294), .ZN(n11730) );
  OR2_X1 U12879 ( .A1(n10267), .A2(n10277), .ZN(n10268) );
  NAND2_X1 U12880 ( .A1(n10350), .A2(n10268), .ZN(n14900) );
  NAND2_X1 U12881 ( .A1(n11686), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10274) );
  OR2_X1 U12882 ( .A1(n10269), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10270) );
  NAND2_X1 U12883 ( .A1(n10269), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10357) );
  AND2_X1 U12884 ( .A1(n10270), .A2(n10357), .ZN(n10366) );
  NAND2_X1 U12885 ( .A1(n11658), .A2(n10366), .ZN(n10273) );
  NAND2_X1 U12886 ( .A1(n11642), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10272) );
  OR2_X1 U12887 ( .A1(n11605), .A2(n9326), .ZN(n10271) );
  NAND4_X1 U12888 ( .A1(n10274), .A2(n10273), .A3(n10272), .A4(n10271), .ZN(
        n13293) );
  AOI22_X1 U12889 ( .A1(n13650), .A2(n13293), .B1(n13295), .B2(n13470), .ZN(
        n10280) );
  INV_X1 U12890 ( .A(n13296), .ZN(n11399) );
  AND2_X1 U12891 ( .A1(n14887), .A2(n11399), .ZN(n10275) );
  XNOR2_X1 U12892 ( .A(n10354), .B(n10277), .ZN(n10278) );
  NAND2_X1 U12893 ( .A1(n10278), .A2(n13521), .ZN(n10279) );
  OAI211_X1 U12894 ( .C1(n14900), .C2(n13647), .A(n10280), .B(n10279), .ZN(
        n14903) );
  NAND2_X1 U12895 ( .A1(n14903), .A2(n13441), .ZN(n10286) );
  INV_X1 U12896 ( .A(n10281), .ZN(n10336) );
  OAI22_X1 U12897 ( .A1(n13441), .A2(n9242), .B1(n10336), .B2(n15592), .ZN(
        n10284) );
  INV_X1 U12898 ( .A(n10296), .ZN(n10282) );
  INV_X1 U12899 ( .A(n11417), .ZN(n14902) );
  OAI211_X1 U12900 ( .C1(n10282), .C2(n14902), .A(n10936), .B(n10367), .ZN(
        n14901) );
  NOR2_X1 U12901 ( .A1(n14901), .A2(n13550), .ZN(n10283) );
  AOI211_X1 U12902 ( .C1(n14557), .C2(n11417), .A(n10284), .B(n10283), .ZN(
        n10285) );
  OAI211_X1 U12903 ( .C1(n14900), .C2(n15596), .A(n10286), .B(n10285), .ZN(
        P2_U3256) );
  NAND2_X1 U12904 ( .A1(n10288), .A2(n10287), .ZN(n10289) );
  NAND2_X1 U12905 ( .A1(n10290), .A2(n10289), .ZN(n14894) );
  AOI22_X1 U12906 ( .A1(n13650), .A2(n13294), .B1(n13296), .B2(n13470), .ZN(
        n10294) );
  XNOR2_X1 U12907 ( .A(n10291), .B(n11732), .ZN(n10292) );
  NAND2_X1 U12908 ( .A1(n10292), .A2(n13521), .ZN(n10293) );
  OAI211_X1 U12909 ( .C1(n14894), .C2(n13647), .A(n10294), .B(n10293), .ZN(
        n14896) );
  NAND2_X1 U12910 ( .A1(n14896), .A2(n13441), .ZN(n10300) );
  OAI22_X1 U12911 ( .A1(n13441), .A2(n9173), .B1(n10295), .B2(n15592), .ZN(
        n10298) );
  OAI211_X1 U12912 ( .C1(n6809), .C2(n7056), .A(n10936), .B(n10296), .ZN(
        n14895) );
  NOR2_X1 U12913 ( .A1(n14895), .A2(n13550), .ZN(n10297) );
  AOI211_X1 U12914 ( .C1(n14557), .C2(n11411), .A(n10298), .B(n10297), .ZN(
        n10299) );
  OAI211_X1 U12915 ( .C1(n14894), .C2(n15596), .A(n10300), .B(n10299), .ZN(
        P2_U3257) );
  AOI21_X1 U12916 ( .B1(n10301), .B2(n12224), .A(n14656), .ZN(n10303) );
  AND2_X1 U12917 ( .A1(n10303), .A2(n10302), .ZN(n14749) );
  NAND2_X1 U12918 ( .A1(n13832), .A2(n14082), .ZN(n14747) );
  INV_X1 U12919 ( .A(n14747), .ZN(n10306) );
  AOI21_X1 U12920 ( .B1(n14744), .B2(n14663), .A(n14661), .ZN(n10304) );
  NAND2_X1 U12921 ( .A1(n10304), .A2(n10420), .ZN(n14748) );
  NAND2_X1 U12922 ( .A1(n13830), .A2(n14079), .ZN(n14746) );
  AOI21_X1 U12923 ( .B1(n14748), .B2(n14746), .A(n14114), .ZN(n10305) );
  NOR3_X1 U12924 ( .A1(n14749), .A2(n10306), .A3(n10305), .ZN(n10313) );
  OAI21_X1 U12925 ( .B1(n10308), .B2(n12224), .A(n10307), .ZN(n14751) );
  NOR2_X1 U12926 ( .A1(n7080), .A2(n14156), .ZN(n10311) );
  OAI22_X1 U12927 ( .A1(n14668), .A2(n10309), .B1(n10845), .B2(n14665), .ZN(
        n10310) );
  AOI211_X1 U12928 ( .C1(n14751), .C2(n14188), .A(n10311), .B(n10310), .ZN(
        n10312) );
  OAI21_X1 U12929 ( .B1(n10313), .B2(n14678), .A(n10312), .ZN(P1_U3283) );
  NAND2_X1 U12930 ( .A1(n12720), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10314) );
  OAI21_X1 U12931 ( .B1(n12487), .B2(n12720), .A(n10314), .ZN(P3_U3521) );
  NOR2_X1 U12932 ( .A1(n10933), .A2(n10315), .ZN(n10317) );
  XOR2_X1 U12933 ( .A(n11063), .B(n10543), .Z(n10318) );
  NAND2_X1 U12934 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n10318), .ZN(n10544) );
  OAI211_X1 U12935 ( .C1(n10318), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14837), 
        .B(n10544), .ZN(n10326) );
  NAND2_X1 U12936 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n11074)
         );
  INV_X1 U12937 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10320) );
  OAI21_X1 U12938 ( .B1(n10321), .B2(n10320), .A(n10319), .ZN(n10550) );
  XNOR2_X1 U12939 ( .A(n10550), .B(n10327), .ZN(n10322) );
  NAND2_X1 U12940 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10322), .ZN(n10551) );
  OAI211_X1 U12941 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n10322), .A(n14843), 
        .B(n10551), .ZN(n10323) );
  NAND2_X1 U12942 ( .A1(n11074), .A2(n10323), .ZN(n10324) );
  AOI21_X1 U12943 ( .B1(n14835), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n10324), 
        .ZN(n10325) );
  OAI211_X1 U12944 ( .C1(n14765), .C2(n10327), .A(n10326), .B(n10325), .ZN(
        P2_U3229) );
  INV_X1 U12945 ( .A(n10328), .ZN(n10330) );
  NAND2_X1 U12946 ( .A1(n10330), .A2(n10329), .ZN(n10331) );
  XNOR2_X1 U12947 ( .A(n11417), .B(n11995), .ZN(n10561) );
  NAND2_X1 U12948 ( .A1(n13294), .A2(n10208), .ZN(n10560) );
  XNOR2_X1 U12949 ( .A(n10561), .B(n10560), .ZN(n10332) );
  AND3_X1 U12950 ( .A1(n10333), .A2(n10332), .A3(n10331), .ZN(n10334) );
  OAI21_X1 U12951 ( .B1(n10559), .B2(n10334), .A(n13249), .ZN(n10340) );
  INV_X1 U12952 ( .A(n10335), .ZN(n10338) );
  INV_X1 U12953 ( .A(n13293), .ZN(n11421) );
  OAI22_X1 U12954 ( .A1(n13258), .A2(n11421), .B1(n13270), .B2(n10336), .ZN(
        n10337) );
  AOI211_X1 U12955 ( .C1(n13244), .C2(n13295), .A(n10338), .B(n10337), .ZN(
        n10339) );
  OAI211_X1 U12956 ( .C1(n14902), .C2(n13242), .A(n10340), .B(n10339), .ZN(
        P2_U3203) );
  INV_X1 U12957 ( .A(n10487), .ZN(n10348) );
  OAI21_X1 U12958 ( .B1(n10342), .B2(n10341), .A(n10596), .ZN(n10343) );
  NAND2_X1 U12959 ( .A1(n10343), .A2(n12436), .ZN(n10347) );
  OAI22_X1 U12960 ( .A1(n10501), .A2(n12442), .B1(n10723), .B2(n12368), .ZN(
        n10344) );
  AOI211_X1 U12961 ( .C1(n12456), .C2(n15165), .A(n10345), .B(n10344), .ZN(
        n10346) );
  OAI211_X1 U12962 ( .C1(n10348), .C2(n12418), .A(n10347), .B(n10346), .ZN(
        P3_U3167) );
  NAND2_X1 U12963 ( .A1(n11417), .A2(n13294), .ZN(n10349) );
  NAND2_X1 U12964 ( .A1(n10351), .A2(n6652), .ZN(n10353) );
  AOI22_X1 U12965 ( .A1(n11683), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n11490), 
        .B2(n14816), .ZN(n10352) );
  XOR2_X1 U12966 ( .A(n13293), .B(n11424), .Z(n11733) );
  XNOR2_X1 U12967 ( .A(n10512), .B(n11733), .ZN(n14907) );
  NAND2_X1 U12968 ( .A1(n10354), .A2(n11730), .ZN(n10356) );
  OR2_X1 U12969 ( .A1(n11417), .A2(n11419), .ZN(n10355) );
  XNOR2_X1 U12970 ( .A(n10520), .B(n11733), .ZN(n10364) );
  NAND2_X1 U12971 ( .A1(n11686), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10362) );
  NAND2_X1 U12972 ( .A1(n11642), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10361) );
  NAND2_X1 U12973 ( .A1(n10357), .A2(n15532), .ZN(n10358) );
  AND2_X1 U12974 ( .A1(n10522), .A2(n10358), .ZN(n10656) );
  NAND2_X1 U12975 ( .A1(n11658), .A2(n10656), .ZN(n10360) );
  OR2_X1 U12976 ( .A1(n11605), .A2(n9830), .ZN(n10359) );
  NAND4_X1 U12977 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n13292) );
  INV_X1 U12978 ( .A(n13292), .ZN(n11433) );
  OAI22_X1 U12979 ( .A1(n11419), .A2(n13538), .B1(n11433), .B2(n13540), .ZN(
        n10363) );
  AOI21_X1 U12980 ( .B1(n10364), .B2(n13521), .A(n10363), .ZN(n10365) );
  OAI21_X1 U12981 ( .B1(n14907), .B2(n13647), .A(n10365), .ZN(n14911) );
  NAND2_X1 U12982 ( .A1(n14911), .A2(n13441), .ZN(n10372) );
  INV_X1 U12983 ( .A(n10366), .ZN(n10564) );
  OAI22_X1 U12984 ( .A1(n13441), .A2(n9326), .B1(n10564), .B2(n15592), .ZN(
        n10370) );
  OAI211_X1 U12985 ( .C1(n14910), .C2(n10368), .A(n10936), .B(n10534), .ZN(
        n14908) );
  NOR2_X1 U12986 ( .A1(n14908), .A2(n13550), .ZN(n10369) );
  AOI211_X1 U12987 ( .C1(n14557), .C2(n11424), .A(n10370), .B(n10369), .ZN(
        n10371) );
  OAI211_X1 U12988 ( .C1(n14907), .C2(n15596), .A(n10372), .B(n10371), .ZN(
        P2_U3255) );
  INV_X1 U12989 ( .A(n14985), .ZN(n10389) );
  INV_X1 U12990 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U12991 ( .A1(n10389), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n10376), 
        .B2(n14985), .ZN(n14970) );
  INV_X1 U12992 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10377) );
  AOI21_X1 U12993 ( .B1(n10378), .B2(n10377), .A(n10699), .ZN(n10396) );
  INV_X1 U12994 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15205) );
  AOI22_X1 U12995 ( .A1(n10389), .A2(n15205), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n14985), .ZN(n14973) );
  OR2_X1 U12996 ( .A1(n10380), .A2(n10379), .ZN(n10382) );
  NAND2_X1 U12997 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10383), .ZN(n10690) );
  OAI21_X1 U12998 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10383), .A(n10690), .ZN(
        n10394) );
  NAND2_X1 U12999 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10587) );
  NAND2_X1 U13000 ( .A1(n15095), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n10384) );
  OAI211_X1 U13001 ( .C1(n15092), .C2(n10689), .A(n10587), .B(n10384), .ZN(
        n10393) );
  MUX2_X1 U13002 ( .A(n10376), .B(n15205), .S(n12758), .Z(n10390) );
  XNOR2_X1 U13003 ( .A(n10390), .B(n14985), .ZN(n14981) );
  OR2_X1 U13004 ( .A1(n10386), .A2(n10385), .ZN(n10388) );
  MUX2_X1 U13005 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12758), .Z(n10679) );
  XNOR2_X1 U13006 ( .A(n10679), .B(n10689), .ZN(n10681) );
  XOR2_X1 U13007 ( .A(n10680), .B(n10681), .Z(n10391) );
  NOR2_X1 U13008 ( .A1(n10391), .A2(n15077), .ZN(n10392) );
  AOI211_X1 U13009 ( .C1(n15087), .C2(n10394), .A(n10393), .B(n10392), .ZN(
        n10395) );
  OAI21_X1 U13010 ( .B1(n10396), .B2(n15102), .A(n10395), .ZN(P3_U3189) );
  INV_X1 U13011 ( .A(n12868), .ZN(n15119) );
  NAND2_X1 U13012 ( .A1(n15144), .A2(n15119), .ZN(n10397) );
  NAND2_X1 U13013 ( .A1(n10398), .A2(n12557), .ZN(n10476) );
  NAND2_X1 U13014 ( .A1(n10476), .A2(n12559), .ZN(n10399) );
  NAND2_X1 U13015 ( .A1(n10399), .A2(n12500), .ZN(n10401) );
  NAND3_X1 U13016 ( .A1(n10476), .A2(n12559), .A3(n7009), .ZN(n10400) );
  AND2_X1 U13017 ( .A1(n10401), .A2(n10400), .ZN(n15173) );
  AND2_X1 U13018 ( .A1(n10480), .A2(n10402), .ZN(n10403) );
  NAND2_X1 U13019 ( .A1(n10481), .A2(n10403), .ZN(n10404) );
  AOI21_X1 U13020 ( .B1(n10404), .B2(n12500), .A(n15132), .ZN(n10408) );
  OAI22_X1 U13021 ( .A1(n10405), .A2(n15134), .B1(n12575), .B2(n15136), .ZN(
        n10406) );
  AOI21_X1 U13022 ( .B1(n10408), .B2(n10407), .A(n10406), .ZN(n15170) );
  MUX2_X1 U13023 ( .A(n15170), .B(n10376), .S(n15146), .Z(n10412) );
  AOI22_X1 U13024 ( .A1(n14528), .A2(n10410), .B1(n15140), .B2(n10409), .ZN(
        n10411) );
  OAI211_X1 U13025 ( .C1(n13002), .C2(n15173), .A(n10412), .B(n10411), .ZN(
        P3_U3227) );
  OAI211_X1 U13026 ( .C1(n10414), .C2(n12225), .A(n10413), .B(n14144), .ZN(
        n10416) );
  AOI22_X1 U13027 ( .A1(n14082), .A2(n13831), .B1(n13829), .B2(n14079), .ZN(
        n10415) );
  NAND2_X1 U13028 ( .A1(n10416), .A2(n10415), .ZN(n14610) );
  INV_X1 U13029 ( .A(n14610), .ZN(n10427) );
  OAI21_X1 U13030 ( .B1(n10419), .B2(n10418), .A(n10417), .ZN(n14612) );
  NAND2_X1 U13031 ( .A1(n14607), .A2(n10420), .ZN(n10421) );
  NAND2_X1 U13032 ( .A1(n10421), .A2(n14176), .ZN(n10422) );
  OR2_X1 U13033 ( .A1(n10576), .A2(n10422), .ZN(n14608) );
  OAI22_X1 U13034 ( .A1(n14668), .A2(n9399), .B1(n14605), .B2(n14665), .ZN(
        n10423) );
  AOI21_X1 U13035 ( .B1(n14607), .B2(n14670), .A(n10423), .ZN(n10424) );
  OAI21_X1 U13036 ( .B1(n14608), .B2(n14673), .A(n10424), .ZN(n10425) );
  AOI21_X1 U13037 ( .B1(n14612), .B2(n14188), .A(n10425), .ZN(n10426) );
  OAI21_X1 U13038 ( .B1(n14678), .B2(n10427), .A(n10426), .ZN(P1_U3282) );
  AOI22_X1 U13039 ( .A1(n12067), .A2(n12326), .B1(n12323), .B2(n13833), .ZN(
        n10428) );
  XNOR2_X1 U13040 ( .A(n10428), .B(n12324), .ZN(n10618) );
  AOI22_X1 U13041 ( .A1(n12067), .A2(n12323), .B1(n12322), .B2(n13833), .ZN(
        n10617) );
  XNOR2_X1 U13042 ( .A(n10618), .B(n10617), .ZN(n10436) );
  INV_X1 U13043 ( .A(n10429), .ZN(n10432) );
  AOI21_X1 U13044 ( .B1(n10436), .B2(n10435), .A(n10619), .ZN(n10442) );
  AOI22_X1 U13045 ( .A1(n14587), .A2(n10437), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10438) );
  OAI21_X1 U13046 ( .B1(n14606), .B2(n10439), .A(n10438), .ZN(n10440) );
  AOI21_X1 U13047 ( .B1(n12067), .B2(n14602), .A(n10440), .ZN(n10441) );
  OAI21_X1 U13048 ( .B1(n10442), .B2(n14598), .A(n10441), .ZN(P1_U3221) );
  XNOR2_X1 U13049 ( .A(n10443), .B(n11727), .ZN(n10452) );
  INV_X1 U13050 ( .A(n10452), .ZN(n14884) );
  OAI211_X1 U13051 ( .C1(n14881), .C2(n10445), .A(n10444), .B(n10936), .ZN(
        n14880) );
  AOI22_X1 U13052 ( .A1(n14557), .A2(n11392), .B1(n14555), .B2(n10446), .ZN(
        n10447) );
  OAI21_X1 U13053 ( .B1(n14880), .B2(n13550), .A(n10447), .ZN(n10454) );
  XNOR2_X1 U13054 ( .A(n10448), .B(n11727), .ZN(n10450) );
  OAI22_X1 U13055 ( .A1(n11384), .A2(n13538), .B1(n11399), .B2(n13540), .ZN(
        n10449) );
  AOI21_X1 U13056 ( .B1(n10450), .B2(n13521), .A(n10449), .ZN(n10451) );
  OAI21_X1 U13057 ( .B1(n10452), .B2(n13647), .A(n10451), .ZN(n14882) );
  MUX2_X1 U13058 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n14882), .S(n13441), .Z(
        n10453) );
  AOI211_X1 U13059 ( .C1(n14884), .C2(n10497), .A(n10454), .B(n10453), .ZN(
        n10455) );
  INV_X1 U13060 ( .A(n10455), .ZN(P2_U3259) );
  OAI21_X1 U13061 ( .B1(n10457), .B2(n11725), .A(n10456), .ZN(n14869) );
  AOI21_X1 U13062 ( .B1(n10458), .B2(n11370), .A(n13459), .ZN(n10460) );
  NAND2_X1 U13063 ( .A1(n10460), .A2(n10459), .ZN(n14865) );
  AOI22_X1 U13064 ( .A1(n14557), .A2(n11370), .B1(n10461), .B2(n14555), .ZN(
        n10462) );
  OAI21_X1 U13065 ( .B1(n13550), .B2(n14865), .A(n10462), .ZN(n10471) );
  NAND3_X1 U13066 ( .A1(n10464), .A2(n11725), .A3(n10463), .ZN(n10465) );
  NAND2_X1 U13067 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  NAND2_X1 U13068 ( .A1(n10467), .A2(n13521), .ZN(n10469) );
  AOI22_X1 U13069 ( .A1(n13650), .A2(n13298), .B1(n13300), .B2(n13470), .ZN(
        n10468) );
  NAND2_X1 U13070 ( .A1(n10469), .A2(n10468), .ZN(n14867) );
  MUX2_X1 U13071 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n14867), .S(n13441), .Z(
        n10470) );
  AOI211_X1 U13072 ( .C1(n14563), .C2(n14869), .A(n10471), .B(n10470), .ZN(
        n10472) );
  INV_X1 U13073 ( .A(n10472), .ZN(P2_U3261) );
  NAND2_X1 U13074 ( .A1(n10473), .A2(n13135), .ZN(n10474) );
  OAI211_X1 U13075 ( .C1(n10475), .C2(n12350), .A(n10474), .B(n12697), .ZN(
        P3_U3272) );
  OAI21_X1 U13076 ( .B1(n10398), .B2(n12557), .A(n10476), .ZN(n15166) );
  INV_X1 U13077 ( .A(n15166), .ZN(n10490) );
  NAND2_X1 U13078 ( .A1(n10503), .A2(n10477), .ZN(n10479) );
  NAND2_X1 U13079 ( .A1(n10479), .A2(n10478), .ZN(n10484) );
  AND2_X1 U13080 ( .A1(n10481), .A2(n10480), .ZN(n10482) );
  OAI21_X1 U13081 ( .B1(n10484), .B2(n10483), .A(n10482), .ZN(n10485) );
  AOI222_X1 U13082 ( .A1(n12987), .A2(n10485), .B1(n12714), .B2(n12990), .C1(
        n12716), .C2(n12993), .ZN(n15168) );
  MUX2_X1 U13083 ( .A(n10486), .B(n15168), .S(n15144), .Z(n10489) );
  AOI22_X1 U13084 ( .A1(n14528), .A2(n15165), .B1(n15140), .B2(n10487), .ZN(
        n10488) );
  OAI211_X1 U13085 ( .C1(n13002), .C2(n10490), .A(n10489), .B(n10488), .ZN(
        P3_U3228) );
  AOI22_X1 U13086 ( .A1(n14557), .A2(n13164), .B1(n14555), .B2(n13165), .ZN(
        n10491) );
  OAI21_X1 U13087 ( .B1(n13550), .B2(n10492), .A(n10491), .ZN(n10495) );
  MUX2_X1 U13088 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10493), .S(n13441), .Z(
        n10494) );
  AOI211_X1 U13089 ( .C1(n10497), .C2(n10496), .A(n10495), .B(n10494), .ZN(
        n10498) );
  INV_X1 U13090 ( .A(n10498), .ZN(P2_U3262) );
  OAI21_X1 U13091 ( .B1(n10500), .B2(n12507), .A(n10499), .ZN(n15157) );
  INV_X1 U13092 ( .A(n15157), .ZN(n10510) );
  OAI22_X1 U13093 ( .A1(n15135), .A2(n15134), .B1(n10501), .B2(n15136), .ZN(
        n10507) );
  NAND2_X1 U13094 ( .A1(n15116), .A2(n10502), .ZN(n10505) );
  INV_X1 U13095 ( .A(n10503), .ZN(n10504) );
  AOI211_X1 U13096 ( .C1(n12507), .C2(n10505), .A(n15132), .B(n10504), .ZN(
        n10506) );
  AOI211_X1 U13097 ( .C1(n15119), .C2(n15157), .A(n10507), .B(n10506), .ZN(
        n15159) );
  MUX2_X1 U13098 ( .A(n9545), .B(n15159), .S(n15144), .Z(n10509) );
  AOI22_X1 U13099 ( .A1(n14528), .A2(n15155), .B1(n15140), .B2(n7740), .ZN(
        n10508) );
  OAI211_X1 U13100 ( .C1(n10510), .C2(n12848), .A(n10509), .B(n10508), .ZN(
        P3_U3230) );
  OR2_X1 U13101 ( .A1(n11424), .A2(n13293), .ZN(n10511) );
  NAND2_X1 U13102 ( .A1(n10512), .A2(n10511), .ZN(n10514) );
  NAND2_X1 U13103 ( .A1(n11424), .A2(n13293), .ZN(n10513) );
  NAND2_X1 U13104 ( .A1(n10514), .A2(n10513), .ZN(n10778) );
  NAND2_X1 U13105 ( .A1(n10515), .A2(n6652), .ZN(n10518) );
  AOI22_X1 U13106 ( .A1(n11683), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11490), 
        .B2(n10516), .ZN(n10517) );
  XNOR2_X1 U13107 ( .A(n14918), .B(n13292), .ZN(n11734) );
  XNOR2_X1 U13108 ( .A(n10778), .B(n11734), .ZN(n14916) );
  INV_X1 U13109 ( .A(n14916), .ZN(n10542) );
  NAND2_X1 U13110 ( .A1(n14916), .A2(n14873), .ZN(n10533) );
  NAND2_X1 U13111 ( .A1(n11424), .A2(n11421), .ZN(n10519) );
  XNOR2_X1 U13112 ( .A(n10747), .B(n11734), .ZN(n10531) );
  NAND2_X1 U13113 ( .A1(n11686), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10527) );
  AND2_X1 U13114 ( .A1(n10522), .A2(n10521), .ZN(n10523) );
  NOR2_X1 U13115 ( .A1(n10760), .A2(n10523), .ZN(n14554) );
  NAND2_X1 U13116 ( .A1(n11658), .A2(n14554), .ZN(n10526) );
  NAND2_X1 U13117 ( .A1(n11642), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10525) );
  OR2_X1 U13118 ( .A1(n11605), .A2(n9832), .ZN(n10524) );
  NAND4_X1 U13119 ( .A1(n10527), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(
        n13291) );
  NAND2_X1 U13120 ( .A1(n13650), .A2(n13291), .ZN(n10529) );
  NAND2_X1 U13121 ( .A1(n13293), .A2(n13470), .ZN(n10528) );
  AND2_X1 U13122 ( .A1(n10529), .A2(n10528), .ZN(n10659) );
  INV_X1 U13123 ( .A(n10659), .ZN(n10530) );
  AOI21_X1 U13124 ( .B1(n10531), .B2(n13521), .A(n10530), .ZN(n10532) );
  NAND2_X1 U13125 ( .A1(n10533), .A2(n10532), .ZN(n14922) );
  NAND2_X1 U13126 ( .A1(n14922), .A2(n13441), .ZN(n10541) );
  NAND2_X1 U13127 ( .A1(n10534), .A2(n14918), .ZN(n10535) );
  NAND2_X1 U13128 ( .A1(n10535), .A2(n10936), .ZN(n10536) );
  NOR2_X1 U13129 ( .A1(n6810), .A2(n10536), .ZN(n14920) );
  INV_X1 U13130 ( .A(n14918), .ZN(n10538) );
  AOI22_X1 U13131 ( .A1(n14556), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10656), 
        .B2(n14555), .ZN(n10537) );
  OAI21_X1 U13132 ( .B1(n10538), .B2(n13528), .A(n10537), .ZN(n10539) );
  AOI21_X1 U13133 ( .B1(n14920), .B2(n15590), .A(n10539), .ZN(n10540) );
  OAI211_X1 U13134 ( .C1(n10542), .C2(n15596), .A(n10541), .B(n10540), .ZN(
        P2_U3254) );
  NAND2_X1 U13135 ( .A1(n11063), .A2(n10543), .ZN(n10545) );
  NAND2_X1 U13136 ( .A1(n10545), .A2(n10544), .ZN(n10549) );
  INV_X1 U13137 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10547) );
  NAND2_X1 U13138 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n11170), .ZN(n13321) );
  INV_X1 U13139 ( .A(n13321), .ZN(n10546) );
  AOI21_X1 U13140 ( .B1(n10547), .B2(n13327), .A(n10546), .ZN(n10548) );
  NAND2_X1 U13141 ( .A1(n10548), .A2(n10549), .ZN(n13320) );
  OAI211_X1 U13142 ( .C1(n10549), .C2(n10548), .A(n14837), .B(n13320), .ZN(
        n10558) );
  NAND2_X1 U13143 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n11202)
         );
  NAND2_X1 U13144 ( .A1(n11063), .A2(n10550), .ZN(n10552) );
  NAND2_X1 U13145 ( .A1(n10552), .A2(n10551), .ZN(n10554) );
  XNOR2_X1 U13146 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13327), .ZN(n10553) );
  NAND2_X1 U13147 ( .A1(n10553), .A2(n10554), .ZN(n13325) );
  OAI211_X1 U13148 ( .C1(n10554), .C2(n10553), .A(n14843), .B(n13325), .ZN(
        n10555) );
  NAND2_X1 U13149 ( .A1(n11202), .A2(n10555), .ZN(n10556) );
  AOI21_X1 U13150 ( .B1(n14835), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n10556), 
        .ZN(n10557) );
  OAI211_X1 U13151 ( .C1(n14765), .C2(n13327), .A(n10558), .B(n10557), .ZN(
        P2_U3230) );
  XNOR2_X1 U13152 ( .A(n11424), .B(n12012), .ZN(n10650) );
  NAND2_X1 U13153 ( .A1(n13293), .A2(n13459), .ZN(n10652) );
  XNOR2_X1 U13154 ( .A(n10650), .B(n10652), .ZN(n10562) );
  OAI211_X1 U13155 ( .C1(n10563), .C2(n10562), .A(n10651), .B(n13249), .ZN(
        n10567) );
  AND2_X1 U13156 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14815) );
  OAI22_X1 U13157 ( .A1(n13258), .A2(n11433), .B1(n10564), .B2(n13270), .ZN(
        n10565) );
  AOI211_X1 U13158 ( .C1(n13244), .C2(n13294), .A(n14815), .B(n10565), .ZN(
        n10566) );
  OAI211_X1 U13159 ( .C1(n14910), .C2(n13242), .A(n10567), .B(n10566), .ZN(
        P2_U3189) );
  OAI211_X1 U13160 ( .C1(n10569), .C2(n12226), .A(n10568), .B(n14144), .ZN(
        n10572) );
  NAND2_X1 U13161 ( .A1(n13830), .A2(n14082), .ZN(n10571) );
  NAND2_X1 U13162 ( .A1(n13828), .A2(n14079), .ZN(n10570) );
  AND2_X1 U13163 ( .A1(n10571), .A2(n10570), .ZN(n11130) );
  NAND2_X1 U13164 ( .A1(n10572), .A2(n11130), .ZN(n10813) );
  INV_X1 U13165 ( .A(n10813), .ZN(n10583) );
  OAI21_X1 U13166 ( .B1(n10575), .B2(n10574), .A(n10573), .ZN(n10815) );
  OR2_X1 U13167 ( .A1(n11135), .A2(n10576), .ZN(n10577) );
  AND3_X1 U13168 ( .A1(n10641), .A2(n10577), .A3(n14176), .ZN(n10814) );
  NAND2_X1 U13169 ( .A1(n10814), .A2(n14165), .ZN(n10580) );
  INV_X1 U13170 ( .A(n10578), .ZN(n11132) );
  AOI22_X1 U13171 ( .A1(n14678), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11132), 
        .B2(n14180), .ZN(n10579) );
  OAI211_X1 U13172 ( .C1(n11135), .C2(n14156), .A(n10580), .B(n10579), .ZN(
        n10581) );
  AOI21_X1 U13173 ( .B1(n10815), .B2(n14188), .A(n10581), .ZN(n10582) );
  OAI21_X1 U13174 ( .B1(n14678), .B2(n10583), .A(n10582), .ZN(P1_U3281) );
  OAI222_X1 U13175 ( .A1(P1_U3086), .A2(n12206), .B1(n14330), .B2(n11523), 
        .C1(n10584), .C2(n14332), .ZN(P1_U3334) );
  OAI222_X1 U13176 ( .A1(n13693), .A2(n10585), .B1(P2_U3088), .B2(n11750), 
        .C1(n11317), .C2(n11523), .ZN(P2_U3306) );
  NOR2_X1 U13177 ( .A1(n10723), .A2(n10592), .ZN(n10598) );
  NOR2_X1 U13178 ( .A1(n10586), .A2(n10598), .ZN(n10799) );
  XNOR2_X1 U13179 ( .A(n12568), .B(n11886), .ZN(n10798) );
  INV_X1 U13180 ( .A(n10798), .ZN(n10597) );
  XNOR2_X1 U13181 ( .A(n10799), .B(n10597), .ZN(n10591) );
  AOI22_X1 U13182 ( .A1(n12714), .A2(n11899), .B1(n12440), .B2(n12712), .ZN(
        n10588) );
  OAI211_X1 U13183 ( .C1(n12446), .C2(n15177), .A(n10588), .B(n10587), .ZN(
        n10589) );
  AOI21_X1 U13184 ( .B1(n10729), .B2(n12451), .A(n10589), .ZN(n10590) );
  OAI21_X1 U13185 ( .B1(n10591), .B2(n12459), .A(n10590), .ZN(P3_U3153) );
  XNOR2_X1 U13186 ( .A(n15194), .B(n11886), .ZN(n10732) );
  XNOR2_X1 U13187 ( .A(n10732), .B(n12711), .ZN(n10609) );
  XNOR2_X1 U13188 ( .A(n15183), .B(n11886), .ZN(n10601) );
  XNOR2_X1 U13189 ( .A(n10601), .B(n12712), .ZN(n10599) );
  NAND2_X1 U13190 ( .A1(n10723), .A2(n10592), .ZN(n10593) );
  AND4_X1 U13191 ( .A1(n10798), .A2(n10599), .A3(n10594), .A4(n10593), .ZN(
        n10595) );
  INV_X1 U13192 ( .A(n10599), .ZN(n10800) );
  OAI21_X1 U13193 ( .B1(n12575), .B2(n10800), .A(n10597), .ZN(n10604) );
  NAND2_X1 U13194 ( .A1(n10599), .A2(n10598), .ZN(n10600) );
  NAND2_X1 U13195 ( .A1(n10798), .A2(n10600), .ZN(n10603) );
  INV_X1 U13196 ( .A(n10601), .ZN(n10602) );
  AOI22_X1 U13197 ( .A1(n10604), .A2(n10603), .B1(n10602), .B2(n12712), .ZN(
        n10605) );
  INV_X1 U13198 ( .A(n10609), .ZN(n10606) );
  INV_X1 U13199 ( .A(n10737), .ZN(n10607) );
  AOI21_X1 U13200 ( .B1(n10609), .B2(n10608), .A(n10607), .ZN(n10615) );
  INV_X1 U13201 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10610) );
  NOR2_X1 U13202 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10610), .ZN(n15020) );
  OAI22_X1 U13203 ( .A1(n10611), .A2(n12442), .B1(n11028), .B2(n12368), .ZN(
        n10612) );
  AOI211_X1 U13204 ( .C1(n12456), .C2(n15194), .A(n15020), .B(n10612), .ZN(
        n10614) );
  NAND2_X1 U13205 ( .A1(n12451), .A2(n10874), .ZN(n10613) );
  OAI211_X1 U13206 ( .C1(n10615), .C2(n12459), .A(n10614), .B(n10613), .ZN(
        P3_U3171) );
  INV_X1 U13207 ( .A(n10616), .ZN(n13804) );
  NAND2_X1 U13208 ( .A1(n14671), .A2(n14743), .ZN(n14736) );
  NAND2_X1 U13209 ( .A1(n14671), .A2(n12326), .ZN(n10621) );
  NAND2_X1 U13210 ( .A1(n13832), .A2(n12323), .ZN(n10620) );
  NAND2_X1 U13211 ( .A1(n10621), .A2(n10620), .ZN(n10622) );
  XNOR2_X1 U13212 ( .A(n10622), .B(n12324), .ZN(n10834) );
  AND2_X1 U13213 ( .A1(n13832), .A2(n12322), .ZN(n10623) );
  AOI21_X1 U13214 ( .B1(n14671), .B2(n12323), .A(n10623), .ZN(n10835) );
  XNOR2_X1 U13215 ( .A(n10834), .B(n10835), .ZN(n10624) );
  OAI211_X1 U13216 ( .C1(n10625), .C2(n10624), .A(n10838), .B(n14585), .ZN(
        n10631) );
  INV_X1 U13217 ( .A(n14666), .ZN(n10629) );
  NAND2_X1 U13218 ( .A1(n13833), .A2(n14082), .ZN(n10627) );
  NAND2_X1 U13219 ( .A1(n13831), .A2(n14079), .ZN(n10626) );
  AND2_X1 U13220 ( .A1(n10627), .A2(n10626), .ZN(n14737) );
  OAI22_X1 U13221 ( .A1(n13808), .A2(n14737), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13925), .ZN(n10628) );
  AOI21_X1 U13222 ( .B1(n13806), .B2(n10629), .A(n10628), .ZN(n10630) );
  OAI211_X1 U13223 ( .C1(n13804), .C2(n14736), .A(n10631), .B(n10630), .ZN(
        P1_U3231) );
  INV_X1 U13224 ( .A(n10632), .ZN(n10633) );
  AOI21_X1 U13225 ( .B1(n10633), .B2(n10639), .A(n14656), .ZN(n10637) );
  NAND2_X1 U13226 ( .A1(n13829), .A2(n14082), .ZN(n10635) );
  NAND2_X1 U13227 ( .A1(n13827), .A2(n14079), .ZN(n10634) );
  NAND2_X1 U13228 ( .A1(n10635), .A2(n10634), .ZN(n11254) );
  AOI21_X1 U13229 ( .B1(n10637), .B2(n10636), .A(n11254), .ZN(n10911) );
  OAI21_X1 U13230 ( .B1(n10640), .B2(n10639), .A(n10638), .ZN(n10913) );
  AOI21_X1 U13231 ( .B1(n10641), .B2(n12092), .A(n14661), .ZN(n10642) );
  NAND2_X1 U13232 ( .A1(n10642), .A2(n10826), .ZN(n10910) );
  NAND2_X1 U13233 ( .A1(n14678), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10643) );
  OAI21_X1 U13234 ( .B1(n14665), .B2(n11251), .A(n10643), .ZN(n10644) );
  AOI21_X1 U13235 ( .B1(n12092), .B2(n14670), .A(n10644), .ZN(n10645) );
  OAI21_X1 U13236 ( .B1(n10910), .B2(n14673), .A(n10645), .ZN(n10646) );
  AOI21_X1 U13237 ( .B1(n10913), .B2(n14188), .A(n10646), .ZN(n10647) );
  OAI21_X1 U13238 ( .B1(n10911), .B2(n14678), .A(n10647), .ZN(P1_U3280) );
  OAI222_X1 U13239 ( .A1(P1_U3086), .A2(n10649), .B1(n14330), .B2(n12262), 
        .C1(n10648), .C2(n14332), .ZN(P1_U3335) );
  XNOR2_X1 U13240 ( .A(n14918), .B(n11995), .ZN(n10654) );
  NAND2_X1 U13241 ( .A1(n13292), .A2(n10208), .ZN(n10653) );
  NOR2_X1 U13242 ( .A1(n10654), .A2(n10653), .ZN(n10854) );
  NOR2_X1 U13243 ( .A1(n10854), .A2(n6811), .ZN(n10655) );
  XNOR2_X1 U13244 ( .A(n10855), .B(n10655), .ZN(n10662) );
  NAND2_X1 U13245 ( .A1(n13219), .A2(n10656), .ZN(n10657) );
  OAI211_X1 U13246 ( .C1(n13217), .C2(n10659), .A(n10658), .B(n10657), .ZN(
        n10660) );
  AOI21_X1 U13247 ( .B1(n14918), .B2(n13273), .A(n10660), .ZN(n10661) );
  OAI21_X1 U13248 ( .B1(n10662), .B2(n13275), .A(n10661), .ZN(P2_U3208) );
  OAI21_X1 U13249 ( .B1(n10664), .B2(n10669), .A(n10663), .ZN(n10665) );
  NOR2_X1 U13250 ( .A1(n10670), .A2(n10665), .ZN(n10666) );
  XNOR2_X1 U13251 ( .A(n10670), .B(n10665), .ZN(n14639) );
  NOR2_X1 U13252 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14639), .ZN(n14638) );
  NOR2_X1 U13253 ( .A1(n10666), .A2(n14638), .ZN(n10882) );
  XNOR2_X1 U13254 ( .A(n10887), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n10881) );
  XNOR2_X1 U13255 ( .A(n10882), .B(n10881), .ZN(n10678) );
  NAND2_X1 U13256 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13744)
         );
  AOI21_X1 U13257 ( .B1(n10669), .B2(n10668), .A(n10667), .ZN(n10671) );
  NOR2_X1 U13258 ( .A1(n10670), .A2(n10671), .ZN(n10672) );
  XOR2_X1 U13259 ( .A(n14646), .B(n10671), .Z(n14641) );
  NOR2_X1 U13260 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14641), .ZN(n14640) );
  NOR2_X1 U13261 ( .A1(n10672), .A2(n14640), .ZN(n10884) );
  XNOR2_X1 U13262 ( .A(n10880), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10886) );
  XNOR2_X1 U13263 ( .A(n10884), .B(n10886), .ZN(n10673) );
  NAND2_X1 U13264 ( .A1(n13966), .A2(n10673), .ZN(n10674) );
  NAND2_X1 U13265 ( .A1(n13744), .A2(n10674), .ZN(n10676) );
  NOR2_X1 U13266 ( .A1(n14647), .A2(n10887), .ZN(n10675) );
  AOI211_X1 U13267 ( .C1(n13929), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n10676), 
        .B(n10675), .ZN(n10677) );
  OAI21_X1 U13268 ( .B1(n10678), .B2(n14645), .A(n10677), .ZN(P1_U3259) );
  MUX2_X1 U13269 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12758), .Z(n10682) );
  OR2_X1 U13270 ( .A1(n10682), .A2(n10701), .ZN(n10683) );
  OAI22_X1 U13271 ( .A1(n10681), .A2(n10680), .B1(n10679), .B2(n10689), .ZN(
        n14998) );
  XNOR2_X1 U13272 ( .A(n10682), .B(n15000), .ZN(n14997) );
  NAND2_X1 U13273 ( .A1(n14998), .A2(n14997), .ZN(n14996) );
  NAND2_X1 U13274 ( .A1(n10683), .A2(n14996), .ZN(n15016) );
  INV_X1 U13275 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15012) );
  INV_X1 U13276 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15211) );
  MUX2_X1 U13277 ( .A(n15012), .B(n15211), .S(n12758), .Z(n10684) );
  OR2_X1 U13278 ( .A1(n10684), .A2(n10702), .ZN(n15013) );
  NAND2_X1 U13279 ( .A1(n10684), .A2(n10702), .ZN(n15014) );
  INV_X1 U13280 ( .A(n15014), .ZN(n10685) );
  AOI21_X1 U13281 ( .B1(n15016), .B2(n15013), .A(n10685), .ZN(n10687) );
  MUX2_X1 U13282 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12758), .Z(n12740) );
  XNOR2_X1 U13283 ( .A(n12740), .B(n12722), .ZN(n10686) );
  NOR2_X1 U13284 ( .A1(n10687), .A2(n10686), .ZN(n12741) );
  AOI21_X1 U13285 ( .B1(n10687), .B2(n10686), .A(n12741), .ZN(n10713) );
  INV_X1 U13286 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15208) );
  AOI22_X1 U13287 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10701), .B1(n15000), 
        .B2(n15208), .ZN(n14995) );
  NAND2_X1 U13288 ( .A1(n10689), .A2(n10688), .ZN(n10691) );
  NAND2_X1 U13289 ( .A1(n15017), .A2(n10692), .ZN(n10693) );
  NAND2_X1 U13290 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15022), .ZN(n15021) );
  NAND2_X1 U13291 ( .A1(n10693), .A2(n15021), .ZN(n10695) );
  MUX2_X1 U13292 ( .A(n15499), .B(P3_REG1_REG_10__SCAN_IN), .S(n12774), .Z(
        n10694) );
  NAND2_X1 U13293 ( .A1(n10695), .A2(n10694), .ZN(n12773) );
  OAI21_X1 U13294 ( .B1(n10695), .B2(n10694), .A(n12773), .ZN(n10696) );
  NAND2_X1 U13295 ( .A1(n10696), .A2(n15087), .ZN(n10712) );
  INV_X1 U13296 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13297 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n15000), .B1(n10701), 
        .B2(n10700), .ZN(n14991) );
  NOR2_X1 U13298 ( .A1(n14992), .A2(n14991), .ZN(n14990) );
  NOR2_X1 U13299 ( .A1(n10702), .A2(n10703), .ZN(n10704) );
  INV_X1 U13300 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10929) );
  MUX2_X1 U13301 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n10929), .S(n12774), .Z(
        n10705) );
  AOI21_X1 U13302 ( .B1(n6814), .B2(n10705), .A(n12721), .ZN(n10709) );
  NAND2_X1 U13303 ( .A1(n15095), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n10708) );
  INV_X1 U13304 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n10706) );
  NOR2_X1 U13305 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10706), .ZN(n10740) );
  INV_X1 U13306 ( .A(n10740), .ZN(n10707) );
  OAI211_X1 U13307 ( .C1(n15102), .C2(n10709), .A(n10708), .B(n10707), .ZN(
        n10710) );
  AOI21_X1 U13308 ( .B1(n12774), .B2(n14999), .A(n10710), .ZN(n10711) );
  OAI211_X1 U13309 ( .C1(n10713), .C2(n15077), .A(n10712), .B(n10711), .ZN(
        P3_U3192) );
  NAND2_X1 U13310 ( .A1(n10398), .A2(n10714), .ZN(n10716) );
  NAND2_X1 U13311 ( .A1(n10716), .A2(n10715), .ZN(n10717) );
  OR2_X1 U13312 ( .A1(n10717), .A2(n10720), .ZN(n10718) );
  NAND2_X1 U13313 ( .A1(n6819), .A2(n10718), .ZN(n10725) );
  INV_X1 U13314 ( .A(n10725), .ZN(n15178) );
  XNOR2_X1 U13315 ( .A(n10719), .B(n10720), .ZN(n10721) );
  NAND2_X1 U13316 ( .A1(n10721), .A2(n12987), .ZN(n10727) );
  NAND2_X1 U13317 ( .A1(n12712), .A2(n12990), .ZN(n10722) );
  OAI21_X1 U13318 ( .B1(n10723), .B2(n15134), .A(n10722), .ZN(n10724) );
  AOI21_X1 U13319 ( .B1(n10725), .B2(n15119), .A(n10724), .ZN(n10726) );
  NAND2_X1 U13320 ( .A1(n10727), .A2(n10726), .ZN(n15180) );
  MUX2_X1 U13321 ( .A(n15180), .B(P3_REG2_REG_7__SCAN_IN), .S(n15146), .Z(
        n10728) );
  INV_X1 U13322 ( .A(n10728), .ZN(n10731) );
  AOI22_X1 U13323 ( .A1(n14528), .A2(n12534), .B1(n15140), .B2(n10729), .ZN(
        n10730) );
  OAI211_X1 U13324 ( .C1(n15178), .C2(n12848), .A(n10731), .B(n10730), .ZN(
        P3_U3226) );
  INV_X1 U13325 ( .A(n10925), .ZN(n10746) );
  INV_X1 U13326 ( .A(n10732), .ZN(n10734) );
  NAND2_X1 U13327 ( .A1(n10734), .A2(n10733), .ZN(n10735) );
  AND2_X1 U13328 ( .A1(n10737), .A2(n10735), .ZN(n10739) );
  XNOR2_X1 U13329 ( .A(n10926), .B(n11886), .ZN(n11026) );
  XNOR2_X1 U13330 ( .A(n11026), .B(n11028), .ZN(n10738) );
  AND2_X1 U13331 ( .A1(n10738), .A2(n10735), .ZN(n10736) );
  NAND2_X1 U13332 ( .A1(n10737), .A2(n10736), .ZN(n11030) );
  OAI211_X1 U13333 ( .C1(n10739), .C2(n10738), .A(n12436), .B(n11030), .ZN(
        n10745) );
  INV_X1 U13334 ( .A(n12676), .ZN(n12657) );
  NAND2_X1 U13335 ( .A1(n12711), .A2(n12657), .ZN(n12581) );
  NOR2_X1 U13336 ( .A1(n12581), .A2(n10802), .ZN(n10920) );
  AOI21_X1 U13337 ( .B1(n12456), .B2(n10926), .A(n10740), .ZN(n10741) );
  OAI21_X1 U13338 ( .B1(n10742), .B2(n12368), .A(n10741), .ZN(n10743) );
  AOI21_X1 U13339 ( .B1(n10920), .B2(n12416), .A(n10743), .ZN(n10744) );
  OAI211_X1 U13340 ( .C1(n10746), .C2(n12418), .A(n10745), .B(n10744), .ZN(
        P3_U3157) );
  NAND2_X1 U13341 ( .A1(n14918), .A2(n11433), .ZN(n10748) );
  NAND2_X1 U13342 ( .A1(n10749), .A2(n6652), .ZN(n10751) );
  AOI22_X1 U13343 ( .A1(n11683), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11490), 
        .B2(n13309), .ZN(n10750) );
  INV_X1 U13344 ( .A(n13291), .ZN(n11435) );
  OR2_X1 U13345 ( .A1(n14558), .A2(n11435), .ZN(n10754) );
  NAND2_X1 U13346 ( .A1(n14558), .A2(n11435), .ZN(n10752) );
  NAND2_X1 U13347 ( .A1(n10754), .A2(n10752), .ZN(n14559) );
  INV_X1 U13348 ( .A(n14559), .ZN(n10753) );
  NAND2_X1 U13349 ( .A1(n10755), .A2(n6652), .ZN(n10758) );
  INV_X1 U13350 ( .A(n10756), .ZN(n14830) );
  AOI22_X1 U13351 ( .A1(n11683), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n14830), 
        .B2(n11490), .ZN(n10757) );
  NAND2_X1 U13352 ( .A1(n11642), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10765) );
  INV_X1 U13353 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10759) );
  OR2_X1 U13354 ( .A1(n9466), .A2(n10759), .ZN(n10764) );
  NAND2_X1 U13355 ( .A1(n10760), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10767) );
  OR2_X1 U13356 ( .A1(n10760), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10761) );
  AND2_X1 U13357 ( .A1(n10767), .A2(n10761), .ZN(n10782) );
  NAND2_X1 U13358 ( .A1(n11658), .A2(n10782), .ZN(n10763) );
  OR2_X1 U13359 ( .A1(n11605), .A2(n9833), .ZN(n10762) );
  NAND4_X1 U13360 ( .A1(n10765), .A2(n10764), .A3(n10763), .A4(n10762), .ZN(
        n13290) );
  XNOR2_X1 U13361 ( .A(n11443), .B(n13290), .ZN(n11735) );
  XNOR2_X1 U13362 ( .A(n11013), .B(n11735), .ZN(n10775) );
  INV_X1 U13363 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U13364 ( .A1(n10767), .A2(n10766), .ZN(n10768) );
  AND2_X1 U13365 ( .A1(n10955), .A2(n10768), .ZN(n11020) );
  NAND2_X1 U13366 ( .A1(n11020), .A2(n11658), .ZN(n10773) );
  NAND2_X1 U13367 ( .A1(n11642), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10772) );
  INV_X1 U13368 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n15535) );
  OR2_X1 U13369 ( .A1(n9466), .A2(n15535), .ZN(n10771) );
  INV_X1 U13370 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10769) );
  OR2_X1 U13371 ( .A1(n11605), .A2(n10769), .ZN(n10770) );
  OAI22_X1 U13372 ( .A1(n11435), .A2(n13538), .B1(n11452), .B2(n13540), .ZN(
        n10902) );
  INV_X1 U13373 ( .A(n10902), .ZN(n10774) );
  OAI21_X1 U13374 ( .B1(n10775), .B2(n14548), .A(n10774), .ZN(n14567) );
  INV_X1 U13375 ( .A(n14567), .ZN(n10787) );
  AND2_X1 U13376 ( .A1(n14918), .A2(n13292), .ZN(n10777) );
  OR2_X1 U13377 ( .A1(n14918), .A2(n13292), .ZN(n10776) );
  NOR2_X1 U13378 ( .A1(n14558), .A2(n13291), .ZN(n10779) );
  NAND2_X1 U13379 ( .A1(n14558), .A2(n13291), .ZN(n10780) );
  XNOR2_X1 U13380 ( .A(n11010), .B(n11735), .ZN(n14569) );
  INV_X1 U13381 ( .A(n14561), .ZN(n10781) );
  OAI211_X1 U13382 ( .C1(n10781), .C2(n7075), .A(n10936), .B(n11019), .ZN(
        n14566) );
  INV_X1 U13383 ( .A(n10782), .ZN(n10904) );
  OAI22_X1 U13384 ( .A1(n13441), .A2(n9833), .B1(n10904), .B2(n15592), .ZN(
        n10783) );
  AOI21_X1 U13385 ( .B1(n11443), .B2(n14557), .A(n10783), .ZN(n10784) );
  OAI21_X1 U13386 ( .B1(n14566), .B2(n13550), .A(n10784), .ZN(n10785) );
  AOI21_X1 U13387 ( .B1(n14569), .B2(n14563), .A(n10785), .ZN(n10786) );
  OAI21_X1 U13388 ( .B1(n10787), .B2(n14556), .A(n10786), .ZN(P2_U3252) );
  INV_X1 U13389 ( .A(n10802), .ZN(n10791) );
  NAND2_X1 U13390 ( .A1(n10981), .A2(n10788), .ZN(n10869) );
  OAI21_X1 U13391 ( .B1(n10788), .B2(n10981), .A(n10869), .ZN(n10789) );
  INV_X1 U13392 ( .A(n10789), .ZN(n10790) );
  OAI222_X1 U13393 ( .A1(n15134), .A2(n12575), .B1(n12581), .B2(n10791), .C1(
        n10790), .C2(n15132), .ZN(n15184) );
  INV_X1 U13394 ( .A(n15184), .ZN(n10797) );
  OAI21_X1 U13395 ( .B1(n10793), .B2(n12572), .A(n10792), .ZN(n15186) );
  AOI22_X1 U13396 ( .A1(n14528), .A2(n10803), .B1(n15140), .B2(n10807), .ZN(
        n10794) );
  OAI21_X1 U13397 ( .B1(n10700), .B2(n15144), .A(n10794), .ZN(n10795) );
  AOI21_X1 U13398 ( .B1(n15186), .B2(n15141), .A(n10795), .ZN(n10796) );
  OAI21_X1 U13399 ( .B1(n10797), .B2(n15146), .A(n10796), .ZN(P3_U3225) );
  MUX2_X1 U13400 ( .A(n12575), .B(n10799), .S(n10798), .Z(n10801) );
  XNOR2_X1 U13401 ( .A(n10801), .B(n10800), .ZN(n10809) );
  NAND2_X1 U13402 ( .A1(n12416), .A2(n10802), .ZN(n10805) );
  AOI22_X1 U13403 ( .A1(n12713), .A2(n11899), .B1(n12456), .B2(n10803), .ZN(
        n10804) );
  NAND2_X1 U13404 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15007) );
  OAI211_X1 U13405 ( .C1(n12581), .C2(n10805), .A(n10804), .B(n15007), .ZN(
        n10806) );
  AOI21_X1 U13406 ( .B1(n10807), .B2(n12451), .A(n10806), .ZN(n10808) );
  OAI21_X1 U13407 ( .B1(n10809), .B2(n12459), .A(n10808), .ZN(P3_U3161) );
  NAND2_X1 U13408 ( .A1(n8669), .A2(n10810), .ZN(n10811) );
  NAND2_X1 U13409 ( .A1(n10812), .A2(n10811), .ZN(n11541) );
  OAI222_X1 U13410 ( .A1(n13693), .A2(n15395), .B1(P2_U3088), .B2(n9569), .C1(
        n11317), .C2(n11541), .ZN(P2_U3305) );
  AOI211_X1 U13411 ( .C1(n14752), .C2(n10815), .A(n10814), .B(n10813), .ZN(
        n10818) );
  INV_X1 U13412 ( .A(n14318), .ZN(n14304) );
  AOI22_X1 U13413 ( .A1(n12082), .A2(n14304), .B1(P1_REG0_REG_12__SCAN_IN), 
        .B2(n14753), .ZN(n10816) );
  OAI21_X1 U13414 ( .B1(n10818), .B2(n14753), .A(n10816), .ZN(P1_U3495) );
  AOI22_X1 U13415 ( .A1(n12082), .A2(n14245), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n14761), .ZN(n10817) );
  OAI21_X1 U13416 ( .B1(n10818), .B2(n14761), .A(n10817), .ZN(P1_U3540) );
  OAI211_X1 U13417 ( .C1(n10820), .C2(n12209), .A(n10819), .B(n14144), .ZN(
        n10824) );
  NAND2_X1 U13418 ( .A1(n13828), .A2(n14082), .ZN(n10822) );
  NAND2_X1 U13419 ( .A1(n13826), .A2(n14079), .ZN(n10821) );
  NAND2_X1 U13420 ( .A1(n10822), .A2(n10821), .ZN(n14588) );
  INV_X1 U13421 ( .A(n14588), .ZN(n10823) );
  NAND2_X1 U13422 ( .A1(n10824), .A2(n10823), .ZN(n10970) );
  INV_X1 U13423 ( .A(n10970), .ZN(n10833) );
  AOI21_X1 U13424 ( .B1(n12209), .B2(n10825), .A(n6798), .ZN(n10971) );
  AOI21_X1 U13425 ( .B1(n14584), .B2(n10826), .A(n14661), .ZN(n10827) );
  NAND2_X1 U13426 ( .A1(n10827), .A2(n6785), .ZN(n10967) );
  AOI22_X1 U13427 ( .A1(n14678), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n10828), 
        .B2(n14180), .ZN(n10830) );
  NAND2_X1 U13428 ( .A1(n14584), .A2(n14670), .ZN(n10829) );
  OAI211_X1 U13429 ( .C1(n10967), .C2(n14673), .A(n10830), .B(n10829), .ZN(
        n10831) );
  AOI21_X1 U13430 ( .B1(n10971), .B2(n14188), .A(n10831), .ZN(n10832) );
  OAI21_X1 U13431 ( .B1(n14678), .B2(n10833), .A(n10832), .ZN(P1_U3279) );
  INV_X1 U13432 ( .A(n10835), .ZN(n10836) );
  NAND2_X1 U13433 ( .A1(n10834), .A2(n10836), .ZN(n10837) );
  AND2_X1 U13434 ( .A1(n13831), .A2(n12322), .ZN(n10839) );
  AOI21_X1 U13435 ( .B1(n14744), .B2(n12323), .A(n10839), .ZN(n11115) );
  AOI22_X1 U13436 ( .A1(n14744), .A2(n12326), .B1(n12323), .B2(n13831), .ZN(
        n10840) );
  XNOR2_X1 U13437 ( .A(n10840), .B(n12324), .ZN(n11114) );
  XOR2_X1 U13438 ( .A(n11115), .B(n11114), .Z(n10841) );
  OAI211_X1 U13439 ( .C1(n10842), .C2(n10841), .A(n11119), .B(n14585), .ZN(
        n10849) );
  INV_X1 U13440 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10843) );
  OAI22_X1 U13441 ( .A1(n14593), .A2(n10844), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10843), .ZN(n10847) );
  NOR2_X1 U13442 ( .A1(n14606), .A2(n10845), .ZN(n10846) );
  AOI211_X1 U13443 ( .C1(n13789), .C2(n13832), .A(n10847), .B(n10846), .ZN(
        n10848) );
  OAI211_X1 U13444 ( .C1(n7080), .C2(n13792), .A(n10849), .B(n10848), .ZN(
        P1_U3217) );
  INV_X1 U13445 ( .A(n11555), .ZN(n10853) );
  NAND2_X1 U13446 ( .A1(n14323), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n10850) );
  OAI211_X1 U13447 ( .C1(n10853), .C2(n14330), .A(n10850), .B(n12260), .ZN(
        P1_U3332) );
  NAND2_X1 U13448 ( .A1(n13676), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n10852) );
  OR2_X1 U13449 ( .A1(n10851), .A2(P2_U3088), .ZN(n11770) );
  OAI211_X1 U13450 ( .C1(n10853), .C2(n11317), .A(n10852), .B(n11770), .ZN(
        P2_U3304) );
  XNOR2_X1 U13451 ( .A(n14558), .B(n12012), .ZN(n10859) );
  INV_X1 U13452 ( .A(n10859), .ZN(n10857) );
  AND2_X1 U13453 ( .A1(n13291), .A2(n13459), .ZN(n10858) );
  INV_X1 U13454 ( .A(n10858), .ZN(n10856) );
  NAND2_X1 U13455 ( .A1(n10857), .A2(n10856), .ZN(n10946) );
  NAND2_X1 U13456 ( .A1(n10859), .A2(n10858), .ZN(n10939) );
  AND2_X1 U13457 ( .A1(n10946), .A2(n10939), .ZN(n10860) );
  NAND2_X1 U13458 ( .A1(n10942), .A2(n10860), .ZN(n10899) );
  OAI21_X1 U13459 ( .B1(n10942), .B2(n10860), .A(n10899), .ZN(n10861) );
  NAND2_X1 U13460 ( .A1(n10861), .A2(n13249), .ZN(n10866) );
  NAND2_X1 U13461 ( .A1(n13650), .A2(n13290), .ZN(n10863) );
  NAND2_X1 U13462 ( .A1(n13292), .A2(n13470), .ZN(n10862) );
  AND2_X1 U13463 ( .A1(n10863), .A2(n10862), .ZN(n14550) );
  NAND2_X1 U13464 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n13307)
         );
  OAI21_X1 U13465 ( .B1(n13217), .B2(n14550), .A(n13307), .ZN(n10864) );
  AOI21_X1 U13466 ( .B1(n14554), .B2(n13219), .A(n10864), .ZN(n10865) );
  OAI211_X1 U13467 ( .C1(n14573), .C2(n13242), .A(n10866), .B(n10865), .ZN(
        P2_U3196) );
  XNOR2_X1 U13468 ( .A(n10867), .B(n7117), .ZN(n15190) );
  NAND2_X1 U13469 ( .A1(n10869), .A2(n10868), .ZN(n10870) );
  INV_X1 U13470 ( .A(n10870), .ZN(n10871) );
  OR2_X1 U13471 ( .A1(n10870), .A2(n12579), .ZN(n10918) );
  OAI211_X1 U13472 ( .C1(n10871), .C2(n7117), .A(n12987), .B(n10918), .ZN(
        n10873) );
  AOI22_X1 U13473 ( .A1(n12710), .A2(n12990), .B1(n12993), .B2(n12712), .ZN(
        n10872) );
  OAI211_X1 U13474 ( .C1(n12868), .C2(n15190), .A(n10873), .B(n10872), .ZN(
        n15191) );
  NAND2_X1 U13475 ( .A1(n15191), .A2(n15144), .ZN(n10879) );
  INV_X1 U13476 ( .A(n15194), .ZN(n10876) );
  INV_X1 U13477 ( .A(n10874), .ZN(n10875) );
  OAI22_X1 U13478 ( .A1(n10876), .A2(n12998), .B1(n10875), .B2(n15108), .ZN(
        n10877) );
  AOI21_X1 U13479 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15146), .A(n10877), .ZN(
        n10878) );
  OAI211_X1 U13480 ( .C1(n15190), .C2(n12848), .A(n10879), .B(n10878), .ZN(
        P3_U3224) );
  XNOR2_X1 U13481 ( .A(n11051), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U13482 ( .A1(n10882), .A2(n10881), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n10880), .ZN(n11044) );
  XOR2_X1 U13483 ( .A(n11046), .B(n11044), .Z(n10894) );
  NAND2_X1 U13484 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13757)
         );
  XNOR2_X1 U13485 ( .A(n10883), .B(n14271), .ZN(n10889) );
  INV_X1 U13486 ( .A(n10884), .ZN(n10885) );
  OAI22_X1 U13487 ( .A1(n15418), .A2(n10887), .B1(n10886), .B2(n10885), .ZN(
        n10888) );
  NAND2_X1 U13488 ( .A1(n10889), .A2(n10888), .ZN(n11050) );
  OAI211_X1 U13489 ( .C1(n10889), .C2(n10888), .A(n13966), .B(n11050), .ZN(
        n10890) );
  NAND2_X1 U13490 ( .A1(n13757), .A2(n10890), .ZN(n10892) );
  NOR2_X1 U13491 ( .A1(n14647), .A2(n11051), .ZN(n10891) );
  AOI211_X1 U13492 ( .C1(n13929), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n10892), 
        .B(n10891), .ZN(n10893) );
  OAI21_X1 U13493 ( .B1(n10894), .B2(n14645), .A(n10893), .ZN(P1_U3260) );
  INV_X1 U13494 ( .A(n10895), .ZN(n10896) );
  OAI222_X1 U13495 ( .A1(P3_U3151), .A2(n10898), .B1(n12350), .B2(n10897), 
        .C1(n11060), .C2(n10896), .ZN(P3_U3271) );
  NAND2_X1 U13496 ( .A1(n10899), .A2(n10946), .ZN(n10901) );
  XNOR2_X1 U13497 ( .A(n11443), .B(n11995), .ZN(n10943) );
  NAND2_X1 U13498 ( .A1(n13290), .A2(n13459), .ZN(n10948) );
  XNOR2_X1 U13499 ( .A(n10943), .B(n10948), .ZN(n10900) );
  XNOR2_X1 U13500 ( .A(n10901), .B(n10900), .ZN(n10907) );
  AOI22_X1 U13501 ( .A1(n13268), .A2(n10902), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10903) );
  OAI21_X1 U13502 ( .B1(n10904), .B2(n13270), .A(n10903), .ZN(n10905) );
  AOI21_X1 U13503 ( .B1(n11443), .B2(n13273), .A(n10905), .ZN(n10906) );
  OAI21_X1 U13504 ( .B1(n10907), .B2(n13275), .A(n10906), .ZN(P2_U3206) );
  AOI22_X1 U13505 ( .A1(n10908), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n13676), .ZN(n10909) );
  OAI21_X1 U13506 ( .B1(n11573), .B2(n11317), .A(n10909), .ZN(P2_U3303) );
  INV_X1 U13507 ( .A(n12092), .ZN(n11257) );
  OAI211_X1 U13508 ( .C1(n11257), .C2(n14731), .A(n10911), .B(n10910), .ZN(
        n10912) );
  AOI21_X1 U13509 ( .B1(n14752), .B2(n10913), .A(n10912), .ZN(n10916) );
  NAND2_X1 U13510 ( .A1(n14761), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10914) );
  OAI21_X1 U13511 ( .B1(n10916), .B2(n14761), .A(n10914), .ZN(P1_U3541) );
  NAND2_X1 U13512 ( .A1(n14753), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10915) );
  OAI21_X1 U13513 ( .B1(n10916), .B2(n14753), .A(n10915), .ZN(P1_U3498) );
  NAND2_X1 U13514 ( .A1(n10918), .A2(n10917), .ZN(n10919) );
  XNOR2_X1 U13515 ( .A(n10919), .B(n12505), .ZN(n10922) );
  AOI21_X1 U13516 ( .B1(n12990), .B2(n12709), .A(n10920), .ZN(n10921) );
  OAI21_X1 U13517 ( .B1(n10922), .B2(n15132), .A(n10921), .ZN(n11001) );
  INV_X1 U13518 ( .A(n11002), .ZN(n10924) );
  AND2_X1 U13519 ( .A1(n10923), .A2(n12505), .ZN(n11000) );
  OR3_X1 U13520 ( .A1(n10924), .A2(n13002), .A3(n11000), .ZN(n10928) );
  AOI22_X1 U13521 ( .A1(n14528), .A2(n10926), .B1(n15140), .B2(n10925), .ZN(
        n10927) );
  OAI211_X1 U13522 ( .C1(n15144), .C2(n10929), .A(n10928), .B(n10927), .ZN(
        n10930) );
  AOI21_X1 U13523 ( .B1(n11001), .B2(n15144), .A(n10930), .ZN(n10931) );
  INV_X1 U13524 ( .A(n10931), .ZN(P3_U3223) );
  NAND2_X1 U13525 ( .A1(n10932), .A2(n6652), .ZN(n10935) );
  AOI22_X1 U13526 ( .A1(n11683), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n11490), 
        .B2(n10933), .ZN(n10934) );
  INV_X1 U13527 ( .A(n13643), .ZN(n11023) );
  NOR2_X1 U13528 ( .A1(n11452), .A2(n10936), .ZN(n10938) );
  XNOR2_X1 U13529 ( .A(n13643), .B(n12012), .ZN(n10937) );
  NOR2_X1 U13530 ( .A1(n10937), .A2(n10938), .ZN(n11068) );
  AOI21_X1 U13531 ( .B1(n10938), .B2(n10937), .A(n11068), .ZN(n10952) );
  INV_X1 U13532 ( .A(n10946), .ZN(n10949) );
  INV_X1 U13533 ( .A(n10948), .ZN(n10945) );
  INV_X1 U13534 ( .A(n10943), .ZN(n10944) );
  OAI21_X1 U13535 ( .B1(n10946), .B2(n10945), .A(n10944), .ZN(n10947) );
  OAI21_X1 U13536 ( .B1(n10949), .B2(n10948), .A(n10947), .ZN(n10950) );
  OAI21_X1 U13537 ( .B1(n10952), .B2(n10951), .A(n6837), .ZN(n10953) );
  NAND2_X1 U13538 ( .A1(n10953), .A2(n13249), .ZN(n10964) );
  AND2_X1 U13539 ( .A1(n10955), .A2(n10954), .ZN(n10956) );
  OR2_X1 U13540 ( .A1(n10956), .A2(n11075), .ZN(n11218) );
  AOI22_X1 U13541 ( .A1(n11686), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n10957), 
        .B2(P2_REG2_REG_15__SCAN_IN), .ZN(n10959) );
  NAND2_X1 U13542 ( .A1(n11642), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n10958) );
  INV_X1 U13543 ( .A(n13288), .ZN(n11167) );
  INV_X1 U13544 ( .A(n11020), .ZN(n10960) );
  OAI22_X1 U13545 ( .A1(n13258), .A2(n11167), .B1(n13270), .B2(n10960), .ZN(
        n10961) );
  AOI211_X1 U13546 ( .C1(n13244), .C2(n13290), .A(n10962), .B(n10961), .ZN(
        n10963) );
  OAI211_X1 U13547 ( .C1(n11023), .C2(n13242), .A(n10964), .B(n10963), .ZN(
        P2_U3187) );
  OAI222_X1 U13548 ( .A1(P1_U3086), .A2(n10966), .B1(n14330), .B2(n11573), 
        .C1(n10965), .C2(n14332), .ZN(P1_U3331) );
  INV_X1 U13549 ( .A(n14584), .ZN(n10968) );
  OAI21_X1 U13550 ( .B1(n10968), .B2(n14731), .A(n10967), .ZN(n10969) );
  AOI211_X1 U13551 ( .C1(n10971), .C2(n14752), .A(n10970), .B(n10969), .ZN(
        n10974) );
  NAND2_X1 U13552 ( .A1(n14753), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10972) );
  OAI21_X1 U13553 ( .B1(n10974), .B2(n14753), .A(n10972), .ZN(P1_U3501) );
  NAND2_X1 U13554 ( .A1(n14761), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10973) );
  OAI21_X1 U13555 ( .B1(n10974), .B2(n14761), .A(n10973), .ZN(P1_U3542) );
  INV_X1 U13556 ( .A(n10975), .ZN(n10976) );
  AOI21_X1 U13557 ( .B1(n12511), .B2(n10977), .A(n10976), .ZN(n14539) );
  INV_X1 U13558 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n15498) );
  INV_X1 U13559 ( .A(n10978), .ZN(n11033) );
  OAI22_X1 U13560 ( .A1(n15144), .A2(n15498), .B1(n11033), .B2(n15108), .ZN(
        n10979) );
  AOI21_X1 U13561 ( .B1(n14528), .B2(n11037), .A(n10979), .ZN(n10989) );
  NAND2_X1 U13562 ( .A1(n10981), .A2(n10980), .ZN(n10983) );
  AND2_X1 U13563 ( .A1(n10983), .A2(n10982), .ZN(n10984) );
  XNOR2_X1 U13564 ( .A(n10984), .B(n12511), .ZN(n10987) );
  OR2_X1 U13565 ( .A1(n11028), .A2(n15134), .ZN(n10986) );
  NAND2_X1 U13566 ( .A1(n11235), .A2(n12990), .ZN(n10985) );
  AND2_X1 U13567 ( .A1(n10986), .A2(n10985), .ZN(n11034) );
  OAI21_X1 U13568 ( .B1(n10987), .B2(n15132), .A(n11034), .ZN(n14540) );
  NAND2_X1 U13569 ( .A1(n14540), .A2(n15144), .ZN(n10988) );
  OAI211_X1 U13570 ( .C1(n14539), .C2(n13002), .A(n10989), .B(n10988), .ZN(
        P3_U3222) );
  XNOR2_X1 U13571 ( .A(n10990), .B(n12234), .ZN(n11106) );
  INV_X1 U13572 ( .A(n11106), .ZN(n10999) );
  OAI211_X1 U13573 ( .C1(n10992), .C2(n12234), .A(n10991), .B(n14144), .ZN(
        n10993) );
  AOI22_X1 U13574 ( .A1(n13825), .A2(n14079), .B1(n13827), .B2(n14082), .ZN(
        n13809) );
  NAND2_X1 U13575 ( .A1(n10993), .A2(n13809), .ZN(n11104) );
  INV_X1 U13576 ( .A(n11098), .ZN(n10994) );
  AOI211_X1 U13577 ( .C1(n13815), .C2(n6785), .A(n14661), .B(n10994), .ZN(
        n11105) );
  NAND2_X1 U13578 ( .A1(n11105), .A2(n14165), .ZN(n10996) );
  AOI22_X1 U13579 ( .A1(n14678), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13805), 
        .B2(n14180), .ZN(n10995) );
  OAI211_X1 U13580 ( .C1(n8817), .C2(n14156), .A(n10996), .B(n10995), .ZN(
        n10997) );
  AOI21_X1 U13581 ( .B1(n14668), .B2(n11104), .A(n10997), .ZN(n10998) );
  OAI21_X1 U13582 ( .B1(n14167), .B2(n10999), .A(n10998), .ZN(P1_U3278) );
  INV_X1 U13583 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11004) );
  NOR2_X1 U13584 ( .A1(n11000), .A2(n15172), .ZN(n11003) );
  AOI21_X1 U13585 ( .B1(n11003), .B2(n11002), .A(n11001), .ZN(n11006) );
  MUX2_X1 U13586 ( .A(n11004), .B(n11006), .S(n15197), .Z(n11005) );
  OAI21_X1 U13587 ( .B1(n13131), .B2(n11008), .A(n11005), .ZN(P3_U3420) );
  INV_X1 U13588 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15499) );
  MUX2_X1 U13589 ( .A(n15499), .B(n11006), .S(n15213), .Z(n11007) );
  OAI21_X1 U13590 ( .B1(n13073), .B2(n11008), .A(n11007), .ZN(P3_U3469) );
  XNOR2_X1 U13591 ( .A(n13643), .B(n11452), .ZN(n11738) );
  NAND2_X1 U13592 ( .A1(n11009), .A2(n7075), .ZN(n11011) );
  XOR2_X1 U13593 ( .A(n11738), .B(n11182), .Z(n13645) );
  INV_X1 U13594 ( .A(n13290), .ZN(n11445) );
  NAND2_X1 U13595 ( .A1(n11443), .A2(n11445), .ZN(n11012) );
  OR2_X1 U13596 ( .A1(n11443), .A2(n11445), .ZN(n11014) );
  INV_X1 U13597 ( .A(n11166), .ZN(n11015) );
  AOI21_X1 U13598 ( .B1(n11738), .B2(n11016), .A(n11015), .ZN(n11017) );
  OAI222_X1 U13599 ( .A1(n13540), .A2(n11167), .B1(n13538), .B2(n11445), .C1(
        n14548), .C2(n11017), .ZN(n13641) );
  OR2_X1 U13600 ( .A1(n13643), .A2(n11019), .ZN(n11217) );
  INV_X1 U13601 ( .A(n11217), .ZN(n11018) );
  AOI211_X1 U13602 ( .C1(n13643), .C2(n11019), .A(n13459), .B(n11018), .ZN(
        n13642) );
  NAND2_X1 U13603 ( .A1(n13642), .A2(n15590), .ZN(n11022) );
  AOI22_X1 U13604 ( .A1(n14556), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11020), 
        .B2(n14555), .ZN(n11021) );
  OAI211_X1 U13605 ( .C1(n11023), .C2(n13528), .A(n11022), .B(n11021), .ZN(
        n11024) );
  AOI21_X1 U13606 ( .B1(n13641), .B2(n13441), .A(n11024), .ZN(n11025) );
  OAI21_X1 U13607 ( .B1(n13496), .B2(n13645), .A(n11025), .ZN(P2_U3251) );
  INV_X1 U13608 ( .A(n11026), .ZN(n11027) );
  OR2_X1 U13609 ( .A1(n11028), .A2(n11027), .ZN(n11029) );
  INV_X1 U13610 ( .A(n11138), .ZN(n11031) );
  AOI21_X1 U13611 ( .B1(n12709), .B2(n11032), .A(n11031), .ZN(n11039) );
  NOR2_X1 U13612 ( .A1(n12418), .A2(n11033), .ZN(n11036) );
  NAND2_X1 U13613 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(P3_U3151), .ZN(n15032)
         );
  OAI21_X1 U13614 ( .B1(n11034), .B2(n12454), .A(n15032), .ZN(n11035) );
  AOI211_X1 U13615 ( .C1(n12456), .C2(n11037), .A(n11036), .B(n11035), .ZN(
        n11038) );
  OAI21_X1 U13616 ( .B1(n11039), .B2(n12459), .A(n11038), .ZN(P3_U3176) );
  INV_X1 U13617 ( .A(n11040), .ZN(n11042) );
  OAI222_X1 U13618 ( .A1(P3_U3151), .A2(n11043), .B1(n11060), .B2(n11042), 
        .C1(n11041), .C2(n12350), .ZN(P3_U3270) );
  INV_X1 U13619 ( .A(n11044), .ZN(n11045) );
  NAND2_X1 U13620 ( .A1(n11046), .A2(n11045), .ZN(n11047) );
  OAI21_X1 U13621 ( .B1(n11048), .B2(n11051), .A(n11047), .ZN(n13958) );
  XNOR2_X1 U13622 ( .A(n11057), .B(n13958), .ZN(n11049) );
  NAND2_X1 U13623 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11049), .ZN(n13961) );
  OAI211_X1 U13624 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n11049), .A(n13963), 
        .B(n13961), .ZN(n11056) );
  NAND2_X1 U13625 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13785)
         );
  OAI21_X1 U13626 ( .B1(n14271), .B2(n11051), .A(n11050), .ZN(n13954) );
  XNOR2_X1 U13627 ( .A(n13954), .B(n11057), .ZN(n11052) );
  NAND2_X1 U13628 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n11052), .ZN(n13956) );
  OAI211_X1 U13629 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11052), .A(n13966), 
        .B(n13956), .ZN(n11053) );
  NAND2_X1 U13630 ( .A1(n13785), .A2(n11053), .ZN(n11054) );
  AOI21_X1 U13631 ( .B1(n13929), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11054), 
        .ZN(n11055) );
  OAI211_X1 U13632 ( .C1(n14647), .C2(n11057), .A(n11056), .B(n11055), .ZN(
        P1_U3261) );
  INV_X1 U13633 ( .A(n11058), .ZN(n11059) );
  OAI222_X1 U13634 ( .A1(P3_U3151), .A2(n11061), .B1(n12350), .B2(n15444), 
        .C1(n11060), .C2(n11059), .ZN(P3_U3269) );
  NAND2_X1 U13635 ( .A1(n11062), .A2(n6652), .ZN(n11065) );
  AOI22_X1 U13636 ( .A1(n11683), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n11490), 
        .B2(n11063), .ZN(n11064) );
  INV_X1 U13637 ( .A(n13637), .ZN(n11221) );
  AND2_X1 U13638 ( .A1(n13288), .A2(n13459), .ZN(n11067) );
  XNOR2_X1 U13639 ( .A(n13637), .B(n12012), .ZN(n11066) );
  NOR2_X1 U13640 ( .A1(n11066), .A2(n11067), .ZN(n11197) );
  AOI21_X1 U13641 ( .B1(n11067), .B2(n11066), .A(n11197), .ZN(n11072) );
  INV_X1 U13642 ( .A(n11068), .ZN(n11069) );
  OAI21_X1 U13643 ( .B1(n11072), .B2(n11071), .A(n11198), .ZN(n11073) );
  NAND2_X1 U13644 ( .A1(n11073), .A2(n13249), .ZN(n11082) );
  INV_X1 U13645 ( .A(n11452), .ZN(n13289) );
  INV_X1 U13646 ( .A(n11074), .ZN(n11080) );
  NOR2_X1 U13647 ( .A1(n11075), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11076) );
  OR2_X1 U13648 ( .A1(n11173), .A2(n11076), .ZN(n11203) );
  AOI22_X1 U13649 ( .A1(n11642), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n11686), 
        .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n11078) );
  OR2_X1 U13650 ( .A1(n11605), .A2(n10547), .ZN(n11077) );
  OAI211_X1 U13651 ( .C1(n11203), .C2(n11551), .A(n11078), .B(n11077), .ZN(
        n13287) );
  INV_X1 U13652 ( .A(n13287), .ZN(n11273) );
  OAI22_X1 U13653 ( .A1(n13258), .A2(n11273), .B1(n13270), .B2(n11218), .ZN(
        n11079) );
  AOI211_X1 U13654 ( .C1(n13244), .C2(n13289), .A(n11080), .B(n11079), .ZN(
        n11081) );
  OAI211_X1 U13655 ( .C1(n11221), .C2(n13242), .A(n11082), .B(n11081), .ZN(
        P2_U3213) );
  XOR2_X1 U13656 ( .A(n12512), .B(n11083), .Z(n11086) );
  NAND2_X1 U13657 ( .A1(n12992), .A2(n12990), .ZN(n11085) );
  NAND2_X1 U13658 ( .A1(n12709), .A2(n12993), .ZN(n11084) );
  NAND2_X1 U13659 ( .A1(n11085), .A2(n11084), .ZN(n11141) );
  AOI21_X1 U13660 ( .B1(n11086), .B2(n12987), .A(n11141), .ZN(n14534) );
  XNOR2_X1 U13661 ( .A(n11087), .B(n12512), .ZN(n14537) );
  NOR2_X1 U13662 ( .A1(n14535), .A2(n12998), .ZN(n11091) );
  INV_X1 U13663 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11089) );
  INV_X1 U13664 ( .A(n11088), .ZN(n11143) );
  OAI22_X1 U13665 ( .A1(n15144), .A2(n11089), .B1(n11143), .B2(n15108), .ZN(
        n11090) );
  AOI211_X1 U13666 ( .C1(n14537), .C2(n15141), .A(n11091), .B(n11090), .ZN(
        n11092) );
  OAI21_X1 U13667 ( .B1(n14534), .B2(n15146), .A(n11092), .ZN(P3_U3221) );
  OAI21_X1 U13668 ( .B1(n6794), .B2(n7556), .A(n11093), .ZN(n11094) );
  AOI222_X1 U13669 ( .A1(n14144), .A2(n11094), .B1(n13824), .B2(n14079), .C1(
        n13826), .C2(n14082), .ZN(n14278) );
  OAI21_X1 U13670 ( .B1(n11096), .B2(n12230), .A(n11095), .ZN(n14274) );
  INV_X1 U13671 ( .A(n14276), .ZN(n13751) );
  INV_X1 U13672 ( .A(n11157), .ZN(n11097) );
  AOI211_X1 U13673 ( .C1(n14276), .C2(n11098), .A(n14661), .B(n11097), .ZN(
        n14275) );
  NAND2_X1 U13674 ( .A1(n14275), .A2(n14165), .ZN(n11101) );
  INV_X1 U13675 ( .A(n13746), .ZN(n11099) );
  AOI22_X1 U13676 ( .A1(n14678), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11099), 
        .B2(n14180), .ZN(n11100) );
  OAI211_X1 U13677 ( .C1(n13751), .C2(n14156), .A(n11101), .B(n11100), .ZN(
        n11102) );
  AOI21_X1 U13678 ( .B1(n14188), .B2(n14274), .A(n11102), .ZN(n11103) );
  OAI21_X1 U13679 ( .B1(n14278), .B2(n14678), .A(n11103), .ZN(P1_U3277) );
  AOI211_X1 U13680 ( .C1(n11106), .C2(n14752), .A(n11105), .B(n11104), .ZN(
        n11108) );
  MUX2_X1 U13681 ( .A(n15452), .B(n11108), .S(n14755), .Z(n11107) );
  OAI21_X1 U13682 ( .B1(n8817), .B2(n14318), .A(n11107), .ZN(P1_U3504) );
  MUX2_X1 U13683 ( .A(n11109), .B(n11108), .S(n14764), .Z(n11110) );
  OAI21_X1 U13684 ( .B1(n8817), .B2(n14273), .A(n11110), .ZN(P1_U3543) );
  INV_X1 U13685 ( .A(n11111), .ZN(n11113) );
  OAI222_X1 U13686 ( .A1(P3_U3151), .A2(n12758), .B1(n11060), .B2(n11113), 
        .C1(n11112), .C2(n12350), .ZN(P3_U3268) );
  INV_X1 U13687 ( .A(n11114), .ZN(n11117) );
  AOI22_X1 U13688 ( .A1(n14607), .A2(n12326), .B1(n12323), .B2(n13830), .ZN(
        n11120) );
  XNOR2_X1 U13689 ( .A(n11120), .B(n12324), .ZN(n11122) );
  AOI22_X1 U13690 ( .A1(n14607), .A2(n12323), .B1(n12322), .B2(n13830), .ZN(
        n11121) );
  XNOR2_X1 U13691 ( .A(n11122), .B(n11121), .ZN(n14597) );
  NAND2_X1 U13692 ( .A1(n12082), .A2(n12326), .ZN(n11124) );
  NAND2_X1 U13693 ( .A1(n13829), .A2(n12323), .ZN(n11123) );
  NAND2_X1 U13694 ( .A1(n11124), .A2(n11123), .ZN(n11125) );
  XNOR2_X1 U13695 ( .A(n11125), .B(n12324), .ZN(n11242) );
  AND2_X1 U13696 ( .A1(n13829), .A2(n12322), .ZN(n11126) );
  AOI21_X1 U13697 ( .B1(n12082), .B2(n12323), .A(n11126), .ZN(n11245) );
  XNOR2_X1 U13698 ( .A(n11242), .B(n11245), .ZN(n11127) );
  NAND2_X1 U13699 ( .A1(n11128), .A2(n11127), .ZN(n11243) );
  OAI211_X1 U13700 ( .C1(n11128), .C2(n11127), .A(n11243), .B(n14585), .ZN(
        n11134) );
  OAI22_X1 U13701 ( .A1(n13808), .A2(n11130), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11129), .ZN(n11131) );
  AOI21_X1 U13702 ( .B1(n13806), .B2(n11132), .A(n11131), .ZN(n11133) );
  OAI211_X1 U13703 ( .C1(n11135), .C2(n13792), .A(n11134), .B(n11133), .ZN(
        P1_U3224) );
  XNOR2_X1 U13704 ( .A(n11136), .B(n11895), .ZN(n11231) );
  XNOR2_X1 U13705 ( .A(n11231), .B(n11235), .ZN(n11140) );
  NAND2_X1 U13706 ( .A1(n11138), .A2(n11137), .ZN(n11139) );
  NAND2_X1 U13707 ( .A1(n11139), .A2(n11140), .ZN(n11233) );
  OAI21_X1 U13708 ( .B1(n11140), .B2(n11139), .A(n11233), .ZN(n11146) );
  NOR2_X1 U13709 ( .A1(n14535), .A2(n12446), .ZN(n11145) );
  NAND2_X1 U13710 ( .A1(n11141), .A2(n12416), .ZN(n11142) );
  NAND2_X1 U13711 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n15052)
         );
  OAI211_X1 U13712 ( .C1(n12418), .C2(n11143), .A(n11142), .B(n15052), .ZN(
        n11144) );
  AOI211_X1 U13713 ( .C1(n11146), .C2(n12436), .A(n11145), .B(n11144), .ZN(
        n11147) );
  INV_X1 U13714 ( .A(n11147), .ZN(P3_U3164) );
  XNOR2_X1 U13715 ( .A(n11148), .B(n12599), .ZN(n13070) );
  INV_X1 U13716 ( .A(n13070), .ZN(n11155) );
  AOI21_X1 U13717 ( .B1(n12599), .B2(n11150), .A(n11149), .ZN(n11151) );
  OAI222_X1 U13718 ( .A1(n15136), .A2(n11297), .B1(n15134), .B2(n11230), .C1(
        n15132), .C2(n11151), .ZN(n13069) );
  AOI22_X1 U13719 ( .A1(n15146), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15140), 
        .B2(n11239), .ZN(n11152) );
  OAI21_X1 U13720 ( .B1(n13130), .B2(n12998), .A(n11152), .ZN(n11153) );
  AOI21_X1 U13721 ( .B1(n13069), .B2(n15144), .A(n11153), .ZN(n11154) );
  OAI21_X1 U13722 ( .B1(n13002), .B2(n11155), .A(n11154), .ZN(P3_U3220) );
  XNOR2_X1 U13723 ( .A(n13761), .B(n13745), .ZN(n12232) );
  XOR2_X1 U13724 ( .A(n12232), .B(n11156), .Z(n14266) );
  AOI211_X1 U13725 ( .C1(n13761), .C2(n11157), .A(n14661), .B(n11287), .ZN(
        n14268) );
  INV_X1 U13726 ( .A(n13761), .ZN(n14319) );
  AOI22_X1 U13727 ( .A1(n14678), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n13756), 
        .B2(n14180), .ZN(n11158) );
  OAI21_X1 U13728 ( .B1(n14319), .B2(n14156), .A(n11158), .ZN(n11159) );
  AOI21_X1 U13729 ( .B1(n14268), .B2(n14165), .A(n11159), .ZN(n11164) );
  XNOR2_X1 U13730 ( .A(n11160), .B(n12232), .ZN(n11161) );
  NOR2_X1 U13731 ( .A1(n11161), .A2(n14656), .ZN(n14269) );
  AND2_X1 U13732 ( .A1(n13825), .A2(n14082), .ZN(n11162) );
  AOI21_X1 U13733 ( .B1(n13823), .B2(n14079), .A(n11162), .ZN(n13759) );
  INV_X1 U13734 ( .A(n13759), .ZN(n14267) );
  OAI21_X1 U13735 ( .B1(n14269), .B2(n14267), .A(n14668), .ZN(n11163) );
  OAI211_X1 U13736 ( .C1(n14266), .C2(n14167), .A(n11164), .B(n11163), .ZN(
        P1_U3276) );
  NAND2_X1 U13737 ( .A1(n13643), .A2(n11452), .ZN(n11165) );
  NAND2_X1 U13738 ( .A1(n11166), .A2(n11165), .ZN(n11223) );
  XNOR2_X1 U13739 ( .A(n13637), .B(n13288), .ZN(n11740) );
  INV_X1 U13740 ( .A(n11740), .ZN(n11222) );
  OR2_X1 U13741 ( .A1(n13637), .A2(n11167), .ZN(n11168) );
  NAND2_X1 U13742 ( .A1(n11169), .A2(n6652), .ZN(n11172) );
  AOI22_X1 U13743 ( .A1(n11683), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n11490), 
        .B2(n11170), .ZN(n11171) );
  XNOR2_X1 U13744 ( .A(n13632), .B(n13287), .ZN(n11737) );
  XNOR2_X1 U13745 ( .A(n11258), .B(n11186), .ZN(n11180) );
  OR2_X1 U13746 ( .A1(n11173), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11174) );
  AND2_X1 U13747 ( .A1(n11265), .A2(n11174), .ZN(n13207) );
  NAND2_X1 U13748 ( .A1(n13207), .A2(n11658), .ZN(n11179) );
  INV_X1 U13749 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13318) );
  NAND2_X1 U13750 ( .A1(n11642), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n11176) );
  NAND2_X1 U13751 ( .A1(n11686), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n11175) );
  OAI211_X1 U13752 ( .C1(n13318), .C2(n11605), .A(n11176), .B(n11175), .ZN(
        n11177) );
  INV_X1 U13753 ( .A(n11177), .ZN(n11178) );
  AOI222_X1 U13754 ( .A1(n13521), .A2(n11180), .B1(n13286), .B2(n13650), .C1(
        n13288), .C2(n13470), .ZN(n13634) );
  NOR2_X1 U13755 ( .A1(n13643), .A2(n13289), .ZN(n11181) );
  NAND2_X1 U13756 ( .A1(n13643), .A2(n13289), .ZN(n11183) );
  NOR2_X1 U13757 ( .A1(n13637), .A2(n13288), .ZN(n11185) );
  OAI21_X1 U13758 ( .B1(n11187), .B2(n11186), .A(n11276), .ZN(n13635) );
  NAND2_X1 U13759 ( .A1(n15599), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11188) );
  OAI21_X1 U13760 ( .B1(n15592), .B2(n11203), .A(n11188), .ZN(n11189) );
  AOI21_X1 U13761 ( .B1(n13632), .B2(n14557), .A(n11189), .ZN(n11192) );
  AOI21_X1 U13762 ( .B1(n11215), .B2(n13632), .A(n13459), .ZN(n11190) );
  AND2_X1 U13763 ( .A1(n11190), .A2(n6787), .ZN(n13631) );
  NAND2_X1 U13764 ( .A1(n13631), .A2(n15590), .ZN(n11191) );
  OAI211_X1 U13765 ( .C1(n13635), .C2(n13496), .A(n11192), .B(n11191), .ZN(
        n11193) );
  INV_X1 U13766 ( .A(n11193), .ZN(n11194) );
  OAI21_X1 U13767 ( .B1(n13634), .B2(n14556), .A(n11194), .ZN(P2_U3249) );
  INV_X1 U13768 ( .A(n13632), .ZN(n11208) );
  AND2_X1 U13769 ( .A1(n13287), .A2(n13459), .ZN(n11196) );
  XNOR2_X1 U13770 ( .A(n13632), .B(n12012), .ZN(n11195) );
  NOR2_X1 U13771 ( .A1(n11195), .A2(n11196), .ZN(n11969) );
  AOI21_X1 U13772 ( .B1(n11196), .B2(n11195), .A(n11969), .ZN(n11200) );
  OAI21_X1 U13773 ( .B1(n11200), .B2(n11199), .A(n11971), .ZN(n11201) );
  NAND2_X1 U13774 ( .A1(n11201), .A2(n13249), .ZN(n11207) );
  INV_X1 U13775 ( .A(n11202), .ZN(n11205) );
  OAI22_X1 U13776 ( .A1(n13258), .A2(n13539), .B1(n13270), .B2(n11203), .ZN(
        n11204) );
  AOI211_X1 U13777 ( .C1(n13244), .C2(n13288), .A(n11205), .B(n11204), .ZN(
        n11206) );
  OAI211_X1 U13778 ( .C1(n11208), .C2(n13242), .A(n11207), .B(n11206), .ZN(
        P2_U3198) );
  INV_X1 U13779 ( .A(n11587), .ZN(n11213) );
  OAI222_X1 U13780 ( .A1(n13693), .A2(n11211), .B1(n11317), .B2(n11213), .C1(
        n11210), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U13781 ( .A1(n14332), .A2(n11214), .B1(n14330), .B2(n11213), .C1(
        P1_U3086), .C2(n11212), .ZN(P1_U3330) );
  XNOR2_X1 U13782 ( .A(n6807), .B(n11740), .ZN(n13640) );
  INV_X1 U13783 ( .A(n11215), .ZN(n11216) );
  AOI211_X1 U13784 ( .C1(n13637), .C2(n11217), .A(n13459), .B(n11216), .ZN(
        n13636) );
  INV_X1 U13785 ( .A(n11218), .ZN(n11219) );
  AOI22_X1 U13786 ( .A1(n15599), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11219), 
        .B2(n14555), .ZN(n11220) );
  OAI21_X1 U13787 ( .B1(n11221), .B2(n13528), .A(n11220), .ZN(n11228) );
  AOI21_X1 U13788 ( .B1(n11223), .B2(n11222), .A(n14548), .ZN(n11226) );
  OAI22_X1 U13789 ( .A1(n11273), .A2(n13540), .B1(n11452), .B2(n13538), .ZN(
        n11224) );
  AOI21_X1 U13790 ( .B1(n11226), .B2(n11225), .A(n11224), .ZN(n13639) );
  NOR2_X1 U13791 ( .A1(n13639), .A2(n15599), .ZN(n11227) );
  AOI211_X1 U13792 ( .C1(n13636), .C2(n15590), .A(n11228), .B(n11227), .ZN(
        n11229) );
  OAI21_X1 U13793 ( .B1(n13640), .B2(n13496), .A(n11229), .ZN(P2_U3250) );
  NAND2_X1 U13794 ( .A1(n11231), .A2(n11230), .ZN(n11232) );
  NAND2_X1 U13795 ( .A1(n11233), .A2(n11232), .ZN(n11296) );
  XNOR2_X1 U13796 ( .A(n13130), .B(n11886), .ZN(n11295) );
  XNOR2_X1 U13797 ( .A(n11295), .B(n11303), .ZN(n11234) );
  XNOR2_X1 U13798 ( .A(n11296), .B(n11234), .ZN(n11241) );
  AOI22_X1 U13799 ( .A1(n11899), .A2(n11235), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11236) );
  OAI21_X1 U13800 ( .B1(n11297), .B2(n12368), .A(n11236), .ZN(n11238) );
  NOR2_X1 U13801 ( .A1(n13130), .A2(n12446), .ZN(n11237) );
  AOI211_X1 U13802 ( .C1(n11239), .C2(n12451), .A(n11238), .B(n11237), .ZN(
        n11240) );
  OAI21_X1 U13803 ( .B1(n11241), .B2(n12459), .A(n11240), .ZN(P3_U3174) );
  INV_X1 U13804 ( .A(n11242), .ZN(n11244) );
  AND2_X1 U13805 ( .A1(n13828), .A2(n12322), .ZN(n11246) );
  AOI21_X1 U13806 ( .B1(n12092), .B2(n12323), .A(n11246), .ZN(n11776) );
  AOI22_X1 U13807 ( .A1(n12092), .A2(n12326), .B1(n12323), .B2(n13828), .ZN(
        n11247) );
  XNOR2_X1 U13808 ( .A(n11247), .B(n12324), .ZN(n11775) );
  XOR2_X1 U13809 ( .A(n11776), .B(n11775), .Z(n11248) );
  OAI211_X1 U13810 ( .C1(n11249), .C2(n11248), .A(n11780), .B(n14585), .ZN(
        n11256) );
  INV_X1 U13811 ( .A(n11250), .ZN(n11253) );
  NOR2_X1 U13812 ( .A1(n14606), .A2(n11251), .ZN(n11252) );
  AOI211_X1 U13813 ( .C1(n14587), .C2(n11254), .A(n11253), .B(n11252), .ZN(
        n11255) );
  OAI211_X1 U13814 ( .C1(n11257), .C2(n13792), .A(n11256), .B(n11255), .ZN(
        P1_U3234) );
  OR2_X1 U13815 ( .A1(n13632), .A2(n11273), .ZN(n11259) );
  NAND2_X1 U13816 ( .A1(n11260), .A2(n11259), .ZN(n11934) );
  NAND2_X1 U13817 ( .A1(n11261), .A2(n6652), .ZN(n11263) );
  INV_X1 U13818 ( .A(n13328), .ZN(n14840) );
  AOI22_X1 U13819 ( .A1(n11683), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n14840), 
        .B2(n11490), .ZN(n11262) );
  XNOR2_X1 U13820 ( .A(n13627), .B(n13539), .ZN(n11905) );
  XNOR2_X1 U13821 ( .A(n11934), .B(n11905), .ZN(n11274) );
  NAND2_X1 U13822 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  NAND2_X1 U13823 ( .A1(n11494), .A2(n11266), .ZN(n13546) );
  OR2_X1 U13824 ( .A1(n13546), .A2(n11551), .ZN(n11272) );
  INV_X1 U13825 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U13826 ( .A1(n11642), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n11268) );
  INV_X1 U13827 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13547) );
  OR2_X1 U13828 ( .A1(n11605), .A2(n13547), .ZN(n11267) );
  OAI211_X1 U13829 ( .C1(n9466), .C2(n11269), .A(n11268), .B(n11267), .ZN(
        n11270) );
  INV_X1 U13830 ( .A(n11270), .ZN(n11271) );
  NAND2_X1 U13831 ( .A1(n11272), .A2(n11271), .ZN(n13285) );
  INV_X1 U13832 ( .A(n13285), .ZN(n13174) );
  OAI22_X1 U13833 ( .A1(n13174), .A2(n13540), .B1(n11273), .B2(n13538), .ZN(
        n13206) );
  AOI21_X1 U13834 ( .B1(n11274), .B2(n13521), .A(n13206), .ZN(n13629) );
  NAND2_X1 U13835 ( .A1(n13632), .A2(n13287), .ZN(n11275) );
  XNOR2_X1 U13836 ( .A(n11906), .B(n11905), .ZN(n13630) );
  INV_X1 U13837 ( .A(n13630), .ZN(n11282) );
  NAND2_X1 U13838 ( .A1(n6787), .A2(n13627), .ZN(n11277) );
  NAND2_X1 U13839 ( .A1(n11277), .A2(n10936), .ZN(n11278) );
  NOR2_X1 U13840 ( .A1(n6788), .A2(n11278), .ZN(n13626) );
  NAND2_X1 U13841 ( .A1(n13626), .A2(n15590), .ZN(n11280) );
  AOI22_X1 U13842 ( .A1(n15599), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13207), 
        .B2(n14555), .ZN(n11279) );
  OAI211_X1 U13843 ( .C1(n7062), .C2(n13528), .A(n11280), .B(n11279), .ZN(
        n11281) );
  AOI21_X1 U13844 ( .B1(n11282), .B2(n14563), .A(n11281), .ZN(n11283) );
  OAI21_X1 U13845 ( .B1(n15599), .B2(n13629), .A(n11283), .ZN(P2_U3248) );
  XNOR2_X1 U13846 ( .A(n11284), .B(n6876), .ZN(n11285) );
  OAI22_X1 U13847 ( .A1(n11285), .A2(n14656), .B1(n13745), .B2(n14170), .ZN(
        n14262) );
  INV_X1 U13848 ( .A(n14262), .ZN(n11294) );
  XNOR2_X1 U13849 ( .A(n11286), .B(n6876), .ZN(n14264) );
  OAI211_X1 U13850 ( .C1(n11287), .C2(n14314), .A(n14175), .B(n14176), .ZN(
        n14259) );
  NOR2_X1 U13851 ( .A1(n14183), .A2(n14261), .ZN(n11290) );
  OAI22_X1 U13852 ( .A1(n14668), .A2(n11288), .B1(n13786), .B2(n14665), .ZN(
        n11289) );
  AOI211_X1 U13853 ( .C1(n11807), .C2(n14670), .A(n11290), .B(n11289), .ZN(
        n11291) );
  OAI21_X1 U13854 ( .B1(n14259), .B2(n14673), .A(n11291), .ZN(n11292) );
  AOI21_X1 U13855 ( .B1(n14264), .B2(n14188), .A(n11292), .ZN(n11293) );
  OAI21_X1 U13856 ( .B1(n11294), .B2(n14678), .A(n11293), .ZN(P1_U3275) );
  XNOR2_X1 U13857 ( .A(n13066), .B(n11886), .ZN(n11299) );
  INV_X1 U13858 ( .A(n11299), .ZN(n11298) );
  NAND2_X1 U13859 ( .A1(n11298), .A2(n11297), .ZN(n11309) );
  NAND2_X1 U13860 ( .A1(n11299), .A2(n12708), .ZN(n11307) );
  NAND2_X1 U13861 ( .A1(n11309), .A2(n11307), .ZN(n11300) );
  XNOR2_X1 U13862 ( .A(n11308), .B(n11300), .ZN(n11306) );
  AOI22_X1 U13863 ( .A1(n12440), .A2(n12991), .B1(P3_REG3_REG_14__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11302) );
  NAND2_X1 U13864 ( .A1(n12451), .A2(n12996), .ZN(n11301) );
  OAI211_X1 U13865 ( .C1(n11303), .C2(n12442), .A(n11302), .B(n11301), .ZN(
        n11304) );
  AOI21_X1 U13866 ( .B1(n12456), .B2(n13066), .A(n11304), .ZN(n11305) );
  OAI21_X1 U13867 ( .B1(n11306), .B2(n12459), .A(n11305), .ZN(P3_U3155) );
  XNOR2_X1 U13868 ( .A(n11311), .B(n11886), .ZN(n11857) );
  XNOR2_X1 U13869 ( .A(n11857), .B(n12991), .ZN(n11310) );
  XNOR2_X1 U13870 ( .A(n11856), .B(n11310), .ZN(n11315) );
  AOI22_X1 U13871 ( .A1(n12708), .A2(n12993), .B1(n12990), .B2(n12946), .ZN(
        n12975) );
  INV_X1 U13872 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n14467) );
  OAI22_X1 U13873 ( .A1(n12975), .A2(n12454), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14467), .ZN(n11313) );
  INV_X1 U13874 ( .A(n11311), .ZN(n13125) );
  NOR2_X1 U13875 ( .A1(n13125), .A2(n12446), .ZN(n11312) );
  AOI211_X1 U13876 ( .C1(n12980), .C2(n12451), .A(n11313), .B(n11312), .ZN(
        n11314) );
  OAI21_X1 U13877 ( .B1(n11315), .B2(n12459), .A(n11314), .ZN(P3_U3181) );
  INV_X1 U13878 ( .A(n11651), .ZN(n11967) );
  OAI222_X1 U13879 ( .A1(n11318), .A2(P2_U3088), .B1(n11317), .B2(n11967), 
        .C1(n11316), .C2(n13693), .ZN(P2_U3301) );
  OAI222_X1 U13880 ( .A1(n12350), .A2(n7396), .B1(n11060), .B2(n11320), .C1(
        n11319), .C2(P3_U3151), .ZN(P3_U3267) );
  NAND2_X1 U13881 ( .A1(n11323), .A2(n11380), .ZN(n11326) );
  NAND2_X1 U13882 ( .A1(n11326), .A2(n11325), .ZN(n11341) );
  INV_X1 U13883 ( .A(n11327), .ZN(n11328) );
  OR2_X1 U13884 ( .A1(n11759), .A2(n11328), .ZN(n11333) );
  NAND3_X1 U13885 ( .A1(n11330), .A2(n11329), .A3(n11333), .ZN(n11335) );
  OAI211_X1 U13886 ( .C1(n11333), .C2(n11332), .A(n11380), .B(n11331), .ZN(
        n11334) );
  NAND2_X1 U13887 ( .A1(n11335), .A2(n11334), .ZN(n11340) );
  NAND2_X1 U13888 ( .A1(n11341), .A2(n11340), .ZN(n11339) );
  NAND2_X1 U13889 ( .A1(n11380), .A2(n13179), .ZN(n11336) );
  NAND2_X1 U13890 ( .A1(n11339), .A2(n11338), .ZN(n11345) );
  INV_X1 U13891 ( .A(n11340), .ZN(n11343) );
  INV_X1 U13892 ( .A(n11341), .ZN(n11342) );
  NAND2_X1 U13893 ( .A1(n11343), .A2(n11342), .ZN(n11344) );
  NAND2_X1 U13894 ( .A1(n11345), .A2(n11344), .ZN(n11352) );
  NAND2_X1 U13895 ( .A1(n11516), .A2(n13246), .ZN(n11347) );
  NAND2_X1 U13896 ( .A1(n11348), .A2(n11347), .ZN(n11351) );
  AOI22_X1 U13897 ( .A1(n11716), .A2(n13246), .B1(n11346), .B2(n11516), .ZN(
        n11349) );
  AOI21_X1 U13898 ( .B1(n11352), .B2(n11351), .A(n11349), .ZN(n11350) );
  INV_X1 U13899 ( .A(n11350), .ZN(n11353) );
  OR2_X1 U13900 ( .A1(n6655), .A2(n11354), .ZN(n11356) );
  NAND2_X1 U13901 ( .A1(n6655), .A2(n13300), .ZN(n11355) );
  NAND2_X1 U13902 ( .A1(n11356), .A2(n11355), .ZN(n11362) );
  NAND2_X1 U13903 ( .A1(n11361), .A2(n11362), .ZN(n11360) );
  NAND2_X1 U13904 ( .A1(n6655), .A2(n13164), .ZN(n11357) );
  OAI21_X1 U13905 ( .B1(n6655), .B2(n11358), .A(n11357), .ZN(n11359) );
  NAND2_X1 U13906 ( .A1(n11360), .A2(n11359), .ZN(n11366) );
  NAND2_X1 U13907 ( .A1(n11364), .A2(n11363), .ZN(n11365) );
  NAND2_X1 U13908 ( .A1(n11366), .A2(n11365), .ZN(n11374) );
  OR2_X1 U13909 ( .A1(n6655), .A2(n11367), .ZN(n11369) );
  NAND2_X1 U13910 ( .A1(n11370), .A2(n6655), .ZN(n11368) );
  NAND2_X1 U13911 ( .A1(n11369), .A2(n11368), .ZN(n11375) );
  NAND2_X1 U13912 ( .A1(n11374), .A2(n11375), .ZN(n11373) );
  AOI22_X1 U13913 ( .A1(n11716), .A2(n11370), .B1(n13299), .B2(n6655), .ZN(
        n11371) );
  NAND2_X1 U13914 ( .A1(n11373), .A2(n11372), .ZN(n11379) );
  INV_X1 U13915 ( .A(n11374), .ZN(n11377) );
  NAND2_X1 U13916 ( .A1(n11379), .A2(n11378), .ZN(n11386) );
  NAND2_X1 U13917 ( .A1(n14874), .A2(n11692), .ZN(n11382) );
  INV_X1 U13918 ( .A(n11716), .ZN(n11516) );
  NAND2_X1 U13919 ( .A1(n11516), .A2(n13298), .ZN(n11381) );
  NAND2_X1 U13920 ( .A1(n11382), .A2(n11381), .ZN(n11387) );
  NAND2_X1 U13921 ( .A1(n14874), .A2(n11516), .ZN(n11383) );
  OAI21_X1 U13922 ( .B1(n11384), .B2(n6655), .A(n11383), .ZN(n11385) );
  INV_X1 U13923 ( .A(n11387), .ZN(n11388) );
  NAND2_X1 U13924 ( .A1(n11392), .A2(n6655), .ZN(n11391) );
  OR2_X1 U13925 ( .A1(n6655), .A2(n11389), .ZN(n11390) );
  NAND2_X1 U13926 ( .A1(n11391), .A2(n11390), .ZN(n11394) );
  AOI22_X1 U13927 ( .A1(n11392), .A2(n11692), .B1(n13297), .B2(n6655), .ZN(
        n11393) );
  NAND2_X1 U13928 ( .A1(n14887), .A2(n11692), .ZN(n11397) );
  NAND2_X1 U13929 ( .A1(n11693), .A2(n13296), .ZN(n11396) );
  NAND2_X1 U13930 ( .A1(n11397), .A2(n11396), .ZN(n11403) );
  NAND2_X1 U13931 ( .A1(n14887), .A2(n11693), .ZN(n11398) );
  OAI21_X1 U13932 ( .B1(n11399), .B2(n11693), .A(n11398), .ZN(n11400) );
  NAND2_X1 U13933 ( .A1(n11401), .A2(n11400), .ZN(n11407) );
  INV_X1 U13934 ( .A(n11402), .ZN(n11405) );
  INV_X1 U13935 ( .A(n11403), .ZN(n11404) );
  NAND2_X1 U13936 ( .A1(n11405), .A2(n11404), .ZN(n11406) );
  NAND2_X1 U13937 ( .A1(n11411), .A2(n11693), .ZN(n11410) );
  OR2_X1 U13938 ( .A1(n11693), .A2(n11408), .ZN(n11409) );
  NAND2_X1 U13939 ( .A1(n11410), .A2(n11409), .ZN(n11413) );
  AOI22_X1 U13940 ( .A1(n11411), .A2(n11692), .B1(n13295), .B2(n11693), .ZN(
        n11412) );
  NAND2_X1 U13941 ( .A1(n11417), .A2(n11692), .ZN(n11416) );
  NAND2_X1 U13942 ( .A1(n11693), .A2(n13294), .ZN(n11415) );
  NAND2_X1 U13943 ( .A1(n11417), .A2(n6655), .ZN(n11418) );
  OAI21_X1 U13944 ( .B1(n11419), .B2(n6655), .A(n11418), .ZN(n11420) );
  NAND2_X1 U13945 ( .A1(n11424), .A2(n11693), .ZN(n11423) );
  OR2_X1 U13946 ( .A1(n11693), .A2(n11421), .ZN(n11422) );
  NAND2_X1 U13947 ( .A1(n11423), .A2(n11422), .ZN(n11426) );
  AOI22_X1 U13948 ( .A1(n11424), .A2(n11692), .B1(n13293), .B2(n6655), .ZN(
        n11425) );
  AOI21_X1 U13949 ( .B1(n11427), .B2(n11426), .A(n11425), .ZN(n11429) );
  NOR2_X1 U13950 ( .A1(n11427), .A2(n11426), .ZN(n11428) );
  NAND2_X1 U13951 ( .A1(n14918), .A2(n11692), .ZN(n11431) );
  NAND2_X1 U13952 ( .A1(n11693), .A2(n13292), .ZN(n11430) );
  NAND2_X1 U13953 ( .A1(n14918), .A2(n11693), .ZN(n11432) );
  OAI21_X1 U13954 ( .B1(n11433), .B2(n11693), .A(n11432), .ZN(n11434) );
  NAND2_X1 U13955 ( .A1(n14558), .A2(n11693), .ZN(n11437) );
  OR2_X1 U13956 ( .A1(n11693), .A2(n11435), .ZN(n11436) );
  AOI22_X1 U13957 ( .A1(n14558), .A2(n11692), .B1(n13291), .B2(n11693), .ZN(
        n11438) );
  INV_X1 U13958 ( .A(n11438), .ZN(n11439) );
  NAND2_X1 U13959 ( .A1(n11443), .A2(n11692), .ZN(n11442) );
  NAND2_X1 U13960 ( .A1(n11693), .A2(n13290), .ZN(n11441) );
  NAND2_X1 U13961 ( .A1(n11442), .A2(n11441), .ZN(n11447) );
  NAND2_X1 U13962 ( .A1(n11443), .A2(n11693), .ZN(n11444) );
  OAI21_X1 U13963 ( .B1(n11445), .B2(n11693), .A(n11444), .ZN(n11446) );
  INV_X1 U13964 ( .A(n11447), .ZN(n11448) );
  NAND2_X1 U13965 ( .A1(n13643), .A2(n11693), .ZN(n11450) );
  OR2_X1 U13966 ( .A1(n11693), .A2(n11452), .ZN(n11449) );
  NAND2_X1 U13967 ( .A1(n11450), .A2(n11449), .ZN(n11456) );
  NAND2_X1 U13968 ( .A1(n11455), .A2(n11456), .ZN(n11454) );
  NAND2_X1 U13969 ( .A1(n13643), .A2(n11716), .ZN(n11451) );
  OAI21_X1 U13970 ( .B1(n11452), .B2(n11699), .A(n11451), .ZN(n11453) );
  NAND2_X1 U13971 ( .A1(n11454), .A2(n11453), .ZN(n11460) );
  INV_X1 U13972 ( .A(n11455), .ZN(n11458) );
  INV_X1 U13973 ( .A(n11456), .ZN(n11457) );
  NAND2_X1 U13974 ( .A1(n11458), .A2(n11457), .ZN(n11459) );
  NAND2_X1 U13975 ( .A1(n13637), .A2(n11716), .ZN(n11462) );
  NAND2_X1 U13976 ( .A1(n13288), .A2(n11693), .ZN(n11461) );
  AOI22_X1 U13977 ( .A1(n13637), .A2(n11693), .B1(n11716), .B2(n13288), .ZN(
        n11463) );
  AOI22_X1 U13978 ( .A1(n13627), .A2(n11693), .B1(n11716), .B2(n13286), .ZN(
        n11466) );
  NAND2_X1 U13979 ( .A1(n13627), .A2(n11692), .ZN(n11465) );
  NAND2_X1 U13980 ( .A1(n13286), .A2(n6655), .ZN(n11464) );
  NAND2_X1 U13981 ( .A1(n11465), .A2(n11464), .ZN(n11477) );
  NAND2_X1 U13982 ( .A1(n11466), .A2(n11477), .ZN(n11475) );
  NAND2_X1 U13983 ( .A1(n13632), .A2(n11693), .ZN(n11468) );
  NAND2_X1 U13984 ( .A1(n13287), .A2(n11716), .ZN(n11467) );
  NAND2_X1 U13985 ( .A1(n11468), .A2(n11467), .ZN(n11473) );
  INV_X1 U13986 ( .A(n11473), .ZN(n11471) );
  AND2_X1 U13987 ( .A1(n13287), .A2(n11693), .ZN(n11469) );
  AOI21_X1 U13988 ( .B1(n13632), .B2(n11699), .A(n11469), .ZN(n11474) );
  INV_X1 U13989 ( .A(n11474), .ZN(n11470) );
  NAND2_X1 U13990 ( .A1(n11471), .A2(n11470), .ZN(n11472) );
  AND2_X1 U13991 ( .A1(n11475), .A2(n11472), .ZN(n11480) );
  NOR2_X1 U13992 ( .A1(n13627), .A2(n13286), .ZN(n11478) );
  NAND3_X1 U13993 ( .A1(n11475), .A2(n11474), .A3(n11473), .ZN(n11476) );
  OAI21_X1 U13994 ( .B1(n11478), .B2(n11477), .A(n11476), .ZN(n11479) );
  NAND2_X1 U13995 ( .A1(n11481), .A2(n6652), .ZN(n11483) );
  AOI22_X1 U13996 ( .A1(n11683), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n13340), 
        .B2(n11490), .ZN(n11482) );
  NAND2_X2 U13997 ( .A1(n11483), .A2(n11482), .ZN(n13553) );
  AND2_X1 U13998 ( .A1(n13285), .A2(n11716), .ZN(n11484) );
  AOI21_X1 U13999 ( .B1(n13553), .B2(n6655), .A(n11484), .ZN(n11485) );
  NAND2_X1 U14000 ( .A1(n11489), .A2(n6652), .ZN(n11492) );
  AOI22_X1 U14001 ( .A1(n11748), .A2(n11490), .B1(n11683), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n11491) );
  INV_X1 U14002 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n11493) );
  NAND2_X1 U14003 ( .A1(n11494), .A2(n11493), .ZN(n11495) );
  AND2_X1 U14004 ( .A1(n11529), .A2(n11495), .ZN(n13526) );
  NAND2_X1 U14005 ( .A1(n13526), .A2(n11658), .ZN(n11501) );
  INV_X1 U14006 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n11498) );
  NAND2_X1 U14007 ( .A1(n11642), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U14008 ( .A1(n11686), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n11496) );
  OAI211_X1 U14009 ( .C1(n11498), .C2(n11605), .A(n11497), .B(n11496), .ZN(
        n11499) );
  INV_X1 U14010 ( .A(n11499), .ZN(n11500) );
  OAI22_X1 U14011 ( .A1(n13529), .A2(n6655), .B1(n13541), .B2(n11699), .ZN(
        n11504) );
  NAND2_X1 U14012 ( .A1(n11503), .A2(n11504), .ZN(n11508) );
  AOI22_X1 U14013 ( .A1(n13616), .A2(n6655), .B1(n11716), .B2(n13284), .ZN(
        n11502) );
  INV_X1 U14014 ( .A(n11503), .ZN(n11506) );
  INV_X1 U14015 ( .A(n11504), .ZN(n11505) );
  INV_X1 U14016 ( .A(n11519), .ZN(n11522) );
  NAND2_X1 U14017 ( .A1(n11683), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n11509) );
  XNOR2_X1 U14018 ( .A(n11529), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13509) );
  NAND2_X1 U14019 ( .A1(n13509), .A2(n11658), .ZN(n11515) );
  INV_X1 U14020 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n15522) );
  NAND2_X1 U14021 ( .A1(n10957), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n11512) );
  NAND2_X1 U14022 ( .A1(n11642), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n11511) );
  OAI211_X1 U14023 ( .C1(n9466), .C2(n15522), .A(n11512), .B(n11511), .ZN(
        n11513) );
  INV_X1 U14024 ( .A(n11513), .ZN(n11514) );
  NAND2_X1 U14025 ( .A1(n11515), .A2(n11514), .ZN(n13283) );
  AOI22_X1 U14026 ( .A1(n13611), .A2(n11516), .B1(n11716), .B2(n13283), .ZN(
        n11518) );
  INV_X1 U14027 ( .A(n11518), .ZN(n11521) );
  INV_X1 U14028 ( .A(n13611), .ZN(n13512) );
  OAI22_X1 U14029 ( .A1(n13512), .A2(n11693), .B1(n13190), .B2(n11699), .ZN(
        n11517) );
  OR2_X1 U14030 ( .A1(n11523), .A2(n11572), .ZN(n11525) );
  NAND2_X1 U14031 ( .A1(n11683), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14032 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n11526) );
  INV_X1 U14033 ( .A(n11544), .ZN(n11531) );
  INV_X1 U14034 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n11528) );
  INV_X1 U14035 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n11527) );
  OAI21_X1 U14036 ( .B1(n11529), .B2(n11528), .A(n11527), .ZN(n11530) );
  NAND2_X1 U14037 ( .A1(n11531), .A2(n11530), .ZN(n13490) );
  OR2_X1 U14038 ( .A1(n13490), .A2(n11551), .ZN(n11537) );
  INV_X1 U14039 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n11534) );
  NAND2_X1 U14040 ( .A1(n10957), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U14041 ( .A1(n11686), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n11532) );
  OAI211_X1 U14042 ( .C1(n9858), .C2(n11534), .A(n11533), .B(n11532), .ZN(
        n11535) );
  INV_X1 U14043 ( .A(n11535), .ZN(n11536) );
  OAI22_X1 U14044 ( .A1(n13493), .A2(n6655), .B1(n13236), .B2(n11699), .ZN(
        n11539) );
  INV_X1 U14045 ( .A(n11539), .ZN(n11540) );
  AOI22_X1 U14046 ( .A1(n13606), .A2(n6655), .B1(n11716), .B2(n13471), .ZN(
        n11538) );
  NAND2_X1 U14047 ( .A1(n11683), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n11542) );
  NOR2_X1 U14048 ( .A1(n11544), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n11545) );
  OR2_X1 U14049 ( .A1(n11558), .A2(n11545), .ZN(n13477) );
  INV_X1 U14050 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n11548) );
  NAND2_X1 U14051 ( .A1(n11686), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U14052 ( .A1(n11642), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n11546) );
  OAI211_X1 U14053 ( .C1(n11605), .C2(n11548), .A(n11547), .B(n11546), .ZN(
        n11549) );
  INV_X1 U14054 ( .A(n11549), .ZN(n11550) );
  OAI21_X1 U14055 ( .B1(n13477), .B2(n11551), .A(n11550), .ZN(n13282) );
  AOI22_X1 U14056 ( .A1(n13601), .A2(n6655), .B1(n11699), .B2(n13282), .ZN(
        n11552) );
  AOI22_X1 U14057 ( .A1(n13601), .A2(n11699), .B1(n13282), .B2(n6655), .ZN(
        n11554) );
  INV_X1 U14058 ( .A(n11552), .ZN(n11553) );
  NAND2_X1 U14059 ( .A1(n11555), .A2(n6652), .ZN(n11557) );
  NAND2_X1 U14060 ( .A1(n11683), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11556) );
  OR2_X1 U14061 ( .A1(n11558), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n11559) );
  NAND2_X1 U14062 ( .A1(n13461), .A2(n11658), .ZN(n11565) );
  INV_X1 U14063 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n11562) );
  NAND2_X1 U14064 ( .A1(n10957), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U14065 ( .A1(n11686), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n11560) );
  OAI211_X1 U14066 ( .C1(n9858), .C2(n11562), .A(n11561), .B(n11560), .ZN(
        n11563) );
  INV_X1 U14067 ( .A(n11563), .ZN(n11564) );
  OAI22_X1 U14068 ( .A1(n13463), .A2(n11693), .B1(n13237), .B2(n11699), .ZN(
        n11567) );
  OAI22_X1 U14069 ( .A1(n13463), .A2(n11699), .B1(n13237), .B2(n11693), .ZN(
        n11566) );
  INV_X1 U14070 ( .A(n11566), .ZN(n11570) );
  OR2_X1 U14071 ( .A1(n11573), .A2(n11572), .ZN(n11575) );
  NAND2_X1 U14072 ( .A1(n11683), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n11574) );
  NAND2_X1 U14073 ( .A1(n11686), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U14074 ( .A1(n11642), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n11579) );
  INV_X1 U14075 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13216) );
  AOI21_X1 U14076 ( .B1(n13216), .B2(n11576), .A(n11590), .ZN(n13438) );
  NAND2_X1 U14077 ( .A1(n11658), .A2(n13438), .ZN(n11578) );
  INV_X1 U14078 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13440) );
  OR2_X1 U14079 ( .A1(n11605), .A2(n13440), .ZN(n11577) );
  NAND4_X1 U14080 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n13422) );
  AOI22_X1 U14081 ( .A1(n13588), .A2(n6655), .B1(n11699), .B2(n13422), .ZN(
        n11583) );
  INV_X1 U14082 ( .A(n11583), .ZN(n11582) );
  AOI22_X1 U14083 ( .A1(n13588), .A2(n11699), .B1(n13422), .B2(n11693), .ZN(
        n11581) );
  AOI21_X1 U14084 ( .B1(n11584), .B2(n11582), .A(n11581), .ZN(n11586) );
  NAND2_X1 U14085 ( .A1(n11587), .A2(n6652), .ZN(n11589) );
  NAND2_X1 U14086 ( .A1(n11683), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n11588) );
  NAND2_X1 U14087 ( .A1(n9574), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14088 ( .A1(n11590), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n11654) );
  OAI21_X1 U14089 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n11590), .A(n11654), 
        .ZN(n11591) );
  INV_X1 U14090 ( .A(n11591), .ZN(n13414) );
  NAND2_X1 U14091 ( .A1(n11658), .A2(n13414), .ZN(n11596) );
  INV_X1 U14092 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n11592) );
  OR2_X1 U14093 ( .A1(n9466), .A2(n11592), .ZN(n11595) );
  INV_X1 U14094 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n11593) );
  OR2_X1 U14095 ( .A1(n11605), .A2(n11593), .ZN(n11594) );
  OAI22_X1 U14096 ( .A1(n13416), .A2(n6655), .B1(n13267), .B2(n11699), .ZN(
        n11669) );
  NAND2_X1 U14097 ( .A1(n13690), .A2(n6652), .ZN(n11600) );
  NAND2_X1 U14098 ( .A1(n11683), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n11599) );
  NAND2_X1 U14099 ( .A1(n11686), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n11609) );
  NAND2_X1 U14100 ( .A1(n9574), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n11608) );
  INV_X1 U14101 ( .A(n11654), .ZN(n11601) );
  INV_X1 U14102 ( .A(n11628), .ZN(n11630) );
  INV_X1 U14103 ( .A(n11602), .ZN(n11656) );
  INV_X1 U14104 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13150) );
  NAND2_X1 U14105 ( .A1(n11656), .A2(n13150), .ZN(n11603) );
  NAND2_X1 U14106 ( .A1(n11658), .A2(n13391), .ZN(n11607) );
  INV_X1 U14107 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n11604) );
  OR2_X1 U14108 ( .A1(n11605), .A2(n11604), .ZN(n11606) );
  NAND4_X1 U14109 ( .A1(n11609), .A2(n11608), .A3(n11607), .A4(n11606), .ZN(
        n13280) );
  AOI22_X1 U14110 ( .A1(n13573), .A2(n11692), .B1(n13280), .B2(n6655), .ZN(
        n11675) );
  NAND2_X1 U14111 ( .A1(n13573), .A2(n11693), .ZN(n11611) );
  OR2_X1 U14112 ( .A1(n11693), .A2(n13266), .ZN(n11610) );
  NAND2_X1 U14113 ( .A1(n11611), .A2(n11610), .ZN(n11674) );
  XNOR2_X1 U14114 ( .A(n11614), .B(SI_30_), .ZN(n11681) );
  INV_X1 U14115 ( .A(n11614), .ZN(n11615) );
  INV_X1 U14116 ( .A(SI_30_), .ZN(n12464) );
  MUX2_X1 U14117 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6643), .Z(n11616) );
  XNOR2_X1 U14118 ( .A(n11616), .B(SI_31_), .ZN(n11617) );
  XNOR2_X1 U14119 ( .A(n11618), .B(n11617), .ZN(n12194) );
  NAND2_X1 U14120 ( .A1(n12194), .A2(n6652), .ZN(n11621) );
  NAND2_X1 U14121 ( .A1(n11683), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n11620) );
  INV_X1 U14122 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n11624) );
  NAND2_X1 U14123 ( .A1(n10957), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n11623) );
  NAND2_X1 U14124 ( .A1(n11686), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n11622) );
  OAI211_X1 U14125 ( .C1(n9858), .C2(n11624), .A(n11623), .B(n11622), .ZN(
        n13354) );
  NAND2_X1 U14126 ( .A1(n11698), .A2(n13354), .ZN(n11625) );
  NAND2_X1 U14127 ( .A1(n13686), .A2(n6652), .ZN(n11627) );
  NAND2_X1 U14128 ( .A1(n11683), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n11626) );
  NAND2_X1 U14129 ( .A1(n9574), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n11637) );
  INV_X1 U14130 ( .A(n11643), .ZN(n11926) );
  INV_X1 U14131 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11629) );
  NAND2_X1 U14132 ( .A1(n11630), .A2(n11629), .ZN(n11631) );
  NAND2_X1 U14133 ( .A1(n11658), .A2(n12016), .ZN(n11636) );
  INV_X1 U14134 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n11632) );
  OR2_X1 U14135 ( .A1(n9466), .A2(n11632), .ZN(n11635) );
  INV_X1 U14136 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n11633) );
  OR2_X1 U14137 ( .A1(n11605), .A2(n11633), .ZN(n11634) );
  NOR2_X1 U14138 ( .A1(n11693), .A2(n11930), .ZN(n11638) );
  AOI21_X1 U14139 ( .B1(n13567), .B2(n11693), .A(n11638), .ZN(n11679) );
  NAND2_X1 U14140 ( .A1(n13567), .A2(n11716), .ZN(n11640) );
  NAND2_X1 U14141 ( .A1(n6655), .A2(n13279), .ZN(n11639) );
  NAND2_X1 U14142 ( .A1(n11640), .A2(n11639), .ZN(n11678) );
  NAND2_X1 U14143 ( .A1(n11683), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11641) );
  NAND2_X1 U14144 ( .A1(n11686), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14145 ( .A1(n11642), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n11646) );
  NAND2_X1 U14146 ( .A1(n11658), .A2(n11643), .ZN(n11645) );
  INV_X1 U14147 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n11927) );
  OR2_X1 U14148 ( .A1(n11605), .A2(n11927), .ZN(n11644) );
  NAND4_X1 U14149 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n13278) );
  AND2_X1 U14150 ( .A1(n11693), .A2(n13278), .ZN(n11648) );
  AOI21_X1 U14151 ( .B1(n13564), .B2(n11699), .A(n11648), .ZN(n11697) );
  NAND2_X1 U14152 ( .A1(n13564), .A2(n6655), .ZN(n11650) );
  NAND2_X1 U14153 ( .A1(n11699), .A2(n13278), .ZN(n11649) );
  NAND2_X1 U14154 ( .A1(n11650), .A2(n11649), .ZN(n11696) );
  AOI21_X1 U14155 ( .B1(n11675), .B2(n11674), .A(n11676), .ZN(n11673) );
  NAND2_X1 U14156 ( .A1(n11651), .A2(n6652), .ZN(n11653) );
  NAND2_X1 U14157 ( .A1(n11683), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n11652) );
  NAND2_X1 U14158 ( .A1(n11642), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n11663) );
  INV_X1 U14159 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n11655) );
  NAND2_X1 U14160 ( .A1(n11655), .A2(n11654), .ZN(n11657) );
  NAND2_X1 U14161 ( .A1(n11658), .A2(n13405), .ZN(n11662) );
  INV_X1 U14162 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n15350) );
  OR2_X1 U14163 ( .A1(n9466), .A2(n15350), .ZN(n11661) );
  INV_X1 U14164 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n11659) );
  OR2_X1 U14165 ( .A1(n11605), .A2(n11659), .ZN(n11660) );
  NOR2_X1 U14166 ( .A1(n11693), .A2(n11944), .ZN(n11664) );
  AOI21_X1 U14167 ( .B1(n13579), .B2(n11693), .A(n11664), .ZN(n11672) );
  NAND2_X1 U14168 ( .A1(n13579), .A2(n11716), .ZN(n11666) );
  NAND2_X1 U14169 ( .A1(n11693), .A2(n13423), .ZN(n11665) );
  NAND2_X1 U14170 ( .A1(n11666), .A2(n11665), .ZN(n11671) );
  OR2_X1 U14171 ( .A1(n11672), .A2(n11671), .ZN(n11667) );
  AOI22_X1 U14172 ( .A1(n13584), .A2(n11693), .B1(n11699), .B2(n13281), .ZN(
        n11668) );
  AOI21_X1 U14173 ( .B1(n11670), .B2(n11669), .A(n11668), .ZN(n11708) );
  OR3_X1 U14174 ( .A1(n11676), .A2(n11675), .A3(n11674), .ZN(n11705) );
  NAND4_X1 U14175 ( .A1(n11747), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11704) );
  INV_X1 U14176 ( .A(n11681), .ZN(n11682) );
  NAND2_X1 U14177 ( .A1(n12266), .A2(n6652), .ZN(n11685) );
  NAND2_X1 U14178 ( .A1(n11683), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11684) );
  INV_X1 U14179 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13362) );
  NAND2_X1 U14180 ( .A1(n11642), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n11688) );
  NAND2_X1 U14181 ( .A1(n11686), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11687) );
  OAI211_X1 U14182 ( .C1(n11605), .C2(n13362), .A(n11688), .B(n11687), .ZN(
        n13277) );
  NAND2_X1 U14183 ( .A1(n6655), .A2(n13354), .ZN(n11712) );
  OR2_X1 U14184 ( .A1(n11690), .A2(n15591), .ZN(n11754) );
  NAND4_X1 U14185 ( .A1(n11712), .A2(n11757), .A3(n11754), .A4(n11764), .ZN(
        n11691) );
  AOI22_X1 U14186 ( .A1(n13365), .A2(n11692), .B1(n13277), .B2(n11691), .ZN(
        n11711) );
  NAND2_X1 U14187 ( .A1(n13365), .A2(n11693), .ZN(n11695) );
  NAND2_X1 U14188 ( .A1(n11699), .A2(n13277), .ZN(n11694) );
  NAND2_X1 U14189 ( .A1(n11695), .A2(n11694), .ZN(n11710) );
  OAI22_X1 U14190 ( .A1(n11711), .A2(n11710), .B1(n11697), .B2(n11696), .ZN(
        n11702) );
  NAND2_X1 U14191 ( .A1(n11699), .A2(n13354), .ZN(n11700) );
  OAI211_X1 U14192 ( .C1(n13558), .C2(n11699), .A(n11700), .B(n11713), .ZN(
        n11701) );
  NAND2_X1 U14193 ( .A1(n11702), .A2(n11701), .ZN(n11703) );
  NAND3_X1 U14194 ( .A1(n11705), .A2(n11704), .A3(n11703), .ZN(n11706) );
  NOR2_X1 U14195 ( .A1(n7572), .A2(n11706), .ZN(n11707) );
  OAI21_X1 U14196 ( .B1(n11709), .B2(n11708), .A(n11707), .ZN(n11719) );
  NAND2_X1 U14197 ( .A1(n11711), .A2(n11710), .ZN(n11718) );
  INV_X1 U14198 ( .A(n11712), .ZN(n11715) );
  INV_X1 U14199 ( .A(n11713), .ZN(n11714) );
  AOI211_X1 U14200 ( .C1(n11716), .C2(n11698), .A(n11715), .B(n11714), .ZN(
        n11717) );
  NAND2_X1 U14201 ( .A1(n13567), .A2(n13279), .ZN(n11922) );
  OR2_X1 U14202 ( .A1(n13567), .A2(n13279), .ZN(n11720) );
  XNOR2_X1 U14203 ( .A(n13573), .B(n13266), .ZN(n13387) );
  XNOR2_X1 U14204 ( .A(n13579), .B(n11944), .ZN(n13401) );
  XNOR2_X1 U14205 ( .A(n13584), .B(n13281), .ZN(n13417) );
  XNOR2_X1 U14206 ( .A(n13601), .B(n13451), .ZN(n13467) );
  NOR2_X1 U14207 ( .A1(n13606), .A2(n13471), .ZN(n11913) );
  AND2_X1 U14208 ( .A1(n13606), .A2(n13471), .ZN(n11912) );
  NOR2_X1 U14209 ( .A1(n11913), .A2(n11912), .ZN(n13494) );
  XNOR2_X1 U14210 ( .A(n13611), .B(n13190), .ZN(n13505) );
  XNOR2_X1 U14211 ( .A(n13616), .B(n13284), .ZN(n13517) );
  OAI21_X1 U14212 ( .B1(n13302), .B2(n13654), .A(n11721), .ZN(n15595) );
  NAND4_X1 U14213 ( .A1(n11722), .A2(n15591), .A3(n15595), .A4(n9570), .ZN(
        n11724) );
  NOR4_X1 U14214 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11729) );
  NAND4_X1 U14215 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11731) );
  NOR4_X1 U14216 ( .A1(n14559), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n11736) );
  NAND4_X1 U14217 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11739) );
  NOR3_X1 U14218 ( .A1(n11905), .A2(n11739), .A3(n11738), .ZN(n11741) );
  XNOR2_X1 U14219 ( .A(n13553), .B(n13285), .ZN(n13536) );
  NAND4_X1 U14220 ( .A1(n13517), .A2(n11741), .A3(n13536), .A4(n11740), .ZN(
        n11742) );
  NOR4_X1 U14221 ( .A1(n13467), .A2(n13494), .A3(n13505), .A4(n11742), .ZN(
        n11743) );
  XNOR2_X1 U14222 ( .A(n13596), .B(n13469), .ZN(n13453) );
  XNOR2_X1 U14223 ( .A(n13588), .B(n13422), .ZN(n11917) );
  NAND4_X1 U14224 ( .A1(n13417), .A2(n11743), .A3(n13453), .A4(n11917), .ZN(
        n11744) );
  NOR4_X1 U14225 ( .A1(n13372), .A2(n13387), .A3(n13401), .A4(n11744), .ZN(
        n11746) );
  XNOR2_X1 U14226 ( .A(n13365), .B(n13277), .ZN(n11745) );
  XNOR2_X1 U14227 ( .A(n13564), .B(n13278), .ZN(n11950) );
  NAND4_X1 U14228 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11950), .ZN(
        n11749) );
  XNOR2_X1 U14229 ( .A(n11749), .B(n11748), .ZN(n11751) );
  NAND2_X1 U14230 ( .A1(n11751), .A2(n11750), .ZN(n11755) );
  NAND2_X1 U14231 ( .A1(n11761), .A2(n11753), .ZN(n11763) );
  OAI211_X1 U14232 ( .C1(n13349), .C2(n11756), .A(n11755), .B(n11754), .ZN(
        n11762) );
  NAND2_X1 U14233 ( .A1(n13349), .A2(n11757), .ZN(n11758) );
  OAI211_X1 U14234 ( .C1(n11759), .C2(n9581), .A(n11764), .B(n11758), .ZN(
        n11760) );
  AOI22_X1 U14235 ( .A1(n11763), .A2(n11762), .B1(n11761), .B2(n11760), .ZN(
        n11771) );
  INV_X1 U14236 ( .A(n11764), .ZN(n11765) );
  NAND4_X1 U14237 ( .A1(n11767), .A2(n11766), .A3(n11765), .A4(n13470), .ZN(
        n11768) );
  OAI211_X1 U14238 ( .C1(n9581), .C2(n11770), .A(n11768), .B(P2_B_REG_SCAN_IN), 
        .ZN(n11769) );
  OAI21_X1 U14239 ( .B1(n11771), .B2(n11770), .A(n11769), .ZN(P2_U3328) );
  NAND2_X1 U14240 ( .A1(n14584), .A2(n12326), .ZN(n11773) );
  NAND2_X1 U14241 ( .A1(n13827), .A2(n12323), .ZN(n11772) );
  NAND2_X1 U14242 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  XNOR2_X1 U14243 ( .A(n11774), .B(n12324), .ZN(n11781) );
  INV_X1 U14244 ( .A(n11781), .ZN(n11783) );
  AOI22_X1 U14245 ( .A1(n14584), .A2(n12323), .B1(n12322), .B2(n13827), .ZN(
        n11782) );
  INV_X1 U14246 ( .A(n11776), .ZN(n11777) );
  XOR2_X1 U14247 ( .A(n11782), .B(n11781), .Z(n14582) );
  NAND2_X1 U14248 ( .A1(n13815), .A2(n12326), .ZN(n11785) );
  NAND2_X1 U14249 ( .A1(n13826), .A2(n12323), .ZN(n11784) );
  NAND2_X1 U14250 ( .A1(n11785), .A2(n11784), .ZN(n11786) );
  XNOR2_X1 U14251 ( .A(n11786), .B(n12324), .ZN(n11787) );
  AOI22_X1 U14252 ( .A1(n13815), .A2(n12323), .B1(n12322), .B2(n13826), .ZN(
        n13811) );
  AND2_X1 U14253 ( .A1(n11788), .A2(n11787), .ZN(n11789) );
  AOI22_X1 U14254 ( .A1(n14276), .A2(n12323), .B1(n12322), .B2(n13825), .ZN(
        n11792) );
  AOI22_X1 U14255 ( .A1(n14276), .A2(n12326), .B1(n12323), .B2(n13825), .ZN(
        n11790) );
  XNOR2_X1 U14256 ( .A(n11790), .B(n12324), .ZN(n11791) );
  XOR2_X1 U14257 ( .A(n11792), .B(n11791), .Z(n13742) );
  NAND2_X1 U14258 ( .A1(n13761), .A2(n12326), .ZN(n11795) );
  NAND2_X1 U14259 ( .A1(n13824), .A2(n12323), .ZN(n11794) );
  NAND2_X1 U14260 ( .A1(n11795), .A2(n11794), .ZN(n11796) );
  XNOR2_X1 U14261 ( .A(n11796), .B(n12324), .ZN(n11799) );
  NAND2_X1 U14262 ( .A1(n13761), .A2(n12323), .ZN(n11798) );
  NAND2_X1 U14263 ( .A1(n13824), .A2(n12322), .ZN(n11797) );
  NAND2_X1 U14264 ( .A1(n11798), .A2(n11797), .ZN(n11800) );
  NAND2_X1 U14265 ( .A1(n11799), .A2(n11800), .ZN(n13752) );
  INV_X1 U14266 ( .A(n11799), .ZN(n11802) );
  INV_X1 U14267 ( .A(n11800), .ZN(n11801) );
  NAND2_X1 U14268 ( .A1(n11802), .A2(n11801), .ZN(n13753) );
  NAND2_X1 U14269 ( .A1(n11803), .A2(n13753), .ZN(n13782) );
  NAND2_X1 U14270 ( .A1(n11807), .A2(n12326), .ZN(n11805) );
  NAND2_X1 U14271 ( .A1(n13823), .A2(n12323), .ZN(n11804) );
  NAND2_X1 U14272 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  XNOR2_X1 U14273 ( .A(n11806), .B(n12324), .ZN(n11813) );
  AOI22_X1 U14274 ( .A1(n11807), .A2(n12323), .B1(n12322), .B2(n13823), .ZN(
        n11814) );
  XNOR2_X1 U14275 ( .A(n11813), .B(n11814), .ZN(n13783) );
  NAND2_X1 U14276 ( .A1(n14185), .A2(n12326), .ZN(n11809) );
  NAND2_X1 U14277 ( .A1(n13822), .A2(n12323), .ZN(n11808) );
  NAND2_X1 U14278 ( .A1(n11809), .A2(n11808), .ZN(n11810) );
  XNOR2_X1 U14279 ( .A(n11810), .B(n12324), .ZN(n11819) );
  AND2_X1 U14280 ( .A1(n13822), .A2(n12322), .ZN(n11812) );
  AOI21_X1 U14281 ( .B1(n14185), .B2(n6648), .A(n11812), .ZN(n11817) );
  XNOR2_X1 U14282 ( .A(n11819), .B(n11817), .ZN(n13717) );
  INV_X1 U14283 ( .A(n11813), .ZN(n11815) );
  NAND2_X1 U14284 ( .A1(n11815), .A2(n11814), .ZN(n13715) );
  INV_X1 U14285 ( .A(n11817), .ZN(n11818) );
  NAND2_X1 U14286 ( .A1(n11819), .A2(n11818), .ZN(n11820) );
  AND2_X1 U14287 ( .A1(n13821), .A2(n12322), .ZN(n11821) );
  AOI21_X1 U14288 ( .B1(n14248), .B2(n12323), .A(n11821), .ZN(n11824) );
  AOI22_X1 U14289 ( .A1(n14248), .A2(n12326), .B1(n12323), .B2(n13821), .ZN(
        n11822) );
  XNOR2_X1 U14290 ( .A(n11822), .B(n12324), .ZN(n11823) );
  XOR2_X1 U14291 ( .A(n11824), .B(n11823), .Z(n13775) );
  INV_X1 U14292 ( .A(n11823), .ZN(n11826) );
  INV_X1 U14293 ( .A(n11824), .ZN(n11825) );
  NAND2_X1 U14294 ( .A1(n11826), .A2(n11825), .ZN(n11827) );
  NAND2_X1 U14295 ( .A1(n14303), .A2(n12326), .ZN(n11829) );
  NAND2_X1 U14296 ( .A1(n13820), .A2(n6648), .ZN(n11828) );
  NAND2_X1 U14297 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  XNOR2_X1 U14298 ( .A(n11830), .B(n12295), .ZN(n11833) );
  AND2_X1 U14299 ( .A1(n13820), .A2(n12322), .ZN(n11831) );
  AOI21_X1 U14300 ( .B1(n14303), .B2(n12323), .A(n11831), .ZN(n11832) );
  NAND2_X1 U14301 ( .A1(n11833), .A2(n11832), .ZN(n11846) );
  OAI21_X1 U14302 ( .B1(n11833), .B2(n11832), .A(n11846), .ZN(n13723) );
  INV_X1 U14303 ( .A(n11846), .ZN(n11844) );
  OAI22_X1 U14304 ( .A1(n14234), .A2(n11834), .B1(n13724), .B2(n11836), .ZN(
        n11835) );
  XNOR2_X1 U14305 ( .A(n11835), .B(n12295), .ZN(n11839) );
  OR2_X1 U14306 ( .A1(n14234), .A2(n11836), .ZN(n11838) );
  NAND2_X1 U14307 ( .A1(n13819), .A2(n12322), .ZN(n11837) );
  AND2_X1 U14308 ( .A1(n11838), .A2(n11837), .ZN(n11840) );
  NAND2_X1 U14309 ( .A1(n11839), .A2(n11840), .ZN(n13702) );
  INV_X1 U14310 ( .A(n11839), .ZN(n11842) );
  INV_X1 U14311 ( .A(n11840), .ZN(n11841) );
  NAND2_X1 U14312 ( .A1(n11842), .A2(n11841), .ZN(n11843) );
  NOR3_X1 U14313 ( .A1(n7573), .A2(n11844), .A3(n11845), .ZN(n11849) );
  INV_X1 U14314 ( .A(n11845), .ZN(n11847) );
  OR2_X1 U14315 ( .A1(n13723), .A2(n11847), .ZN(n12278) );
  OR2_X1 U14316 ( .A1(n12268), .A2(n12278), .ZN(n11848) );
  OR2_X1 U14317 ( .A1(n11847), .A2(n11846), .ZN(n12279) );
  NAND2_X1 U14318 ( .A1(n11848), .A2(n12279), .ZN(n13705) );
  OAI21_X1 U14319 ( .B1(n11849), .B2(n13705), .A(n14585), .ZN(n11854) );
  INV_X1 U14320 ( .A(n11850), .ZN(n14128) );
  AOI22_X1 U14321 ( .A1(n13820), .A2(n14082), .B1(n14079), .B2(n14081), .ZN(
        n14232) );
  INV_X1 U14322 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n11851) );
  OAI22_X1 U14323 ( .A1(n14232), .A2(n13808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11851), .ZN(n11852) );
  AOI21_X1 U14324 ( .B1(n14128), .B2(n13806), .A(n11852), .ZN(n11853) );
  OAI211_X1 U14325 ( .C1(n13792), .C2(n14234), .A(n11854), .B(n11853), .ZN(
        P1_U3235) );
  NAND2_X1 U14326 ( .A1(n11857), .A2(n12991), .ZN(n11855) );
  NAND2_X1 U14327 ( .A1(n11856), .A2(n11855), .ZN(n11861) );
  INV_X1 U14328 ( .A(n11857), .ZN(n11859) );
  NAND2_X1 U14329 ( .A1(n11859), .A2(n11858), .ZN(n11860) );
  XNOR2_X1 U14330 ( .A(n12399), .B(n11895), .ZN(n11863) );
  XNOR2_X1 U14331 ( .A(n11863), .B(n12405), .ZN(n12396) );
  INV_X1 U14332 ( .A(n11863), .ZN(n11864) );
  NAND2_X1 U14333 ( .A1(n11864), .A2(n12946), .ZN(n11865) );
  XNOR2_X1 U14334 ( .A(n13052), .B(n11895), .ZN(n11866) );
  XNOR2_X1 U14335 ( .A(n11866), .B(n12707), .ZN(n12402) );
  NAND2_X1 U14336 ( .A1(n12403), .A2(n12402), .ZN(n12401) );
  INV_X1 U14337 ( .A(n11866), .ZN(n11867) );
  NAND2_X1 U14338 ( .A1(n11867), .A2(n12707), .ZN(n11868) );
  NAND2_X1 U14339 ( .A1(n12401), .A2(n11868), .ZN(n12439) );
  XNOR2_X1 U14340 ( .A(n11869), .B(n11886), .ZN(n11870) );
  XNOR2_X1 U14341 ( .A(n11870), .B(n12918), .ZN(n12438) );
  NAND2_X1 U14342 ( .A1(n12439), .A2(n12438), .ZN(n12437) );
  INV_X1 U14343 ( .A(n12918), .ZN(n12947) );
  NAND2_X1 U14344 ( .A1(n11870), .A2(n12947), .ZN(n11871) );
  NAND2_X1 U14345 ( .A1(n12437), .A2(n11871), .ZN(n12367) );
  XNOR2_X1 U14346 ( .A(n13112), .B(n11895), .ZN(n11872) );
  XNOR2_X1 U14347 ( .A(n11872), .B(n12931), .ZN(n12366) );
  NAND2_X1 U14348 ( .A1(n12367), .A2(n12366), .ZN(n12365) );
  NAND2_X1 U14349 ( .A1(n11872), .A2(n12899), .ZN(n11873) );
  NAND2_X1 U14350 ( .A1(n12365), .A2(n11873), .ZN(n12425) );
  XNOR2_X1 U14351 ( .A(n12905), .B(n11895), .ZN(n11874) );
  XNOR2_X1 U14352 ( .A(n11874), .B(n12706), .ZN(n12424) );
  INV_X1 U14353 ( .A(n11874), .ZN(n11875) );
  NAND2_X1 U14354 ( .A1(n11875), .A2(n12706), .ZN(n11876) );
  XNOR2_X1 U14355 ( .A(n11877), .B(n11895), .ZN(n11879) );
  XNOR2_X1 U14356 ( .A(n11879), .B(n11878), .ZN(n12376) );
  XNOR2_X1 U14357 ( .A(n11880), .B(n11886), .ZN(n11881) );
  INV_X1 U14358 ( .A(n11881), .ZN(n11882) );
  AND2_X1 U14359 ( .A1(n11883), .A2(n11882), .ZN(n11884) );
  XNOR2_X1 U14360 ( .A(n13021), .B(n11895), .ZN(n12413) );
  XNOR2_X1 U14361 ( .A(n12651), .B(n11886), .ZN(n12409) );
  INV_X1 U14362 ( .A(n12409), .ZN(n11887) );
  OAI22_X1 U14363 ( .A1(n12413), .A2(n12412), .B1(n12650), .B2(n11887), .ZN(
        n11891) );
  OAI21_X1 U14364 ( .B1(n12409), .B2(n12704), .A(n12703), .ZN(n11889) );
  NOR2_X1 U14365 ( .A1(n12704), .A2(n12703), .ZN(n11888) );
  AOI22_X1 U14366 ( .A1(n12413), .A2(n11889), .B1(n11888), .B2(n11887), .ZN(
        n11890) );
  XNOR2_X1 U14367 ( .A(n13091), .B(n11895), .ZN(n11892) );
  XNOR2_X1 U14368 ( .A(n11892), .B(n12656), .ZN(n12383) );
  INV_X1 U14369 ( .A(n11892), .ZN(n11893) );
  XNOR2_X1 U14370 ( .A(n13087), .B(n11895), .ZN(n11894) );
  XNOR2_X1 U14371 ( .A(n11894), .B(n12702), .ZN(n12448) );
  XNOR2_X1 U14372 ( .A(n12822), .B(n11895), .ZN(n11896) );
  XNOR2_X1 U14373 ( .A(n11896), .B(n12701), .ZN(n12352) );
  XNOR2_X1 U14374 ( .A(n12800), .B(n11895), .ZN(n11897) );
  XNOR2_X1 U14375 ( .A(n11898), .B(n11897), .ZN(n11904) );
  AOI22_X1 U14376 ( .A1(n12701), .A2(n11899), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11900) );
  OAI21_X1 U14377 ( .B1(n12803), .B2(n12368), .A(n11900), .ZN(n11902) );
  NOR2_X1 U14378 ( .A1(n13080), .A2(n12446), .ZN(n11901) );
  AOI211_X1 U14379 ( .C1(n12807), .C2(n12451), .A(n11902), .B(n11901), .ZN(
        n11903) );
  OAI21_X1 U14380 ( .B1(n11904), .B2(n12459), .A(n11903), .ZN(P3_U3160) );
  NAND2_X1 U14381 ( .A1(n11906), .A2(n11905), .ZN(n11908) );
  NAND2_X1 U14382 ( .A1(n13627), .A2(n13286), .ZN(n11907) );
  OR2_X1 U14383 ( .A1(n13553), .A2(n13285), .ZN(n11909) );
  OR2_X1 U14384 ( .A1(n13529), .A2(n13541), .ZN(n11910) );
  NAND2_X1 U14385 ( .A1(n13611), .A2(n13283), .ZN(n11911) );
  INV_X1 U14386 ( .A(n11913), .ZN(n11914) );
  INV_X1 U14387 ( .A(n13467), .ZN(n13473) );
  NAND2_X1 U14388 ( .A1(n13463), .A2(n13237), .ZN(n11915) );
  NAND2_X1 U14389 ( .A1(n13588), .A2(n13422), .ZN(n11918) );
  NAND2_X1 U14390 ( .A1(n13416), .A2(n13267), .ZN(n11919) );
  NAND2_X1 U14391 ( .A1(n13579), .A2(n13423), .ZN(n11921) );
  NOR2_X1 U14392 ( .A1(n13579), .A2(n13423), .ZN(n11920) );
  NAND2_X1 U14393 ( .A1(n13388), .A2(n13387), .ZN(n13571) );
  OAI21_X1 U14394 ( .B1(n13390), .B2(n13266), .A(n13571), .ZN(n13373) );
  NAND2_X1 U14395 ( .A1(n13373), .A2(n13372), .ZN(n13371) );
  INV_X1 U14396 ( .A(n13553), .ZN(n13623) );
  AND2_X1 U14397 ( .A1(n13508), .A2(n13493), .ZN(n13488) );
  NAND2_X1 U14398 ( .A1(n13390), .A2(n13404), .ZN(n13389) );
  AOI21_X1 U14399 ( .B1(n13564), .B2(n13377), .A(n13459), .ZN(n11925) );
  OAI22_X1 U14400 ( .A1(n13441), .A2(n11927), .B1(n11926), .B2(n15592), .ZN(
        n11929) );
  NOR2_X1 U14401 ( .A1(n7057), .A2(n13528), .ZN(n11928) );
  AOI211_X1 U14402 ( .C1(n15590), .C2(n13563), .A(n11929), .B(n11928), .ZN(
        n11957) );
  NOR2_X1 U14403 ( .A1(n13567), .A2(n11930), .ZN(n11931) );
  XNOR2_X1 U14404 ( .A(n11950), .B(n11931), .ZN(n11955) );
  NOR2_X1 U14405 ( .A1(n13627), .A2(n13539), .ZN(n11933) );
  NAND2_X1 U14406 ( .A1(n13627), .A2(n13539), .ZN(n11932) );
  AND2_X1 U14407 ( .A1(n13553), .A2(n13174), .ZN(n11935) );
  OR2_X1 U14408 ( .A1(n13553), .A2(n13174), .ZN(n11936) );
  NAND2_X1 U14409 ( .A1(n13501), .A2(n13500), .ZN(n11938) );
  NAND2_X1 U14410 ( .A1(n13611), .A2(n13190), .ZN(n11937) );
  NOR2_X1 U14411 ( .A1(n13493), .A2(n13471), .ZN(n11940) );
  NAND2_X1 U14412 ( .A1(n13493), .A2(n13471), .ZN(n11939) );
  NAND2_X1 U14413 ( .A1(n13449), .A2(n13453), .ZN(n11942) );
  NAND2_X1 U14414 ( .A1(n13463), .A2(n13469), .ZN(n11941) );
  INV_X1 U14415 ( .A(n13422), .ZN(n13450) );
  NAND2_X1 U14416 ( .A1(n13588), .A2(n13450), .ZN(n13418) );
  OR2_X1 U14417 ( .A1(n13416), .A2(n13281), .ZN(n11943) );
  NAND2_X1 U14418 ( .A1(n13421), .A2(n11943), .ZN(n13397) );
  NAND2_X1 U14419 ( .A1(n7065), .A2(n13423), .ZN(n11946) );
  AND2_X1 U14420 ( .A1(n13579), .A2(n11944), .ZN(n11945) );
  NAND2_X1 U14421 ( .A1(n13573), .A2(n13266), .ZN(n11947) );
  NOR2_X1 U14422 ( .A1(n13691), .A2(n11948), .ZN(n11949) );
  NOR2_X1 U14423 ( .A1(n13540), .A2(n11949), .ZN(n13355) );
  AOI22_X1 U14424 ( .A1(n13470), .A2(n13279), .B1(n13355), .B2(n13277), .ZN(
        n11954) );
  INV_X1 U14425 ( .A(n13372), .ZN(n11952) );
  NAND4_X1 U14426 ( .A1(n11923), .A2(n13367), .A3(n13521), .A4(n11952), .ZN(
        n11953) );
  NAND2_X1 U14427 ( .A1(n13562), .A2(n13441), .ZN(n11956) );
  OAI211_X1 U14428 ( .C1(n13565), .C2(n13496), .A(n11957), .B(n11956), .ZN(
        P2_U3236) );
  OAI21_X1 U14429 ( .B1(n11960), .B2(n11959), .A(n11958), .ZN(n11961) );
  NAND2_X1 U14430 ( .A1(n11961), .A2(n14585), .ZN(n11966) );
  OAI22_X1 U14431 ( .A1(n11962), .A2(n14594), .B1(n14593), .B2(n6649), .ZN(
        n11963) );
  AOI21_X1 U14432 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n11964), .A(n11963), .ZN(
        n11965) );
  OAI211_X1 U14433 ( .C1(n14714), .C2(n13792), .A(n11966), .B(n11965), .ZN(
        P1_U3237) );
  OAI222_X1 U14434 ( .A1(P1_U3086), .A2(n11968), .B1(n14330), .B2(n11967), 
        .C1(n15349), .C2(n14332), .ZN(P1_U3329) );
  INV_X1 U14435 ( .A(n11969), .ZN(n11970) );
  AND2_X1 U14436 ( .A1(n13286), .A2(n13459), .ZN(n11973) );
  XNOR2_X1 U14437 ( .A(n13627), .B(n12012), .ZN(n11972) );
  NOR2_X1 U14438 ( .A1(n11972), .A2(n11973), .ZN(n11974) );
  AOI21_X1 U14439 ( .B1(n11973), .B2(n11972), .A(n11974), .ZN(n13202) );
  XNOR2_X1 U14440 ( .A(n13553), .B(n12012), .ZN(n11976) );
  NAND2_X1 U14441 ( .A1(n13285), .A2(n13459), .ZN(n11975) );
  XNOR2_X1 U14442 ( .A(n11976), .B(n11975), .ZN(n13255) );
  INV_X1 U14443 ( .A(n11975), .ZN(n11977) );
  NOR2_X1 U14444 ( .A1(n13541), .A2(n10936), .ZN(n11979) );
  XNOR2_X1 U14445 ( .A(n13529), .B(n11995), .ZN(n11978) );
  NOR2_X1 U14446 ( .A1(n11978), .A2(n11979), .ZN(n11980) );
  AOI21_X1 U14447 ( .B1(n11979), .B2(n11978), .A(n11980), .ZN(n13171) );
  INV_X1 U14448 ( .A(n11980), .ZN(n11981) );
  NAND2_X1 U14449 ( .A1(n13170), .A2(n11981), .ZN(n13227) );
  XNOR2_X1 U14450 ( .A(n13611), .B(n12012), .ZN(n11983) );
  AND2_X1 U14451 ( .A1(n13283), .A2(n13459), .ZN(n11982) );
  NOR2_X1 U14452 ( .A1(n11983), .A2(n11982), .ZN(n13223) );
  NAND2_X1 U14453 ( .A1(n11983), .A2(n11982), .ZN(n13224) );
  XNOR2_X1 U14454 ( .A(n13606), .B(n12012), .ZN(n11984) );
  NAND2_X1 U14455 ( .A1(n13471), .A2(n13459), .ZN(n11985) );
  XNOR2_X1 U14456 ( .A(n11984), .B(n11985), .ZN(n13188) );
  NAND2_X1 U14457 ( .A1(n13189), .A2(n13188), .ZN(n13187) );
  INV_X1 U14458 ( .A(n11985), .ZN(n11986) );
  NAND2_X1 U14459 ( .A1(n11984), .A2(n11986), .ZN(n11987) );
  NAND2_X1 U14460 ( .A1(n13187), .A2(n11987), .ZN(n11988) );
  XNOR2_X1 U14461 ( .A(n13601), .B(n11995), .ZN(n11989) );
  XNOR2_X1 U14462 ( .A(n11988), .B(n11989), .ZN(n13233) );
  NOR2_X1 U14463 ( .A1(n13451), .A2(n10936), .ZN(n13235) );
  NAND2_X1 U14464 ( .A1(n13233), .A2(n13235), .ZN(n13234) );
  INV_X1 U14465 ( .A(n11988), .ZN(n11990) );
  NAND2_X1 U14466 ( .A1(n13234), .A2(n7562), .ZN(n11993) );
  XNOR2_X1 U14467 ( .A(n13463), .B(n12012), .ZN(n11991) );
  XNOR2_X1 U14468 ( .A(n11993), .B(n11991), .ZN(n13154) );
  NOR2_X1 U14469 ( .A1(n13237), .A2(n10936), .ZN(n13156) );
  NAND2_X1 U14470 ( .A1(n13154), .A2(n13156), .ZN(n13155) );
  INV_X1 U14471 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U14472 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  NAND2_X1 U14473 ( .A1(n13155), .A2(n11994), .ZN(n13212) );
  XNOR2_X1 U14474 ( .A(n13588), .B(n11995), .ZN(n11997) );
  NAND2_X1 U14475 ( .A1(n13422), .A2(n13459), .ZN(n11996) );
  NOR2_X1 U14476 ( .A1(n11997), .A2(n11996), .ZN(n11998) );
  AOI21_X1 U14477 ( .B1(n11997), .B2(n11996), .A(n11998), .ZN(n13214) );
  NAND2_X1 U14478 ( .A1(n13212), .A2(n13214), .ZN(n13213) );
  INV_X1 U14479 ( .A(n11998), .ZN(n11999) );
  NAND2_X1 U14480 ( .A1(n13213), .A2(n11999), .ZN(n13195) );
  XNOR2_X1 U14481 ( .A(n13416), .B(n12012), .ZN(n12001) );
  OR2_X1 U14482 ( .A1(n13267), .A2(n10936), .ZN(n12000) );
  NOR2_X1 U14483 ( .A1(n12001), .A2(n12000), .ZN(n12002) );
  AOI21_X1 U14484 ( .B1(n12001), .B2(n12000), .A(n12002), .ZN(n13197) );
  NAND2_X1 U14485 ( .A1(n13195), .A2(n13197), .ZN(n13196) );
  INV_X1 U14486 ( .A(n12002), .ZN(n12003) );
  XNOR2_X1 U14487 ( .A(n13579), .B(n12012), .ZN(n12004) );
  NAND2_X1 U14488 ( .A1(n13423), .A2(n13459), .ZN(n12005) );
  XOR2_X1 U14489 ( .A(n12004), .B(n12005), .Z(n13265) );
  INV_X1 U14490 ( .A(n12004), .ZN(n12006) );
  NAND2_X1 U14491 ( .A1(n12006), .A2(n12005), .ZN(n12007) );
  XNOR2_X1 U14492 ( .A(n13573), .B(n12012), .ZN(n12009) );
  AND2_X1 U14493 ( .A1(n13280), .A2(n13459), .ZN(n12008) );
  NAND2_X1 U14494 ( .A1(n12009), .A2(n12008), .ZN(n12010) );
  OAI21_X1 U14495 ( .B1(n12009), .B2(n12008), .A(n12010), .ZN(n13146) );
  NAND2_X1 U14496 ( .A1(n13148), .A2(n12010), .ZN(n12015) );
  NAND2_X1 U14497 ( .A1(n13279), .A2(n13459), .ZN(n12011) );
  XNOR2_X1 U14498 ( .A(n12012), .B(n12011), .ZN(n12013) );
  XNOR2_X1 U14499 ( .A(n13567), .B(n12013), .ZN(n12014) );
  XNOR2_X1 U14500 ( .A(n12015), .B(n12014), .ZN(n12021) );
  INV_X1 U14501 ( .A(n12016), .ZN(n13375) );
  INV_X1 U14502 ( .A(n13278), .ZN(n12017) );
  OAI22_X1 U14503 ( .A1(n13266), .A2(n13538), .B1(n12017), .B2(n13540), .ZN(
        n13369) );
  AOI22_X1 U14504 ( .A1(n13268), .A2(n13369), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12018) );
  OAI21_X1 U14505 ( .B1(n13375), .B2(n13270), .A(n12018), .ZN(n12019) );
  AOI21_X1 U14506 ( .B1(n13567), .B2(n13273), .A(n12019), .ZN(n12020) );
  OAI21_X1 U14507 ( .B1(n12021), .B2(n13275), .A(n12020), .ZN(P2_U3192) );
  NAND2_X1 U14508 ( .A1(n12023), .A2(n14114), .ZN(n12024) );
  NAND2_X1 U14509 ( .A1(n14114), .A2(n12025), .ZN(n12026) );
  NAND3_X1 U14510 ( .A1(n12027), .A2(n12205), .A3(n12026), .ZN(n12028) );
  MUX2_X1 U14511 ( .A(n14081), .B(n14110), .S(n12152), .Z(n12148) );
  NAND2_X1 U14512 ( .A1(n12032), .A2(n12029), .ZN(n12031) );
  INV_X1 U14513 ( .A(n12032), .ZN(n12033) );
  AND2_X1 U14514 ( .A1(n9350), .A2(n12152), .ZN(n12036) );
  NOR2_X1 U14515 ( .A1(n9350), .A2(n12152), .ZN(n12035) );
  MUX2_X1 U14516 ( .A(n12039), .B(n12038), .S(n12066), .Z(n12040) );
  MUX2_X1 U14517 ( .A(n12042), .B(n12041), .S(n12066), .Z(n12043) );
  NAND2_X1 U14518 ( .A1(n12044), .A2(n12043), .ZN(n12049) );
  INV_X1 U14519 ( .A(n14722), .ZN(n12045) );
  MUX2_X1 U14520 ( .A(n12046), .B(n12045), .S(n12066), .Z(n12048) );
  MUX2_X1 U14521 ( .A(n14722), .B(n13837), .S(n12066), .Z(n12047) );
  OAI21_X1 U14522 ( .B1(n12049), .B2(n12048), .A(n12047), .ZN(n12051) );
  NAND2_X1 U14523 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  MUX2_X1 U14524 ( .A(n12052), .B(n13836), .S(n12066), .Z(n12054) );
  MUX2_X1 U14525 ( .A(n12052), .B(n13836), .S(n12152), .Z(n12053) );
  INV_X1 U14526 ( .A(n12054), .ZN(n12055) );
  MUX2_X1 U14527 ( .A(n13835), .B(n12056), .S(n12066), .Z(n12060) );
  NAND2_X1 U14528 ( .A1(n12059), .A2(n12060), .ZN(n12058) );
  MUX2_X1 U14529 ( .A(n12056), .B(n13835), .S(n12066), .Z(n12057) );
  INV_X1 U14530 ( .A(n12059), .ZN(n12062) );
  INV_X1 U14531 ( .A(n12060), .ZN(n12061) );
  MUX2_X1 U14532 ( .A(n13834), .B(n12064), .S(n12152), .Z(n12063) );
  MUX2_X1 U14533 ( .A(n13834), .B(n12064), .S(n12066), .Z(n12065) );
  MUX2_X1 U14534 ( .A(n13833), .B(n12067), .S(n12066), .Z(n12069) );
  MUX2_X1 U14535 ( .A(n13833), .B(n12067), .S(n12152), .Z(n12068) );
  MUX2_X1 U14536 ( .A(n13832), .B(n14671), .S(n12152), .Z(n12071) );
  MUX2_X1 U14537 ( .A(n13832), .B(n14671), .S(n12066), .Z(n12070) );
  MUX2_X1 U14538 ( .A(n13831), .B(n14744), .S(n12066), .Z(n12074) );
  MUX2_X1 U14539 ( .A(n13831), .B(n14744), .S(n12152), .Z(n12072) );
  INV_X1 U14540 ( .A(n12074), .ZN(n12075) );
  MUX2_X1 U14541 ( .A(n13830), .B(n14607), .S(n12152), .Z(n12076) );
  NAND2_X1 U14542 ( .A1(n12077), .A2(n12076), .ZN(n12079) );
  MUX2_X1 U14543 ( .A(n13830), .B(n14607), .S(n12066), .Z(n12078) );
  NAND2_X1 U14544 ( .A1(n12079), .A2(n12078), .ZN(n12080) );
  MUX2_X1 U14545 ( .A(n13829), .B(n12082), .S(n12066), .Z(n12084) );
  MUX2_X1 U14546 ( .A(n13829), .B(n12082), .S(n12152), .Z(n12083) );
  INV_X1 U14547 ( .A(n12084), .ZN(n12085) );
  MUX2_X1 U14548 ( .A(n13828), .B(n12092), .S(n12152), .Z(n12094) );
  NAND2_X1 U14549 ( .A1(n13828), .A2(n12152), .ZN(n12087) );
  NAND2_X1 U14550 ( .A1(n12092), .A2(n12066), .ZN(n12086) );
  NAND3_X1 U14551 ( .A1(n12094), .A2(n12087), .A3(n12086), .ZN(n12088) );
  NAND2_X1 U14552 ( .A1(n12103), .A2(n12089), .ZN(n12096) );
  NAND2_X1 U14553 ( .A1(n12090), .A2(n12152), .ZN(n12091) );
  OAI21_X1 U14554 ( .B1(n12092), .B2(n12152), .A(n12091), .ZN(n12093) );
  NOR2_X1 U14555 ( .A1(n12094), .A2(n12093), .ZN(n12095) );
  AOI22_X1 U14556 ( .A1(n12096), .A2(n12066), .B1(n12209), .B2(n12095), .ZN(
        n12100) );
  NAND2_X1 U14557 ( .A1(n12102), .A2(n12097), .ZN(n12098) );
  NAND2_X1 U14558 ( .A1(n12098), .A2(n12152), .ZN(n12099) );
  NAND3_X1 U14559 ( .A1(n12101), .A2(n12100), .A3(n12099), .ZN(n12111) );
  MUX2_X1 U14560 ( .A(n12103), .B(n12102), .S(n12066), .Z(n12110) );
  MUX2_X1 U14561 ( .A(n12104), .B(n13751), .S(n12066), .Z(n12115) );
  AND2_X1 U14562 ( .A1(n13825), .A2(n12066), .ZN(n12105) );
  AOI21_X1 U14563 ( .B1(n14276), .B2(n12152), .A(n12105), .ZN(n12106) );
  NAND3_X1 U14564 ( .A1(n12108), .A2(n12107), .A3(n12106), .ZN(n12116) );
  OAI21_X1 U14565 ( .B1(n12232), .B2(n12115), .A(n12116), .ZN(n12109) );
  AND2_X1 U14566 ( .A1(n13824), .A2(n12152), .ZN(n12113) );
  OAI21_X1 U14567 ( .B1(n12152), .B2(n13824), .A(n13761), .ZN(n12112) );
  OAI21_X1 U14568 ( .B1(n12113), .B2(n13761), .A(n12112), .ZN(n12114) );
  OAI21_X1 U14569 ( .B1(n12116), .B2(n12115), .A(n12114), .ZN(n12117) );
  INV_X1 U14570 ( .A(n12119), .ZN(n12122) );
  INV_X1 U14571 ( .A(n12120), .ZN(n12121) );
  MUX2_X1 U14572 ( .A(n12122), .B(n12121), .S(n12152), .Z(n12123) );
  MUX2_X1 U14573 ( .A(n12125), .B(n12124), .S(n12152), .Z(n12126) );
  MUX2_X1 U14574 ( .A(n14248), .B(n13821), .S(n12152), .Z(n12130) );
  NAND2_X1 U14575 ( .A1(n12129), .A2(n12130), .ZN(n12128) );
  MUX2_X1 U14576 ( .A(n14248), .B(n13821), .S(n12066), .Z(n12127) );
  NAND2_X1 U14577 ( .A1(n12128), .A2(n12127), .ZN(n12134) );
  INV_X1 U14578 ( .A(n12129), .ZN(n12132) );
  INV_X1 U14579 ( .A(n12130), .ZN(n12131) );
  NAND2_X1 U14580 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  MUX2_X1 U14581 ( .A(n13820), .B(n14303), .S(n12152), .Z(n12136) );
  MUX2_X1 U14582 ( .A(n13820), .B(n14303), .S(n12066), .Z(n12135) );
  INV_X1 U14583 ( .A(n12136), .ZN(n12137) );
  INV_X1 U14584 ( .A(n14234), .ZN(n12138) );
  MUX2_X1 U14585 ( .A(n13819), .B(n12138), .S(n12066), .Z(n12141) );
  MUX2_X1 U14586 ( .A(n13724), .B(n14234), .S(n12152), .Z(n12139) );
  INV_X1 U14587 ( .A(n12140), .ZN(n12143) );
  NAND2_X1 U14588 ( .A1(n12143), .A2(n6723), .ZN(n12147) );
  NAND2_X1 U14589 ( .A1(n12147), .A2(n12148), .ZN(n12145) );
  MUX2_X1 U14590 ( .A(n14081), .B(n14110), .S(n12066), .Z(n12144) );
  NAND2_X1 U14591 ( .A1(n12145), .A2(n12144), .ZN(n12146) );
  MUX2_X1 U14592 ( .A(n14061), .B(n14094), .S(n12066), .Z(n12151) );
  MUX2_X1 U14593 ( .A(n14091), .B(n12149), .S(n12066), .Z(n12150) );
  MUX2_X1 U14594 ( .A(n14080), .B(n14067), .S(n12152), .Z(n12154) );
  MUX2_X1 U14595 ( .A(n14080), .B(n14067), .S(n12066), .Z(n12153) );
  INV_X1 U14596 ( .A(n12153), .ZN(n12156) );
  MUX2_X1 U14597 ( .A(n14060), .B(n14049), .S(n12066), .Z(n12160) );
  NAND2_X1 U14598 ( .A1(n12159), .A2(n12160), .ZN(n12158) );
  MUX2_X1 U14599 ( .A(n14049), .B(n14060), .S(n12066), .Z(n12157) );
  NAND2_X1 U14600 ( .A1(n12158), .A2(n12157), .ZN(n12164) );
  INV_X1 U14601 ( .A(n12159), .ZN(n12162) );
  INV_X1 U14602 ( .A(n12160), .ZN(n12161) );
  NAND2_X1 U14603 ( .A1(n12162), .A2(n12161), .ZN(n12163) );
  NAND2_X1 U14604 ( .A1(n12164), .A2(n12163), .ZN(n12167) );
  MUX2_X1 U14605 ( .A(n14032), .B(n14042), .S(n12066), .Z(n12168) );
  NAND2_X1 U14606 ( .A1(n12167), .A2(n12168), .ZN(n12166) );
  MUX2_X1 U14607 ( .A(n14042), .B(n14032), .S(n12066), .Z(n12165) );
  NAND2_X1 U14608 ( .A1(n12166), .A2(n12165), .ZN(n12172) );
  INV_X1 U14609 ( .A(n12167), .ZN(n12170) );
  INV_X1 U14610 ( .A(n12168), .ZN(n12169) );
  NAND2_X1 U14611 ( .A1(n12170), .A2(n12169), .ZN(n12171) );
  MUX2_X1 U14612 ( .A(n13818), .B(n14200), .S(n12066), .Z(n12174) );
  MUX2_X1 U14613 ( .A(n13818), .B(n14200), .S(n12152), .Z(n12173) );
  MUX2_X1 U14614 ( .A(n14002), .B(n13992), .S(n12152), .Z(n12176) );
  MUX2_X1 U14615 ( .A(n14002), .B(n13992), .S(n12066), .Z(n12175) );
  INV_X1 U14616 ( .A(n12176), .ZN(n12177) );
  INV_X1 U14617 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U14618 ( .A1(n12178), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12181) );
  INV_X1 U14619 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14193) );
  OR2_X1 U14620 ( .A1(n12179), .A2(n14193), .ZN(n12180) );
  OAI211_X1 U14621 ( .C1(n6650), .C2(n12182), .A(n12181), .B(n12180), .ZN(
        n13975) );
  OAI21_X1 U14622 ( .B1(n13975), .B2(n12183), .A(n13817), .ZN(n12184) );
  INV_X1 U14623 ( .A(n12184), .ZN(n12187) );
  NAND2_X1 U14624 ( .A1(n12266), .A2(n12195), .ZN(n12186) );
  NAND2_X1 U14625 ( .A1(n12196), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12185) );
  MUX2_X1 U14626 ( .A(n12187), .B(n13985), .S(n12066), .Z(n12192) );
  INV_X1 U14627 ( .A(n13817), .ZN(n12191) );
  INV_X1 U14628 ( .A(n12188), .ZN(n12189) );
  AOI21_X1 U14629 ( .B1(n13975), .B2(n12066), .A(n12189), .ZN(n12190) );
  OAI22_X1 U14630 ( .A1(n14288), .A2(n12066), .B1(n12191), .B2(n12190), .ZN(
        n12193) );
  NAND2_X1 U14631 ( .A1(n12194), .A2(n12195), .ZN(n12198) );
  NAND2_X1 U14632 ( .A1(n12196), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12197) );
  INV_X1 U14633 ( .A(n13975), .ZN(n12203) );
  XNOR2_X1 U14634 ( .A(n12202), .B(n12203), .ZN(n12246) );
  OAI21_X1 U14635 ( .B1(n12201), .B2(n12200), .A(n12199), .ZN(n12248) );
  NOR3_X1 U14636 ( .A1(n12208), .A2(n12246), .A3(n12248), .ZN(n12255) );
  MUX2_X1 U14637 ( .A(n12202), .B(n13975), .S(n12066), .Z(n12204) );
  INV_X1 U14638 ( .A(n12247), .ZN(n12207) );
  NAND2_X1 U14639 ( .A1(n12206), .A2(n12205), .ZN(n12251) );
  AND3_X1 U14640 ( .A1(n12208), .A2(n12207), .A3(n7560), .ZN(n12254) );
  INV_X1 U14641 ( .A(n12246), .ZN(n12244) );
  INV_X1 U14642 ( .A(n12209), .ZN(n12231) );
  NOR3_X1 U14643 ( .A1(n12212), .A2(n12211), .A3(n12210), .ZN(n12215) );
  NAND4_X1 U14644 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n12217) );
  NOR2_X1 U14645 ( .A1(n12218), .A2(n12217), .ZN(n12221) );
  NAND4_X1 U14646 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(
        n12223) );
  NOR2_X1 U14647 ( .A1(n12224), .A2(n12223), .ZN(n12227) );
  NAND4_X1 U14648 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12229) );
  NOR4_X1 U14649 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12233) );
  NAND4_X1 U14650 ( .A1(n14168), .A2(n6876), .A3(n12234), .A4(n12233), .ZN(
        n12235) );
  NOR4_X1 U14651 ( .A1(n14126), .A2(n14142), .A3(n14157), .A4(n12235), .ZN(
        n12236) );
  NAND4_X1 U14652 ( .A1(n12237), .A2(n12236), .A3(n14083), .A4(n14106), .ZN(
        n12238) );
  NOR4_X1 U14653 ( .A1(n12240), .A2(n14021), .A3(n12239), .A4(n12238), .ZN(
        n12243) );
  XNOR2_X1 U14654 ( .A(n13985), .B(n13817), .ZN(n12242) );
  NAND4_X1 U14655 ( .A1(n12244), .A2(n12243), .A3(n12242), .A4(n12241), .ZN(
        n12245) );
  XNOR2_X1 U14656 ( .A(n12245), .B(n8775), .ZN(n12252) );
  NAND2_X1 U14657 ( .A1(n12246), .A2(n7560), .ZN(n12249) );
  MUX2_X1 U14658 ( .A(n12249), .B(n12248), .S(n12247), .Z(n12250) );
  OAI21_X1 U14659 ( .B1(n12252), .B2(n12251), .A(n12250), .ZN(n12253) );
  NOR3_X1 U14660 ( .A1(n12255), .A2(n12254), .A3(n12253), .ZN(n12261) );
  NAND3_X1 U14661 ( .A1(n12257), .A2(n12256), .A3(n14082), .ZN(n12258) );
  OAI211_X1 U14662 ( .C1(n14335), .C2(n12260), .A(n12258), .B(P1_B_REG_SCAN_IN), .ZN(n12259) );
  OAI21_X1 U14663 ( .B1(n12261), .B2(n12260), .A(n12259), .ZN(P1_U3242) );
  OAI222_X1 U14664 ( .A1(n13693), .A2(n12263), .B1(P2_U3088), .B2(n6656), .C1(
        n11317), .C2(n12262), .ZN(P2_U3307) );
  INV_X1 U14665 ( .A(n13686), .ZN(n12264) );
  OAI222_X1 U14666 ( .A1(n14332), .A2(n12265), .B1(n14330), .B2(n12264), .C1(
        P1_U3086), .C2(n8816), .ZN(P1_U3327) );
  INV_X1 U14667 ( .A(n12266), .ZN(n12335) );
  INV_X1 U14668 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12346) );
  OAI222_X1 U14669 ( .A1(n11317), .A2(n12335), .B1(P2_U3088), .B2(n12267), 
        .C1(n12346), .C2(n13693), .ZN(P2_U3297) );
  NAND2_X1 U14670 ( .A1(n14110), .A2(n12326), .ZN(n12270) );
  NAND2_X1 U14671 ( .A1(n14081), .A2(n12323), .ZN(n12269) );
  NAND2_X1 U14672 ( .A1(n12270), .A2(n12269), .ZN(n12271) );
  XNOR2_X1 U14673 ( .A(n12271), .B(n12295), .ZN(n12273) );
  AND2_X1 U14674 ( .A1(n14081), .A2(n12322), .ZN(n12272) );
  AOI21_X1 U14675 ( .B1(n14110), .B2(n12323), .A(n12272), .ZN(n12274) );
  NAND2_X1 U14676 ( .A1(n12273), .A2(n12274), .ZN(n13764) );
  INV_X1 U14677 ( .A(n12273), .ZN(n12276) );
  INV_X1 U14678 ( .A(n12274), .ZN(n12275) );
  NAND2_X1 U14679 ( .A1(n12276), .A2(n12275), .ZN(n12277) );
  INV_X1 U14680 ( .A(n13703), .ZN(n12281) );
  AND2_X1 U14681 ( .A1(n12279), .A2(n13702), .ZN(n12280) );
  AND2_X1 U14682 ( .A1(n13706), .A2(n13764), .ZN(n12282) );
  NAND2_X1 U14683 ( .A1(n13707), .A2(n12282), .ZN(n12292) );
  NAND2_X1 U14684 ( .A1(n14094), .A2(n12326), .ZN(n12284) );
  NAND2_X1 U14685 ( .A1(n14061), .A2(n6648), .ZN(n12283) );
  NAND2_X1 U14686 ( .A1(n12284), .A2(n12283), .ZN(n12285) );
  XNOR2_X1 U14687 ( .A(n12285), .B(n12295), .ZN(n12287) );
  AND2_X1 U14688 ( .A1(n14061), .A2(n12322), .ZN(n12286) );
  AOI21_X1 U14689 ( .B1(n14094), .B2(n12323), .A(n12286), .ZN(n12288) );
  NAND2_X1 U14690 ( .A1(n12287), .A2(n12288), .ZN(n13734) );
  INV_X1 U14691 ( .A(n12287), .ZN(n12290) );
  INV_X1 U14692 ( .A(n12288), .ZN(n12289) );
  NAND2_X1 U14693 ( .A1(n12290), .A2(n12289), .ZN(n12291) );
  NAND2_X1 U14694 ( .A1(n12292), .A2(n13765), .ZN(n13731) );
  NAND2_X1 U14695 ( .A1(n13731), .A2(n13734), .ZN(n12303) );
  NAND2_X1 U14696 ( .A1(n14067), .A2(n12326), .ZN(n12294) );
  NAND2_X1 U14697 ( .A1(n14080), .A2(n12323), .ZN(n12293) );
  NAND2_X1 U14698 ( .A1(n12294), .A2(n12293), .ZN(n12296) );
  XNOR2_X1 U14699 ( .A(n12296), .B(n12295), .ZN(n12298) );
  AND2_X1 U14700 ( .A1(n14080), .A2(n12322), .ZN(n12297) );
  AOI21_X1 U14701 ( .B1(n14067), .B2(n12323), .A(n12297), .ZN(n12299) );
  NAND2_X1 U14702 ( .A1(n12298), .A2(n12299), .ZN(n12304) );
  INV_X1 U14703 ( .A(n12298), .ZN(n12301) );
  INV_X1 U14704 ( .A(n12299), .ZN(n12300) );
  NAND2_X1 U14705 ( .A1(n12301), .A2(n12300), .ZN(n12302) );
  AND2_X1 U14706 ( .A1(n12304), .A2(n12302), .ZN(n13732) );
  NAND2_X1 U14707 ( .A1(n12303), .A2(n13732), .ZN(n13736) );
  NAND2_X1 U14708 ( .A1(n14049), .A2(n12326), .ZN(n12306) );
  NAND2_X1 U14709 ( .A1(n14060), .A2(n12323), .ZN(n12305) );
  NAND2_X1 U14710 ( .A1(n12306), .A2(n12305), .ZN(n12307) );
  XNOR2_X1 U14711 ( .A(n12307), .B(n12324), .ZN(n12311) );
  NAND2_X1 U14712 ( .A1(n14049), .A2(n12323), .ZN(n12309) );
  NAND2_X1 U14713 ( .A1(n14060), .A2(n12322), .ZN(n12308) );
  NAND2_X1 U14714 ( .A1(n12309), .A2(n12308), .ZN(n12310) );
  NOR2_X1 U14715 ( .A1(n12311), .A2(n12310), .ZN(n12312) );
  AOI21_X1 U14716 ( .B1(n12311), .B2(n12310), .A(n12312), .ZN(n13795) );
  INV_X1 U14717 ( .A(n12312), .ZN(n12313) );
  NAND2_X1 U14718 ( .A1(n14032), .A2(n12326), .ZN(n12315) );
  NAND2_X1 U14719 ( .A1(n14042), .A2(n12323), .ZN(n12314) );
  NAND2_X1 U14720 ( .A1(n12315), .A2(n12314), .ZN(n12316) );
  XNOR2_X1 U14721 ( .A(n12316), .B(n12324), .ZN(n12320) );
  NAND2_X1 U14722 ( .A1(n14032), .A2(n6648), .ZN(n12318) );
  NAND2_X1 U14723 ( .A1(n14042), .A2(n12322), .ZN(n12317) );
  NAND2_X1 U14724 ( .A1(n12318), .A2(n12317), .ZN(n12319) );
  NOR2_X1 U14725 ( .A1(n12320), .A2(n12319), .ZN(n12321) );
  AOI21_X1 U14726 ( .B1(n12320), .B2(n12319), .A(n12321), .ZN(n13696) );
  AOI22_X1 U14727 ( .A1(n14200), .A2(n6648), .B1(n12322), .B2(n13818), .ZN(
        n12325) );
  XNOR2_X1 U14728 ( .A(n12325), .B(n12324), .ZN(n12328) );
  AOI22_X1 U14729 ( .A1(n14200), .A2(n12326), .B1(n6648), .B2(n13818), .ZN(
        n12327) );
  XNOR2_X1 U14730 ( .A(n12328), .B(n12327), .ZN(n12329) );
  AOI22_X1 U14731 ( .A1(n13789), .A2(n14042), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12331) );
  NAND2_X1 U14732 ( .A1(n13797), .A2(n14002), .ZN(n12330) );
  OAI211_X1 U14733 ( .C1(n14606), .C2(n14012), .A(n12331), .B(n12330), .ZN(
        n12332) );
  AOI21_X1 U14734 ( .B1(n14200), .B2(n14602), .A(n12332), .ZN(n12333) );
  OAI21_X1 U14735 ( .B1(n12334), .B2(n14598), .A(n12333), .ZN(P1_U3220) );
  INV_X1 U14736 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15473) );
  OAI222_X1 U14737 ( .A1(n14330), .A2(n12335), .B1(P1_U3086), .B2(n8220), .C1(
        n15473), .C2(n14332), .ZN(P1_U3325) );
  INV_X1 U14738 ( .A(n12336), .ZN(n12341) );
  NOR2_X1 U14739 ( .A1(n12337), .A2(n15108), .ZN(n12795) );
  AOI21_X1 U14740 ( .B1(n15146), .B2(P3_REG2_REG_29__SCAN_IN), .A(n12795), 
        .ZN(n12338) );
  OAI21_X1 U14741 ( .B1(n12339), .B2(n12998), .A(n12338), .ZN(n12340) );
  AOI21_X1 U14742 ( .B1(n12341), .B2(n15141), .A(n12340), .ZN(n12342) );
  OAI21_X1 U14743 ( .B1(n12343), .B2(n15146), .A(n12342), .ZN(P3_U3204) );
  NAND2_X1 U14744 ( .A1(n14326), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12344) );
  NAND2_X1 U14745 ( .A1(n12345), .A2(n12344), .ZN(n12474) );
  NAND2_X1 U14746 ( .A1(n15473), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12475) );
  NAND2_X1 U14747 ( .A1(n12346), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12347) );
  AND2_X1 U14748 ( .A1(n12475), .A2(n12347), .ZN(n12473) );
  INV_X1 U14749 ( .A(n12473), .ZN(n12348) );
  XNOR2_X1 U14750 ( .A(n12474), .B(n12348), .ZN(n12463) );
  INV_X1 U14751 ( .A(n12463), .ZN(n12349) );
  OAI222_X1 U14752 ( .A1(n12350), .A2(n12464), .B1(n11060), .B2(n12349), .C1(
        n7706), .C2(P3_U3151), .ZN(P3_U3265) );
  XOR2_X1 U14753 ( .A(n12352), .B(n12351), .Z(n12359) );
  OAI22_X1 U14754 ( .A1(n12354), .A2(n15136), .B1(n12353), .B2(n15134), .ZN(
        n12818) );
  INV_X1 U14755 ( .A(n12818), .ZN(n12356) );
  AOI22_X1 U14756 ( .A1(n12823), .A2(n12451), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12355) );
  OAI21_X1 U14757 ( .B1(n12356), .B2(n12454), .A(n12355), .ZN(n12357) );
  AOI21_X1 U14758 ( .B1(n12822), .B2(n12456), .A(n12357), .ZN(n12358) );
  OAI21_X1 U14759 ( .B1(n12359), .B2(n12459), .A(n12358), .ZN(P3_U3154) );
  XNOR2_X1 U14760 ( .A(n12410), .B(n12409), .ZN(n12411) );
  XNOR2_X1 U14761 ( .A(n12411), .B(n12650), .ZN(n12364) );
  AOI22_X1 U14762 ( .A1(n12703), .A2(n12990), .B1(n12993), .B2(n12705), .ZN(
        n12867) );
  INV_X1 U14763 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12360) );
  OAI22_X1 U14764 ( .A1(n12867), .A2(n12454), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12360), .ZN(n12362) );
  NOR2_X1 U14765 ( .A1(n13096), .A2(n12446), .ZN(n12361) );
  AOI211_X1 U14766 ( .C1(n12871), .C2(n12451), .A(n12362), .B(n12361), .ZN(
        n12363) );
  OAI21_X1 U14767 ( .B1(n12364), .B2(n12459), .A(n12363), .ZN(P3_U3156) );
  OAI211_X1 U14768 ( .C1(n12367), .C2(n12366), .A(n12365), .B(n12436), .ZN(
        n12374) );
  OR2_X1 U14769 ( .A1(n12921), .A2(n12368), .ZN(n12369) );
  NAND2_X1 U14770 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12768)
         );
  OAI211_X1 U14771 ( .C1(n12442), .C2(n12918), .A(n12369), .B(n12768), .ZN(
        n12370) );
  INV_X1 U14772 ( .A(n12370), .ZN(n12373) );
  OR2_X1 U14773 ( .A1(n13112), .A2(n12446), .ZN(n12372) );
  NAND2_X1 U14774 ( .A1(n12451), .A2(n12922), .ZN(n12371) );
  NAND4_X1 U14775 ( .A1(n12374), .A2(n12373), .A3(n12372), .A4(n12371), .ZN(
        P3_U3159) );
  AOI21_X1 U14776 ( .B1(n12376), .B2(n12375), .A(n6724), .ZN(n12381) );
  AOI22_X1 U14777 ( .A1(n12706), .A2(n12993), .B1(n12990), .B2(n12705), .ZN(
        n12888) );
  INV_X1 U14778 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12377) );
  OAI22_X1 U14779 ( .A1(n12888), .A2(n12454), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12377), .ZN(n12379) );
  NOR2_X1 U14780 ( .A1(n13104), .A2(n12446), .ZN(n12378) );
  AOI211_X1 U14781 ( .C1(n12892), .C2(n12451), .A(n12379), .B(n12378), .ZN(
        n12380) );
  OAI21_X1 U14782 ( .B1(n12381), .B2(n12459), .A(n12380), .ZN(P3_U3163) );
  XOR2_X1 U14783 ( .A(n12383), .B(n12382), .Z(n12388) );
  AOI22_X1 U14784 ( .A1(n12702), .A2(n12990), .B1(n12993), .B2(n12703), .ZN(
        n12842) );
  OAI22_X1 U14785 ( .A1(n12842), .A2(n12454), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12384), .ZN(n12386) );
  NOR2_X1 U14786 ( .A1(n13091), .A2(n12446), .ZN(n12385) );
  AOI211_X1 U14787 ( .C1(n12844), .C2(n12451), .A(n12386), .B(n12385), .ZN(
        n12387) );
  OAI21_X1 U14788 ( .B1(n12388), .B2(n12459), .A(n12387), .ZN(P3_U3165) );
  INV_X1 U14789 ( .A(n12969), .ZN(n12392) );
  OR2_X1 U14790 ( .A1(n12930), .A2(n15136), .ZN(n12390) );
  NAND2_X1 U14791 ( .A1(n12991), .A2(n12993), .ZN(n12389) );
  NAND2_X1 U14792 ( .A1(n12390), .A2(n12389), .ZN(n12962) );
  AOI22_X1 U14793 ( .A1(n12962), .A2(n12416), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12391) );
  OAI21_X1 U14794 ( .B1(n12392), .B2(n12418), .A(n12391), .ZN(n12398) );
  INV_X1 U14795 ( .A(n12393), .ZN(n12394) );
  AOI211_X1 U14796 ( .C1(n12396), .C2(n12395), .A(n12459), .B(n12394), .ZN(
        n12397) );
  AOI211_X1 U14797 ( .C1(n12456), .C2(n12399), .A(n12398), .B(n12397), .ZN(
        n12400) );
  INV_X1 U14798 ( .A(n12400), .ZN(P3_U3166) );
  INV_X1 U14799 ( .A(n13052), .ZN(n12957) );
  OAI211_X1 U14800 ( .C1(n12403), .C2(n12402), .A(n12401), .B(n12436), .ZN(
        n12408) );
  AOI22_X1 U14801 ( .A1(n12947), .A2(n12440), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12404) );
  OAI21_X1 U14802 ( .B1(n12405), .B2(n12442), .A(n12404), .ZN(n12406) );
  AOI21_X1 U14803 ( .B1(n12955), .B2(n12451), .A(n12406), .ZN(n12407) );
  OAI211_X1 U14804 ( .C1(n12957), .C2(n12446), .A(n12408), .B(n12407), .ZN(
        P3_U3168) );
  OAI22_X1 U14805 ( .A1(n12411), .A2(n12704), .B1(n12410), .B2(n12409), .ZN(
        n12415) );
  XNOR2_X1 U14806 ( .A(n12413), .B(n12412), .ZN(n12414) );
  XNOR2_X1 U14807 ( .A(n12415), .B(n12414), .ZN(n12422) );
  INV_X1 U14808 ( .A(n12856), .ZN(n12419) );
  OAI22_X1 U14809 ( .A1(n12656), .A2(n15136), .B1(n12650), .B2(n15134), .ZN(
        n12852) );
  AOI22_X1 U14810 ( .A1(n12852), .A2(n12416), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12417) );
  OAI21_X1 U14811 ( .B1(n12419), .B2(n12418), .A(n12417), .ZN(n12420) );
  AOI21_X1 U14812 ( .B1(n13021), .B2(n12456), .A(n12420), .ZN(n12421) );
  OAI21_X1 U14813 ( .B1(n12422), .B2(n12459), .A(n12421), .ZN(P3_U3169) );
  OAI211_X1 U14814 ( .C1(n12425), .C2(n12424), .A(n12423), .B(n12436), .ZN(
        n12429) );
  AOI22_X1 U14815 ( .A1(n12440), .A2(n12898), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12426) );
  OAI21_X1 U14816 ( .B1(n12931), .B2(n12442), .A(n12426), .ZN(n12427) );
  AOI21_X1 U14817 ( .B1(n12901), .B2(n12451), .A(n12427), .ZN(n12428) );
  OAI211_X1 U14818 ( .C1(n13108), .C2(n12446), .A(n12429), .B(n12428), .ZN(
        P3_U3173) );
  XNOR2_X1 U14819 ( .A(n12430), .B(n12705), .ZN(n12435) );
  AOI22_X1 U14820 ( .A1(n12704), .A2(n12990), .B1(n12993), .B2(n12898), .ZN(
        n12878) );
  OAI22_X1 U14821 ( .A1(n12878), .A2(n12454), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12431), .ZN(n12433) );
  NOR2_X1 U14822 ( .A1(n13100), .A2(n12446), .ZN(n12432) );
  AOI211_X1 U14823 ( .C1(n12882), .C2(n12451), .A(n12433), .B(n12432), .ZN(
        n12434) );
  OAI21_X1 U14824 ( .B1(n12435), .B2(n12459), .A(n12434), .ZN(P3_U3175) );
  OAI211_X1 U14825 ( .C1(n12439), .C2(n12438), .A(n12437), .B(n12436), .ZN(
        n12445) );
  AOI22_X1 U14826 ( .A1(n12440), .A2(n12899), .B1(P3_REG3_REG_18__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12441) );
  OAI21_X1 U14827 ( .B1(n12930), .B2(n12442), .A(n12441), .ZN(n12443) );
  AOI21_X1 U14828 ( .B1(n12940), .B2(n12451), .A(n12443), .ZN(n12444) );
  OAI211_X1 U14829 ( .C1(n13116), .C2(n12446), .A(n12445), .B(n12444), .ZN(
        P3_U3178) );
  XOR2_X1 U14830 ( .A(n12448), .B(n12447), .Z(n12460) );
  OR2_X1 U14831 ( .A1(n12802), .A2(n15136), .ZN(n12450) );
  OR2_X1 U14832 ( .A1(n12656), .A2(n15134), .ZN(n12449) );
  AND2_X1 U14833 ( .A1(n12450), .A2(n12449), .ZN(n12829) );
  NAND2_X1 U14834 ( .A1(n12833), .A2(n12451), .ZN(n12453) );
  NAND2_X1 U14835 ( .A1(P3_U3151), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n12452)
         );
  OAI211_X1 U14836 ( .C1(n12829), .C2(n12454), .A(n12453), .B(n12452), .ZN(
        n12455) );
  AOI21_X1 U14837 ( .B1(n12457), .B2(n12456), .A(n12455), .ZN(n12458) );
  OAI21_X1 U14838 ( .B1(n12460), .B2(n12459), .A(n12458), .ZN(P3_U3180) );
  INV_X1 U14839 ( .A(n12461), .ZN(n12679) );
  NOR2_X1 U14840 ( .A1(n12462), .A2(n12679), .ZN(n12490) );
  NAND2_X1 U14841 ( .A1(n12463), .A2(n12480), .ZN(n12466) );
  OR2_X1 U14842 ( .A1(n7882), .A2(n12464), .ZN(n12465) );
  NAND2_X1 U14843 ( .A1(n12466), .A2(n12465), .ZN(n14532) );
  INV_X1 U14844 ( .A(n14532), .ZN(n12486) );
  NAND2_X1 U14845 ( .A1(n12467), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12470) );
  NAND2_X1 U14846 ( .A1(n8083), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12469) );
  NAND2_X1 U14847 ( .A1(n8058), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12468) );
  AND3_X1 U14848 ( .A1(n12470), .A2(n12469), .A3(n12468), .ZN(n12471) );
  INV_X1 U14849 ( .A(n12794), .ZN(n12699) );
  NAND2_X1 U14850 ( .A1(n12474), .A2(n12473), .ZN(n12476) );
  NAND2_X1 U14851 ( .A1(n12476), .A2(n12475), .ZN(n12479) );
  INV_X1 U14852 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12477) );
  XNOR2_X1 U14853 ( .A(n12477), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12478) );
  XNOR2_X1 U14854 ( .A(n12479), .B(n12478), .ZN(n13136) );
  NAND2_X1 U14855 ( .A1(n13136), .A2(n12480), .ZN(n12482) );
  INV_X1 U14856 ( .A(SI_31_), .ZN(n13141) );
  OR2_X1 U14857 ( .A1(n7882), .A2(n13141), .ZN(n12481) );
  NAND2_X1 U14858 ( .A1(n12482), .A2(n12481), .ZN(n12493) );
  OR2_X1 U14859 ( .A1(n12493), .A2(n12794), .ZN(n12527) );
  NAND2_X1 U14860 ( .A1(n14532), .A2(n12487), .ZN(n12483) );
  NAND2_X1 U14861 ( .A1(n12527), .A2(n12483), .ZN(n12524) );
  INV_X1 U14862 ( .A(n12484), .ZN(n12485) );
  NOR2_X1 U14863 ( .A1(n12524), .A2(n12485), .ZN(n12677) );
  OAI21_X1 U14864 ( .B1(n12486), .B2(n12699), .A(n12677), .ZN(n12489) );
  NOR2_X1 U14865 ( .A1(n14532), .A2(n12487), .ZN(n12494) );
  NOR2_X1 U14866 ( .A1(n12494), .A2(n12794), .ZN(n12488) );
  OAI22_X1 U14867 ( .A1(n12490), .A2(n12489), .B1(n13076), .B2(n12488), .ZN(
        n12491) );
  XNOR2_X1 U14868 ( .A(n12491), .B(n12525), .ZN(n12689) );
  INV_X1 U14869 ( .A(n12492), .ZN(n12688) );
  NAND2_X1 U14870 ( .A1(n12493), .A2(n12794), .ZN(n12496) );
  INV_X1 U14871 ( .A(n12494), .ZN(n12495) );
  AND2_X1 U14872 ( .A1(n12496), .A2(n12495), .ZN(n12681) );
  INV_X1 U14873 ( .A(n12681), .ZN(n12523) );
  INV_X1 U14874 ( .A(n12816), .ZN(n12668) );
  INV_X1 U14875 ( .A(n12665), .ZN(n12497) );
  NAND2_X1 U14876 ( .A1(n8127), .A2(n12499), .ZN(n12640) );
  AND2_X1 U14877 ( .A1(n12557), .A2(n12500), .ZN(n12504) );
  NOR2_X1 U14878 ( .A1(n12502), .A2(n12501), .ZN(n12503) );
  INV_X1 U14879 ( .A(n15139), .ZN(n15130) );
  NAND4_X1 U14880 ( .A1(n12504), .A2(n12579), .A3(n12503), .A4(n15130), .ZN(
        n12510) );
  NOR2_X1 U14881 ( .A1(n12568), .A2(n12505), .ZN(n12508) );
  NAND4_X1 U14882 ( .A1(n12508), .A2(n12507), .A3(n12506), .A4(n12572), .ZN(
        n12509) );
  NOR2_X1 U14883 ( .A1(n12510), .A2(n12509), .ZN(n12513) );
  INV_X1 U14884 ( .A(n12511), .ZN(n12587) );
  NAND4_X1 U14885 ( .A1(n12513), .A2(n12512), .A3(n12599), .A4(n12587), .ZN(
        n12514) );
  NOR2_X1 U14886 ( .A1(n12514), .A2(n12988), .ZN(n12515) );
  NAND4_X1 U14887 ( .A1(n12936), .A2(n12978), .A3(n12965), .A4(n12515), .ZN(
        n12516) );
  NOR4_X1 U14888 ( .A1(n12890), .A2(n12917), .A3(n12517), .A4(n12516), .ZN(
        n12518) );
  NAND4_X1 U14889 ( .A1(n12863), .A2(n8004), .A3(n12881), .A4(n12518), .ZN(
        n12519) );
  NOR4_X1 U14890 ( .A1(n12832), .A2(n12840), .A3(n12854), .A4(n12519), .ZN(
        n12520) );
  NAND4_X1 U14891 ( .A1(n12521), .A2(n12668), .A3(n12800), .A4(n12520), .ZN(
        n12522) );
  NOR3_X1 U14892 ( .A1(n12524), .A2(n12523), .A3(n12522), .ZN(n12526) );
  XNOR2_X1 U14893 ( .A(n12526), .B(n12525), .ZN(n12685) );
  INV_X1 U14894 ( .A(n12527), .ZN(n12682) );
  OAI21_X1 U14895 ( .B1(n12529), .B2(n12676), .A(n12528), .ZN(n12675) );
  AOI21_X1 U14896 ( .B1(n12531), .B2(n12530), .A(n12672), .ZN(n12533) );
  MUX2_X1 U14897 ( .A(n12657), .B(n12533), .S(n12532), .Z(n12663) );
  OR2_X1 U14898 ( .A1(n12534), .A2(n12657), .ZN(n12574) );
  NAND3_X1 U14899 ( .A1(n12539), .A2(n12536), .A3(n12535), .ZN(n12537) );
  NAND2_X1 U14900 ( .A1(n12537), .A2(n12676), .ZN(n12538) );
  NAND2_X1 U14901 ( .A1(n15114), .A2(n12538), .ZN(n12544) );
  NAND2_X1 U14902 ( .A1(n12539), .A2(n12672), .ZN(n12540) );
  AOI21_X1 U14903 ( .B1(n12542), .B2(n12541), .A(n12540), .ZN(n12543) );
  AOI21_X1 U14904 ( .B1(n15104), .B2(n12544), .A(n12543), .ZN(n12553) );
  NAND2_X1 U14905 ( .A1(n12550), .A2(n12545), .ZN(n12548) );
  NAND2_X1 U14906 ( .A1(n12549), .A2(n12546), .ZN(n12547) );
  MUX2_X1 U14907 ( .A(n12548), .B(n12547), .S(n12676), .Z(n12552) );
  MUX2_X1 U14908 ( .A(n12550), .B(n12549), .S(n12657), .Z(n12551) );
  OAI211_X1 U14909 ( .C1(n12553), .C2(n12552), .A(n8097), .B(n12551), .ZN(
        n12558) );
  MUX2_X1 U14910 ( .A(n12555), .B(n12554), .S(n12676), .Z(n12556) );
  NAND3_X1 U14911 ( .A1(n12558), .A2(n12557), .A3(n12556), .ZN(n12562) );
  NAND2_X1 U14912 ( .A1(n12571), .A2(n12559), .ZN(n12560) );
  NAND2_X1 U14913 ( .A1(n12560), .A2(n12672), .ZN(n12561) );
  NAND2_X1 U14914 ( .A1(n12562), .A2(n12561), .ZN(n12566) );
  AOI21_X1 U14915 ( .B1(n12565), .B2(n12563), .A(n12672), .ZN(n12564) );
  AOI21_X1 U14916 ( .B1(n12566), .B2(n12565), .A(n12564), .ZN(n12569) );
  OAI22_X1 U14917 ( .A1(n12569), .A2(n12568), .B1(n12567), .B2(n12676), .ZN(
        n12570) );
  OAI21_X1 U14918 ( .B1(n12672), .B2(n12571), .A(n12570), .ZN(n12573) );
  OAI211_X1 U14919 ( .C1(n12575), .C2(n12574), .A(n12573), .B(n12572), .ZN(
        n12580) );
  NAND2_X1 U14920 ( .A1(n12712), .A2(n15183), .ZN(n12577) );
  MUX2_X1 U14921 ( .A(n12577), .B(n12576), .S(n12676), .Z(n12578) );
  NAND3_X1 U14922 ( .A1(n12580), .A2(n12579), .A3(n12578), .ZN(n12584) );
  MUX2_X1 U14923 ( .A(n12711), .B(n12657), .S(n15194), .Z(n12582) );
  NAND2_X1 U14924 ( .A1(n12582), .A2(n12581), .ZN(n12583) );
  NAND2_X1 U14925 ( .A1(n12584), .A2(n12583), .ZN(n12591) );
  MUX2_X1 U14926 ( .A(n12586), .B(n12585), .S(n12657), .Z(n12588) );
  NAND2_X1 U14927 ( .A1(n12588), .A2(n12587), .ZN(n12589) );
  AOI21_X1 U14928 ( .B1(n12591), .B2(n12590), .A(n12589), .ZN(n12601) );
  NAND2_X1 U14929 ( .A1(n12709), .A2(n14538), .ZN(n12592) );
  NAND2_X1 U14930 ( .A1(n12597), .A2(n12592), .ZN(n12595) );
  NAND2_X1 U14931 ( .A1(n12596), .A2(n12593), .ZN(n12594) );
  MUX2_X1 U14932 ( .A(n12595), .B(n12594), .S(n12676), .Z(n12600) );
  MUX2_X1 U14933 ( .A(n12597), .B(n12596), .S(n12657), .Z(n12598) );
  OAI211_X1 U14934 ( .C1(n12601), .C2(n12600), .A(n12599), .B(n12598), .ZN(
        n12605) );
  INV_X1 U14935 ( .A(n12988), .ZN(n12985) );
  MUX2_X1 U14936 ( .A(n12603), .B(n12602), .S(n12672), .Z(n12604) );
  NAND4_X1 U14937 ( .A1(n12605), .A2(n12978), .A3(n12985), .A4(n12604), .ZN(
        n12613) );
  INV_X1 U14938 ( .A(n12606), .ZN(n12607) );
  NAND2_X1 U14939 ( .A1(n12978), .A2(n12607), .ZN(n12609) );
  NAND3_X1 U14940 ( .A1(n12609), .A2(n12608), .A3(n12618), .ZN(n12610) );
  NAND2_X1 U14941 ( .A1(n12610), .A2(n12676), .ZN(n12612) );
  INV_X1 U14942 ( .A(n12615), .ZN(n12611) );
  AOI21_X1 U14943 ( .B1(n12613), .B2(n12612), .A(n12611), .ZN(n12620) );
  INV_X1 U14944 ( .A(n12910), .ZN(n12614) );
  NAND2_X1 U14945 ( .A1(n12978), .A2(n12614), .ZN(n12616) );
  NAND3_X1 U14946 ( .A1(n12616), .A2(n12615), .A3(n12964), .ZN(n12617) );
  AND2_X1 U14947 ( .A1(n12617), .A2(n12657), .ZN(n12619) );
  OAI22_X1 U14948 ( .A1(n12620), .A2(n12619), .B1(n12618), .B2(n12676), .ZN(
        n12621) );
  NAND3_X1 U14949 ( .A1(n12621), .A2(n12936), .A3(n12953), .ZN(n12632) );
  NAND2_X1 U14950 ( .A1(n12936), .A2(n12622), .ZN(n12623) );
  NAND3_X1 U14951 ( .A1(n12623), .A2(n12633), .A3(n12624), .ZN(n12629) );
  INV_X1 U14952 ( .A(n12624), .ZN(n12627) );
  OAI211_X1 U14953 ( .C1(n12627), .C2(n12626), .A(n12634), .B(n12625), .ZN(
        n12628) );
  MUX2_X1 U14954 ( .A(n12629), .B(n12628), .S(n12657), .Z(n12630) );
  INV_X1 U14955 ( .A(n12630), .ZN(n12631) );
  NAND2_X1 U14956 ( .A1(n12632), .A2(n12631), .ZN(n12636) );
  MUX2_X1 U14957 ( .A(n12634), .B(n12633), .S(n12672), .Z(n12635) );
  NAND3_X1 U14958 ( .A1(n12636), .A2(n8004), .A3(n12635), .ZN(n12641) );
  MUX2_X1 U14959 ( .A(n12638), .B(n12637), .S(n12676), .Z(n12639) );
  NAND3_X1 U14960 ( .A1(n12641), .A2(n12640), .A3(n12639), .ZN(n12645) );
  MUX2_X1 U14961 ( .A(n12643), .B(n12642), .S(n12657), .Z(n12644) );
  NAND3_X1 U14962 ( .A1(n12645), .A2(n12881), .A3(n12644), .ZN(n12649) );
  MUX2_X1 U14963 ( .A(n12647), .B(n12646), .S(n12676), .Z(n12648) );
  NAND3_X1 U14964 ( .A1(n12649), .A2(n12863), .A3(n12648), .ZN(n12653) );
  NAND3_X1 U14965 ( .A1(n12651), .A2(n12650), .A3(n12657), .ZN(n12652) );
  AOI21_X1 U14966 ( .B1(n12653), .B2(n12652), .A(n12854), .ZN(n12654) );
  OR2_X1 U14967 ( .A1(n12654), .A2(n12840), .ZN(n12662) );
  INV_X1 U14968 ( .A(n12655), .ZN(n12659) );
  NOR2_X1 U14969 ( .A1(n12845), .A2(n12656), .ZN(n12658) );
  MUX2_X1 U14970 ( .A(n12659), .B(n12658), .S(n12657), .Z(n12660) );
  NOR2_X1 U14971 ( .A1(n12832), .A2(n12660), .ZN(n12661) );
  OAI211_X1 U14972 ( .C1(n12663), .C2(n12662), .A(n12661), .B(n12668), .ZN(
        n12670) );
  INV_X1 U14973 ( .A(n12664), .ZN(n12666) );
  NAND2_X1 U14974 ( .A1(n12668), .A2(n12667), .ZN(n12669) );
  OAI211_X1 U14975 ( .C1(n12672), .C2(n12671), .A(n12670), .B(n12669), .ZN(
        n12673) );
  NAND2_X1 U14976 ( .A1(n12673), .A2(n12800), .ZN(n12674) );
  MUX2_X1 U14977 ( .A(n12676), .B(n12675), .S(n12674), .Z(n12678) );
  OAI21_X1 U14978 ( .B1(n12679), .B2(n12678), .A(n12677), .ZN(n12680) );
  OAI21_X1 U14979 ( .B1(n12682), .B2(n12681), .A(n12680), .ZN(n12683) );
  MUX2_X1 U14980 ( .A(n12692), .B(n15137), .S(n12683), .Z(n12684) );
  OAI21_X1 U14981 ( .B1(n12686), .B2(n12685), .A(n12684), .ZN(n12687) );
  AOI21_X1 U14982 ( .B1(n12689), .B2(n12688), .A(n12687), .ZN(n12698) );
  INV_X1 U14983 ( .A(n12690), .ZN(n12691) );
  NOR4_X1 U14984 ( .A1(n15134), .A2(n12693), .A3(n12692), .A4(n12691), .ZN(
        n12696) );
  OAI21_X1 U14985 ( .B1(n12697), .B2(n12694), .A(P3_B_REG_SCAN_IN), .ZN(n12695) );
  OAI22_X1 U14986 ( .A1(n12698), .A2(n12697), .B1(n12696), .B2(n12695), .ZN(
        P3_U3296) );
  MUX2_X1 U14987 ( .A(n12699), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12720), .Z(
        P3_U3522) );
  MUX2_X1 U14988 ( .A(n12700), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12720), .Z(
        P3_U3520) );
  MUX2_X1 U14989 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12701), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14990 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12702), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14991 ( .A(n12703), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12720), .Z(
        P3_U3515) );
  MUX2_X1 U14992 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12704), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14993 ( .A(n12705), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12720), .Z(
        P3_U3513) );
  MUX2_X1 U14994 ( .A(n12898), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12720), .Z(
        P3_U3512) );
  MUX2_X1 U14995 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12706), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14996 ( .A(n12899), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12720), .Z(
        P3_U3510) );
  MUX2_X1 U14997 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12947), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14998 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12707), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14999 ( .A(n12946), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12720), .Z(
        P3_U3507) );
  MUX2_X1 U15000 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12708), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15001 ( .A(n12992), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12720), .Z(
        P3_U3504) );
  MUX2_X1 U15002 ( .A(n12709), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12720), .Z(
        P3_U3502) );
  MUX2_X1 U15003 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12710), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15004 ( .A(n12711), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12720), .Z(
        P3_U3500) );
  MUX2_X1 U15005 ( .A(n12712), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12720), .Z(
        P3_U3499) );
  MUX2_X1 U15006 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12713), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15007 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12714), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15008 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12715), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15009 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12716), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15010 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12717), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15011 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12718), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15012 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12719), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15013 ( .A(n15125), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12720), .Z(
        P3_U3491) );
  XNOR2_X1 U15014 ( .A(n12769), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12737) );
  INV_X1 U15015 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14464) );
  INV_X1 U15016 ( .A(n15071), .ZN(n12749) );
  NOR2_X1 U15017 ( .A1(n12775), .A2(n12723), .ZN(n12724) );
  MUX2_X1 U15018 ( .A(n11089), .B(P3_REG2_REG_12__SCAN_IN), .S(n15051), .Z(
        n15046) );
  NAND2_X1 U15019 ( .A1(n15051), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12726) );
  NOR2_X1 U15020 ( .A1(n12749), .A2(n12727), .ZN(n12728) );
  INV_X1 U15021 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15066) );
  INV_X1 U15022 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12729) );
  OR2_X1 U15023 ( .A1(n12751), .A2(n12729), .ZN(n12754) );
  NAND2_X1 U15024 ( .A1(n12751), .A2(n12729), .ZN(n12730) );
  NAND2_X1 U15025 ( .A1(n12754), .A2(n12730), .ZN(n15083) );
  XNOR2_X1 U15026 ( .A(n14470), .B(n12732), .ZN(n14463) );
  AND2_X1 U15027 ( .A1(n14470), .A2(n12732), .ZN(n12733) );
  NAND2_X1 U15028 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12772), .ZN(n12734) );
  OAI21_X1 U15029 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12772), .A(n12734), 
        .ZN(n14491) );
  INV_X1 U15030 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n15481) );
  INV_X1 U15031 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U15032 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14511), .B1(n12770), 
        .B2(n12738), .ZN(n14521) );
  XOR2_X1 U15033 ( .A(n12737), .B(n12736), .Z(n12792) );
  XNOR2_X1 U15034 ( .A(n12769), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12788) );
  MUX2_X1 U15035 ( .A(n12737), .B(n12788), .S(n12758), .Z(n12766) );
  INV_X1 U15036 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13050) );
  MUX2_X1 U15037 ( .A(n12738), .B(n13050), .S(n12758), .Z(n14516) );
  MUX2_X1 U15038 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12758), .Z(n12761) );
  AND2_X1 U15039 ( .A1(n12761), .A2(n12785), .ZN(n12762) );
  MUX2_X1 U15040 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12758), .Z(n12739) );
  AND2_X1 U15041 ( .A1(n12739), .A2(n12772), .ZN(n14481) );
  MUX2_X1 U15042 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12758), .Z(n12747) );
  INV_X1 U15043 ( .A(n12747), .ZN(n12748) );
  INV_X1 U15044 ( .A(n15051), .ZN(n12778) );
  MUX2_X1 U15045 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12758), .Z(n12745) );
  INV_X1 U15046 ( .A(n12745), .ZN(n12746) );
  MUX2_X1 U15047 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12758), .Z(n12743) );
  INV_X1 U15048 ( .A(n12743), .ZN(n12744) );
  INV_X1 U15049 ( .A(n12740), .ZN(n12742) );
  XNOR2_X1 U15050 ( .A(n12743), .B(n15031), .ZN(n15037) );
  XNOR2_X1 U15051 ( .A(n12745), .B(n12778), .ZN(n15059) );
  OAI21_X1 U15052 ( .B1(n12778), .B2(n12746), .A(n15058), .ZN(n15075) );
  XNOR2_X1 U15053 ( .A(n12747), .B(n15071), .ZN(n15076) );
  NOR2_X1 U15054 ( .A1(n15075), .A2(n15076), .ZN(n15074) );
  INV_X1 U15055 ( .A(n15083), .ZN(n12753) );
  INV_X1 U15056 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12750) );
  OR2_X1 U15057 ( .A1(n12751), .A2(n12750), .ZN(n12781) );
  NAND2_X1 U15058 ( .A1(n12751), .A2(n12750), .ZN(n12752) );
  AND2_X1 U15059 ( .A1(n12781), .A2(n12752), .ZN(n15085) );
  MUX2_X1 U15060 ( .A(n12753), .B(n15085), .S(n12758), .Z(n15098) );
  MUX2_X1 U15061 ( .A(n12754), .B(n12781), .S(n12758), .Z(n12755) );
  AOI21_X1 U15062 ( .B1(n14470), .B2(n12756), .A(n12757), .ZN(n14474) );
  INV_X1 U15063 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13063) );
  MUX2_X1 U15064 ( .A(n14464), .B(n13063), .S(n12758), .Z(n14473) );
  AND2_X1 U15065 ( .A1(n14474), .A2(n14473), .ZN(n14476) );
  NOR2_X1 U15066 ( .A1(n12757), .A2(n14476), .ZN(n14485) );
  INV_X1 U15067 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12771) );
  MUX2_X1 U15068 ( .A(n6859), .B(n12771), .S(n12758), .Z(n12759) );
  NAND2_X1 U15069 ( .A1(n12759), .A2(n14480), .ZN(n14483) );
  INV_X1 U15070 ( .A(n12762), .ZN(n12760) );
  OAI21_X1 U15071 ( .B1(n12761), .B2(n12785), .A(n12760), .ZN(n14501) );
  NAND2_X1 U15072 ( .A1(n14516), .A2(n14517), .ZN(n14515) );
  NAND2_X1 U15073 ( .A1(n14511), .A2(n12763), .ZN(n12764) );
  NAND2_X1 U15074 ( .A1(n14515), .A2(n12764), .ZN(n12765) );
  XOR2_X1 U15075 ( .A(n12766), .B(n12765), .Z(n12790) );
  NAND2_X1 U15076 ( .A1(n15095), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12767) );
  OAI211_X1 U15077 ( .C1(n15092), .C2(n12769), .A(n12768), .B(n12767), .ZN(
        n12789) );
  AOI22_X1 U15078 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12770), .B1(n14511), 
        .B2(n13050), .ZN(n14514) );
  NAND2_X1 U15079 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12772), .ZN(n12784) );
  AOI22_X1 U15080 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12772), .B1(n14480), 
        .B2(n12771), .ZN(n14488) );
  INV_X1 U15081 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n15434) );
  OAI21_X1 U15082 ( .B1(n12774), .B2(n15499), .A(n12773), .ZN(n12776) );
  NAND2_X1 U15083 ( .A1(n15031), .A2(n12776), .ZN(n12777) );
  XNOR2_X1 U15084 ( .A(n12776), .B(n12775), .ZN(n15030) );
  NAND2_X1 U15085 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15030), .ZN(n15029) );
  MUX2_X1 U15086 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n15434), .S(n15051), .Z(
        n15049) );
  NAND2_X1 U15087 ( .A1(n15071), .A2(n12779), .ZN(n12780) );
  NAND2_X1 U15088 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n15068), .ZN(n15067) );
  NAND2_X1 U15089 ( .A1(n14470), .A2(n12782), .ZN(n12783) );
  NAND2_X1 U15090 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14466), .ZN(n14465) );
  NAND2_X1 U15091 ( .A1(n12783), .A2(n14465), .ZN(n14487) );
  NAND2_X1 U15092 ( .A1(n14488), .A2(n14487), .ZN(n14486) );
  NAND2_X1 U15093 ( .A1(n12784), .A2(n14486), .ZN(n12786) );
  NAND2_X1 U15094 ( .A1(n12785), .A2(n12786), .ZN(n12787) );
  XNOR2_X1 U15095 ( .A(n14497), .B(n12786), .ZN(n14499) );
  NAND2_X1 U15096 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14499), .ZN(n14498) );
  NAND2_X1 U15097 ( .A1(n12787), .A2(n14498), .ZN(n14513) );
  NAND2_X1 U15098 ( .A1(n14514), .A2(n14513), .ZN(n14512) );
  OAI21_X1 U15099 ( .B1(n12792), .B2(n15102), .A(n12791), .ZN(P3_U3201) );
  AOI21_X1 U15100 ( .B1(n14531), .B2(n15144), .A(n12795), .ZN(n14530) );
  NAND2_X1 U15101 ( .A1(n15146), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12796) );
  OAI211_X1 U15102 ( .C1(n13076), .C2(n12998), .A(n14530), .B(n12796), .ZN(
        P3_U3202) );
  INV_X1 U15103 ( .A(n12797), .ZN(n12798) );
  NOR2_X1 U15104 ( .A1(n12814), .A2(n12798), .ZN(n12799) );
  XNOR2_X1 U15105 ( .A(n12799), .B(n12800), .ZN(n13006) );
  AOI21_X1 U15106 ( .B1(n12801), .B2(n12800), .A(n15132), .ZN(n12806) );
  OAI22_X1 U15107 ( .A1(n12803), .A2(n15136), .B1(n12802), .B2(n15134), .ZN(
        n12804) );
  AOI21_X1 U15108 ( .B1(n12806), .B2(n12805), .A(n12804), .ZN(n13005) );
  INV_X1 U15109 ( .A(n13005), .ZN(n12810) );
  AOI22_X1 U15110 ( .A1(n12807), .A2(n15140), .B1(n15146), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12808) );
  OAI21_X1 U15111 ( .B1(n13080), .B2(n12998), .A(n12808), .ZN(n12809) );
  AOI21_X1 U15112 ( .B1(n12810), .B2(n15144), .A(n12809), .ZN(n12811) );
  OAI21_X1 U15113 ( .B1(n13002), .B2(n13006), .A(n12811), .ZN(P3_U3205) );
  AND2_X1 U15114 ( .A1(n12812), .A2(n12816), .ZN(n12813) );
  OR2_X2 U15115 ( .A1(n12814), .A2(n12813), .ZN(n13010) );
  INV_X1 U15116 ( .A(n13010), .ZN(n12821) );
  OAI21_X1 U15117 ( .B1(n12817), .B2(n12816), .A(n12815), .ZN(n12819) );
  AOI21_X1 U15118 ( .B1(n12819), .B2(n12987), .A(n12818), .ZN(n12820) );
  OAI21_X1 U15119 ( .B1(n12868), .B2(n12821), .A(n12820), .ZN(n13009) );
  NAND2_X1 U15120 ( .A1(n13010), .A2(n12874), .ZN(n12825) );
  AOI22_X1 U15121 ( .A1(n12823), .A2(n15140), .B1(n15146), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12824) );
  OAI211_X1 U15122 ( .C1(n8131), .C2(n12998), .A(n12825), .B(n12824), .ZN(
        n12826) );
  AOI21_X1 U15123 ( .B1(n13009), .B2(n15144), .A(n12826), .ZN(n12827) );
  INV_X1 U15124 ( .A(n12827), .ZN(P3_U3206) );
  XNOR2_X1 U15125 ( .A(n12828), .B(n12832), .ZN(n12830) );
  OAI21_X1 U15126 ( .B1(n12830), .B2(n15132), .A(n12829), .ZN(n13013) );
  INV_X1 U15127 ( .A(n13013), .ZN(n12837) );
  XOR2_X1 U15128 ( .A(n12832), .B(n12831), .Z(n13014) );
  AOI22_X1 U15129 ( .A1(n12833), .A2(n15140), .B1(n15146), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12834) );
  OAI21_X1 U15130 ( .B1(n13087), .B2(n12998), .A(n12834), .ZN(n12835) );
  AOI21_X1 U15131 ( .B1(n13014), .B2(n15141), .A(n12835), .ZN(n12836) );
  OAI21_X1 U15132 ( .B1(n12837), .B2(n15146), .A(n12836), .ZN(P3_U3207) );
  XNOR2_X1 U15133 ( .A(n12838), .B(n12840), .ZN(n13017) );
  OAI211_X1 U15134 ( .C1(n12841), .C2(n12840), .A(n12839), .B(n12987), .ZN(
        n12843) );
  OAI211_X1 U15135 ( .C1(n12868), .C2(n13017), .A(n12843), .B(n12842), .ZN(
        n13018) );
  AOI22_X1 U15136 ( .A1(n12844), .A2(n15140), .B1(n15146), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12847) );
  NAND2_X1 U15137 ( .A1(n12845), .A2(n14528), .ZN(n12846) );
  OAI211_X1 U15138 ( .C1(n13017), .C2(n12848), .A(n12847), .B(n12846), .ZN(
        n12849) );
  AOI21_X1 U15139 ( .B1(n13018), .B2(n15144), .A(n12849), .ZN(n12850) );
  INV_X1 U15140 ( .A(n12850), .ZN(P3_U3208) );
  XNOR2_X1 U15141 ( .A(n12851), .B(n12854), .ZN(n12853) );
  AOI21_X1 U15142 ( .B1(n12853), .B2(n12987), .A(n12852), .ZN(n13023) );
  AOI21_X1 U15143 ( .B1(n12855), .B2(n12854), .A(n6731), .ZN(n13024) );
  INV_X1 U15144 ( .A(n13024), .ZN(n12860) );
  AOI22_X1 U15145 ( .A1(n15146), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15140), 
        .B2(n12856), .ZN(n12857) );
  OAI21_X1 U15146 ( .B1(n12858), .B2(n12998), .A(n12857), .ZN(n12859) );
  AOI21_X1 U15147 ( .B1(n12860), .B2(n15141), .A(n12859), .ZN(n12861) );
  OAI21_X1 U15148 ( .B1(n13023), .B2(n15146), .A(n12861), .ZN(P3_U3209) );
  XNOR2_X1 U15149 ( .A(n12862), .B(n12863), .ZN(n12870) );
  OR2_X1 U15150 ( .A1(n12864), .A2(n12863), .ZN(n12865) );
  NAND2_X1 U15151 ( .A1(n12866), .A2(n12865), .ZN(n13025) );
  OAI21_X1 U15152 ( .B1(n13025), .B2(n12868), .A(n12867), .ZN(n12869) );
  AOI21_X1 U15153 ( .B1(n12870), .B2(n12987), .A(n12869), .ZN(n13027) );
  INV_X1 U15154 ( .A(n13025), .ZN(n12875) );
  AOI22_X1 U15155 ( .A1(n15146), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15140), 
        .B2(n12871), .ZN(n12872) );
  OAI21_X1 U15156 ( .B1(n13096), .B2(n12998), .A(n12872), .ZN(n12873) );
  AOI21_X1 U15157 ( .B1(n12875), .B2(n12874), .A(n12873), .ZN(n12876) );
  OAI21_X1 U15158 ( .B1(n13027), .B2(n15146), .A(n12876), .ZN(P3_U3210) );
  XNOR2_X1 U15159 ( .A(n12877), .B(n12881), .ZN(n12879) );
  OAI21_X1 U15160 ( .B1(n12879), .B2(n15132), .A(n12878), .ZN(n13030) );
  INV_X1 U15161 ( .A(n13030), .ZN(n12886) );
  XOR2_X1 U15162 ( .A(n12881), .B(n12880), .Z(n13031) );
  AOI22_X1 U15163 ( .A1(n15146), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15140), 
        .B2(n12882), .ZN(n12883) );
  OAI21_X1 U15164 ( .B1(n13100), .B2(n12998), .A(n12883), .ZN(n12884) );
  AOI21_X1 U15165 ( .B1(n13031), .B2(n15141), .A(n12884), .ZN(n12885) );
  OAI21_X1 U15166 ( .B1(n12886), .B2(n15146), .A(n12885), .ZN(P3_U3211) );
  XNOR2_X1 U15167 ( .A(n12887), .B(n12890), .ZN(n12889) );
  OAI21_X1 U15168 ( .B1(n12889), .B2(n15132), .A(n12888), .ZN(n13034) );
  INV_X1 U15169 ( .A(n13034), .ZN(n12896) );
  XNOR2_X1 U15170 ( .A(n12891), .B(n12890), .ZN(n13035) );
  AOI22_X1 U15171 ( .A1(n15146), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15140), 
        .B2(n12892), .ZN(n12893) );
  OAI21_X1 U15172 ( .B1(n13104), .B2(n12998), .A(n12893), .ZN(n12894) );
  AOI21_X1 U15173 ( .B1(n13035), .B2(n15141), .A(n12894), .ZN(n12895) );
  OAI21_X1 U15174 ( .B1(n12896), .B2(n15146), .A(n12895), .ZN(P3_U3212) );
  XNOR2_X1 U15175 ( .A(n12897), .B(n8004), .ZN(n12900) );
  AOI222_X1 U15176 ( .A1(n12987), .A2(n12900), .B1(n12899), .B2(n12993), .C1(
        n12898), .C2(n12990), .ZN(n13041) );
  INV_X1 U15177 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12903) );
  INV_X1 U15178 ( .A(n12901), .ZN(n12902) );
  OAI22_X1 U15179 ( .A1(n15144), .A2(n12903), .B1(n12902), .B2(n15108), .ZN(
        n12904) );
  AOI21_X1 U15180 ( .B1(n12905), .B2(n14528), .A(n12904), .ZN(n12909) );
  NAND2_X1 U15181 ( .A1(n12907), .A2(n12906), .ZN(n13038) );
  NAND3_X1 U15182 ( .A1(n13039), .A2(n13038), .A3(n15141), .ZN(n12908) );
  OAI211_X1 U15183 ( .C1(n13041), .C2(n15146), .A(n12909), .B(n12908), .ZN(
        P3_U3213) );
  NAND2_X1 U15184 ( .A1(n12911), .A2(n12910), .ZN(n12979) );
  NAND2_X1 U15185 ( .A1(n12979), .A2(n12912), .ZN(n12914) );
  AND2_X1 U15186 ( .A1(n12914), .A2(n12913), .ZN(n12915) );
  XNOR2_X1 U15187 ( .A(n12915), .B(n12917), .ZN(n13045) );
  INV_X1 U15188 ( .A(n13045), .ZN(n12926) );
  OAI211_X1 U15189 ( .C1(n6808), .C2(n12917), .A(n12916), .B(n12987), .ZN(
        n12920) );
  OR2_X1 U15190 ( .A1(n12918), .A2(n15134), .ZN(n12919) );
  OAI211_X1 U15191 ( .C1(n12921), .C2(n15136), .A(n12920), .B(n12919), .ZN(
        n13044) );
  AOI22_X1 U15192 ( .A1(n15146), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15140), 
        .B2(n12922), .ZN(n12923) );
  OAI21_X1 U15193 ( .B1(n13112), .B2(n12998), .A(n12923), .ZN(n12924) );
  AOI21_X1 U15194 ( .B1(n13044), .B2(n15144), .A(n12924), .ZN(n12925) );
  OAI21_X1 U15195 ( .B1(n13002), .B2(n12926), .A(n12925), .ZN(P3_U3214) );
  AOI21_X1 U15196 ( .B1(n12936), .B2(n12928), .A(n12927), .ZN(n12929) );
  OAI222_X1 U15197 ( .A1(n15136), .A2(n12931), .B1(n15134), .B2(n12930), .C1(
        n15132), .C2(n12929), .ZN(n13048) );
  INV_X1 U15198 ( .A(n13048), .ZN(n12944) );
  NAND2_X1 U15199 ( .A1(n12979), .A2(n12932), .ZN(n12935) );
  AND2_X1 U15200 ( .A1(n12935), .A2(n12933), .ZN(n12939) );
  AND2_X1 U15201 ( .A1(n12935), .A2(n12934), .ZN(n12952) );
  AOI21_X1 U15202 ( .B1(n12952), .B2(n12937), .A(n12936), .ZN(n12938) );
  NOR2_X1 U15203 ( .A1(n12939), .A2(n12938), .ZN(n13049) );
  AOI22_X1 U15204 ( .A1(n15146), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15140), 
        .B2(n12940), .ZN(n12941) );
  OAI21_X1 U15205 ( .B1(n13116), .B2(n12998), .A(n12941), .ZN(n12942) );
  AOI21_X1 U15206 ( .B1(n13049), .B2(n15141), .A(n12942), .ZN(n12943) );
  OAI21_X1 U15207 ( .B1(n12944), .B2(n15146), .A(n12943), .ZN(P3_U3215) );
  XNOR2_X1 U15208 ( .A(n12945), .B(n12953), .ZN(n12948) );
  AOI222_X1 U15209 ( .A1(n12987), .A2(n12948), .B1(n12947), .B2(n12990), .C1(
        n12946), .C2(n12993), .ZN(n13055) );
  NAND2_X1 U15210 ( .A1(n12979), .A2(n12949), .ZN(n12951) );
  NAND2_X1 U15211 ( .A1(n12951), .A2(n12950), .ZN(n12954) );
  OAI21_X1 U15212 ( .B1(n12954), .B2(n12953), .A(n12952), .ZN(n13053) );
  AOI22_X1 U15213 ( .A1(n15146), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15140), 
        .B2(n12955), .ZN(n12956) );
  OAI21_X1 U15214 ( .B1(n12957), .B2(n12998), .A(n12956), .ZN(n12958) );
  AOI21_X1 U15215 ( .B1(n13053), .B2(n15141), .A(n12958), .ZN(n12959) );
  OAI21_X1 U15216 ( .B1(n13055), .B2(n15146), .A(n12959), .ZN(P3_U3216) );
  INV_X1 U15217 ( .A(n12965), .ZN(n12960) );
  XNOR2_X1 U15218 ( .A(n12961), .B(n12960), .ZN(n12963) );
  AOI21_X1 U15219 ( .B1(n12963), .B2(n12987), .A(n12962), .ZN(n13058) );
  NAND2_X1 U15220 ( .A1(n12979), .A2(n12978), .ZN(n12977) );
  NAND2_X1 U15221 ( .A1(n12977), .A2(n12964), .ZN(n12966) );
  NAND2_X1 U15222 ( .A1(n12966), .A2(n12965), .ZN(n12968) );
  OR2_X1 U15223 ( .A1(n12966), .A2(n12965), .ZN(n12967) );
  NAND2_X1 U15224 ( .A1(n12968), .A2(n12967), .ZN(n13056) );
  AOI22_X1 U15225 ( .A1(n15146), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15140), 
        .B2(n12969), .ZN(n12970) );
  OAI21_X1 U15226 ( .B1(n13121), .B2(n12998), .A(n12970), .ZN(n12971) );
  AOI21_X1 U15227 ( .B1(n13056), .B2(n15141), .A(n12971), .ZN(n12972) );
  OAI21_X1 U15228 ( .B1(n13058), .B2(n15146), .A(n12972), .ZN(P3_U3217) );
  NAND2_X1 U15229 ( .A1(n6786), .A2(n12973), .ZN(n12974) );
  XOR2_X1 U15230 ( .A(n12978), .B(n12974), .Z(n12976) );
  OAI21_X1 U15231 ( .B1(n12976), .B2(n15132), .A(n12975), .ZN(n13061) );
  INV_X1 U15232 ( .A(n13061), .ZN(n12984) );
  OAI21_X1 U15233 ( .B1(n12979), .B2(n12978), .A(n12977), .ZN(n13062) );
  AOI22_X1 U15234 ( .A1(n15146), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15140), 
        .B2(n12980), .ZN(n12981) );
  OAI21_X1 U15235 ( .B1(n13125), .B2(n12998), .A(n12981), .ZN(n12982) );
  AOI21_X1 U15236 ( .B1(n13062), .B2(n15141), .A(n12982), .ZN(n12983) );
  OAI21_X1 U15237 ( .B1(n12984), .B2(n15146), .A(n12983), .ZN(P3_U3218) );
  XNOR2_X1 U15238 ( .A(n12986), .B(n12985), .ZN(n13068) );
  OAI211_X1 U15239 ( .C1(n12989), .C2(n12988), .A(n6786), .B(n12987), .ZN(
        n12995) );
  AOI22_X1 U15240 ( .A1(n12993), .A2(n12992), .B1(n12991), .B2(n12990), .ZN(
        n12994) );
  NAND2_X1 U15241 ( .A1(n12995), .A2(n12994), .ZN(n13065) );
  INV_X1 U15242 ( .A(n13066), .ZN(n12999) );
  AOI22_X1 U15243 ( .A1(n15146), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15140), 
        .B2(n12996), .ZN(n12997) );
  OAI21_X1 U15244 ( .B1(n12999), .B2(n12998), .A(n12997), .ZN(n13000) );
  AOI21_X1 U15245 ( .B1(n13065), .B2(n15144), .A(n13000), .ZN(n13001) );
  OAI21_X1 U15246 ( .B1(n13002), .B2(n13068), .A(n13001), .ZN(P3_U3219) );
  NAND2_X1 U15247 ( .A1(n15210), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13004) );
  NAND2_X1 U15248 ( .A1(n14531), .A2(n15213), .ZN(n13003) );
  OAI211_X1 U15249 ( .C1(n13076), .C2(n13073), .A(n13004), .B(n13003), .ZN(
        P3_U3490) );
  MUX2_X1 U15250 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13077), .S(n15213), .Z(
        n13007) );
  INV_X1 U15251 ( .A(n13007), .ZN(n13008) );
  OAI21_X1 U15252 ( .B1(n13080), .B2(n13073), .A(n13008), .ZN(P3_U3487) );
  INV_X1 U15253 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13011) );
  INV_X1 U15254 ( .A(n15189), .ZN(n15156) );
  AOI21_X1 U15255 ( .B1(n15156), .B2(n13010), .A(n13009), .ZN(n13081) );
  MUX2_X1 U15256 ( .A(n13011), .B(n13081), .S(n15213), .Z(n13012) );
  OAI21_X1 U15257 ( .B1(n8131), .B2(n13073), .A(n13012), .ZN(P3_U3486) );
  INV_X1 U15258 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13015) );
  AOI21_X1 U15259 ( .B1(n13014), .B2(n15187), .A(n13013), .ZN(n13084) );
  MUX2_X1 U15260 ( .A(n13015), .B(n13084), .S(n15213), .Z(n13016) );
  OAI21_X1 U15261 ( .B1(n13087), .B2(n13073), .A(n13016), .ZN(P3_U3485) );
  INV_X1 U15262 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n15417) );
  INV_X1 U15263 ( .A(n13017), .ZN(n13019) );
  AOI21_X1 U15264 ( .B1(n15156), .B2(n13019), .A(n13018), .ZN(n13088) );
  MUX2_X1 U15265 ( .A(n15417), .B(n13088), .S(n15213), .Z(n13020) );
  OAI21_X1 U15266 ( .B1(n13091), .B2(n13073), .A(n13020), .ZN(P3_U3484) );
  NAND2_X1 U15267 ( .A1(n13021), .A2(n15193), .ZN(n13022) );
  OAI211_X1 U15268 ( .C1(n15172), .C2(n13024), .A(n13023), .B(n13022), .ZN(
        n13092) );
  MUX2_X1 U15269 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13092), .S(n15213), .Z(
        P3_U3483) );
  INV_X1 U15270 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13028) );
  OR2_X1 U15271 ( .A1(n13025), .A2(n15189), .ZN(n13026) );
  AND2_X1 U15272 ( .A1(n13027), .A2(n13026), .ZN(n13093) );
  MUX2_X1 U15273 ( .A(n13028), .B(n13093), .S(n15213), .Z(n13029) );
  OAI21_X1 U15274 ( .B1(n13096), .B2(n13073), .A(n13029), .ZN(P3_U3482) );
  INV_X1 U15275 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13032) );
  AOI21_X1 U15276 ( .B1(n15187), .B2(n13031), .A(n13030), .ZN(n13097) );
  MUX2_X1 U15277 ( .A(n13032), .B(n13097), .S(n15213), .Z(n13033) );
  OAI21_X1 U15278 ( .B1(n13100), .B2(n13073), .A(n13033), .ZN(P3_U3481) );
  INV_X1 U15279 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13036) );
  AOI21_X1 U15280 ( .B1(n13035), .B2(n15187), .A(n13034), .ZN(n13101) );
  MUX2_X1 U15281 ( .A(n13036), .B(n13101), .S(n15213), .Z(n13037) );
  OAI21_X1 U15282 ( .B1(n13104), .B2(n13073), .A(n13037), .ZN(P3_U3480) );
  INV_X1 U15283 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13042) );
  NAND3_X1 U15284 ( .A1(n13039), .A2(n13038), .A3(n15187), .ZN(n13040) );
  AND2_X1 U15285 ( .A1(n13041), .A2(n13040), .ZN(n13105) );
  MUX2_X1 U15286 ( .A(n13042), .B(n13105), .S(n15213), .Z(n13043) );
  OAI21_X1 U15287 ( .B1(n13108), .B2(n13073), .A(n13043), .ZN(P3_U3479) );
  INV_X1 U15288 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13046) );
  AOI21_X1 U15289 ( .B1(n15187), .B2(n13045), .A(n13044), .ZN(n13109) );
  MUX2_X1 U15290 ( .A(n13046), .B(n13109), .S(n15213), .Z(n13047) );
  OAI21_X1 U15291 ( .B1(n13073), .B2(n13112), .A(n13047), .ZN(P3_U3478) );
  AOI21_X1 U15292 ( .B1(n13049), .B2(n15187), .A(n13048), .ZN(n13113) );
  MUX2_X1 U15293 ( .A(n13050), .B(n13113), .S(n15213), .Z(n13051) );
  OAI21_X1 U15294 ( .B1(n13116), .B2(n13073), .A(n13051), .ZN(P3_U3477) );
  AOI22_X1 U15295 ( .A1(n13053), .A2(n15187), .B1(n15193), .B2(n13052), .ZN(
        n13054) );
  NAND2_X1 U15296 ( .A1(n13055), .A2(n13054), .ZN(n13117) );
  MUX2_X1 U15297 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13117), .S(n15213), .Z(
        P3_U3476) );
  NAND2_X1 U15298 ( .A1(n13056), .A2(n15187), .ZN(n13057) );
  NAND2_X1 U15299 ( .A1(n13058), .A2(n13057), .ZN(n13118) );
  MUX2_X1 U15300 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13118), .S(n15213), .Z(
        n13059) );
  INV_X1 U15301 ( .A(n13059), .ZN(n13060) );
  OAI21_X1 U15302 ( .B1(n13121), .B2(n13073), .A(n13060), .ZN(P3_U3475) );
  AOI21_X1 U15303 ( .B1(n15187), .B2(n13062), .A(n13061), .ZN(n13122) );
  MUX2_X1 U15304 ( .A(n13063), .B(n13122), .S(n15213), .Z(n13064) );
  OAI21_X1 U15305 ( .B1(n13125), .B2(n13073), .A(n13064), .ZN(P3_U3474) );
  AOI21_X1 U15306 ( .B1(n15193), .B2(n13066), .A(n13065), .ZN(n13067) );
  OAI21_X1 U15307 ( .B1(n15172), .B2(n13068), .A(n13067), .ZN(n13126) );
  MUX2_X1 U15308 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n13126), .S(n15213), .Z(
        P3_U3473) );
  INV_X1 U15309 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13071) );
  AOI21_X1 U15310 ( .B1(n13070), .B2(n15187), .A(n13069), .ZN(n13127) );
  MUX2_X1 U15311 ( .A(n13071), .B(n13127), .S(n15213), .Z(n13072) );
  OAI21_X1 U15312 ( .B1(n13073), .B2(n13130), .A(n13072), .ZN(P3_U3472) );
  INV_X1 U15313 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n15449) );
  NOR2_X1 U15314 ( .A1(n15197), .A2(n15449), .ZN(n13074) );
  AOI21_X1 U15315 ( .B1(n14531), .B2(n15197), .A(n13074), .ZN(n13075) );
  OAI21_X1 U15316 ( .B1(n13076), .B2(n13131), .A(n13075), .ZN(P3_U3458) );
  INV_X1 U15317 ( .A(n13077), .ZN(n13078) );
  OAI21_X1 U15318 ( .B1(n13080), .B2(n13131), .A(n13079), .ZN(P3_U3455) );
  MUX2_X1 U15319 ( .A(n13082), .B(n13081), .S(n15197), .Z(n13083) );
  OAI21_X1 U15320 ( .B1(n8131), .B2(n13131), .A(n13083), .ZN(P3_U3454) );
  MUX2_X1 U15321 ( .A(n13085), .B(n13084), .S(n15197), .Z(n13086) );
  OAI21_X1 U15322 ( .B1(n13087), .B2(n13131), .A(n13086), .ZN(P3_U3453) );
  INV_X1 U15323 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13089) );
  MUX2_X1 U15324 ( .A(n13089), .B(n13088), .S(n15197), .Z(n13090) );
  OAI21_X1 U15325 ( .B1(n13091), .B2(n13131), .A(n13090), .ZN(P3_U3452) );
  MUX2_X1 U15326 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13092), .S(n15197), .Z(
        P3_U3451) );
  INV_X1 U15327 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13094) );
  MUX2_X1 U15328 ( .A(n13094), .B(n13093), .S(n15197), .Z(n13095) );
  OAI21_X1 U15329 ( .B1(n13096), .B2(n13131), .A(n13095), .ZN(P3_U3450) );
  INV_X1 U15330 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13098) );
  MUX2_X1 U15331 ( .A(n13098), .B(n13097), .S(n15197), .Z(n13099) );
  OAI21_X1 U15332 ( .B1(n13100), .B2(n13131), .A(n13099), .ZN(P3_U3449) );
  INV_X1 U15333 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13102) );
  MUX2_X1 U15334 ( .A(n13102), .B(n13101), .S(n15197), .Z(n13103) );
  OAI21_X1 U15335 ( .B1(n13104), .B2(n13131), .A(n13103), .ZN(P3_U3448) );
  INV_X1 U15336 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13106) );
  MUX2_X1 U15337 ( .A(n13106), .B(n13105), .S(n15197), .Z(n13107) );
  OAI21_X1 U15338 ( .B1(n13108), .B2(n13131), .A(n13107), .ZN(P3_U3447) );
  INV_X1 U15339 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13110) );
  MUX2_X1 U15340 ( .A(n13110), .B(n13109), .S(n15197), .Z(n13111) );
  OAI21_X1 U15341 ( .B1(n13131), .B2(n13112), .A(n13111), .ZN(P3_U3446) );
  INV_X1 U15342 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13114) );
  MUX2_X1 U15343 ( .A(n13114), .B(n13113), .S(n15197), .Z(n13115) );
  OAI21_X1 U15344 ( .B1(n13116), .B2(n13131), .A(n13115), .ZN(P3_U3444) );
  MUX2_X1 U15345 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13117), .S(n15197), .Z(
        P3_U3441) );
  MUX2_X1 U15346 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13118), .S(n15197), .Z(
        n13119) );
  INV_X1 U15347 ( .A(n13119), .ZN(n13120) );
  OAI21_X1 U15348 ( .B1(n13121), .B2(n13131), .A(n13120), .ZN(P3_U3438) );
  INV_X1 U15349 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13123) );
  MUX2_X1 U15350 ( .A(n13123), .B(n13122), .S(n15197), .Z(n13124) );
  OAI21_X1 U15351 ( .B1(n13125), .B2(n13131), .A(n13124), .ZN(P3_U3435) );
  MUX2_X1 U15352 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n13126), .S(n15197), .Z(
        P3_U3432) );
  INV_X1 U15353 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13128) );
  MUX2_X1 U15354 ( .A(n13128), .B(n13127), .S(n15197), .Z(n13129) );
  OAI21_X1 U15355 ( .B1(n13131), .B2(n13130), .A(n13129), .ZN(P3_U3429) );
  MUX2_X1 U15356 ( .A(n13132), .B(P3_D_REG_1__SCAN_IN), .S(n13133), .Z(
        P3_U3377) );
  MUX2_X1 U15357 ( .A(n13134), .B(P3_D_REG_0__SCAN_IN), .S(n13133), .Z(
        P3_U3376) );
  NAND2_X1 U15358 ( .A1(n13136), .A2(n13135), .ZN(n13140) );
  OR4_X1 U15359 ( .A1(n13138), .A2(P3_IR_REG_30__SCAN_IN), .A3(n13137), .A4(
        P3_U3151), .ZN(n13139) );
  OAI211_X1 U15360 ( .C1(n13141), .C2(n12350), .A(n13140), .B(n13139), .ZN(
        P3_U3264) );
  OAI222_X1 U15361 ( .A1(P3_U3151), .A2(n13144), .B1(n11060), .B2(n13143), 
        .C1(n13142), .C2(n12350), .ZN(P3_U3266) );
  MUX2_X1 U15362 ( .A(n13145), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AOI21_X1 U15363 ( .B1(n13147), .B2(n13146), .A(n13275), .ZN(n13149) );
  NAND2_X1 U15364 ( .A1(n13149), .A2(n13148), .ZN(n13153) );
  AOI22_X1 U15365 ( .A1(n13650), .A2(n13279), .B1(n13423), .B2(n13470), .ZN(
        n13384) );
  OAI22_X1 U15366 ( .A1(n13217), .A2(n13384), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13150), .ZN(n13151) );
  AOI21_X1 U15367 ( .B1(n13391), .B2(n13219), .A(n13151), .ZN(n13152) );
  OAI211_X1 U15368 ( .C1(n13390), .C2(n13242), .A(n13153), .B(n13152), .ZN(
        P2_U3186) );
  OAI211_X1 U15369 ( .C1(n13154), .C2(n13156), .A(n13155), .B(n13249), .ZN(
        n13160) );
  AOI22_X1 U15370 ( .A1(n13244), .A2(n13282), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13159) );
  AOI22_X1 U15371 ( .A1(n13243), .A2(n13422), .B1(n13219), .B2(n13461), .ZN(
        n13158) );
  NAND2_X1 U15372 ( .A1(n13596), .A2(n13273), .ZN(n13157) );
  NAND4_X1 U15373 ( .A1(n13160), .A2(n13159), .A3(n13158), .A4(n13157), .ZN(
        P2_U3188) );
  OAI211_X1 U15374 ( .C1(n13163), .C2(n13162), .A(n13161), .B(n13249), .ZN(
        n13169) );
  AOI22_X1 U15375 ( .A1(n13244), .A2(n11346), .B1(n13243), .B2(n13299), .ZN(
        n13168) );
  AOI22_X1 U15376 ( .A1(n13273), .A2(n13164), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13167) );
  NAND2_X1 U15377 ( .A1(n13219), .A2(n13165), .ZN(n13166) );
  NAND4_X1 U15378 ( .A1(n13169), .A2(n13168), .A3(n13167), .A4(n13166), .ZN(
        P2_U3190) );
  OAI21_X1 U15379 ( .B1(n13172), .B2(n13171), .A(n13170), .ZN(n13173) );
  NAND2_X1 U15380 ( .A1(n13173), .A2(n13249), .ZN(n13178) );
  OAI22_X1 U15381 ( .A1(n13190), .A2(n13540), .B1(n13174), .B2(n13538), .ZN(
        n13520) );
  INV_X1 U15382 ( .A(n13520), .ZN(n13175) );
  NAND2_X1 U15383 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13352)
         );
  OAI21_X1 U15384 ( .B1(n13175), .B2(n13217), .A(n13352), .ZN(n13176) );
  AOI21_X1 U15385 ( .B1(n13526), .B2(n13219), .A(n13176), .ZN(n13177) );
  OAI211_X1 U15386 ( .C1(n13529), .C2(n13242), .A(n13178), .B(n13177), .ZN(
        P2_U3191) );
  AOI22_X1 U15387 ( .A1(n13244), .A2(n13302), .B1(n13243), .B2(n11346), .ZN(
        n13186) );
  AOI22_X1 U15388 ( .A1(n13273), .A2(n13179), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13245), .ZN(n13185) );
  OAI21_X1 U15389 ( .B1(n13182), .B2(n13181), .A(n13180), .ZN(n13183) );
  NAND2_X1 U15390 ( .A1(n13183), .A2(n13249), .ZN(n13184) );
  NAND3_X1 U15391 ( .A1(n13186), .A2(n13185), .A3(n13184), .ZN(P2_U3194) );
  OAI211_X1 U15392 ( .C1(n13189), .C2(n13188), .A(n13187), .B(n13249), .ZN(
        n13194) );
  OAI22_X1 U15393 ( .A1(n13451), .A2(n13540), .B1(n13190), .B2(n13538), .ZN(
        n13486) );
  AOI22_X1 U15394 ( .A1(n13486), .A2(n13268), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13191) );
  OAI21_X1 U15395 ( .B1(n13490), .B2(n13270), .A(n13191), .ZN(n13192) );
  AOI21_X1 U15396 ( .B1(n13606), .B2(n13273), .A(n13192), .ZN(n13193) );
  NAND2_X1 U15397 ( .A1(n13194), .A2(n13193), .ZN(P2_U3195) );
  OAI211_X1 U15398 ( .C1(n13195), .C2(n13197), .A(n13196), .B(n13249), .ZN(
        n13201) );
  AOI22_X1 U15399 ( .A1(n13244), .A2(n13422), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13200) );
  AOI22_X1 U15400 ( .A1(n13243), .A2(n13423), .B1(n13219), .B2(n13414), .ZN(
        n13199) );
  NAND2_X1 U15401 ( .A1(n13584), .A2(n13273), .ZN(n13198) );
  NAND4_X1 U15402 ( .A1(n13201), .A2(n13200), .A3(n13199), .A4(n13198), .ZN(
        P2_U3197) );
  NOR2_X1 U15403 ( .A1(n13203), .A2(n13202), .ZN(n13204) );
  OAI21_X1 U15404 ( .B1(n13205), .B2(n13204), .A(n13249), .ZN(n13211) );
  AOI22_X1 U15405 ( .A1(n13268), .A2(n13206), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13210) );
  NAND2_X1 U15406 ( .A1(n13627), .A2(n13273), .ZN(n13209) );
  NAND2_X1 U15407 ( .A1(n13219), .A2(n13207), .ZN(n13208) );
  NAND4_X1 U15408 ( .A1(n13211), .A2(n13210), .A3(n13209), .A4(n13208), .ZN(
        P2_U3200) );
  INV_X1 U15409 ( .A(n13588), .ZN(n13222) );
  OAI211_X1 U15410 ( .C1(n13212), .C2(n13214), .A(n13213), .B(n13249), .ZN(
        n13221) );
  NOR2_X1 U15411 ( .A1(n13267), .A2(n13540), .ZN(n13215) );
  AOI21_X1 U15412 ( .B1(n13469), .B2(n13470), .A(n13215), .ZN(n13433) );
  OAI22_X1 U15413 ( .A1(n13433), .A2(n13217), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13216), .ZN(n13218) );
  AOI21_X1 U15414 ( .B1(n13438), .B2(n13219), .A(n13218), .ZN(n13220) );
  OAI211_X1 U15415 ( .C1(n13222), .C2(n13242), .A(n13221), .B(n13220), .ZN(
        P2_U3201) );
  INV_X1 U15416 ( .A(n13223), .ZN(n13225) );
  NAND2_X1 U15417 ( .A1(n13225), .A2(n13224), .ZN(n13226) );
  XNOR2_X1 U15418 ( .A(n13227), .B(n13226), .ZN(n13232) );
  INV_X1 U15419 ( .A(n13509), .ZN(n13229) );
  OAI22_X1 U15420 ( .A1(n13236), .A2(n13540), .B1(n13541), .B2(n13538), .ZN(
        n13502) );
  AOI22_X1 U15421 ( .A1(n13502), .A2(n13268), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13228) );
  OAI21_X1 U15422 ( .B1(n13229), .B2(n13270), .A(n13228), .ZN(n13230) );
  AOI21_X1 U15423 ( .B1(n13611), .B2(n13273), .A(n13230), .ZN(n13231) );
  OAI21_X1 U15424 ( .B1(n13232), .B2(n13275), .A(n13231), .ZN(P2_U3205) );
  OAI211_X1 U15425 ( .C1(n13233), .C2(n13235), .A(n13234), .B(n13249), .ZN(
        n13241) );
  NOR2_X1 U15426 ( .A1(n13257), .A2(n13236), .ZN(n13239) );
  OAI22_X1 U15427 ( .A1(n13258), .A2(n13237), .B1(n13477), .B2(n13270), .ZN(
        n13238) );
  AOI211_X1 U15428 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3088), .A(n13239), 
        .B(n13238), .ZN(n13240) );
  OAI211_X1 U15429 ( .C1(n13481), .C2(n13242), .A(n13241), .B(n13240), .ZN(
        P2_U3207) );
  AOI22_X1 U15430 ( .A1(n13244), .A2(n11323), .B1(n13243), .B2(n13300), .ZN(
        n13254) );
  AOI22_X1 U15431 ( .A1(n13273), .A2(n13246), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n13245), .ZN(n13253) );
  AND3_X1 U15432 ( .A1(n13180), .A2(n13248), .A3(n13247), .ZN(n13250) );
  OAI21_X1 U15433 ( .B1(n13251), .B2(n13250), .A(n13249), .ZN(n13252) );
  NAND3_X1 U15434 ( .A1(n13254), .A2(n13253), .A3(n13252), .ZN(P2_U3209) );
  XNOR2_X1 U15435 ( .A(n13256), .B(n13255), .ZN(n13262) );
  NAND2_X1 U15436 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13323)
         );
  OAI21_X1 U15437 ( .B1(n13257), .B2(n13539), .A(n13323), .ZN(n13260) );
  OAI22_X1 U15438 ( .A1(n13258), .A2(n13541), .B1(n13270), .B2(n13546), .ZN(
        n13259) );
  AOI211_X1 U15439 ( .C1(n13553), .C2(n13273), .A(n13260), .B(n13259), .ZN(
        n13261) );
  OAI21_X1 U15440 ( .B1(n13262), .B2(n13275), .A(n13261), .ZN(P2_U3210) );
  INV_X1 U15441 ( .A(n13405), .ZN(n13271) );
  OAI22_X1 U15442 ( .A1(n13267), .A2(n13538), .B1(n13266), .B2(n13540), .ZN(
        n13398) );
  AOI22_X1 U15443 ( .A1(n13268), .A2(n13398), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13269) );
  OAI21_X1 U15444 ( .B1(n13271), .B2(n13270), .A(n13269), .ZN(n13272) );
  AOI21_X1 U15445 ( .B1(n13579), .B2(n13273), .A(n13272), .ZN(n13274) );
  OAI21_X1 U15446 ( .B1(n13276), .B2(n13275), .A(n13274), .ZN(P2_U3212) );
  MUX2_X1 U15447 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13354), .S(n13301), .Z(
        P2_U3562) );
  MUX2_X1 U15448 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13277), .S(n13301), .Z(
        P2_U3561) );
  MUX2_X1 U15449 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13278), .S(n13301), .Z(
        P2_U3560) );
  MUX2_X1 U15450 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13279), .S(n13301), .Z(
        P2_U3559) );
  MUX2_X1 U15451 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13280), .S(n13301), .Z(
        P2_U3558) );
  MUX2_X1 U15452 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13423), .S(n13301), .Z(
        P2_U3557) );
  MUX2_X1 U15453 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13281), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15454 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13422), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15455 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13469), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15456 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13282), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15457 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13471), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15458 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13283), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15459 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13284), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15460 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13285), .S(n13301), .Z(
        P2_U3549) );
  MUX2_X1 U15461 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13286), .S(n13301), .Z(
        P2_U3548) );
  MUX2_X1 U15462 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13287), .S(n13301), .Z(
        P2_U3547) );
  MUX2_X1 U15463 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13288), .S(n13301), .Z(
        P2_U3546) );
  MUX2_X1 U15464 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13289), .S(n13301), .Z(
        P2_U3545) );
  MUX2_X1 U15465 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13290), .S(n13301), .Z(
        P2_U3544) );
  MUX2_X1 U15466 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13291), .S(n13301), .Z(
        P2_U3543) );
  MUX2_X1 U15467 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13292), .S(n13301), .Z(
        P2_U3542) );
  MUX2_X1 U15468 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13293), .S(n13301), .Z(
        P2_U3541) );
  MUX2_X1 U15469 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13294), .S(n13301), .Z(
        P2_U3540) );
  MUX2_X1 U15470 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13295), .S(n13301), .Z(
        P2_U3539) );
  MUX2_X1 U15471 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13296), .S(n13301), .Z(
        P2_U3538) );
  MUX2_X1 U15472 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13297), .S(n13301), .Z(
        P2_U3537) );
  MUX2_X1 U15473 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13298), .S(n13301), .Z(
        P2_U3536) );
  MUX2_X1 U15474 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13299), .S(n13301), .Z(
        P2_U3535) );
  MUX2_X1 U15475 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13300), .S(n13301), .Z(
        P2_U3534) );
  MUX2_X1 U15476 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n11346), .S(n13301), .Z(
        P2_U3533) );
  MUX2_X1 U15477 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n11323), .S(n13301), .Z(
        P2_U3532) );
  MUX2_X1 U15478 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13302), .S(n13301), .Z(
        P2_U3531) );
  NOR2_X1 U15479 ( .A1(n13304), .A2(n13303), .ZN(n13306) );
  OAI21_X1 U15480 ( .B1(n13306), .B2(n13305), .A(n14843), .ZN(n13317) );
  INV_X1 U15481 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14622) );
  OAI21_X1 U15482 ( .B1(n14823), .B2(n14622), .A(n13307), .ZN(n13308) );
  AOI21_X1 U15483 ( .B1(n13309), .B2(n14841), .A(n13308), .ZN(n13316) );
  AND3_X1 U15484 ( .A1(n13312), .A2(n13311), .A3(n13310), .ZN(n13313) );
  OAI21_X1 U15485 ( .B1(n13314), .B2(n13313), .A(n14837), .ZN(n13315) );
  NAND3_X1 U15486 ( .A1(n13317), .A2(n13316), .A3(n13315), .ZN(P2_U3226) );
  NOR2_X1 U15487 ( .A1(n13328), .A2(n13318), .ZN(n13319) );
  AOI21_X1 U15488 ( .B1(n13318), .B2(n13328), .A(n13319), .ZN(n14838) );
  NAND2_X1 U15489 ( .A1(n13321), .A2(n13320), .ZN(n14839) );
  NAND2_X1 U15490 ( .A1(n14838), .A2(n14839), .ZN(n14836) );
  OAI21_X1 U15491 ( .B1(n13328), .B2(n13318), .A(n14836), .ZN(n13335) );
  XNOR2_X1 U15492 ( .A(n13340), .B(n13335), .ZN(n13322) );
  NOR2_X1 U15493 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13322), .ZN(n13337) );
  AOI21_X1 U15494 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13322), .A(n13337), 
        .ZN(n13334) );
  INV_X1 U15495 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n13324) );
  OAI21_X1 U15496 ( .B1(n14823), .B2(n13324), .A(n13323), .ZN(n13332) );
  INV_X1 U15497 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n15411) );
  XNOR2_X1 U15498 ( .A(n13328), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14845) );
  INV_X1 U15499 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13326) );
  OAI21_X1 U15500 ( .B1(n13327), .B2(n13326), .A(n13325), .ZN(n14844) );
  NAND2_X1 U15501 ( .A1(n14845), .A2(n14844), .ZN(n14842) );
  OAI21_X1 U15502 ( .B1(n13328), .B2(n15411), .A(n14842), .ZN(n13339) );
  XOR2_X1 U15503 ( .A(n13340), .B(n13339), .Z(n13329) );
  NAND2_X1 U15504 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n13329), .ZN(n13342) );
  OAI21_X1 U15505 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n13329), .A(n13342), 
        .ZN(n13330) );
  NOR2_X1 U15506 ( .A1(n13330), .A2(n14798), .ZN(n13331) );
  AOI211_X1 U15507 ( .C1(n14841), .C2(n13340), .A(n13332), .B(n13331), .ZN(
        n13333) );
  OAI21_X1 U15508 ( .B1(n13334), .B2(n14811), .A(n13333), .ZN(P2_U3232) );
  NOR2_X1 U15509 ( .A1(n13340), .A2(n13335), .ZN(n13336) );
  NOR2_X1 U15510 ( .A1(n13337), .A2(n13336), .ZN(n13338) );
  XOR2_X1 U15511 ( .A(n13338), .B(n11498), .Z(n13348) );
  INV_X1 U15512 ( .A(n13348), .ZN(n13346) );
  NAND2_X1 U15513 ( .A1(n13340), .A2(n13339), .ZN(n13341) );
  NAND2_X1 U15514 ( .A1(n13342), .A2(n13341), .ZN(n13344) );
  INV_X1 U15515 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13343) );
  XOR2_X1 U15516 ( .A(n13344), .B(n13343), .Z(n13347) );
  NAND2_X1 U15517 ( .A1(n13347), .A2(n14843), .ZN(n13345) );
  OAI211_X1 U15518 ( .C1(n13346), .C2(n14811), .A(n14765), .B(n13345), .ZN(
        n13351) );
  OAI22_X1 U15519 ( .A1(n13348), .A2(n14811), .B1(n13347), .B2(n14798), .ZN(
        n13350) );
  XNOR2_X1 U15520 ( .A(n13359), .B(n11698), .ZN(n13353) );
  NAND2_X1 U15521 ( .A1(n13353), .A2(n10936), .ZN(n13557) );
  NAND2_X1 U15522 ( .A1(n13355), .A2(n13354), .ZN(n13559) );
  NOR2_X1 U15523 ( .A1(n14556), .A2(n13559), .ZN(n13363) );
  NOR2_X1 U15524 ( .A1(n13558), .A2(n13528), .ZN(n13356) );
  AOI211_X1 U15525 ( .C1(n14556), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13363), 
        .B(n13356), .ZN(n13357) );
  OAI21_X1 U15526 ( .B1(n13557), .B2(n13550), .A(n13357), .ZN(P2_U3234) );
  INV_X1 U15527 ( .A(n13365), .ZN(n13561) );
  INV_X1 U15528 ( .A(n13358), .ZN(n13361) );
  OAI211_X1 U15529 ( .C1(n13561), .C2(n13361), .A(n13360), .B(n10936), .ZN(
        n13560) );
  NOR2_X1 U15530 ( .A1(n13441), .A2(n13362), .ZN(n13364) );
  AOI211_X1 U15531 ( .C1(n13365), .C2(n14557), .A(n13364), .B(n13363), .ZN(
        n13366) );
  OAI21_X1 U15532 ( .B1(n13560), .B2(n13550), .A(n13366), .ZN(P2_U3235) );
  AOI21_X1 U15533 ( .B1(n13372), .B2(n11951), .A(n13368), .ZN(n13370) );
  NOR2_X1 U15534 ( .A1(n13370), .A2(n13369), .ZN(n13569) );
  OAI21_X1 U15535 ( .B1(n13373), .B2(n13372), .A(n13371), .ZN(n13570) );
  NAND2_X1 U15536 ( .A1(n15599), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n13374) );
  OAI21_X1 U15537 ( .B1(n15592), .B2(n13375), .A(n13374), .ZN(n13376) );
  AOI21_X1 U15538 ( .B1(n13567), .B2(n14557), .A(n13376), .ZN(n13380) );
  AOI21_X1 U15539 ( .B1(n13389), .B2(n13567), .A(n13459), .ZN(n13378) );
  NAND2_X1 U15540 ( .A1(n13566), .A2(n15590), .ZN(n13379) );
  OAI211_X1 U15541 ( .C1(n13570), .C2(n13496), .A(n13380), .B(n13379), .ZN(
        n13381) );
  INV_X1 U15542 ( .A(n13381), .ZN(n13382) );
  OAI21_X1 U15543 ( .B1(n15599), .B2(n13569), .A(n13382), .ZN(P2_U3237) );
  XNOR2_X1 U15544 ( .A(n13383), .B(n13387), .ZN(n13386) );
  INV_X1 U15545 ( .A(n13384), .ZN(n13385) );
  AOI21_X1 U15546 ( .B1(n13386), .B2(n13521), .A(n13385), .ZN(n13576) );
  OR2_X1 U15547 ( .A1(n13388), .A2(n13387), .ZN(n13572) );
  NAND3_X1 U15548 ( .A1(n13572), .A2(n13571), .A3(n14563), .ZN(n13396) );
  OAI211_X1 U15549 ( .C1(n13390), .C2(n13404), .A(n10936), .B(n13389), .ZN(
        n13575) );
  AOI22_X1 U15550 ( .A1(n14556), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13391), 
        .B2(n14555), .ZN(n13393) );
  NAND2_X1 U15551 ( .A1(n13573), .A2(n14557), .ZN(n13392) );
  OAI211_X1 U15552 ( .C1(n13575), .C2(n13550), .A(n13393), .B(n13392), .ZN(
        n13394) );
  INV_X1 U15553 ( .A(n13394), .ZN(n13395) );
  OAI211_X1 U15554 ( .C1(n15599), .C2(n13576), .A(n13396), .B(n13395), .ZN(
        P2_U3238) );
  XOR2_X1 U15555 ( .A(n13401), .B(n13397), .Z(n13399) );
  AOI21_X1 U15556 ( .B1(n13399), .B2(n13521), .A(n13398), .ZN(n13581) );
  XOR2_X1 U15557 ( .A(n13401), .B(n13400), .Z(n13582) );
  INV_X1 U15558 ( .A(n13582), .ZN(n13409) );
  NAND2_X1 U15559 ( .A1(n13579), .A2(n13412), .ZN(n13402) );
  NAND2_X1 U15560 ( .A1(n13402), .A2(n10936), .ZN(n13403) );
  NOR2_X1 U15561 ( .A1(n13404), .A2(n13403), .ZN(n13578) );
  NAND2_X1 U15562 ( .A1(n13578), .A2(n15590), .ZN(n13407) );
  AOI22_X1 U15563 ( .A1(n14556), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13405), 
        .B2(n14555), .ZN(n13406) );
  OAI211_X1 U15564 ( .C1(n7065), .C2(n13528), .A(n13407), .B(n13406), .ZN(
        n13408) );
  AOI21_X1 U15565 ( .B1(n13409), .B2(n14563), .A(n13408), .ZN(n13410) );
  OAI21_X1 U15566 ( .B1(n15599), .B2(n13581), .A(n13410), .ZN(P2_U3239) );
  XOR2_X1 U15567 ( .A(n13417), .B(n13411), .Z(n13587) );
  INV_X1 U15568 ( .A(n13412), .ZN(n13413) );
  AOI211_X1 U15569 ( .C1(n13584), .C2(n7069), .A(n13459), .B(n13413), .ZN(
        n13583) );
  AOI22_X1 U15570 ( .A1(n14556), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13414), 
        .B2(n14555), .ZN(n13415) );
  OAI21_X1 U15571 ( .B1(n13416), .B2(n13528), .A(n13415), .ZN(n13426) );
  INV_X1 U15572 ( .A(n13417), .ZN(n13419) );
  NAND3_X1 U15573 ( .A1(n13432), .A2(n13419), .A3(n13418), .ZN(n13420) );
  NAND2_X1 U15574 ( .A1(n13421), .A2(n13420), .ZN(n13424) );
  AOI222_X1 U15575 ( .A1(n13521), .A2(n13424), .B1(n13423), .B2(n13650), .C1(
        n13422), .C2(n13470), .ZN(n13586) );
  NOR2_X1 U15576 ( .A1(n13586), .A2(n14556), .ZN(n13425) );
  AOI211_X1 U15577 ( .C1(n13583), .C2(n15590), .A(n13426), .B(n13425), .ZN(
        n13427) );
  OAI21_X1 U15578 ( .B1(n13587), .B2(n13496), .A(n13427), .ZN(P2_U3240) );
  OAI21_X1 U15579 ( .B1(n6773), .B2(n13429), .A(n13428), .ZN(n13591) );
  OR2_X1 U15580 ( .A1(n13591), .A2(n13647), .ZN(n13437) );
  NAND2_X1 U15581 ( .A1(n13430), .A2(n13429), .ZN(n13431) );
  NAND2_X1 U15582 ( .A1(n13432), .A2(n13431), .ZN(n13435) );
  INV_X1 U15583 ( .A(n13433), .ZN(n13434) );
  AOI21_X1 U15584 ( .B1(n13435), .B2(n13521), .A(n13434), .ZN(n13436) );
  NAND2_X1 U15585 ( .A1(n13437), .A2(n13436), .ZN(n13592) );
  NAND2_X1 U15586 ( .A1(n13592), .A2(n13441), .ZN(n13448) );
  INV_X1 U15587 ( .A(n13438), .ZN(n13439) );
  OAI22_X1 U15588 ( .A1(n13441), .A2(n13440), .B1(n13439), .B2(n15592), .ZN(
        n13446) );
  NAND2_X1 U15589 ( .A1(n13588), .A2(n13457), .ZN(n13442) );
  NAND2_X1 U15590 ( .A1(n13442), .A2(n10936), .ZN(n13444) );
  OR2_X1 U15591 ( .A1(n13444), .A2(n13443), .ZN(n13589) );
  NOR2_X1 U15592 ( .A1(n13589), .A2(n13550), .ZN(n13445) );
  AOI211_X1 U15593 ( .C1(n14557), .C2(n13588), .A(n13446), .B(n13445), .ZN(
        n13447) );
  OAI211_X1 U15594 ( .C1(n13591), .C2(n15596), .A(n13448), .B(n13447), .ZN(
        P2_U3241) );
  XOR2_X1 U15595 ( .A(n13449), .B(n13453), .Z(n13456) );
  OAI22_X1 U15596 ( .A1(n13451), .A2(n13538), .B1(n13450), .B2(n13540), .ZN(
        n13455) );
  XOR2_X1 U15597 ( .A(n13453), .B(n13452), .Z(n13599) );
  NOR2_X1 U15598 ( .A1(n13599), .A2(n13647), .ZN(n13454) );
  AOI211_X1 U15599 ( .C1(n13456), .C2(n13521), .A(n13455), .B(n13454), .ZN(
        n13598) );
  INV_X1 U15600 ( .A(n13475), .ZN(n13460) );
  INV_X1 U15601 ( .A(n13457), .ZN(n13458) );
  AOI211_X1 U15602 ( .C1(n13596), .C2(n13460), .A(n13459), .B(n13458), .ZN(
        n13595) );
  AOI22_X1 U15603 ( .A1(n13461), .A2(n14555), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n15599), .ZN(n13462) );
  OAI21_X1 U15604 ( .B1(n13463), .B2(n13528), .A(n13462), .ZN(n13465) );
  NOR2_X1 U15605 ( .A1(n13599), .A2(n15596), .ZN(n13464) );
  AOI211_X1 U15606 ( .C1(n13595), .C2(n15590), .A(n13465), .B(n13464), .ZN(
        n13466) );
  OAI21_X1 U15607 ( .B1(n13598), .B2(n14556), .A(n13466), .ZN(P2_U3242) );
  XNOR2_X1 U15608 ( .A(n13468), .B(n13467), .ZN(n13472) );
  AOI222_X1 U15609 ( .A1(n13521), .A2(n13472), .B1(n13471), .B2(n13470), .C1(
        n13469), .C2(n13650), .ZN(n13603) );
  XNOR2_X1 U15610 ( .A(n13474), .B(n13473), .ZN(n13604) );
  INV_X1 U15611 ( .A(n13604), .ZN(n13483) );
  OAI21_X1 U15612 ( .B1(n13488), .B2(n13481), .A(n10936), .ZN(n13476) );
  NOR2_X1 U15613 ( .A1(n13476), .A2(n13475), .ZN(n13600) );
  NAND2_X1 U15614 ( .A1(n13600), .A2(n15590), .ZN(n13480) );
  INV_X1 U15615 ( .A(n13477), .ZN(n13478) );
  AOI22_X1 U15616 ( .A1(n13478), .A2(n14555), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n15599), .ZN(n13479) );
  OAI211_X1 U15617 ( .C1(n13481), .C2(n13528), .A(n13480), .B(n13479), .ZN(
        n13482) );
  AOI21_X1 U15618 ( .B1(n13483), .B2(n14563), .A(n13482), .ZN(n13484) );
  OAI21_X1 U15619 ( .B1(n13603), .B2(n14556), .A(n13484), .ZN(P2_U3243) );
  XOR2_X1 U15620 ( .A(n13494), .B(n13485), .Z(n13487) );
  AOI21_X1 U15621 ( .B1(n13487), .B2(n13521), .A(n13486), .ZN(n13608) );
  OAI21_X1 U15622 ( .B1(n13508), .B2(n13493), .A(n10936), .ZN(n13489) );
  NOR2_X1 U15623 ( .A1(n13489), .A2(n13488), .ZN(n13605) );
  INV_X1 U15624 ( .A(n13490), .ZN(n13491) );
  AOI22_X1 U15625 ( .A1(n13491), .A2(n14555), .B1(n15599), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n13492) );
  OAI21_X1 U15626 ( .B1(n13493), .B2(n13528), .A(n13492), .ZN(n13498) );
  XNOR2_X1 U15627 ( .A(n13495), .B(n13494), .ZN(n13609) );
  NOR2_X1 U15628 ( .A1(n13609), .A2(n13496), .ZN(n13497) );
  AOI211_X1 U15629 ( .C1(n13605), .C2(n15590), .A(n13498), .B(n13497), .ZN(
        n13499) );
  OAI21_X1 U15630 ( .B1(n15599), .B2(n13608), .A(n13499), .ZN(P2_U3244) );
  XNOR2_X1 U15631 ( .A(n13501), .B(n13500), .ZN(n13503) );
  AOI21_X1 U15632 ( .B1(n13503), .B2(n13521), .A(n13502), .ZN(n13613) );
  OAI21_X1 U15633 ( .B1(n6796), .B2(n13505), .A(n13504), .ZN(n13614) );
  INV_X1 U15634 ( .A(n13614), .ZN(n13514) );
  NAND2_X1 U15635 ( .A1(n13611), .A2(n13523), .ZN(n13506) );
  NAND2_X1 U15636 ( .A1(n13506), .A2(n10936), .ZN(n13507) );
  NOR2_X1 U15637 ( .A1(n13508), .A2(n13507), .ZN(n13610) );
  NAND2_X1 U15638 ( .A1(n13610), .A2(n15590), .ZN(n13511) );
  AOI22_X1 U15639 ( .A1(n14556), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13509), 
        .B2(n14555), .ZN(n13510) );
  OAI211_X1 U15640 ( .C1(n13512), .C2(n13528), .A(n13511), .B(n13510), .ZN(
        n13513) );
  AOI21_X1 U15641 ( .B1(n13514), .B2(n14563), .A(n13513), .ZN(n13515) );
  OAI21_X1 U15642 ( .B1(n15599), .B2(n13613), .A(n13515), .ZN(P2_U3245) );
  XOR2_X1 U15643 ( .A(n13516), .B(n13517), .Z(n13522) );
  XNOR2_X1 U15644 ( .A(n13518), .B(n13517), .ZN(n13619) );
  NOR2_X1 U15645 ( .A1(n13619), .A2(n13647), .ZN(n13519) );
  AOI211_X1 U15646 ( .C1(n13522), .C2(n13521), .A(n13520), .B(n13519), .ZN(
        n13618) );
  INV_X1 U15647 ( .A(n13548), .ZN(n13525) );
  INV_X1 U15648 ( .A(n13523), .ZN(n13524) );
  AOI211_X1 U15649 ( .C1(n13616), .C2(n13525), .A(n13459), .B(n13524), .ZN(
        n13615) );
  AOI22_X1 U15650 ( .A1(n15599), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13526), 
        .B2(n14555), .ZN(n13527) );
  OAI21_X1 U15651 ( .B1(n13529), .B2(n13528), .A(n13527), .ZN(n13531) );
  NOR2_X1 U15652 ( .A1(n13619), .A2(n15596), .ZN(n13530) );
  AOI211_X1 U15653 ( .C1(n13615), .C2(n15590), .A(n13531), .B(n13530), .ZN(
        n13532) );
  OAI21_X1 U15654 ( .B1(n13618), .B2(n14556), .A(n13532), .ZN(P2_U3246) );
  NAND2_X1 U15655 ( .A1(n13533), .A2(n13536), .ZN(n13534) );
  NAND2_X1 U15656 ( .A1(n13535), .A2(n13534), .ZN(n13620) );
  INV_X1 U15657 ( .A(n13620), .ZN(n13556) );
  XNOR2_X1 U15658 ( .A(n13537), .B(n7276), .ZN(n13545) );
  NAND2_X1 U15659 ( .A1(n13620), .A2(n14873), .ZN(n13544) );
  OAI22_X1 U15660 ( .A1(n13541), .A2(n13540), .B1(n13539), .B2(n13538), .ZN(
        n13542) );
  INV_X1 U15661 ( .A(n13542), .ZN(n13543) );
  OAI211_X1 U15662 ( .C1(n14548), .C2(n13545), .A(n13544), .B(n13543), .ZN(
        n13625) );
  NAND2_X1 U15663 ( .A1(n13625), .A2(n13441), .ZN(n13555) );
  OAI22_X1 U15664 ( .A1(n13441), .A2(n13547), .B1(n13546), .B2(n15592), .ZN(
        n13552) );
  OAI21_X1 U15665 ( .B1(n6788), .B2(n13623), .A(n10936), .ZN(n13549) );
  OR2_X1 U15666 ( .A1(n13549), .A2(n13548), .ZN(n13621) );
  NOR2_X1 U15667 ( .A1(n13621), .A2(n13550), .ZN(n13551) );
  AOI211_X1 U15668 ( .C1(n14557), .C2(n7063), .A(n13552), .B(n13551), .ZN(
        n13554) );
  OAI211_X1 U15669 ( .C1(n13556), .C2(n15596), .A(n13555), .B(n13554), .ZN(
        P2_U3247) );
  OAI211_X1 U15670 ( .C1(n13558), .C2(n14909), .A(n13557), .B(n13559), .ZN(
        n13656) );
  MUX2_X1 U15671 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13656), .S(n14943), .Z(
        P2_U3530) );
  OAI211_X1 U15672 ( .C1(n13561), .C2(n14909), .A(n13560), .B(n13559), .ZN(
        n13657) );
  MUX2_X1 U15673 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13657), .S(n14943), .Z(
        P2_U3529) );
  MUX2_X1 U15674 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13658), .S(n14943), .Z(
        P2_U3528) );
  AOI21_X1 U15675 ( .B1(n14917), .B2(n13567), .A(n13566), .ZN(n13568) );
  OAI211_X1 U15676 ( .C1(n13570), .C2(n14890), .A(n13569), .B(n13568), .ZN(
        n13659) );
  MUX2_X1 U15677 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13659), .S(n14943), .Z(
        P2_U3527) );
  INV_X1 U15678 ( .A(n14890), .ZN(n14870) );
  NAND3_X1 U15679 ( .A1(n13572), .A2(n13571), .A3(n14870), .ZN(n13577) );
  NAND2_X1 U15680 ( .A1(n13573), .A2(n14917), .ZN(n13574) );
  NAND4_X1 U15681 ( .A1(n13577), .A2(n13576), .A3(n13575), .A4(n13574), .ZN(
        n13660) );
  MUX2_X1 U15682 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13660), .S(n14943), .Z(
        P2_U3526) );
  AOI21_X1 U15683 ( .B1(n14917), .B2(n13579), .A(n13578), .ZN(n13580) );
  OAI211_X1 U15684 ( .C1(n13582), .C2(n14890), .A(n13581), .B(n13580), .ZN(
        n13661) );
  MUX2_X1 U15685 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13661), .S(n14943), .Z(
        P2_U3525) );
  AOI21_X1 U15686 ( .B1(n14917), .B2(n13584), .A(n13583), .ZN(n13585) );
  OAI211_X1 U15687 ( .C1(n13587), .C2(n14890), .A(n13586), .B(n13585), .ZN(
        n13662) );
  MUX2_X1 U15688 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13662), .S(n14943), .Z(
        P2_U3524) );
  INV_X1 U15689 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n15359) );
  NAND2_X1 U15690 ( .A1(n13588), .A2(n14917), .ZN(n13590) );
  OAI211_X1 U15691 ( .C1(n13591), .C2(n13655), .A(n13590), .B(n13589), .ZN(
        n13593) );
  NOR2_X1 U15692 ( .A1(n13593), .A2(n13592), .ZN(n13663) );
  MUX2_X1 U15693 ( .A(n15359), .B(n13663), .S(n14943), .Z(n13594) );
  INV_X1 U15694 ( .A(n13594), .ZN(P2_U3523) );
  AOI21_X1 U15695 ( .B1(n14917), .B2(n13596), .A(n13595), .ZN(n13597) );
  OAI211_X1 U15696 ( .C1(n13599), .C2(n13655), .A(n13598), .B(n13597), .ZN(
        n13666) );
  MUX2_X1 U15697 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13666), .S(n14943), .Z(
        P2_U3522) );
  AOI21_X1 U15698 ( .B1(n14917), .B2(n13601), .A(n13600), .ZN(n13602) );
  OAI211_X1 U15699 ( .C1(n14890), .C2(n13604), .A(n13603), .B(n13602), .ZN(
        n13667) );
  MUX2_X1 U15700 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13667), .S(n14943), .Z(
        P2_U3521) );
  AOI21_X1 U15701 ( .B1(n14917), .B2(n13606), .A(n13605), .ZN(n13607) );
  OAI211_X1 U15702 ( .C1(n13609), .C2(n14890), .A(n13608), .B(n13607), .ZN(
        n13668) );
  MUX2_X1 U15703 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13668), .S(n14943), .Z(
        P2_U3520) );
  AOI21_X1 U15704 ( .B1(n14917), .B2(n13611), .A(n13610), .ZN(n13612) );
  OAI211_X1 U15705 ( .C1(n13614), .C2(n14890), .A(n13613), .B(n13612), .ZN(
        n13669) );
  MUX2_X1 U15706 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13669), .S(n14943), .Z(
        P2_U3519) );
  AOI21_X1 U15707 ( .B1(n14917), .B2(n13616), .A(n13615), .ZN(n13617) );
  OAI211_X1 U15708 ( .C1(n13655), .C2(n13619), .A(n13618), .B(n13617), .ZN(
        n13670) );
  MUX2_X1 U15709 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13670), .S(n14943), .Z(
        P2_U3518) );
  NAND2_X1 U15710 ( .A1(n13620), .A2(n14915), .ZN(n13622) );
  OAI211_X1 U15711 ( .C1(n13623), .C2(n14909), .A(n13622), .B(n13621), .ZN(
        n13624) );
  MUX2_X1 U15712 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13671), .S(n14943), .Z(
        P2_U3517) );
  AOI21_X1 U15713 ( .B1(n14917), .B2(n13627), .A(n13626), .ZN(n13628) );
  OAI211_X1 U15714 ( .C1(n13630), .C2(n14890), .A(n13629), .B(n13628), .ZN(
        n13672) );
  MUX2_X1 U15715 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13672), .S(n14943), .Z(
        P2_U3516) );
  AOI21_X1 U15716 ( .B1(n14917), .B2(n13632), .A(n13631), .ZN(n13633) );
  OAI211_X1 U15717 ( .C1(n14890), .C2(n13635), .A(n13634), .B(n13633), .ZN(
        n13673) );
  MUX2_X1 U15718 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13673), .S(n14943), .Z(
        P2_U3515) );
  AOI21_X1 U15719 ( .B1(n14917), .B2(n13637), .A(n13636), .ZN(n13638) );
  OAI211_X1 U15720 ( .C1(n13640), .C2(n14890), .A(n13639), .B(n13638), .ZN(
        n13674) );
  MUX2_X1 U15721 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13674), .S(n14943), .Z(
        P2_U3514) );
  AOI211_X1 U15722 ( .C1(n14917), .C2(n13643), .A(n13642), .B(n13641), .ZN(
        n13644) );
  OAI21_X1 U15723 ( .B1(n14890), .B2(n13645), .A(n13644), .ZN(n13675) );
  MUX2_X1 U15724 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13675), .S(n14943), .Z(
        P2_U3513) );
  MUX2_X1 U15725 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n13646), .S(n14943), .Z(
        P2_U3500) );
  INV_X1 U15726 ( .A(n15595), .ZN(n13649) );
  NAND2_X1 U15727 ( .A1(n13647), .A2(n14548), .ZN(n13648) );
  NAND2_X1 U15728 ( .A1(n13649), .A2(n13648), .ZN(n13652) );
  NAND2_X1 U15729 ( .A1(n13650), .A2(n11323), .ZN(n13651) );
  AND2_X1 U15730 ( .A1(n13652), .A2(n13651), .ZN(n15594) );
  NAND2_X1 U15731 ( .A1(n13654), .A2(n13653), .ZN(n15601) );
  OAI211_X1 U15732 ( .C1(n15595), .C2(n13655), .A(n15594), .B(n15601), .ZN(
        n14858) );
  MUX2_X1 U15733 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n14858), .S(n14943), .Z(
        P2_U3499) );
  MUX2_X1 U15734 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13656), .S(n14925), .Z(
        P2_U3498) );
  MUX2_X1 U15735 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13657), .S(n14925), .Z(
        P2_U3497) );
  MUX2_X1 U15736 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13659), .S(n14925), .Z(
        P2_U3495) );
  MUX2_X1 U15737 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13660), .S(n14925), .Z(
        P2_U3494) );
  MUX2_X1 U15738 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13661), .S(n14925), .Z(
        P2_U3493) );
  MUX2_X1 U15739 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13662), .S(n14925), .Z(
        P2_U3492) );
  INV_X1 U15740 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13664) );
  MUX2_X1 U15741 ( .A(n13664), .B(n13663), .S(n14925), .Z(n13665) );
  INV_X1 U15742 ( .A(n13665), .ZN(P2_U3491) );
  MUX2_X1 U15743 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13666), .S(n14925), .Z(
        P2_U3490) );
  MUX2_X1 U15744 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13667), .S(n14925), .Z(
        P2_U3489) );
  MUX2_X1 U15745 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13668), .S(n14925), .Z(
        P2_U3488) );
  MUX2_X1 U15746 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13669), .S(n14925), .Z(
        P2_U3487) );
  MUX2_X1 U15747 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13670), .S(n14925), .Z(
        P2_U3486) );
  MUX2_X1 U15748 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13671), .S(n14925), .Z(
        P2_U3484) );
  MUX2_X1 U15749 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13672), .S(n14925), .Z(
        P2_U3481) );
  MUX2_X1 U15750 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13673), .S(n14925), .Z(
        P2_U3478) );
  MUX2_X1 U15751 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13674), .S(n14925), .Z(
        P2_U3475) );
  MUX2_X1 U15752 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13675), .S(n14925), .Z(
        P2_U3472) );
  INV_X1 U15753 ( .A(n12194), .ZN(n14325) );
  NAND2_X1 U15754 ( .A1(n13676), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13681) );
  INV_X1 U15755 ( .A(n13677), .ZN(n13679) );
  NAND4_X1 U15756 ( .A1(n13679), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .A4(n13678), .ZN(n13680) );
  OAI211_X1 U15757 ( .C1(n14325), .C2(n11317), .A(n13681), .B(n13680), .ZN(
        P2_U3296) );
  INV_X1 U15758 ( .A(n13682), .ZN(n14327) );
  OAI222_X1 U15759 ( .A1(n11317), .A2(n14327), .B1(P2_U3088), .B2(n13683), 
        .C1(n13684), .C2(n13693), .ZN(P2_U3298) );
  NAND2_X1 U15760 ( .A1(n13686), .A2(n13685), .ZN(n13688) );
  OAI211_X1 U15761 ( .C1(n13693), .C2(n13689), .A(n13688), .B(n13687), .ZN(
        P2_U3299) );
  INV_X1 U15762 ( .A(n13690), .ZN(n14329) );
  OAI222_X1 U15763 ( .A1(n13693), .A2(n13692), .B1(n11317), .B2(n14329), .C1(
        n13691), .C2(P2_U3088), .ZN(P2_U3300) );
  MUX2_X1 U15764 ( .A(n13694), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15765 ( .A(n14033), .ZN(n13700) );
  AOI22_X1 U15766 ( .A1(n13797), .A2(n13818), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13698) );
  OAI21_X1 U15767 ( .B1(n8809), .B2(n14594), .A(n13698), .ZN(n13699) );
  AOI21_X1 U15768 ( .B1(n13700), .B2(n13806), .A(n13699), .ZN(n13701) );
  NAND2_X1 U15769 ( .A1(n14110), .A2(n14743), .ZN(n14225) );
  INV_X1 U15770 ( .A(n13702), .ZN(n13704) );
  NOR3_X1 U15771 ( .A1(n13705), .A2(n13704), .A3(n13703), .ZN(n13708) );
  OAI21_X1 U15772 ( .B1(n13708), .B2(n6715), .A(n14585), .ZN(n13713) );
  INV_X1 U15773 ( .A(n14101), .ZN(n13711) );
  AND2_X1 U15774 ( .A1(n14061), .A2(n14079), .ZN(n13709) );
  AOI21_X1 U15775 ( .B1(n13819), .B2(n14082), .A(n13709), .ZN(n14226) );
  OAI22_X1 U15776 ( .A1(n14226), .A2(n13808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15519), .ZN(n13710) );
  AOI21_X1 U15777 ( .B1(n13711), .B2(n13806), .A(n13710), .ZN(n13712) );
  OAI211_X1 U15778 ( .C1(n13804), .C2(n14225), .A(n13713), .B(n13712), .ZN(
        P1_U3216) );
  AND2_X1 U15779 ( .A1(n13714), .A2(n13715), .ZN(n13718) );
  OAI211_X1 U15780 ( .C1(n13718), .C2(n13717), .A(n14585), .B(n13716), .ZN(
        n13722) );
  NAND2_X1 U15781 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13972)
         );
  OAI21_X1 U15782 ( .B1(n14593), .B2(n14253), .A(n13972), .ZN(n13720) );
  NOR2_X1 U15783 ( .A1(n14606), .A2(n14179), .ZN(n13719) );
  AOI211_X1 U15784 ( .C1(n13789), .C2(n13823), .A(n13720), .B(n13719), .ZN(
        n13721) );
  OAI211_X1 U15785 ( .C1(n14310), .C2(n13792), .A(n13722), .B(n13721), .ZN(
        P1_U3219) );
  AOI21_X1 U15786 ( .B1(n12268), .B2(n13723), .A(n7573), .ZN(n13728) );
  OAI22_X1 U15787 ( .A1(n13724), .A2(n14260), .B1(n14253), .B2(n14170), .ZN(
        n14146) );
  AOI22_X1 U15788 ( .A1(n14146), .A2(n14587), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13725) );
  OAI21_X1 U15789 ( .B1(n14138), .B2(n14606), .A(n13725), .ZN(n13726) );
  AOI21_X1 U15790 ( .B1(n14303), .B2(n14602), .A(n13726), .ZN(n13727) );
  OAI21_X1 U15791 ( .B1(n13728), .B2(n14598), .A(n13727), .ZN(P1_U3223) );
  AOI22_X1 U15792 ( .A1(n13797), .A2(n14060), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13730) );
  NAND2_X1 U15793 ( .A1(n13789), .A2(n14061), .ZN(n13729) );
  OAI211_X1 U15794 ( .C1(n14606), .C2(n14064), .A(n13730), .B(n13729), .ZN(
        n13738) );
  INV_X1 U15795 ( .A(n13732), .ZN(n13733) );
  NAND3_X1 U15796 ( .A1(n13731), .A2(n13734), .A3(n13733), .ZN(n13735) );
  AOI21_X1 U15797 ( .B1(n13736), .B2(n13735), .A(n14598), .ZN(n13737) );
  AOI211_X1 U15798 ( .C1(n14602), .C2(n14067), .A(n13738), .B(n13737), .ZN(
        n13739) );
  INV_X1 U15799 ( .A(n13739), .ZN(P1_U3225) );
  OAI21_X1 U15800 ( .B1(n13742), .B2(n13741), .A(n13740), .ZN(n13743) );
  NAND2_X1 U15801 ( .A1(n13743), .A2(n14585), .ZN(n13750) );
  OAI21_X1 U15802 ( .B1(n14593), .B2(n13745), .A(n13744), .ZN(n13748) );
  NOR2_X1 U15803 ( .A1(n14606), .A2(n13746), .ZN(n13747) );
  AOI211_X1 U15804 ( .C1(n13789), .C2(n13826), .A(n13748), .B(n13747), .ZN(
        n13749) );
  OAI211_X1 U15805 ( .C1(n13751), .C2(n13792), .A(n13750), .B(n13749), .ZN(
        P1_U3226) );
  NAND2_X1 U15806 ( .A1(n13753), .A2(n13752), .ZN(n13754) );
  XNOR2_X1 U15807 ( .A(n13755), .B(n13754), .ZN(n13763) );
  NAND2_X1 U15808 ( .A1(n13806), .A2(n13756), .ZN(n13758) );
  OAI211_X1 U15809 ( .C1(n13759), .C2(n13808), .A(n13758), .B(n13757), .ZN(
        n13760) );
  AOI21_X1 U15810 ( .B1(n13761), .B2(n14602), .A(n13760), .ZN(n13762) );
  OAI21_X1 U15811 ( .B1(n13763), .B2(n14598), .A(n13762), .ZN(P1_U3228) );
  NAND2_X1 U15812 ( .A1(n14094), .A2(n14743), .ZN(n14220) );
  INV_X1 U15813 ( .A(n13764), .ZN(n13766) );
  NOR3_X1 U15814 ( .A1(n6715), .A2(n13766), .A3(n13765), .ZN(n13768) );
  INV_X1 U15815 ( .A(n13731), .ZN(n13767) );
  OAI21_X1 U15816 ( .B1(n13768), .B2(n13767), .A(n14585), .ZN(n13774) );
  INV_X1 U15817 ( .A(n14088), .ZN(n13772) );
  AOI22_X1 U15818 ( .A1(n13797), .A2(n14080), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13769) );
  OAI21_X1 U15819 ( .B1(n13770), .B2(n14594), .A(n13769), .ZN(n13771) );
  AOI21_X1 U15820 ( .B1(n13772), .B2(n13806), .A(n13771), .ZN(n13773) );
  OAI211_X1 U15821 ( .C1(n13804), .C2(n14220), .A(n13774), .B(n13773), .ZN(
        P1_U3229) );
  XNOR2_X1 U15822 ( .A(n13776), .B(n13775), .ZN(n13781) );
  AOI22_X1 U15823 ( .A1(n13820), .A2(n13797), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13778) );
  NAND2_X1 U15824 ( .A1(n13789), .A2(n13822), .ZN(n13777) );
  OAI211_X1 U15825 ( .C1(n14606), .C2(n14153), .A(n13778), .B(n13777), .ZN(
        n13779) );
  AOI21_X1 U15826 ( .B1(n14248), .B2(n14602), .A(n13779), .ZN(n13780) );
  OAI21_X1 U15827 ( .B1(n13781), .B2(n14598), .A(n13780), .ZN(P1_U3233) );
  OAI21_X1 U15828 ( .B1(n13783), .B2(n13782), .A(n13714), .ZN(n13784) );
  NAND2_X1 U15829 ( .A1(n13784), .A2(n14585), .ZN(n13791) );
  OAI21_X1 U15830 ( .B1(n14593), .B2(n14261), .A(n13785), .ZN(n13788) );
  NOR2_X1 U15831 ( .A1(n14606), .A2(n13786), .ZN(n13787) );
  AOI211_X1 U15832 ( .C1(n13789), .C2(n13824), .A(n13788), .B(n13787), .ZN(
        n13790) );
  OAI211_X1 U15833 ( .C1(n14314), .C2(n13792), .A(n13791), .B(n13790), .ZN(
        P1_U3238) );
  NAND2_X1 U15834 ( .A1(n14049), .A2(n14743), .ZN(n14212) );
  OAI21_X1 U15835 ( .B1(n13795), .B2(n13794), .A(n13793), .ZN(n13796) );
  NAND2_X1 U15836 ( .A1(n13796), .A2(n14585), .ZN(n13803) );
  INV_X1 U15837 ( .A(n14044), .ZN(n13801) );
  AOI22_X1 U15838 ( .A1(n13797), .A2(n14042), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13798) );
  OAI21_X1 U15839 ( .B1(n13799), .B2(n14594), .A(n13798), .ZN(n13800) );
  AOI21_X1 U15840 ( .B1(n13801), .B2(n13806), .A(n13800), .ZN(n13802) );
  OAI211_X1 U15841 ( .C1(n13804), .C2(n14212), .A(n13803), .B(n13802), .ZN(
        P1_U3240) );
  NAND2_X1 U15842 ( .A1(n13806), .A2(n13805), .ZN(n13807) );
  NAND2_X1 U15843 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14649)
         );
  OAI211_X1 U15844 ( .C1(n13809), .C2(n13808), .A(n13807), .B(n14649), .ZN(
        n13814) );
  AOI211_X1 U15845 ( .C1(n13812), .C2(n13811), .A(n14598), .B(n6827), .ZN(
        n13813) );
  AOI211_X1 U15846 ( .C1(n14602), .C2(n13815), .A(n13814), .B(n13813), .ZN(
        n13816) );
  INV_X1 U15847 ( .A(n13816), .ZN(P1_U3241) );
  MUX2_X1 U15848 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13975), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15849 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13817), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15850 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14002), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15851 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13818), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15852 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14042), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15853 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14060), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15854 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14080), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15855 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14061), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15856 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14081), .S(n13847), .Z(
        P1_U3583) );
  MUX2_X1 U15857 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13819), .S(n13847), .Z(
        P1_U3582) );
  MUX2_X1 U15858 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13820), .S(n13847), .Z(
        P1_U3581) );
  MUX2_X1 U15859 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13821), .S(n13847), .Z(
        P1_U3580) );
  MUX2_X1 U15860 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13822), .S(n13847), .Z(
        P1_U3579) );
  MUX2_X1 U15861 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13823), .S(n13847), .Z(
        P1_U3578) );
  MUX2_X1 U15862 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13824), .S(n13847), .Z(
        P1_U3577) );
  MUX2_X1 U15863 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13825), .S(n13847), .Z(
        P1_U3576) );
  MUX2_X1 U15864 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13826), .S(n13847), .Z(
        P1_U3575) );
  MUX2_X1 U15865 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13827), .S(n13847), .Z(
        P1_U3574) );
  MUX2_X1 U15866 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13828), .S(n13847), .Z(
        P1_U3573) );
  MUX2_X1 U15867 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13829), .S(n13847), .Z(
        P1_U3572) );
  MUX2_X1 U15868 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13830), .S(n13847), .Z(
        P1_U3571) );
  MUX2_X1 U15869 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13831), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15870 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13832), .S(n13847), .Z(
        P1_U3569) );
  MUX2_X1 U15871 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13833), .S(n13847), .Z(
        P1_U3568) );
  MUX2_X1 U15872 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13834), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15873 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13835), .S(n13847), .Z(
        P1_U3566) );
  MUX2_X1 U15874 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13836), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15875 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13837), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15876 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13838), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15877 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13839), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15878 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9350), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15879 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13841), .S(P1_U4016), .Z(
        P1_U3560) );
  MUX2_X1 U15880 ( .A(n13843), .B(n13842), .S(n6843), .Z(n13848) );
  NAND2_X1 U15881 ( .A1(n13845), .A2(n13844), .ZN(n13846) );
  OAI211_X1 U15882 ( .C1(n13848), .C2(n8816), .A(n13847), .B(n13846), .ZN(
        n13896) );
  AOI22_X1 U15883 ( .A1(n13929), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13864) );
  INV_X1 U15884 ( .A(n13849), .ZN(n13872) );
  MUX2_X1 U15885 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9122), .S(n13861), .Z(
        n13852) );
  NAND3_X1 U15886 ( .A1(n13852), .A2(n13851), .A3(n13850), .ZN(n13853) );
  NAND3_X1 U15887 ( .A1(n13966), .A2(n13872), .A3(n13853), .ZN(n13860) );
  INV_X1 U15888 ( .A(n13875), .ZN(n13858) );
  MUX2_X1 U15889 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9129), .S(n13861), .Z(
        n13856) );
  NAND3_X1 U15890 ( .A1(n13856), .A2(n13855), .A3(n13854), .ZN(n13857) );
  NAND3_X1 U15891 ( .A1(n13963), .A2(n13858), .A3(n13857), .ZN(n13859) );
  OAI211_X1 U15892 ( .C1(n14647), .C2(n13861), .A(n13860), .B(n13859), .ZN(
        n13862) );
  INV_X1 U15893 ( .A(n13862), .ZN(n13863) );
  NAND3_X1 U15894 ( .A1(n13896), .A2(n13864), .A3(n13863), .ZN(P1_U3245) );
  INV_X1 U15895 ( .A(n14647), .ZN(n13943) );
  INV_X1 U15896 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n13866) );
  OAI21_X1 U15897 ( .B1(n14651), .B2(n13866), .A(n13865), .ZN(n13867) );
  AOI21_X1 U15898 ( .B1(n13869), .B2(n13943), .A(n13867), .ZN(n13880) );
  INV_X1 U15899 ( .A(n13868), .ZN(n13871) );
  MUX2_X1 U15900 ( .A(n9125), .B(P1_REG1_REG_3__SCAN_IN), .S(n13869), .Z(
        n13870) );
  NAND3_X1 U15901 ( .A1(n13872), .A2(n13871), .A3(n13870), .ZN(n13873) );
  NAND3_X1 U15902 ( .A1(n13966), .A2(n13883), .A3(n13873), .ZN(n13879) );
  OR3_X1 U15903 ( .A1(n13876), .A2(n13875), .A3(n13874), .ZN(n13877) );
  NAND3_X1 U15904 ( .A1(n13963), .A2(n13888), .A3(n13877), .ZN(n13878) );
  NAND3_X1 U15905 ( .A1(n13880), .A2(n13879), .A3(n13878), .ZN(P1_U3246) );
  AND3_X1 U15906 ( .A1(n13883), .A2(n13882), .A3(n13881), .ZN(n13884) );
  NOR3_X1 U15907 ( .A1(n14643), .A2(n13885), .A3(n13884), .ZN(n13895) );
  AND3_X1 U15908 ( .A1(n13888), .A2(n13887), .A3(n13886), .ZN(n13889) );
  NOR3_X1 U15909 ( .A1(n14645), .A2(n13890), .A3(n13889), .ZN(n13894) );
  OAI21_X1 U15910 ( .B1(n14647), .B2(n13892), .A(n13891), .ZN(n13893) );
  NOR3_X1 U15911 ( .A1(n13895), .A2(n13894), .A3(n13893), .ZN(n13898) );
  NAND2_X1 U15912 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n13929), .ZN(n13897) );
  NAND3_X1 U15913 ( .A1(n13898), .A2(n13897), .A3(n13896), .ZN(P1_U3247) );
  NOR2_X1 U15914 ( .A1(n14647), .A2(n13899), .ZN(n13900) );
  AOI211_X1 U15915 ( .C1(n13929), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n13901), .B(
        n13900), .ZN(n13918) );
  INV_X1 U15916 ( .A(n13902), .ZN(n13905) );
  MUX2_X1 U15917 ( .A(n13903), .B(P1_REG1_REG_7__SCAN_IN), .S(n13910), .Z(
        n13904) );
  NAND2_X1 U15918 ( .A1(n13905), .A2(n13904), .ZN(n13907) );
  OAI211_X1 U15919 ( .C1(n13908), .C2(n13907), .A(n13906), .B(n13966), .ZN(
        n13917) );
  INV_X1 U15920 ( .A(n13909), .ZN(n13912) );
  MUX2_X1 U15921 ( .A(n9205), .B(P1_REG2_REG_7__SCAN_IN), .S(n13910), .Z(
        n13911) );
  NAND2_X1 U15922 ( .A1(n13912), .A2(n13911), .ZN(n13914) );
  OAI211_X1 U15923 ( .C1(n13915), .C2(n13914), .A(n13963), .B(n13913), .ZN(
        n13916) );
  NAND3_X1 U15924 ( .A1(n13918), .A2(n13917), .A3(n13916), .ZN(P1_U3250) );
  INV_X1 U15925 ( .A(n13919), .ZN(n13924) );
  NOR3_X1 U15926 ( .A1(n13922), .A2(n13921), .A3(n13920), .ZN(n13923) );
  OAI21_X1 U15927 ( .B1(n13924), .B2(n13923), .A(n13966), .ZN(n13937) );
  NOR2_X1 U15928 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13925), .ZN(n13928) );
  NOR2_X1 U15929 ( .A1(n14647), .A2(n13926), .ZN(n13927) );
  AOI211_X1 U15930 ( .C1(n13929), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n13928), .B(
        n13927), .ZN(n13936) );
  OR3_X1 U15931 ( .A1(n13932), .A2(n13931), .A3(n13930), .ZN(n13933) );
  NAND3_X1 U15932 ( .A1(n13934), .A2(n13963), .A3(n13933), .ZN(n13935) );
  NAND3_X1 U15933 ( .A1(n13937), .A2(n13936), .A3(n13935), .ZN(P1_U3252) );
  OAI21_X1 U15934 ( .B1(n13940), .B2(n13939), .A(n13938), .ZN(n13941) );
  NAND2_X1 U15935 ( .A1(n13941), .A2(n13966), .ZN(n13953) );
  NAND2_X1 U15936 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14603)
         );
  OAI21_X1 U15937 ( .B1(n14651), .B2(n14356), .A(n14603), .ZN(n13942) );
  AOI21_X1 U15938 ( .B1(n13945), .B2(n13943), .A(n13942), .ZN(n13952) );
  INV_X1 U15939 ( .A(n13944), .ZN(n13947) );
  MUX2_X1 U15940 ( .A(n9399), .B(P1_REG2_REG_11__SCAN_IN), .S(n13945), .Z(
        n13946) );
  NAND2_X1 U15941 ( .A1(n13947), .A2(n13946), .ZN(n13949) );
  OAI211_X1 U15942 ( .C1(n13950), .C2(n13949), .A(n13948), .B(n13963), .ZN(
        n13951) );
  NAND3_X1 U15943 ( .A1(n13953), .A2(n13952), .A3(n13951), .ZN(P1_U3254) );
  INV_X1 U15944 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14458) );
  NAND2_X1 U15945 ( .A1(n13959), .A2(n13954), .ZN(n13955) );
  NAND2_X1 U15946 ( .A1(n13956), .A2(n13955), .ZN(n13957) );
  XOR2_X1 U15947 ( .A(n13957), .B(P1_REG1_REG_19__SCAN_IN), .Z(n13964) );
  NAND2_X1 U15948 ( .A1(n13959), .A2(n13958), .ZN(n13960) );
  NAND2_X1 U15949 ( .A1(n13961), .A2(n13960), .ZN(n13962) );
  XOR2_X1 U15950 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13962), .Z(n13968) );
  AOI22_X1 U15951 ( .A1(n13964), .A2(n13966), .B1(n13963), .B2(n13968), .ZN(
        n13971) );
  INV_X1 U15952 ( .A(n13964), .ZN(n13965) );
  NAND2_X1 U15953 ( .A1(n13966), .A2(n13965), .ZN(n13967) );
  OAI211_X1 U15954 ( .C1(n13968), .C2(n14645), .A(n14647), .B(n13967), .ZN(
        n13969) );
  INV_X1 U15955 ( .A(n13969), .ZN(n13970) );
  MUX2_X1 U15956 ( .A(n13971), .B(n13970), .S(n14114), .Z(n13973) );
  OAI211_X1 U15957 ( .C1(n14458), .C2(n14651), .A(n13973), .B(n13972), .ZN(
        P1_U3262) );
  NAND2_X1 U15958 ( .A1(n14192), .A2(n14165), .ZN(n13977) );
  AND2_X1 U15959 ( .A1(n13975), .A2(n13974), .ZN(n14191) );
  INV_X1 U15960 ( .A(n14191), .ZN(n14195) );
  NOR2_X1 U15961 ( .A1(n14678), .A2(n14195), .ZN(n13983) );
  AOI21_X1 U15962 ( .B1(n14678), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13983), 
        .ZN(n13976) );
  OAI211_X1 U15963 ( .C1(n14284), .C2(n14156), .A(n13977), .B(n13976), .ZN(
        P1_U3263) );
  NAND2_X1 U15964 ( .A1(n13985), .A2(n13978), .ZN(n13979) );
  NAND2_X1 U15965 ( .A1(n13979), .A2(n14176), .ZN(n13981) );
  NOR2_X1 U15966 ( .A1(n14668), .A2(n13982), .ZN(n13984) );
  AOI211_X1 U15967 ( .C1(n13985), .C2(n14670), .A(n13984), .B(n13983), .ZN(
        n13986) );
  OAI21_X1 U15968 ( .B1(n14196), .B2(n14673), .A(n13986), .ZN(P1_U3264) );
  INV_X1 U15969 ( .A(n13987), .ZN(n13999) );
  OAI22_X1 U15970 ( .A1(n13990), .A2(n13989), .B1(n13988), .B2(n14665), .ZN(
        n13991) );
  AOI21_X1 U15971 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14678), .A(n13991), 
        .ZN(n13994) );
  NAND2_X1 U15972 ( .A1(n13992), .A2(n14670), .ZN(n13993) );
  OAI211_X1 U15973 ( .C1(n13995), .C2(n14673), .A(n13994), .B(n13993), .ZN(
        n13996) );
  AOI21_X1 U15974 ( .B1(n13997), .B2(n14188), .A(n13996), .ZN(n13998) );
  OAI21_X1 U15975 ( .B1(n13999), .B2(n14678), .A(n13998), .ZN(P1_U3356) );
  NAND2_X1 U15976 ( .A1(n14001), .A2(n7563), .ZN(n14006) );
  NAND2_X1 U15977 ( .A1(n14002), .A2(n14079), .ZN(n14004) );
  NAND2_X1 U15978 ( .A1(n14042), .A2(n14082), .ZN(n14003) );
  AOI21_X1 U15979 ( .B1(n14009), .B2(n14008), .A(n14007), .ZN(n14010) );
  INV_X1 U15980 ( .A(n14010), .ZN(n14203) );
  NAND2_X1 U15981 ( .A1(n14678), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14011) );
  OAI21_X1 U15982 ( .B1(n14665), .B2(n14012), .A(n14011), .ZN(n14013) );
  AOI21_X1 U15983 ( .B1(n14200), .B2(n14670), .A(n14013), .ZN(n14017) );
  AOI21_X1 U15984 ( .B1(n14030), .B2(n14200), .A(n14661), .ZN(n14015) );
  NAND2_X1 U15985 ( .A1(n14199), .A2(n14165), .ZN(n14016) );
  OAI211_X1 U15986 ( .C1(n14203), .C2(n14167), .A(n14017), .B(n14016), .ZN(
        n14018) );
  INV_X1 U15987 ( .A(n14018), .ZN(n14019) );
  OAI21_X1 U15988 ( .B1(n14678), .B2(n14202), .A(n14019), .ZN(P1_U3265) );
  OAI21_X1 U15989 ( .B1(n14022), .B2(n14021), .A(n14020), .ZN(n14206) );
  INV_X1 U15990 ( .A(n14206), .ZN(n14039) );
  OAI21_X1 U15991 ( .B1(n14025), .B2(n14024), .A(n14023), .ZN(n14028) );
  OAI22_X1 U15992 ( .A1(n14026), .A2(n14260), .B1(n8809), .B2(n14170), .ZN(
        n14027) );
  AOI21_X1 U15993 ( .B1(n14028), .B2(n14144), .A(n14027), .ZN(n14029) );
  OAI21_X1 U15994 ( .B1(n14039), .B2(n14087), .A(n14029), .ZN(n14204) );
  NAND2_X1 U15995 ( .A1(n14204), .A2(n14668), .ZN(n14038) );
  INV_X1 U15996 ( .A(n14030), .ZN(n14031) );
  AOI211_X1 U15997 ( .C1(n14032), .C2(n6689), .A(n14661), .B(n14031), .ZN(
        n14205) );
  NOR2_X1 U15998 ( .A1(n14292), .A2(n14156), .ZN(n14036) );
  OAI22_X1 U15999 ( .A1(n14668), .A2(n14034), .B1(n14033), .B2(n14665), .ZN(
        n14035) );
  AOI211_X1 U16000 ( .C1(n14205), .C2(n14165), .A(n14036), .B(n14035), .ZN(
        n14037) );
  OAI211_X1 U16001 ( .C1(n14039), .C2(n14097), .A(n14038), .B(n14037), .ZN(
        P1_U3266) );
  OAI21_X1 U16002 ( .B1(n14041), .B2(n14050), .A(n14040), .ZN(n14043) );
  AOI222_X1 U16003 ( .A1(n14144), .A2(n14043), .B1(n14042), .B2(n14079), .C1(
        n14080), .C2(n14082), .ZN(n14213) );
  OAI22_X1 U16004 ( .A1(n14668), .A2(n14045), .B1(n14044), .B2(n14665), .ZN(
        n14048) );
  INV_X1 U16005 ( .A(n14065), .ZN(n14046) );
  OAI211_X1 U16006 ( .C1(n7092), .C2(n14046), .A(n6689), .B(n14176), .ZN(
        n14210) );
  NOR2_X1 U16007 ( .A1(n14210), .A2(n14673), .ZN(n14047) );
  AOI211_X1 U16008 ( .C1(n14670), .C2(n14049), .A(n14048), .B(n14047), .ZN(
        n14053) );
  XNOR2_X1 U16009 ( .A(n14051), .B(n14050), .ZN(n14209) );
  NAND2_X1 U16010 ( .A1(n14209), .A2(n14188), .ZN(n14052) );
  OAI211_X1 U16011 ( .C1(n14213), .C2(n14678), .A(n14053), .B(n14052), .ZN(
        P1_U3267) );
  NAND2_X1 U16012 ( .A1(n14054), .A2(n14055), .ZN(n14056) );
  NAND2_X1 U16013 ( .A1(n14056), .A2(n14070), .ZN(n14058) );
  NAND2_X1 U16014 ( .A1(n14058), .A2(n14057), .ZN(n14059) );
  NAND2_X1 U16015 ( .A1(n14059), .A2(n14144), .ZN(n14063) );
  AOI22_X1 U16016 ( .A1(n14082), .A2(n14061), .B1(n14060), .B2(n14079), .ZN(
        n14062) );
  OAI21_X1 U16017 ( .B1(n14064), .B2(n14665), .A(n14215), .ZN(n14074) );
  AOI21_X1 U16018 ( .B1(n14067), .B2(n14090), .A(n14661), .ZN(n14066) );
  NAND2_X1 U16019 ( .A1(n14066), .A2(n14065), .ZN(n14214) );
  AOI22_X1 U16020 ( .A1(n14067), .A2(n14670), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n14678), .ZN(n14068) );
  OAI21_X1 U16021 ( .B1(n14214), .B2(n14673), .A(n14068), .ZN(n14073) );
  OAI21_X1 U16022 ( .B1(n14071), .B2(n14070), .A(n14069), .ZN(n14216) );
  NOR2_X1 U16023 ( .A1(n14216), .A2(n14167), .ZN(n14072) );
  AOI211_X1 U16024 ( .C1(n14668), .C2(n14074), .A(n14073), .B(n14072), .ZN(
        n14075) );
  INV_X1 U16025 ( .A(n14075), .ZN(P1_U3268) );
  INV_X1 U16026 ( .A(n14076), .ZN(n14077) );
  AOI21_X1 U16027 ( .B1(n14083), .B2(n14078), .A(n14077), .ZN(n14222) );
  AOI22_X1 U16028 ( .A1(n14082), .A2(n14081), .B1(n14080), .B2(n14079), .ZN(
        n14086) );
  OAI211_X1 U16029 ( .C1(n14084), .C2(n14083), .A(n14054), .B(n14144), .ZN(
        n14085) );
  OAI211_X1 U16030 ( .C1(n14222), .C2(n14087), .A(n14086), .B(n14085), .ZN(
        n14224) );
  NAND2_X1 U16031 ( .A1(n14224), .A2(n14668), .ZN(n14096) );
  OAI22_X1 U16032 ( .A1(n14668), .A2(n14089), .B1(n14088), .B2(n14665), .ZN(
        n14093) );
  OAI211_X1 U16033 ( .C1(n14091), .C2(n14113), .A(n14090), .B(n14176), .ZN(
        n14219) );
  NOR2_X1 U16034 ( .A1(n14219), .A2(n14673), .ZN(n14092) );
  AOI211_X1 U16035 ( .C1(n14670), .C2(n14094), .A(n14093), .B(n14092), .ZN(
        n14095) );
  OAI211_X1 U16036 ( .C1(n14222), .C2(n14097), .A(n14096), .B(n14095), .ZN(
        P1_U3269) );
  INV_X1 U16037 ( .A(n14098), .ZN(n14099) );
  AOI21_X1 U16038 ( .B1(n14106), .B2(n14100), .A(n14099), .ZN(n14230) );
  INV_X1 U16039 ( .A(n14230), .ZN(n14118) );
  OAI22_X1 U16040 ( .A1(n14668), .A2(n14102), .B1(n14101), .B2(n14665), .ZN(
        n14103) );
  AOI21_X1 U16041 ( .B1(n14110), .B2(n14670), .A(n14103), .ZN(n14117) );
  INV_X1 U16042 ( .A(n14104), .ZN(n14105) );
  NOR2_X1 U16043 ( .A1(n14106), .A2(n14105), .ZN(n14107) );
  NAND2_X1 U16044 ( .A1(n14122), .A2(n14107), .ZN(n14108) );
  AOI21_X1 U16045 ( .B1(n14109), .B2(n14108), .A(n14656), .ZN(n14229) );
  NAND2_X1 U16046 ( .A1(n14110), .A2(n14119), .ZN(n14111) );
  NAND2_X1 U16047 ( .A1(n14111), .A2(n14176), .ZN(n14112) );
  OR2_X1 U16048 ( .A1(n14113), .A2(n14112), .ZN(n14227) );
  OAI21_X1 U16049 ( .B1(n14227), .B2(n14114), .A(n14226), .ZN(n14115) );
  OAI21_X1 U16050 ( .B1(n14229), .B2(n14115), .A(n14668), .ZN(n14116) );
  OAI211_X1 U16051 ( .C1(n14118), .C2(n14167), .A(n14117), .B(n14116), .ZN(
        P1_U3270) );
  OAI211_X1 U16052 ( .C1(n14136), .C2(n14234), .A(n14119), .B(n14176), .ZN(
        n14233) );
  INV_X1 U16053 ( .A(n14233), .ZN(n14124) );
  INV_X1 U16054 ( .A(n14232), .ZN(n14123) );
  NAND2_X1 U16055 ( .A1(n14120), .A2(n14126), .ZN(n14121) );
  AOI21_X1 U16056 ( .B1(n14122), .B2(n14121), .A(n14656), .ZN(n14235) );
  AOI211_X1 U16057 ( .C1(n14124), .C2(n8775), .A(n14123), .B(n14235), .ZN(
        n14132) );
  OAI21_X1 U16058 ( .B1(n14127), .B2(n14126), .A(n14125), .ZN(n14237) );
  AOI22_X1 U16059 ( .A1(n14128), .A2(n14180), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14678), .ZN(n14129) );
  OAI21_X1 U16060 ( .B1(n14234), .B2(n14156), .A(n14129), .ZN(n14130) );
  AOI21_X1 U16061 ( .B1(n14237), .B2(n14188), .A(n14130), .ZN(n14131) );
  OAI21_X1 U16062 ( .B1(n14132), .B2(n14678), .A(n14131), .ZN(P1_U3271) );
  XNOR2_X1 U16063 ( .A(n14134), .B(n14133), .ZN(n14242) );
  NAND2_X1 U16064 ( .A1(n14151), .A2(n14303), .ZN(n14135) );
  NAND2_X1 U16065 ( .A1(n14135), .A2(n14176), .ZN(n14137) );
  OR2_X1 U16066 ( .A1(n14137), .A2(n14136), .ZN(n14239) );
  OAI22_X1 U16067 ( .A1(n14668), .A2(n14139), .B1(n14138), .B2(n14665), .ZN(
        n14140) );
  AOI21_X1 U16068 ( .B1(n14303), .B2(n14670), .A(n14140), .ZN(n14141) );
  OAI21_X1 U16069 ( .B1(n14239), .B2(n14673), .A(n14141), .ZN(n14148) );
  XNOR2_X1 U16070 ( .A(n14143), .B(n14142), .ZN(n14145) );
  NAND2_X1 U16071 ( .A1(n14145), .A2(n14144), .ZN(n14241) );
  INV_X1 U16072 ( .A(n14146), .ZN(n14240) );
  AOI21_X1 U16073 ( .B1(n14241), .B2(n14240), .A(n14678), .ZN(n14147) );
  AOI211_X1 U16074 ( .C1(n14188), .C2(n14242), .A(n14148), .B(n14147), .ZN(
        n14149) );
  INV_X1 U16075 ( .A(n14149), .ZN(P1_U3272) );
  XNOR2_X1 U16076 ( .A(n14150), .B(n7536), .ZN(n14251) );
  INV_X1 U16077 ( .A(n14151), .ZN(n14152) );
  AOI211_X1 U16078 ( .C1(n14248), .C2(n14177), .A(n14661), .B(n14152), .ZN(
        n14247) );
  INV_X1 U16079 ( .A(n14153), .ZN(n14154) );
  AOI22_X1 U16080 ( .A1(n14678), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14154), 
        .B2(n14180), .ZN(n14155) );
  OAI21_X1 U16081 ( .B1(n7082), .B2(n14156), .A(n14155), .ZN(n14164) );
  AOI21_X1 U16082 ( .B1(n14158), .B2(n14157), .A(n14656), .ZN(n14162) );
  OAI22_X1 U16083 ( .A1(n14159), .A2(n14260), .B1(n14261), .B2(n14170), .ZN(
        n14160) );
  AOI21_X1 U16084 ( .B1(n14162), .B2(n14161), .A(n14160), .ZN(n14250) );
  NOR2_X1 U16085 ( .A1(n14250), .A2(n14678), .ZN(n14163) );
  AOI211_X1 U16086 ( .C1(n14247), .C2(n14165), .A(n14164), .B(n14163), .ZN(
        n14166) );
  OAI21_X1 U16087 ( .B1(n14167), .B2(n14251), .A(n14166), .ZN(P1_U3273) );
  XNOR2_X1 U16088 ( .A(n14169), .B(n14168), .ZN(n14172) );
  OAI22_X1 U16089 ( .A1(n14172), .A2(n14656), .B1(n14171), .B2(n14170), .ZN(
        n14254) );
  INV_X1 U16090 ( .A(n14254), .ZN(n14190) );
  OAI21_X1 U16091 ( .B1(n14174), .B2(n8633), .A(n14173), .ZN(n14256) );
  INV_X1 U16092 ( .A(n14175), .ZN(n14178) );
  OAI211_X1 U16093 ( .C1(n14310), .C2(n14178), .A(n14177), .B(n14176), .ZN(
        n14252) );
  INV_X1 U16094 ( .A(n14179), .ZN(n14181) );
  AOI22_X1 U16095 ( .A1(n14678), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14181), 
        .B2(n14180), .ZN(n14182) );
  OAI21_X1 U16096 ( .B1(n14183), .B2(n14253), .A(n14182), .ZN(n14184) );
  AOI21_X1 U16097 ( .B1(n14185), .B2(n14670), .A(n14184), .ZN(n14186) );
  OAI21_X1 U16098 ( .B1(n14252), .B2(n14673), .A(n14186), .ZN(n14187) );
  AOI21_X1 U16099 ( .B1(n14256), .B2(n14188), .A(n14187), .ZN(n14189) );
  OAI21_X1 U16100 ( .B1(n14190), .B2(n14678), .A(n14189), .ZN(P1_U3274) );
  MUX2_X1 U16101 ( .A(n14193), .B(n14281), .S(n14764), .Z(n14194) );
  OAI21_X1 U16102 ( .B1(n14284), .B2(n14273), .A(n14194), .ZN(P1_U3559) );
  NAND2_X1 U16103 ( .A1(n14196), .A2(n14195), .ZN(n14285) );
  MUX2_X1 U16104 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14285), .S(n14764), .Z(
        n14197) );
  INV_X1 U16105 ( .A(n14197), .ZN(n14198) );
  OAI21_X1 U16106 ( .B1(n14288), .B2(n14273), .A(n14198), .ZN(P1_U3558) );
  AOI21_X1 U16107 ( .B1(n14743), .B2(n14200), .A(n14199), .ZN(n14201) );
  OAI211_X1 U16108 ( .C1(n14203), .C2(n14280), .A(n14202), .B(n14201), .ZN(
        n14289) );
  MUX2_X1 U16109 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14289), .S(n14764), .Z(
        P1_U3556) );
  INV_X1 U16110 ( .A(n14221), .ZN(n14716) );
  MUX2_X1 U16111 ( .A(n14207), .B(n14290), .S(n14764), .Z(n14208) );
  OAI21_X1 U16112 ( .B1(n14292), .B2(n14273), .A(n14208), .ZN(P1_U3555) );
  NAND2_X1 U16113 ( .A1(n14209), .A2(n14752), .ZN(n14211) );
  NAND4_X1 U16114 ( .A1(n14213), .A2(n14212), .A3(n14211), .A4(n14210), .ZN(
        n14293) );
  MUX2_X1 U16115 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14293), .S(n14764), .Z(
        P1_U3554) );
  OAI211_X1 U16116 ( .C1(n14216), .C2(n14280), .A(n14215), .B(n14214), .ZN(
        n14294) );
  MUX2_X1 U16117 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14294), .S(n14764), .Z(
        n14217) );
  INV_X1 U16118 ( .A(n14217), .ZN(n14218) );
  OAI21_X1 U16119 ( .B1(n14297), .B2(n14273), .A(n14218), .ZN(P1_U3553) );
  OAI211_X1 U16120 ( .C1(n14222), .C2(n14221), .A(n14220), .B(n14219), .ZN(
        n14223) );
  OR2_X1 U16121 ( .A1(n14224), .A2(n14223), .ZN(n14298) );
  MUX2_X1 U16122 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14298), .S(n14764), .Z(
        P1_U3552) );
  NAND3_X1 U16123 ( .A1(n14227), .A2(n14226), .A3(n14225), .ZN(n14228) );
  AOI211_X1 U16124 ( .C1(n14230), .C2(n14752), .A(n14229), .B(n14228), .ZN(
        n14231) );
  INV_X1 U16125 ( .A(n14231), .ZN(n14299) );
  MUX2_X1 U16126 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14299), .S(n14764), .Z(
        P1_U3551) );
  OAI211_X1 U16127 ( .C1(n14731), .C2(n14234), .A(n14233), .B(n14232), .ZN(
        n14236) );
  AOI211_X1 U16128 ( .C1(n14752), .C2(n14237), .A(n14236), .B(n14235), .ZN(
        n14238) );
  INV_X1 U16129 ( .A(n14238), .ZN(n14300) );
  MUX2_X1 U16130 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14300), .S(n14764), .Z(
        P1_U3550) );
  NAND2_X1 U16131 ( .A1(n14242), .A2(n14752), .ZN(n14243) );
  NAND2_X1 U16132 ( .A1(n7574), .A2(n14243), .ZN(n14301) );
  MUX2_X1 U16133 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14301), .S(n14764), .Z(
        n14244) );
  AOI21_X1 U16134 ( .B1(n14245), .B2(n14303), .A(n14244), .ZN(n14246) );
  INV_X1 U16135 ( .A(n14246), .ZN(P1_U3549) );
  AOI21_X1 U16136 ( .B1(n14743), .B2(n14248), .A(n14247), .ZN(n14249) );
  OAI211_X1 U16137 ( .C1(n14251), .C2(n14280), .A(n14250), .B(n14249), .ZN(
        n14306) );
  MUX2_X1 U16138 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14306), .S(n14764), .Z(
        P1_U3548) );
  INV_X1 U16139 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14257) );
  OAI21_X1 U16140 ( .B1(n14253), .B2(n14260), .A(n14252), .ZN(n14255) );
  AOI211_X1 U16141 ( .C1(n14752), .C2(n14256), .A(n14255), .B(n14254), .ZN(
        n14307) );
  MUX2_X1 U16142 ( .A(n14257), .B(n14307), .S(n14764), .Z(n14258) );
  OAI21_X1 U16143 ( .B1(n14310), .B2(n14273), .A(n14258), .ZN(P1_U3547) );
  INV_X1 U16144 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15345) );
  OAI21_X1 U16145 ( .B1(n14261), .B2(n14260), .A(n14259), .ZN(n14263) );
  AOI211_X1 U16146 ( .C1(n14264), .C2(n14752), .A(n14263), .B(n14262), .ZN(
        n14311) );
  MUX2_X1 U16147 ( .A(n15345), .B(n14311), .S(n14764), .Z(n14265) );
  OAI21_X1 U16148 ( .B1(n14314), .B2(n14273), .A(n14265), .ZN(P1_U3546) );
  NOR2_X1 U16149 ( .A1(n14266), .A2(n14280), .ZN(n14270) );
  NOR4_X1 U16150 ( .A1(n14270), .A2(n14269), .A3(n14268), .A4(n14267), .ZN(
        n14315) );
  MUX2_X1 U16151 ( .A(n14271), .B(n14315), .S(n14764), .Z(n14272) );
  OAI21_X1 U16152 ( .B1(n14319), .B2(n14273), .A(n14272), .ZN(P1_U3545) );
  INV_X1 U16153 ( .A(n14274), .ZN(n14279) );
  AOI21_X1 U16154 ( .B1(n14743), .B2(n14276), .A(n14275), .ZN(n14277) );
  OAI211_X1 U16155 ( .C1(n14280), .C2(n14279), .A(n14278), .B(n14277), .ZN(
        n14320) );
  MUX2_X1 U16156 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14320), .S(n14764), .Z(
        P1_U3544) );
  INV_X1 U16157 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14282) );
  MUX2_X1 U16158 ( .A(n14282), .B(n14281), .S(n14755), .Z(n14283) );
  OAI21_X1 U16159 ( .B1(n14284), .B2(n14318), .A(n14283), .ZN(P1_U3527) );
  MUX2_X1 U16160 ( .A(n14285), .B(P1_REG0_REG_30__SCAN_IN), .S(n14753), .Z(
        n14286) );
  INV_X1 U16161 ( .A(n14286), .ZN(n14287) );
  OAI21_X1 U16162 ( .B1(n14288), .B2(n14318), .A(n14287), .ZN(P1_U3526) );
  MUX2_X1 U16163 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14289), .S(n14755), .Z(
        P1_U3524) );
  OAI21_X1 U16164 ( .B1(n14292), .B2(n14318), .A(n14291), .ZN(P1_U3523) );
  MUX2_X1 U16165 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14293), .S(n14755), .Z(
        P1_U3522) );
  MUX2_X1 U16166 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14294), .S(n14755), .Z(
        n14295) );
  INV_X1 U16167 ( .A(n14295), .ZN(n14296) );
  OAI21_X1 U16168 ( .B1(n14297), .B2(n14318), .A(n14296), .ZN(P1_U3521) );
  MUX2_X1 U16169 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14298), .S(n14755), .Z(
        P1_U3520) );
  MUX2_X1 U16170 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14299), .S(n14755), .Z(
        P1_U3519) );
  MUX2_X1 U16171 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14300), .S(n14755), .Z(
        P1_U3518) );
  MUX2_X1 U16172 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14301), .S(n14755), .Z(
        n14302) );
  AOI21_X1 U16173 ( .B1(n14304), .B2(n14303), .A(n14302), .ZN(n14305) );
  INV_X1 U16174 ( .A(n14305), .ZN(P1_U3517) );
  MUX2_X1 U16175 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14306), .S(n14755), .Z(
        P1_U3516) );
  INV_X1 U16176 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14308) );
  MUX2_X1 U16177 ( .A(n14308), .B(n14307), .S(n14755), .Z(n14309) );
  OAI21_X1 U16178 ( .B1(n14310), .B2(n14318), .A(n14309), .ZN(P1_U3515) );
  INV_X1 U16179 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14312) );
  MUX2_X1 U16180 ( .A(n14312), .B(n14311), .S(n14755), .Z(n14313) );
  OAI21_X1 U16181 ( .B1(n14314), .B2(n14318), .A(n14313), .ZN(P1_U3513) );
  INV_X1 U16182 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14316) );
  MUX2_X1 U16183 ( .A(n14316), .B(n14315), .S(n14755), .Z(n14317) );
  OAI21_X1 U16184 ( .B1(n14319), .B2(n14318), .A(n14317), .ZN(P1_U3510) );
  MUX2_X1 U16185 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14320), .S(n14755), .Z(
        P1_U3507) );
  NOR4_X1 U16186 ( .A1(n14321), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8317), .A4(
        P1_U3086), .ZN(n14322) );
  AOI21_X1 U16187 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14323), .A(n14322), 
        .ZN(n14324) );
  OAI21_X1 U16188 ( .B1(n14325), .B2(n14330), .A(n14324), .ZN(P1_U3324) );
  OAI222_X1 U16189 ( .A1(n14332), .A2(n14331), .B1(n14330), .B2(n14329), .C1(
        P1_U3086), .C2(n6843), .ZN(P1_U3328) );
  MUX2_X1 U16190 ( .A(n14335), .B(n14334), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16191 ( .A(n14336), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16192 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14424) );
  XOR2_X1 U16193 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n14424), .Z(n14365) );
  INV_X1 U16194 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14364) );
  INV_X1 U16195 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14652) );
  NOR2_X1 U16196 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14652), .ZN(n14363) );
  INV_X1 U16197 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14362) );
  XOR2_X1 U16198 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n14362), .Z(n14366) );
  INV_X1 U16199 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15053) );
  XOR2_X1 U16200 ( .A(n15053), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14416) );
  INV_X1 U16201 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14355) );
  INV_X1 U16202 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14353) );
  XOR2_X1 U16203 ( .A(n14353), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14409) );
  INV_X1 U16204 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15009) );
  AOI22_X1 U16205 ( .A1(n14380), .A2(n14337), .B1(P3_ADDR_REG_1__SCAN_IN), 
        .B2(n14379), .ZN(n14377) );
  XNOR2_X1 U16206 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15391), .ZN(n14378) );
  NOR2_X1 U16207 ( .A1(n14340), .A2(n14339), .ZN(n14341) );
  NOR2_X1 U16208 ( .A1(n14344), .A2(n9716), .ZN(n14346) );
  NOR2_X1 U16209 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14392), .ZN(n14345) );
  INV_X1 U16210 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14396) );
  NOR2_X1 U16211 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14396), .ZN(n14347) );
  NOR2_X1 U16212 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14348), .ZN(n14350) );
  XNOR2_X1 U16213 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14348), .ZN(n14402) );
  NOR2_X1 U16214 ( .A1(n14402), .A2(n14403), .ZN(n14349) );
  XOR2_X1 U16215 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n14374) );
  NOR2_X1 U16216 ( .A1(n14375), .A2(n14374), .ZN(n14351) );
  NAND2_X1 U16217 ( .A1(n14409), .A2(n14408), .ZN(n14352) );
  XNOR2_X1 U16218 ( .A(n14355), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n14372) );
  NOR2_X1 U16219 ( .A1(n14373), .A2(n14372), .ZN(n14354) );
  XNOR2_X1 U16220 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n14356), .ZN(n14370) );
  NOR2_X1 U16221 ( .A1(n14371), .A2(n14370), .ZN(n14357) );
  NAND2_X1 U16222 ( .A1(n14416), .A2(n14415), .ZN(n14358) );
  INV_X1 U16223 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14359) );
  NAND2_X1 U16224 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14359), .ZN(n14360) );
  AOI22_X1 U16225 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n15445), .B1(n14368), 
        .B2(n14360), .ZN(n14367) );
  NAND2_X1 U16226 ( .A1(n14366), .A2(n14367), .ZN(n14361) );
  OAI22_X1 U16227 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14364), .B1(n14363), 
        .B2(n14420), .ZN(n14425) );
  XOR2_X1 U16228 ( .A(n14365), .B(n14425), .Z(n14423) );
  INV_X1 U16229 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14418) );
  XOR2_X1 U16230 ( .A(n14367), .B(n14366), .Z(n14631) );
  XOR2_X1 U16231 ( .A(n15445), .B(P3_ADDR_REG_13__SCAN_IN), .Z(n14369) );
  XNOR2_X1 U16232 ( .A(n14369), .B(n14368), .ZN(n14625) );
  XOR2_X1 U16233 ( .A(n14371), .B(n14370), .Z(n14617) );
  XOR2_X1 U16234 ( .A(n14373), .B(n14372), .Z(n14445) );
  XOR2_X1 U16235 ( .A(n14375), .B(n14374), .Z(n14407) );
  XNOR2_X1 U16236 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14376), .ZN(n14389) );
  NAND2_X1 U16237 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14389), .ZN(n14391) );
  XNOR2_X1 U16238 ( .A(n14378), .B(n14377), .ZN(n14385) );
  INV_X1 U16239 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15518) );
  OR2_X1 U16240 ( .A1(n15518), .A2(n14381), .ZN(n14383) );
  AOI21_X1 U16241 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14952), .A(n14380), .ZN(
        n15609) );
  INV_X1 U16242 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15608) );
  NOR2_X1 U16243 ( .A1(n15609), .A2(n15608), .ZN(n15617) );
  NAND2_X1 U16244 ( .A1(n15617), .A2(n15616), .ZN(n14382) );
  NAND2_X1 U16245 ( .A1(n14383), .A2(n14382), .ZN(n14384) );
  NOR2_X1 U16246 ( .A1(n14385), .A2(n14384), .ZN(n14438) );
  XNOR2_X1 U16247 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14386), .ZN(n15613) );
  NAND2_X1 U16248 ( .A1(n15614), .A2(n15613), .ZN(n14387) );
  AOI21_X1 U16249 ( .B1(n14388), .B2(n14387), .A(n15612), .ZN(n15606) );
  XOR2_X1 U16250 ( .A(n14389), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15605) );
  NAND2_X1 U16251 ( .A1(n15606), .A2(n15605), .ZN(n14390) );
  NAND2_X1 U16252 ( .A1(n14391), .A2(n14390), .ZN(n14395) );
  INV_X1 U16253 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14393) );
  XOR2_X1 U16254 ( .A(n14393), .B(n14392), .Z(n14394) );
  XOR2_X1 U16255 ( .A(n14396), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14398) );
  XOR2_X1 U16256 ( .A(n14398), .B(n14397), .Z(n14440) );
  NAND2_X1 U16257 ( .A1(n14399), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14400) );
  NAND2_X1 U16258 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14401), .ZN(n14405) );
  XOR2_X1 U16259 ( .A(n14403), .B(n14402), .Z(n15610) );
  NAND2_X1 U16260 ( .A1(n15611), .A2(n15610), .ZN(n14404) );
  XNOR2_X1 U16261 ( .A(n14409), .B(n14408), .ZN(n14411) );
  NAND2_X1 U16262 ( .A1(n14410), .A2(n14411), .ZN(n14412) );
  NOR2_X1 U16263 ( .A1(n14445), .A2(n14446), .ZN(n14413) );
  INV_X1 U16264 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14822) );
  NAND2_X1 U16265 ( .A1(n14445), .A2(n14446), .ZN(n14444) );
  XNOR2_X1 U16266 ( .A(n14416), .B(n14415), .ZN(n14621) );
  NAND2_X1 U16267 ( .A1(n14620), .A2(n14621), .ZN(n14619) );
  INV_X1 U16268 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14627) );
  NAND2_X1 U16269 ( .A1(n14631), .A2(n14630), .ZN(n14417) );
  XNOR2_X1 U16270 ( .A(n14652), .B(P3_ADDR_REG_15__SCAN_IN), .ZN(n14419) );
  XNOR2_X1 U16271 ( .A(n14420), .B(n14419), .ZN(n14635) );
  OR2_X1 U16272 ( .A1(n14634), .A2(n14635), .ZN(n14422) );
  NAND2_X1 U16273 ( .A1(n14634), .A2(n14635), .ZN(n14633) );
  INV_X1 U16274 ( .A(n14633), .ZN(n14421) );
  INV_X1 U16275 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14432) );
  AND2_X1 U16276 ( .A1(n14424), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n14426) );
  OAI22_X1 U16277 ( .A1(n14426), .A2(n14425), .B1(P3_ADDR_REG_16__SCAN_IN), 
        .B2(n14424), .ZN(n14430) );
  XNOR2_X1 U16278 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14430), .ZN(n14431) );
  XNOR2_X1 U16279 ( .A(n14432), .B(n14431), .ZN(n14428) );
  NOR2_X1 U16280 ( .A1(n14427), .A2(n14428), .ZN(n14449) );
  NOR2_X1 U16281 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n14448), .ZN(n14429) );
  NOR2_X1 U16282 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14430), .ZN(n14434) );
  NOR2_X1 U16283 ( .A1(n14432), .A2(n14431), .ZN(n14433) );
  NOR2_X1 U16284 ( .A1(n14434), .A2(n14433), .ZN(n14455) );
  INV_X1 U16285 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14457) );
  XNOR2_X1 U16286 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n14457), .ZN(n14454) );
  XNOR2_X1 U16287 ( .A(n14455), .B(n14454), .ZN(n14452) );
  XNOR2_X1 U16288 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14451), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16289 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14435) );
  OAI21_X1 U16290 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14435), 
        .ZN(U28) );
  AOI21_X1 U16291 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14436) );
  OAI21_X1 U16292 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14436), 
        .ZN(U29) );
  NOR2_X1 U16293 ( .A1(n14438), .A2(n14437), .ZN(n14439) );
  XOR2_X1 U16294 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n14439), .Z(SUB_1596_U61) );
  XOR2_X1 U16295 ( .A(n14441), .B(n14440), .Z(SUB_1596_U57) );
  XNOR2_X1 U16296 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14442), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16297 ( .A(n14443), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  OAI21_X1 U16298 ( .B1(n14446), .B2(n14445), .A(n14444), .ZN(n14447) );
  XOR2_X1 U16299 ( .A(n14447), .B(n14822), .Z(SUB_1596_U70) );
  NOR2_X1 U16300 ( .A1(n14449), .A2(n14448), .ZN(n14450) );
  XOR2_X1 U16301 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14450), .Z(SUB_1596_U63)
         );
  NOR2_X1 U16302 ( .A1(n14455), .A2(n14454), .ZN(n14456) );
  AOI21_X1 U16303 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14457), .A(n14456), 
        .ZN(n14461) );
  XNOR2_X1 U16304 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n14459) );
  XNOR2_X1 U16305 ( .A(n14459), .B(n14458), .ZN(n14460) );
  AOI21_X1 U16306 ( .B1(n14464), .B2(n14463), .A(n14462), .ZN(n14479) );
  OAI21_X1 U16307 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14466), .A(n14465), 
        .ZN(n14472) );
  NOR2_X1 U16308 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14467), .ZN(n14468) );
  AOI21_X1 U16309 ( .B1(n15095), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n14468), 
        .ZN(n14469) );
  OAI21_X1 U16310 ( .B1(n15092), .B2(n14470), .A(n14469), .ZN(n14471) );
  AOI21_X1 U16311 ( .B1(n14472), .B2(n15087), .A(n14471), .ZN(n14478) );
  NOR2_X1 U16312 ( .A1(n14474), .A2(n14473), .ZN(n14475) );
  OAI21_X1 U16313 ( .B1(n14476), .B2(n14475), .A(n15096), .ZN(n14477) );
  OAI211_X1 U16314 ( .C1(n14479), .C2(n15102), .A(n14478), .B(n14477), .ZN(
        P3_U3197) );
  AOI22_X1 U16315 ( .A1(n14999), .A2(n14480), .B1(n15095), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14496) );
  INV_X1 U16316 ( .A(n14481), .ZN(n14482) );
  NAND2_X1 U16317 ( .A1(n14483), .A2(n14482), .ZN(n14484) );
  XNOR2_X1 U16318 ( .A(n14485), .B(n14484), .ZN(n14490) );
  OAI21_X1 U16319 ( .B1(n14488), .B2(n14487), .A(n14486), .ZN(n14489) );
  AOI22_X1 U16320 ( .A1(n14490), .A2(n15096), .B1(n15087), .B2(n14489), .ZN(
        n14495) );
  NAND2_X1 U16321 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14494)
         );
  OAI221_X1 U16322 ( .B1(n14492), .B2(n6780), .C1(n14492), .C2(n14491), .A(
        n14520), .ZN(n14493) );
  NAND4_X1 U16323 ( .A1(n14496), .A2(n14495), .A3(n14494), .A4(n14493), .ZN(
        P3_U3198) );
  AOI22_X1 U16324 ( .A1(n14999), .A2(n14497), .B1(n15095), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14510) );
  OAI21_X1 U16325 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14499), .A(n14498), 
        .ZN(n14504) );
  AOI211_X1 U16326 ( .C1(n14502), .C2(n14501), .A(n14500), .B(n15077), .ZN(
        n14503) );
  AOI21_X1 U16327 ( .B1(n15087), .B2(n14504), .A(n14503), .ZN(n14509) );
  NAND2_X1 U16328 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14508)
         );
  OAI221_X1 U16329 ( .B1(n14506), .B2(n15481), .C1(n14506), .C2(n14505), .A(
        n14520), .ZN(n14507) );
  NAND4_X1 U16330 ( .A1(n14510), .A2(n14509), .A3(n14508), .A4(n14507), .ZN(
        P3_U3199) );
  AOI22_X1 U16331 ( .A1(n14999), .A2(n14511), .B1(n15095), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14527) );
  OAI21_X1 U16332 ( .B1(n14514), .B2(n14513), .A(n14512), .ZN(n14519) );
  OAI21_X1 U16333 ( .B1(n14517), .B2(n14516), .A(n14515), .ZN(n14518) );
  AOI22_X1 U16334 ( .A1(n14519), .A2(n15087), .B1(n15096), .B2(n14518), .ZN(
        n14526) );
  NAND2_X1 U16335 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n14525)
         );
  OAI221_X1 U16336 ( .B1(n14523), .B2(n14522), .C1(n14523), .C2(n14521), .A(
        n14520), .ZN(n14524) );
  NAND4_X1 U16337 ( .A1(n14527), .A2(n14526), .A3(n14525), .A4(n14524), .ZN(
        P3_U3200) );
  AOI22_X1 U16338 ( .A1(n14532), .A2(n14528), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15146), .ZN(n14529) );
  NAND2_X1 U16339 ( .A1(n14530), .A2(n14529), .ZN(P3_U3203) );
  AOI21_X1 U16340 ( .B1(n14532), .B2(n15193), .A(n14531), .ZN(n14543) );
  INV_X1 U16341 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14533) );
  AOI22_X1 U16342 ( .A1(n15213), .A2(n14543), .B1(n14533), .B2(n15210), .ZN(
        P3_U3489) );
  OAI21_X1 U16343 ( .B1(n15182), .B2(n14535), .A(n14534), .ZN(n14536) );
  AOI21_X1 U16344 ( .B1(n14537), .B2(n15187), .A(n14536), .ZN(n14545) );
  AOI22_X1 U16345 ( .A1(n15213), .A2(n14545), .B1(n15434), .B2(n15210), .ZN(
        P3_U3471) );
  OAI22_X1 U16346 ( .A1(n14539), .A2(n15172), .B1(n14538), .B2(n15182), .ZN(
        n14541) );
  NOR2_X1 U16347 ( .A1(n14541), .A2(n14540), .ZN(n14547) );
  INV_X1 U16348 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14542) );
  AOI22_X1 U16349 ( .A1(n15213), .A2(n14547), .B1(n14542), .B2(n15210), .ZN(
        P3_U3470) );
  INV_X1 U16350 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n15333) );
  AOI22_X1 U16351 ( .A1(n15197), .A2(n14543), .B1(n15333), .B2(n15195), .ZN(
        P3_U3457) );
  INV_X1 U16352 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14544) );
  AOI22_X1 U16353 ( .A1(n15197), .A2(n14545), .B1(n14544), .B2(n15195), .ZN(
        P3_U3426) );
  INV_X1 U16354 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14546) );
  AOI22_X1 U16355 ( .A1(n15197), .A2(n14547), .B1(n14546), .B2(n15195), .ZN(
        P3_U3423) );
  AOI21_X1 U16356 ( .B1(n14549), .B2(n14559), .A(n14548), .ZN(n14553) );
  INV_X1 U16357 ( .A(n14550), .ZN(n14551) );
  AOI21_X1 U16358 ( .B1(n14553), .B2(n14552), .A(n14551), .ZN(n14572) );
  AOI222_X1 U16359 ( .A1(n14558), .A2(n14557), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n14556), .C1(n14555), .C2(n14554), .ZN(n14565) );
  XNOR2_X1 U16360 ( .A(n14560), .B(n14559), .ZN(n14575) );
  OAI211_X1 U16361 ( .C1(n14573), .C2(n6810), .A(n10936), .B(n14561), .ZN(
        n14571) );
  INV_X1 U16362 ( .A(n14571), .ZN(n14562) );
  AOI22_X1 U16363 ( .A1(n14575), .A2(n14563), .B1(n15590), .B2(n14562), .ZN(
        n14564) );
  OAI211_X1 U16364 ( .C1(n15599), .C2(n14572), .A(n14565), .B(n14564), .ZN(
        P2_U3253) );
  OAI21_X1 U16365 ( .B1(n7075), .B2(n14909), .A(n14566), .ZN(n14568) );
  AOI211_X1 U16366 ( .C1(n14870), .C2(n14569), .A(n14568), .B(n14567), .ZN(
        n14577) );
  AOI22_X1 U16367 ( .A1(n14943), .A2(n14577), .B1(n14570), .B2(n14940), .ZN(
        P2_U3512) );
  OAI211_X1 U16368 ( .C1(n14573), .C2(n14909), .A(n14572), .B(n14571), .ZN(
        n14574) );
  AOI21_X1 U16369 ( .B1(n14870), .B2(n14575), .A(n14574), .ZN(n14579) );
  AOI22_X1 U16370 ( .A1(n14943), .A2(n14579), .B1(n14576), .B2(n14940), .ZN(
        P2_U3511) );
  AOI22_X1 U16371 ( .A1(n14925), .A2(n14577), .B1(n10759), .B2(n14923), .ZN(
        P2_U3469) );
  INV_X1 U16372 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14578) );
  AOI22_X1 U16373 ( .A1(n14925), .A2(n14579), .B1(n14578), .B2(n14923), .ZN(
        P2_U3466) );
  AOI21_X1 U16374 ( .B1(n14582), .B2(n14581), .A(n14580), .ZN(n14583) );
  INV_X1 U16375 ( .A(n14583), .ZN(n14586) );
  AOI222_X1 U16376 ( .A1(n14588), .A2(n14587), .B1(n14586), .B2(n14585), .C1(
        n14584), .C2(n14602), .ZN(n14590) );
  OAI211_X1 U16377 ( .C1(n14606), .C2(n14591), .A(n14590), .B(n14589), .ZN(
        P1_U3215) );
  OAI22_X1 U16378 ( .A1(n14595), .A2(n14594), .B1(n14593), .B2(n14592), .ZN(
        n14601) );
  AOI21_X1 U16379 ( .B1(n14597), .B2(n14596), .A(n6799), .ZN(n14599) );
  NOR2_X1 U16380 ( .A1(n14599), .A2(n14598), .ZN(n14600) );
  AOI211_X1 U16381 ( .C1(n14602), .C2(n14607), .A(n14601), .B(n14600), .ZN(
        n14604) );
  OAI211_X1 U16382 ( .C1(n14606), .C2(n14605), .A(n14604), .B(n14603), .ZN(
        P1_U3236) );
  INV_X1 U16383 ( .A(n14607), .ZN(n14609) );
  OAI21_X1 U16384 ( .B1(n14609), .B2(n14731), .A(n14608), .ZN(n14611) );
  AOI211_X1 U16385 ( .C1(n14752), .C2(n14612), .A(n14611), .B(n14610), .ZN(
        n14614) );
  AOI22_X1 U16386 ( .A1(n14764), .A2(n14614), .B1(n8510), .B2(n14761), .ZN(
        P1_U3539) );
  INV_X1 U16387 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14613) );
  AOI22_X1 U16388 ( .A1(n14755), .A2(n14614), .B1(n14613), .B2(n14753), .ZN(
        P1_U3492) );
  AOI21_X1 U16389 ( .B1(n14617), .B2(n14616), .A(n14615), .ZN(n14618) );
  XOR2_X1 U16390 ( .A(n14618), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16391 ( .B1(n14621), .B2(n14620), .A(n14619), .ZN(n14623) );
  XOR2_X1 U16392 ( .A(n14623), .B(n14622), .Z(SUB_1596_U68) );
  OAI21_X1 U16393 ( .B1(n14626), .B2(n14625), .A(n14624), .ZN(n14628) );
  XOR2_X1 U16394 ( .A(n14628), .B(n14627), .Z(SUB_1596_U67) );
  AOI21_X1 U16395 ( .B1(n14631), .B2(n14630), .A(n14629), .ZN(n14632) );
  XOR2_X1 U16396 ( .A(n14632), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  OAI21_X1 U16397 ( .B1(n14635), .B2(n14634), .A(n14633), .ZN(n14636) );
  XNOR2_X1 U16398 ( .A(n14636), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  NOR2_X1 U16399 ( .A1(n6757), .A2(n6670), .ZN(n14637) );
  XOR2_X1 U16400 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14637), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16401 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14639), .A(n14638), 
        .ZN(n14644) );
  AOI21_X1 U16402 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14641), .A(n14640), 
        .ZN(n14642) );
  OAI222_X1 U16403 ( .A1(n14647), .A2(n14646), .B1(n14645), .B2(n14644), .C1(
        n14643), .C2(n14642), .ZN(n14648) );
  INV_X1 U16404 ( .A(n14648), .ZN(n14650) );
  OAI211_X1 U16405 ( .C1(n14652), .C2(n14651), .A(n14650), .B(n14649), .ZN(
        P1_U3258) );
  OAI21_X1 U16406 ( .B1(n14654), .B2(n7361), .A(n14653), .ZN(n14741) );
  INV_X1 U16407 ( .A(n14737), .ZN(n14659) );
  NAND2_X1 U16408 ( .A1(n14655), .A2(n7361), .ZN(n14657) );
  AOI21_X1 U16409 ( .B1(n14658), .B2(n14657), .A(n14656), .ZN(n14739) );
  AOI211_X1 U16410 ( .C1(n14660), .C2(n14741), .A(n14659), .B(n14739), .ZN(
        n14677) );
  AOI21_X1 U16411 ( .B1(n14662), .B2(n14671), .A(n14661), .ZN(n14664) );
  NAND2_X1 U16412 ( .A1(n14664), .A2(n14663), .ZN(n14738) );
  OAI22_X1 U16413 ( .A1(n14668), .A2(n14667), .B1(n14666), .B2(n14665), .ZN(
        n14669) );
  AOI21_X1 U16414 ( .B1(n14671), .B2(n14670), .A(n14669), .ZN(n14672) );
  OAI21_X1 U16415 ( .B1(n14738), .B2(n14673), .A(n14672), .ZN(n14674) );
  AOI21_X1 U16416 ( .B1(n14741), .B2(n14675), .A(n14674), .ZN(n14676) );
  OAI21_X1 U16417 ( .B1(n14678), .B2(n14677), .A(n14676), .ZN(P1_U3284) );
  INV_X1 U16418 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14679) );
  NOR2_X1 U16419 ( .A1(n14706), .A2(n14679), .ZN(P1_U3294) );
  INV_X1 U16420 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15326) );
  NOR2_X1 U16421 ( .A1(n14706), .A2(n15326), .ZN(P1_U3295) );
  INV_X1 U16422 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14680) );
  NOR2_X1 U16423 ( .A1(n14706), .A2(n14680), .ZN(P1_U3296) );
  INV_X1 U16424 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14681) );
  NOR2_X1 U16425 ( .A1(n14706), .A2(n14681), .ZN(P1_U3297) );
  INV_X1 U16426 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14682) );
  NOR2_X1 U16427 ( .A1(n14706), .A2(n14682), .ZN(P1_U3298) );
  INV_X1 U16428 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14683) );
  NOR2_X1 U16429 ( .A1(n14706), .A2(n14683), .ZN(P1_U3299) );
  INV_X1 U16430 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15363) );
  NOR2_X1 U16431 ( .A1(n14706), .A2(n15363), .ZN(P1_U3300) );
  INV_X1 U16432 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14684) );
  NOR2_X1 U16433 ( .A1(n14706), .A2(n14684), .ZN(P1_U3301) );
  INV_X1 U16434 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14685) );
  NOR2_X1 U16435 ( .A1(n14706), .A2(n14685), .ZN(P1_U3302) );
  INV_X1 U16436 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14686) );
  NOR2_X1 U16437 ( .A1(n14706), .A2(n14686), .ZN(P1_U3303) );
  INV_X1 U16438 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14687) );
  NOR2_X1 U16439 ( .A1(n14706), .A2(n14687), .ZN(P1_U3304) );
  INV_X1 U16440 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14688) );
  NOR2_X1 U16441 ( .A1(n14706), .A2(n14688), .ZN(P1_U3305) );
  INV_X1 U16442 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14689) );
  NOR2_X1 U16443 ( .A1(n14706), .A2(n14689), .ZN(P1_U3306) );
  INV_X1 U16444 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14690) );
  NOR2_X1 U16445 ( .A1(n14706), .A2(n14690), .ZN(P1_U3307) );
  INV_X1 U16446 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14691) );
  NOR2_X1 U16447 ( .A1(n14706), .A2(n14691), .ZN(P1_U3308) );
  INV_X1 U16448 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14692) );
  NOR2_X1 U16449 ( .A1(n14706), .A2(n14692), .ZN(P1_U3309) );
  INV_X1 U16450 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14693) );
  NOR2_X1 U16451 ( .A1(n14706), .A2(n14693), .ZN(P1_U3310) );
  INV_X1 U16452 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14694) );
  NOR2_X1 U16453 ( .A1(n14706), .A2(n14694), .ZN(P1_U3311) );
  INV_X1 U16454 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14695) );
  NOR2_X1 U16455 ( .A1(n14706), .A2(n14695), .ZN(P1_U3312) );
  INV_X1 U16456 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14696) );
  NOR2_X1 U16457 ( .A1(n14706), .A2(n14696), .ZN(P1_U3313) );
  INV_X1 U16458 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14697) );
  NOR2_X1 U16459 ( .A1(n14706), .A2(n14697), .ZN(P1_U3314) );
  INV_X1 U16460 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14698) );
  NOR2_X1 U16461 ( .A1(n14706), .A2(n14698), .ZN(P1_U3315) );
  INV_X1 U16462 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14699) );
  NOR2_X1 U16463 ( .A1(n14706), .A2(n14699), .ZN(P1_U3316) );
  INV_X1 U16464 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15463) );
  NOR2_X1 U16465 ( .A1(n14706), .A2(n15463), .ZN(P1_U3317) );
  INV_X1 U16466 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14700) );
  NOR2_X1 U16467 ( .A1(n14706), .A2(n14700), .ZN(P1_U3318) );
  INV_X1 U16468 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14701) );
  NOR2_X1 U16469 ( .A1(n14706), .A2(n14701), .ZN(P1_U3319) );
  INV_X1 U16470 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14702) );
  NOR2_X1 U16471 ( .A1(n14706), .A2(n14702), .ZN(P1_U3320) );
  INV_X1 U16472 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14703) );
  NOR2_X1 U16473 ( .A1(n14706), .A2(n14703), .ZN(P1_U3321) );
  INV_X1 U16474 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14704) );
  NOR2_X1 U16475 ( .A1(n14706), .A2(n14704), .ZN(P1_U3322) );
  INV_X1 U16476 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14705) );
  NOR2_X1 U16477 ( .A1(n14706), .A2(n14705), .ZN(P1_U3323) );
  OAI21_X1 U16478 ( .B1(n14708), .B2(n14731), .A(n14707), .ZN(n14710) );
  AOI211_X1 U16479 ( .C1(n14716), .C2(n14711), .A(n14710), .B(n14709), .ZN(
        n14756) );
  INV_X1 U16480 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14712) );
  AOI22_X1 U16481 ( .A1(n14755), .A2(n14756), .B1(n14712), .B2(n14753), .ZN(
        P1_U3462) );
  OAI21_X1 U16482 ( .B1(n14714), .B2(n14731), .A(n14713), .ZN(n14715) );
  AOI21_X1 U16483 ( .B1(n14717), .B2(n14716), .A(n14715), .ZN(n14718) );
  AND2_X1 U16484 ( .A1(n14719), .A2(n14718), .ZN(n14757) );
  INV_X1 U16485 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14720) );
  AOI22_X1 U16486 ( .A1(n14755), .A2(n14757), .B1(n14720), .B2(n14753), .ZN(
        P1_U3465) );
  AOI21_X1 U16487 ( .B1(n14743), .B2(n14722), .A(n14721), .ZN(n14724) );
  NAND3_X1 U16488 ( .A1(n14725), .A2(n14724), .A3(n14723), .ZN(n14726) );
  AOI21_X1 U16489 ( .B1(n14752), .B2(n14727), .A(n14726), .ZN(n14758) );
  INV_X1 U16490 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14728) );
  AOI22_X1 U16491 ( .A1(n14755), .A2(n14758), .B1(n14728), .B2(n14753), .ZN(
        P1_U3471) );
  OAI211_X1 U16492 ( .C1(n14732), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        n14733) );
  AOI21_X1 U16493 ( .B1(n14752), .B2(n14734), .A(n14733), .ZN(n14759) );
  INV_X1 U16494 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14735) );
  AOI22_X1 U16495 ( .A1(n14755), .A2(n14759), .B1(n14735), .B2(n14753), .ZN(
        P1_U3477) );
  NAND3_X1 U16496 ( .A1(n14738), .A2(n14737), .A3(n14736), .ZN(n14740) );
  AOI211_X1 U16497 ( .C1(n14752), .C2(n14741), .A(n14740), .B(n14739), .ZN(
        n14760) );
  INV_X1 U16498 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14742) );
  AOI22_X1 U16499 ( .A1(n14755), .A2(n14760), .B1(n14742), .B2(n14753), .ZN(
        P1_U3486) );
  NAND2_X1 U16500 ( .A1(n14744), .A2(n14743), .ZN(n14745) );
  NAND4_X1 U16501 ( .A1(n14748), .A2(n14747), .A3(n14746), .A4(n14745), .ZN(
        n14750) );
  AOI211_X1 U16502 ( .C1(n14752), .C2(n14751), .A(n14750), .B(n14749), .ZN(
        n14763) );
  INV_X1 U16503 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14754) );
  AOI22_X1 U16504 ( .A1(n14755), .A2(n14763), .B1(n14754), .B2(n14753), .ZN(
        P1_U3489) );
  AOI22_X1 U16505 ( .A1(n14764), .A2(n14756), .B1(n9093), .B2(n14761), .ZN(
        P1_U3529) );
  AOI22_X1 U16506 ( .A1(n14764), .A2(n14757), .B1(n9122), .B2(n14761), .ZN(
        P1_U3530) );
  AOI22_X1 U16507 ( .A1(n14764), .A2(n14758), .B1(n8399), .B2(n14761), .ZN(
        P1_U3532) );
  AOI22_X1 U16508 ( .A1(n14764), .A2(n14759), .B1(n9198), .B2(n14761), .ZN(
        P1_U3534) );
  AOI22_X1 U16509 ( .A1(n14764), .A2(n14760), .B1(n8478), .B2(n14761), .ZN(
        P1_U3537) );
  AOI22_X1 U16510 ( .A1(n14764), .A2(n14763), .B1(n14762), .B2(n14761), .ZN(
        P1_U3538) );
  NOR2_X1 U16511 ( .A1(n14835), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI22_X1 U16512 ( .A1(n14765), .A2(n9562), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10146), .ZN(n14766) );
  AOI21_X1 U16513 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n14835), .A(n14766), .ZN(
        n14778) );
  AOI211_X1 U16514 ( .C1(n14769), .C2(n14768), .A(n14767), .B(n14798), .ZN(
        n14770) );
  INV_X1 U16515 ( .A(n14770), .ZN(n14777) );
  AND2_X1 U16516 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14775) );
  INV_X1 U16517 ( .A(n14771), .ZN(n14774) );
  INV_X1 U16518 ( .A(n14772), .ZN(n14773) );
  OAI211_X1 U16519 ( .C1(n14775), .C2(n14774), .A(n14837), .B(n14773), .ZN(
        n14776) );
  NAND3_X1 U16520 ( .A1(n14778), .A2(n14777), .A3(n14776), .ZN(P2_U3215) );
  INV_X1 U16521 ( .A(n14779), .ZN(n14795) );
  OAI21_X1 U16522 ( .B1(n14795), .B2(n14780), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14781) );
  OAI21_X1 U16523 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14781), .ZN(n14793) );
  AOI211_X1 U16524 ( .C1(n14784), .C2(n14783), .A(n14782), .B(n14798), .ZN(
        n14785) );
  INV_X1 U16525 ( .A(n14785), .ZN(n14792) );
  AOI211_X1 U16526 ( .C1(n14788), .C2(n14787), .A(n14786), .B(n14811), .ZN(
        n14789) );
  INV_X1 U16527 ( .A(n14789), .ZN(n14791) );
  NAND2_X1 U16528 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n14835), .ZN(n14790) );
  NAND4_X1 U16529 ( .A1(n14793), .A2(n14792), .A3(n14791), .A4(n14790), .ZN(
        P2_U3216) );
  OAI21_X1 U16530 ( .B1(n14795), .B2(n14794), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14796) );
  OAI21_X1 U16531 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14796), .ZN(n14809) );
  AOI211_X1 U16532 ( .C1(n14800), .C2(n14799), .A(n14798), .B(n14797), .ZN(
        n14801) );
  INV_X1 U16533 ( .A(n14801), .ZN(n14808) );
  NAND2_X1 U16534 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n14835), .ZN(n14807) );
  AOI211_X1 U16535 ( .C1(n14804), .C2(n14803), .A(n14811), .B(n14802), .ZN(
        n14805) );
  INV_X1 U16536 ( .A(n14805), .ZN(n14806) );
  NAND4_X1 U16537 ( .A1(n14809), .A2(n14808), .A3(n14807), .A4(n14806), .ZN(
        P2_U3220) );
  AOI211_X1 U16538 ( .C1(n14813), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        n14814) );
  AOI211_X1 U16539 ( .C1(n14841), .C2(n14816), .A(n14815), .B(n14814), .ZN(
        n14821) );
  OAI211_X1 U16540 ( .C1(n14819), .C2(n14818), .A(n14817), .B(n14843), .ZN(
        n14820) );
  OAI211_X1 U16541 ( .C1(n14823), .C2(n14822), .A(n14821), .B(n14820), .ZN(
        P2_U3224) );
  AOI22_X1 U16542 ( .A1(n14835), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14834) );
  OAI211_X1 U16543 ( .C1(n14826), .C2(n14825), .A(n14824), .B(n14843), .ZN(
        n14833) );
  OAI211_X1 U16544 ( .C1(n14829), .C2(n14828), .A(n14827), .B(n14837), .ZN(
        n14832) );
  NAND2_X1 U16545 ( .A1(n14841), .A2(n14830), .ZN(n14831) );
  NAND4_X1 U16546 ( .A1(n14834), .A2(n14833), .A3(n14832), .A4(n14831), .ZN(
        P2_U3227) );
  AOI22_X1 U16547 ( .A1(n14835), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14849) );
  OAI211_X1 U16548 ( .C1(n14839), .C2(n14838), .A(n14837), .B(n14836), .ZN(
        n14848) );
  NAND2_X1 U16549 ( .A1(n14841), .A2(n14840), .ZN(n14847) );
  OAI211_X1 U16550 ( .C1(n14845), .C2(n14844), .A(n14843), .B(n14842), .ZN(
        n14846) );
  NAND4_X1 U16551 ( .A1(n14849), .A2(n14848), .A3(n14847), .A4(n14846), .ZN(
        P2_U3231) );
  AND2_X1 U16552 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14852), .ZN(P2_U3266) );
  AND2_X1 U16553 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14852), .ZN(P2_U3267) );
  AND2_X1 U16554 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14852), .ZN(P2_U3268) );
  AND2_X1 U16555 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14852), .ZN(P2_U3269) );
  AND2_X1 U16556 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14852), .ZN(P2_U3270) );
  INV_X1 U16557 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15459) );
  NOR2_X1 U16558 ( .A1(n14851), .A2(n15459), .ZN(P2_U3271) );
  AND2_X1 U16559 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14852), .ZN(P2_U3272) );
  INV_X1 U16560 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15531) );
  NOR2_X1 U16561 ( .A1(n14851), .A2(n15531), .ZN(P2_U3273) );
  INV_X1 U16562 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15450) );
  NOR2_X1 U16563 ( .A1(n14851), .A2(n15450), .ZN(P2_U3274) );
  AND2_X1 U16564 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14852), .ZN(P2_U3275) );
  AND2_X1 U16565 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14852), .ZN(P2_U3276) );
  AND2_X1 U16566 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14852), .ZN(P2_U3277) );
  AND2_X1 U16567 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14852), .ZN(P2_U3278) );
  AND2_X1 U16568 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14852), .ZN(P2_U3279) );
  AND2_X1 U16569 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14852), .ZN(P2_U3280) );
  AND2_X1 U16570 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14852), .ZN(P2_U3281) );
  AND2_X1 U16571 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14852), .ZN(P2_U3282) );
  AND2_X1 U16572 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14852), .ZN(P2_U3283) );
  INV_X1 U16573 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15377) );
  NOR2_X1 U16574 ( .A1(n14851), .A2(n15377), .ZN(P2_U3284) );
  AND2_X1 U16575 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14852), .ZN(P2_U3285) );
  AND2_X1 U16576 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14852), .ZN(P2_U3286) );
  AND2_X1 U16577 ( .A1(n14852), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3287) );
  AND2_X1 U16578 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14852), .ZN(P2_U3288) );
  AND2_X1 U16579 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14852), .ZN(P2_U3289) );
  INV_X1 U16580 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15502) );
  NOR2_X1 U16581 ( .A1(n14851), .A2(n15502), .ZN(P2_U3290) );
  INV_X1 U16582 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15534) );
  NOR2_X1 U16583 ( .A1(n14851), .A2(n15534), .ZN(P2_U3291) );
  AND2_X1 U16584 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14852), .ZN(P2_U3292) );
  AND2_X1 U16585 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14852), .ZN(P2_U3293) );
  INV_X1 U16586 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15501) );
  NOR2_X1 U16587 ( .A1(n14851), .A2(n15501), .ZN(P2_U3294) );
  AND2_X1 U16588 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14852), .ZN(P2_U3295) );
  AOI21_X1 U16589 ( .B1(n14854), .B2(n14857), .A(n14853), .ZN(P2_U3416) );
  AOI21_X1 U16590 ( .B1(n14857), .B2(n14856), .A(n14855), .ZN(P2_U3417) );
  INV_X1 U16591 ( .A(n14858), .ZN(n14859) );
  AOI22_X1 U16592 ( .A1(n14925), .A2(n14859), .B1(n9465), .B2(n14923), .ZN(
        P2_U3430) );
  OAI21_X1 U16593 ( .B1(n9646), .B2(n14909), .A(n14860), .ZN(n14863) );
  INV_X1 U16594 ( .A(n14861), .ZN(n14862) );
  AOI211_X1 U16595 ( .C1(n14915), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14927) );
  AOI22_X1 U16596 ( .A1(n14925), .A2(n14927), .B1(n9573), .B2(n14923), .ZN(
        P2_U3436) );
  OAI21_X1 U16597 ( .B1(n14866), .B2(n14909), .A(n14865), .ZN(n14868) );
  AOI211_X1 U16598 ( .C1(n14870), .C2(n14869), .A(n14868), .B(n14867), .ZN(
        n14928) );
  INV_X1 U16599 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14871) );
  AOI22_X1 U16600 ( .A1(n14925), .A2(n14928), .B1(n14871), .B2(n14923), .ZN(
        P2_U3442) );
  OAI21_X1 U16601 ( .B1(n14873), .B2(n14915), .A(n14872), .ZN(n14878) );
  NAND2_X1 U16602 ( .A1(n14874), .A2(n14917), .ZN(n14876) );
  INV_X1 U16603 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14879) );
  AOI22_X1 U16604 ( .A1(n14925), .A2(n14930), .B1(n14879), .B2(n14923), .ZN(
        P2_U3445) );
  OAI21_X1 U16605 ( .B1(n14881), .B2(n14909), .A(n14880), .ZN(n14883) );
  AOI211_X1 U16606 ( .C1(n14915), .C2(n14884), .A(n14883), .B(n14882), .ZN(
        n14932) );
  INV_X1 U16607 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14885) );
  AOI22_X1 U16608 ( .A1(n14925), .A2(n14932), .B1(n14885), .B2(n14923), .ZN(
        P2_U3448) );
  AOI21_X1 U16609 ( .B1(n14917), .B2(n14887), .A(n14886), .ZN(n14889) );
  OAI211_X1 U16610 ( .C1(n14891), .C2(n14890), .A(n14889), .B(n14888), .ZN(
        n14892) );
  INV_X1 U16611 ( .A(n14892), .ZN(n14934) );
  INV_X1 U16612 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14893) );
  AOI22_X1 U16613 ( .A1(n14925), .A2(n14934), .B1(n14893), .B2(n14923), .ZN(
        P2_U3451) );
  INV_X1 U16614 ( .A(n14894), .ZN(n14898) );
  OAI21_X1 U16615 ( .B1(n7056), .B2(n14909), .A(n14895), .ZN(n14897) );
  AOI211_X1 U16616 ( .C1(n14915), .C2(n14898), .A(n14897), .B(n14896), .ZN(
        n14936) );
  INV_X1 U16617 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14899) );
  AOI22_X1 U16618 ( .A1(n14925), .A2(n14936), .B1(n14899), .B2(n14923), .ZN(
        P2_U3454) );
  INV_X1 U16619 ( .A(n14900), .ZN(n14905) );
  OAI21_X1 U16620 ( .B1(n14902), .B2(n14909), .A(n14901), .ZN(n14904) );
  AOI211_X1 U16621 ( .C1(n14915), .C2(n14905), .A(n14904), .B(n14903), .ZN(
        n14938) );
  INV_X1 U16622 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14906) );
  AOI22_X1 U16623 ( .A1(n14925), .A2(n14938), .B1(n14906), .B2(n14923), .ZN(
        P2_U3457) );
  INV_X1 U16624 ( .A(n14907), .ZN(n14913) );
  OAI21_X1 U16625 ( .B1(n14910), .B2(n14909), .A(n14908), .ZN(n14912) );
  AOI211_X1 U16626 ( .C1(n14915), .C2(n14913), .A(n14912), .B(n14911), .ZN(
        n14939) );
  INV_X1 U16627 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14914) );
  AOI22_X1 U16628 ( .A1(n14925), .A2(n14939), .B1(n14914), .B2(n14923), .ZN(
        P2_U3460) );
  AND2_X1 U16629 ( .A1(n14916), .A2(n14915), .ZN(n14921) );
  AND2_X1 U16630 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  NOR4_X1 U16631 ( .A1(n14922), .A2(n14921), .A3(n14920), .A4(n14919), .ZN(
        n14942) );
  INV_X1 U16632 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14924) );
  AOI22_X1 U16633 ( .A1(n14925), .A2(n14942), .B1(n14924), .B2(n14923), .ZN(
        P2_U3463) );
  AOI22_X1 U16634 ( .A1(n14943), .A2(n14927), .B1(n14926), .B2(n14940), .ZN(
        P2_U3501) );
  AOI22_X1 U16635 ( .A1(n14943), .A2(n14928), .B1(n15327), .B2(n14940), .ZN(
        P2_U3503) );
  AOI22_X1 U16636 ( .A1(n14943), .A2(n14930), .B1(n14929), .B2(n14940), .ZN(
        P2_U3504) );
  AOI22_X1 U16637 ( .A1(n14943), .A2(n14932), .B1(n14931), .B2(n14940), .ZN(
        P2_U3505) );
  AOI22_X1 U16638 ( .A1(n14943), .A2(n14934), .B1(n14933), .B2(n14940), .ZN(
        P2_U3506) );
  AOI22_X1 U16639 ( .A1(n14943), .A2(n14936), .B1(n14935), .B2(n14940), .ZN(
        P2_U3507) );
  AOI22_X1 U16640 ( .A1(n14943), .A2(n14938), .B1(n14937), .B2(n14940), .ZN(
        P2_U3508) );
  AOI22_X1 U16641 ( .A1(n14943), .A2(n14939), .B1(n9320), .B2(n14940), .ZN(
        P2_U3509) );
  AOI22_X1 U16642 ( .A1(n14943), .A2(n14942), .B1(n14941), .B2(n14940), .ZN(
        P2_U3510) );
  NOR2_X1 U16643 ( .A1(P3_U3897), .A2(n15095), .ZN(P3_U3150) );
  INV_X1 U16644 ( .A(n14944), .ZN(n14945) );
  AOI21_X1 U16645 ( .B1(n14999), .B2(P3_IR_REG_0__SCAN_IN), .A(n14945), .ZN(
        n14951) );
  NOR2_X1 U16646 ( .A1(n14946), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14948) );
  NAND3_X1 U16647 ( .A1(n15102), .A2(n15003), .A3(n15077), .ZN(n14947) );
  OAI21_X1 U16648 ( .B1(n14949), .B2(n14948), .A(n14947), .ZN(n14950) );
  OAI211_X1 U16649 ( .C1(n14952), .C2(n15054), .A(n14951), .B(n14950), .ZN(
        P3_U3182) );
  XNOR2_X1 U16650 ( .A(n14954), .B(n14953), .ZN(n14965) );
  NOR2_X1 U16651 ( .A1(n15092), .A2(n14955), .ZN(n14964) );
  AOI21_X1 U16652 ( .B1(n14958), .B2(n14957), .A(n14956), .ZN(n14962) );
  XOR2_X1 U16653 ( .A(n14960), .B(n14959), .Z(n14961) );
  OAI22_X1 U16654 ( .A1(n14962), .A2(n15102), .B1(n15003), .B2(n14961), .ZN(
        n14963) );
  AOI211_X1 U16655 ( .C1(n14965), .C2(n15096), .A(n14964), .B(n14963), .ZN(
        n14967) );
  OAI211_X1 U16656 ( .C1(n14968), .C2(n15054), .A(n14967), .B(n14966), .ZN(
        P3_U3186) );
  AOI21_X1 U16657 ( .B1(n14971), .B2(n14970), .A(n14969), .ZN(n14977) );
  OAI21_X1 U16658 ( .B1(n14974), .B2(n14973), .A(n14972), .ZN(n14975) );
  INV_X1 U16659 ( .A(n14975), .ZN(n14976) );
  OAI22_X1 U16660 ( .A1(n14977), .A2(n15102), .B1(n15003), .B2(n14976), .ZN(
        n14978) );
  INV_X1 U16661 ( .A(n14978), .ZN(n14984) );
  OAI21_X1 U16662 ( .B1(n14981), .B2(n14980), .A(n14979), .ZN(n14982) );
  NAND2_X1 U16663 ( .A1(n14982), .A2(n15096), .ZN(n14983) );
  OAI211_X1 U16664 ( .C1(n15092), .C2(n14985), .A(n14984), .B(n14983), .ZN(
        n14986) );
  INV_X1 U16665 ( .A(n14986), .ZN(n14988) );
  OAI211_X1 U16666 ( .C1(n14989), .C2(n15054), .A(n14988), .B(n14987), .ZN(
        P3_U3188) );
  AOI21_X1 U16667 ( .B1(n14992), .B2(n14991), .A(n14990), .ZN(n14993) );
  NOR2_X1 U16668 ( .A1(n14993), .A2(n15102), .ZN(n15006) );
  XOR2_X1 U16669 ( .A(n14995), .B(n14994), .Z(n15004) );
  OAI21_X1 U16670 ( .B1(n14998), .B2(n14997), .A(n14996), .ZN(n15001) );
  AOI22_X1 U16671 ( .A1(n15001), .A2(n15096), .B1(n15000), .B2(n14999), .ZN(
        n15002) );
  OAI21_X1 U16672 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n15005) );
  NOR2_X1 U16673 ( .A1(n15006), .A2(n15005), .ZN(n15008) );
  OAI211_X1 U16674 ( .C1(n15009), .C2(n15054), .A(n15008), .B(n15007), .ZN(
        P3_U3190) );
  AOI21_X1 U16675 ( .B1(n15012), .B2(n15011), .A(n15010), .ZN(n15026) );
  NAND2_X1 U16676 ( .A1(n15014), .A2(n15013), .ZN(n15015) );
  XNOR2_X1 U16677 ( .A(n15016), .B(n15015), .ZN(n15018) );
  OAI22_X1 U16678 ( .A1(n15018), .A2(n15077), .B1(n15017), .B2(n15092), .ZN(
        n15019) );
  AOI211_X1 U16679 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15095), .A(n15020), .B(
        n15019), .ZN(n15025) );
  OAI21_X1 U16680 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15022), .A(n15021), .ZN(
        n15023) );
  NAND2_X1 U16681 ( .A1(n15023), .A2(n15087), .ZN(n15024) );
  OAI211_X1 U16682 ( .C1(n15026), .C2(n15102), .A(n15025), .B(n15024), .ZN(
        P3_U3191) );
  AOI21_X1 U16683 ( .B1(n15498), .B2(n15028), .A(n15027), .ZN(n15042) );
  OAI21_X1 U16684 ( .B1(n15030), .B2(P3_REG1_REG_11__SCAN_IN), .A(n15029), 
        .ZN(n15035) );
  NOR2_X1 U16685 ( .A1(n15092), .A2(n15031), .ZN(n15034) );
  OAI21_X1 U16686 ( .B1(n15054), .B2(n15462), .A(n15032), .ZN(n15033) );
  AOI211_X1 U16687 ( .C1(n15035), .C2(n15087), .A(n15034), .B(n15033), .ZN(
        n15041) );
  AOI21_X1 U16688 ( .B1(n15038), .B2(n15037), .A(n15036), .ZN(n15039) );
  OR2_X1 U16689 ( .A1(n15039), .A2(n15077), .ZN(n15040) );
  OAI211_X1 U16690 ( .C1(n15042), .C2(n15102), .A(n15041), .B(n15040), .ZN(
        P3_U3193) );
  INV_X1 U16691 ( .A(n15044), .ZN(n15045) );
  AOI21_X1 U16692 ( .B1(n15047), .B2(n15046), .A(n15045), .ZN(n15063) );
  OAI21_X1 U16693 ( .B1(n15050), .B2(n15049), .A(n15048), .ZN(n15057) );
  NOR2_X1 U16694 ( .A1(n15092), .A2(n15051), .ZN(n15056) );
  OAI21_X1 U16695 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(n15055) );
  AOI211_X1 U16696 ( .C1(n15057), .C2(n15087), .A(n15056), .B(n15055), .ZN(
        n15062) );
  OAI211_X1 U16697 ( .C1(n15060), .C2(n15059), .A(n15058), .B(n15096), .ZN(
        n15061) );
  OAI211_X1 U16698 ( .C1(n15063), .C2(n15102), .A(n15062), .B(n15061), .ZN(
        P3_U3194) );
  AOI21_X1 U16699 ( .B1(n15066), .B2(n15065), .A(n15064), .ZN(n15081) );
  OAI21_X1 U16700 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15068), .A(n15067), 
        .ZN(n15073) );
  AND2_X1 U16701 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n15069) );
  AOI21_X1 U16702 ( .B1(n15095), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15069), 
        .ZN(n15070) );
  OAI21_X1 U16703 ( .B1(n15092), .B2(n15071), .A(n15070), .ZN(n15072) );
  AOI21_X1 U16704 ( .B1(n15073), .B2(n15087), .A(n15072), .ZN(n15080) );
  AOI21_X1 U16705 ( .B1(n15076), .B2(n15075), .A(n15074), .ZN(n15078) );
  OR2_X1 U16706 ( .A1(n15078), .A2(n15077), .ZN(n15079) );
  OAI211_X1 U16707 ( .C1(n15081), .C2(n15102), .A(n15080), .B(n15079), .ZN(
        P3_U3195) );
  AOI21_X1 U16708 ( .B1(n6791), .B2(n15083), .A(n15082), .ZN(n15103) );
  OAI21_X1 U16709 ( .B1(n15086), .B2(n15085), .A(n15084), .ZN(n15088) );
  AND2_X1 U16710 ( .A1(n15088), .A2(n15087), .ZN(n15094) );
  NAND2_X1 U16711 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n15090)
         );
  OAI21_X1 U16712 ( .B1(n15092), .B2(n15091), .A(n15090), .ZN(n15093) );
  AOI211_X1 U16713 ( .C1(P3_ADDR_REG_14__SCAN_IN), .C2(n15095), .A(n15094), 
        .B(n15093), .ZN(n15101) );
  OAI211_X1 U16714 ( .C1(n15099), .C2(n15098), .A(n15097), .B(n15096), .ZN(
        n15100) );
  OAI211_X1 U16715 ( .C1(n15103), .C2(n15102), .A(n15101), .B(n15100), .ZN(
        P3_U3196) );
  OAI21_X1 U16716 ( .B1(n15105), .B2(n15114), .A(n15104), .ZN(n15153) );
  NOR2_X1 U16717 ( .A1(n15106), .A2(n15182), .ZN(n15152) );
  INV_X1 U16718 ( .A(n15152), .ZN(n15110) );
  INV_X1 U16719 ( .A(n15137), .ZN(n15109) );
  OAI22_X1 U16720 ( .A1(n15110), .A2(n15109), .B1(n15108), .B2(n15107), .ZN(
        n15121) );
  OAI22_X1 U16721 ( .A1(n15112), .A2(n15134), .B1(n15111), .B2(n15136), .ZN(
        n15118) );
  NAND3_X1 U16722 ( .A1(n15127), .A2(n15114), .A3(n15113), .ZN(n15115) );
  AOI21_X1 U16723 ( .B1(n15116), .B2(n15115), .A(n15132), .ZN(n15117) );
  AOI211_X1 U16724 ( .C1(n15119), .C2(n15153), .A(n15118), .B(n15117), .ZN(
        n15120) );
  INV_X1 U16725 ( .A(n15120), .ZN(n15151) );
  AOI211_X1 U16726 ( .C1(n15122), .C2(n15153), .A(n15121), .B(n15151), .ZN(
        n15123) );
  AOI22_X1 U16727 ( .A1(n15146), .A2(n9524), .B1(n15123), .B2(n15144), .ZN(
        P3_U3231) );
  NOR2_X1 U16728 ( .A1(n15124), .A2(n15182), .ZN(n15148) );
  INV_X1 U16729 ( .A(n15125), .ZN(n15133) );
  INV_X1 U16730 ( .A(n15126), .ZN(n15129) );
  INV_X1 U16731 ( .A(n15127), .ZN(n15128) );
  AOI21_X1 U16732 ( .B1(n15130), .B2(n15129), .A(n15128), .ZN(n15131) );
  OAI222_X1 U16733 ( .A1(n15136), .A2(n15135), .B1(n15134), .B2(n15133), .C1(
        n15132), .C2(n15131), .ZN(n15147) );
  AOI21_X1 U16734 ( .B1(n15148), .B2(n15137), .A(n15147), .ZN(n15145) );
  XNOR2_X1 U16735 ( .A(n15139), .B(n15138), .ZN(n15149) );
  AOI22_X1 U16736 ( .A1(n15149), .A2(n15141), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15140), .ZN(n15142) );
  OAI221_X1 U16737 ( .B1(n15146), .B2(n15145), .C1(n15144), .C2(n15143), .A(
        n15142), .ZN(P3_U3232) );
  AOI211_X1 U16738 ( .C1(n15187), .C2(n15149), .A(n15148), .B(n15147), .ZN(
        n15198) );
  INV_X1 U16739 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15150) );
  AOI22_X1 U16740 ( .A1(n15197), .A2(n15198), .B1(n15150), .B2(n15195), .ZN(
        P3_U3393) );
  AOI211_X1 U16741 ( .C1(n15156), .C2(n15153), .A(n15152), .B(n15151), .ZN(
        n15199) );
  INV_X1 U16742 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U16743 ( .A1(n15197), .A2(n15199), .B1(n15154), .B2(n15195), .ZN(
        P3_U3396) );
  AOI22_X1 U16744 ( .A1(n15157), .A2(n15156), .B1(n15193), .B2(n15155), .ZN(
        n15158) );
  AND2_X1 U16745 ( .A1(n15159), .A2(n15158), .ZN(n15200) );
  INV_X1 U16746 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U16747 ( .A1(n15197), .A2(n15200), .B1(n15403), .B2(n15195), .ZN(
        P3_U3399) );
  OAI22_X1 U16748 ( .A1(n15161), .A2(n15189), .B1(n15182), .B2(n15160), .ZN(
        n15162) );
  NOR2_X1 U16749 ( .A1(n15163), .A2(n15162), .ZN(n15202) );
  INV_X1 U16750 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U16751 ( .A1(n15197), .A2(n15202), .B1(n15164), .B2(n15195), .ZN(
        P3_U3402) );
  AOI22_X1 U16752 ( .A1(n15166), .A2(n15187), .B1(n15193), .B2(n15165), .ZN(
        n15167) );
  AND2_X1 U16753 ( .A1(n15168), .A2(n15167), .ZN(n15204) );
  INV_X1 U16754 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U16755 ( .A1(n15197), .A2(n15204), .B1(n15169), .B2(n15195), .ZN(
        P3_U3405) );
  INV_X1 U16756 ( .A(n15170), .ZN(n15175) );
  OAI22_X1 U16757 ( .A1(n15173), .A2(n15172), .B1(n15171), .B2(n15182), .ZN(
        n15174) );
  NOR2_X1 U16758 ( .A1(n15175), .A2(n15174), .ZN(n15206) );
  INV_X1 U16759 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15176) );
  AOI22_X1 U16760 ( .A1(n15197), .A2(n15206), .B1(n15176), .B2(n15195), .ZN(
        P3_U3408) );
  OAI22_X1 U16761 ( .A1(n15178), .A2(n15189), .B1(n15182), .B2(n15177), .ZN(
        n15179) );
  NOR2_X1 U16762 ( .A1(n15180), .A2(n15179), .ZN(n15207) );
  INV_X1 U16763 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15181) );
  AOI22_X1 U16764 ( .A1(n15197), .A2(n15207), .B1(n15181), .B2(n15195), .ZN(
        P3_U3411) );
  NOR2_X1 U16765 ( .A1(n15183), .A2(n15182), .ZN(n15185) );
  AOI211_X1 U16766 ( .C1(n15187), .C2(n15186), .A(n15185), .B(n15184), .ZN(
        n15209) );
  INV_X1 U16767 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15188) );
  AOI22_X1 U16768 ( .A1(n15197), .A2(n15209), .B1(n15188), .B2(n15195), .ZN(
        P3_U3414) );
  NOR2_X1 U16769 ( .A1(n15190), .A2(n15189), .ZN(n15192) );
  AOI211_X1 U16770 ( .C1(n15194), .C2(n15193), .A(n15192), .B(n15191), .ZN(
        n15212) );
  INV_X1 U16771 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15196) );
  AOI22_X1 U16772 ( .A1(n15197), .A2(n15212), .B1(n15196), .B2(n15195), .ZN(
        P3_U3417) );
  AOI22_X1 U16773 ( .A1(n15213), .A2(n15198), .B1(n9507), .B2(n15210), .ZN(
        P3_U3460) );
  AOI22_X1 U16774 ( .A1(n15213), .A2(n15199), .B1(n9527), .B2(n15210), .ZN(
        P3_U3461) );
  AOI22_X1 U16775 ( .A1(n15213), .A2(n15200), .B1(n9709), .B2(n15210), .ZN(
        P3_U3462) );
  AOI22_X1 U16776 ( .A1(n15213), .A2(n15202), .B1(n15201), .B2(n15210), .ZN(
        P3_U3463) );
  INV_X1 U16777 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15203) );
  AOI22_X1 U16778 ( .A1(n15213), .A2(n15204), .B1(n15203), .B2(n15210), .ZN(
        P3_U3464) );
  AOI22_X1 U16779 ( .A1(n15213), .A2(n15206), .B1(n15205), .B2(n15210), .ZN(
        P3_U3465) );
  INV_X1 U16780 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15351) );
  AOI22_X1 U16781 ( .A1(n15213), .A2(n15207), .B1(n15351), .B2(n15210), .ZN(
        P3_U3466) );
  AOI22_X1 U16782 ( .A1(n15213), .A2(n15209), .B1(n15208), .B2(n15210), .ZN(
        P3_U3467) );
  AOI22_X1 U16783 ( .A1(n15213), .A2(n15212), .B1(n15211), .B2(n15210), .ZN(
        P3_U3468) );
  OAI22_X1 U16784 ( .A1(P3_REG0_REG_28__SCAN_IN), .A2(keyinput52), .B1(
        keyinput36), .B2(P2_REG1_REG_4__SCAN_IN), .ZN(n15214) );
  AOI221_X1 U16785 ( .B1(P3_REG0_REG_28__SCAN_IN), .B2(keyinput52), .C1(
        P2_REG1_REG_4__SCAN_IN), .C2(keyinput36), .A(n15214), .ZN(n15221) );
  OAI22_X1 U16786 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput34), .B1(
        keyinput111), .B2(P2_REG3_REG_14__SCAN_IN), .ZN(n15215) );
  AOI221_X1 U16787 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput34), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput111), .A(n15215), .ZN(n15220) );
  OAI22_X1 U16788 ( .A1(P3_REG0_REG_30__SCAN_IN), .A2(keyinput32), .B1(
        keyinput28), .B2(P1_D_REG_30__SCAN_IN), .ZN(n15216) );
  AOI221_X1 U16789 ( .B1(P3_REG0_REG_30__SCAN_IN), .B2(keyinput32), .C1(
        P1_D_REG_30__SCAN_IN), .C2(keyinput28), .A(n15216), .ZN(n15219) );
  OAI22_X1 U16790 ( .A1(P3_REG0_REG_3__SCAN_IN), .A2(keyinput11), .B1(
        P2_REG2_REG_26__SCAN_IN), .B2(keyinput22), .ZN(n15217) );
  AOI221_X1 U16791 ( .B1(P3_REG0_REG_3__SCAN_IN), .B2(keyinput11), .C1(
        keyinput22), .C2(P2_REG2_REG_26__SCAN_IN), .A(n15217), .ZN(n15218) );
  NAND4_X1 U16792 ( .A1(n15221), .A2(n15220), .A3(n15219), .A4(n15218), .ZN(
        n15249) );
  OAI22_X1 U16793 ( .A1(P3_REG2_REG_15__SCAN_IN), .A2(keyinput14), .B1(
        P1_REG1_REG_14__SCAN_IN), .B2(keyinput83), .ZN(n15222) );
  AOI221_X1 U16794 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(keyinput14), .C1(
        keyinput83), .C2(P1_REG1_REG_14__SCAN_IN), .A(n15222), .ZN(n15229) );
  OAI22_X1 U16795 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput91), .B1(
        P3_DATAO_REG_12__SCAN_IN), .B2(keyinput109), .ZN(n15223) );
  AOI221_X1 U16796 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput91), .C1(
        keyinput109), .C2(P3_DATAO_REG_12__SCAN_IN), .A(n15223), .ZN(n15228)
         );
  OAI22_X1 U16797 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput3), .B1(
        P3_ADDR_REG_1__SCAN_IN), .B2(keyinput125), .ZN(n15224) );
  AOI221_X1 U16798 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput3), .C1(keyinput125), .C2(P3_ADDR_REG_1__SCAN_IN), .A(n15224), .ZN(n15227) );
  OAI22_X1 U16799 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(keyinput63), .B1(
        P2_REG1_REG_17__SCAN_IN), .B2(keyinput2), .ZN(n15225) );
  AOI221_X1 U16800 ( .B1(P3_IR_REG_12__SCAN_IN), .B2(keyinput63), .C1(
        keyinput2), .C2(P2_REG1_REG_17__SCAN_IN), .A(n15225), .ZN(n15226) );
  NAND4_X1 U16801 ( .A1(n15229), .A2(n15228), .A3(n15227), .A4(n15226), .ZN(
        n15248) );
  OAI22_X1 U16802 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(keyinput48), .B1(
        keyinput29), .B2(SI_12_), .ZN(n15230) );
  AOI221_X1 U16803 ( .B1(P3_IR_REG_19__SCAN_IN), .B2(keyinput48), .C1(SI_12_), 
        .C2(keyinput29), .A(n15230), .ZN(n15237) );
  OAI22_X1 U16804 ( .A1(P3_D_REG_31__SCAN_IN), .A2(keyinput50), .B1(keyinput8), 
        .B2(P1_REG1_REG_29__SCAN_IN), .ZN(n15231) );
  AOI221_X1 U16805 ( .B1(P3_D_REG_31__SCAN_IN), .B2(keyinput50), .C1(
        P1_REG1_REG_29__SCAN_IN), .C2(keyinput8), .A(n15231), .ZN(n15236) );
  OAI22_X1 U16806 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput41), .B1(
        keyinput47), .B2(P1_IR_REG_7__SCAN_IN), .ZN(n15232) );
  AOI221_X1 U16807 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput41), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput47), .A(n15232), .ZN(n15235) );
  OAI22_X1 U16808 ( .A1(P2_D_REG_10__SCAN_IN), .A2(keyinput124), .B1(
        keyinput59), .B2(P1_D_REG_25__SCAN_IN), .ZN(n15233) );
  AOI221_X1 U16809 ( .B1(P2_D_REG_10__SCAN_IN), .B2(keyinput124), .C1(
        P1_D_REG_25__SCAN_IN), .C2(keyinput59), .A(n15233), .ZN(n15234) );
  NAND4_X1 U16810 ( .A1(n15237), .A2(n15236), .A3(n15235), .A4(n15234), .ZN(
        n15247) );
  OAI22_X1 U16811 ( .A1(P3_D_REG_2__SCAN_IN), .A2(keyinput35), .B1(keyinput110), .B2(P3_ADDR_REG_2__SCAN_IN), .ZN(n15238) );
  AOI221_X1 U16812 ( .B1(P3_D_REG_2__SCAN_IN), .B2(keyinput35), .C1(
        P3_ADDR_REG_2__SCAN_IN), .C2(keyinput110), .A(n15238), .ZN(n15245) );
  OAI22_X1 U16813 ( .A1(P2_REG0_REG_28__SCAN_IN), .A2(keyinput13), .B1(
        keyinput56), .B2(P2_REG1_REG_24__SCAN_IN), .ZN(n15239) );
  AOI221_X1 U16814 ( .B1(P2_REG0_REG_28__SCAN_IN), .B2(keyinput13), .C1(
        P2_REG1_REG_24__SCAN_IN), .C2(keyinput56), .A(n15239), .ZN(n15244) );
  OAI22_X1 U16815 ( .A1(SI_10_), .A2(keyinput96), .B1(keyinput9), .B2(
        P1_D_REG_2__SCAN_IN), .ZN(n15240) );
  AOI221_X1 U16816 ( .B1(SI_10_), .B2(keyinput96), .C1(P1_D_REG_2__SCAN_IN), 
        .C2(keyinput9), .A(n15240), .ZN(n15243) );
  OAI22_X1 U16817 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(keyinput90), .B1(
        keyinput6), .B2(P2_REG2_REG_22__SCAN_IN), .ZN(n15241) );
  AOI221_X1 U16818 ( .B1(P1_DATAO_REG_22__SCAN_IN), .B2(keyinput90), .C1(
        P2_REG2_REG_22__SCAN_IN), .C2(keyinput6), .A(n15241), .ZN(n15242) );
  NAND4_X1 U16819 ( .A1(n15245), .A2(n15244), .A3(n15243), .A4(n15242), .ZN(
        n15246) );
  NOR4_X1 U16820 ( .A1(n15249), .A2(n15248), .A3(n15247), .A4(n15246), .ZN(
        n15589) );
  AOI22_X1 U16821 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(keyinput149), .B1(
        P3_D_REG_14__SCAN_IN), .B2(keyinput194), .ZN(n15250) );
  OAI221_X1 U16822 ( .B1(P2_IR_REG_5__SCAN_IN), .B2(keyinput149), .C1(
        P3_D_REG_14__SCAN_IN), .C2(keyinput194), .A(n15250), .ZN(n15257) );
  AOI22_X1 U16823 ( .A1(SI_5_), .A2(keyinput240), .B1(SI_24_), .B2(keyinput200), .ZN(n15251) );
  OAI221_X1 U16824 ( .B1(SI_5_), .B2(keyinput240), .C1(SI_24_), .C2(
        keyinput200), .A(n15251), .ZN(n15256) );
  AOI22_X1 U16825 ( .A1(P2_D_REG_3__SCAN_IN), .A2(keyinput243), .B1(
        P3_IR_REG_15__SCAN_IN), .B2(keyinput220), .ZN(n15252) );
  OAI221_X1 U16826 ( .B1(P2_D_REG_3__SCAN_IN), .B2(keyinput243), .C1(
        P3_IR_REG_15__SCAN_IN), .C2(keyinput220), .A(n15252), .ZN(n15255) );
  AOI22_X1 U16827 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(keyinput254), .B1(
        P3_IR_REG_23__SCAN_IN), .B2(keyinput143), .ZN(n15253) );
  OAI221_X1 U16828 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(keyinput254), .C1(
        P3_IR_REG_23__SCAN_IN), .C2(keyinput143), .A(n15253), .ZN(n15254) );
  NOR4_X1 U16829 ( .A1(n15257), .A2(n15256), .A3(n15255), .A4(n15254), .ZN(
        n15285) );
  AOI22_X1 U16830 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(keyinput144), .B1(
        P1_IR_REG_28__SCAN_IN), .B2(keyinput147), .ZN(n15258) );
  OAI221_X1 U16831 ( .B1(P1_REG2_REG_21__SCAN_IN), .B2(keyinput144), .C1(
        P1_IR_REG_28__SCAN_IN), .C2(keyinput147), .A(n15258), .ZN(n15265) );
  AOI22_X1 U16832 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput239), .B1(
        P2_IR_REG_2__SCAN_IN), .B2(keyinput216), .ZN(n15259) );
  OAI221_X1 U16833 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput239), .C1(
        P2_IR_REG_2__SCAN_IN), .C2(keyinput216), .A(n15259), .ZN(n15264) );
  AOI22_X1 U16834 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(keyinput206), .B1(SI_18_), 
        .B2(keyinput248), .ZN(n15260) );
  OAI221_X1 U16835 ( .B1(P2_IR_REG_20__SCAN_IN), .B2(keyinput206), .C1(SI_18_), 
        .C2(keyinput248), .A(n15260), .ZN(n15263) );
  AOI22_X1 U16836 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(keyinput148), .B1(
        P3_IR_REG_19__SCAN_IN), .B2(keyinput176), .ZN(n15261) );
  OAI221_X1 U16837 ( .B1(P2_REG0_REG_14__SCAN_IN), .B2(keyinput148), .C1(
        P3_IR_REG_19__SCAN_IN), .C2(keyinput176), .A(n15261), .ZN(n15262) );
  NOR4_X1 U16838 ( .A1(n15265), .A2(n15264), .A3(n15263), .A4(n15262), .ZN(
        n15284) );
  AOI22_X1 U16839 ( .A1(P3_REG2_REG_30__SCAN_IN), .A2(keyinput166), .B1(
        P3_REG1_REG_3__SCAN_IN), .B2(keyinput204), .ZN(n15266) );
  OAI221_X1 U16840 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(keyinput166), .C1(
        P3_REG1_REG_3__SCAN_IN), .C2(keyinput204), .A(n15266), .ZN(n15273) );
  AOI22_X1 U16841 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(keyinput195), .B1(
        P3_REG0_REG_5__SCAN_IN), .B2(keyinput165), .ZN(n15267) );
  OAI221_X1 U16842 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(keyinput195), .C1(
        P3_REG0_REG_5__SCAN_IN), .C2(keyinput165), .A(n15267), .ZN(n15272) );
  AOI22_X1 U16843 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(keyinput211), .B1(
        P2_D_REG_10__SCAN_IN), .B2(keyinput252), .ZN(n15268) );
  OAI221_X1 U16844 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(keyinput211), .C1(
        P2_D_REG_10__SCAN_IN), .C2(keyinput252), .A(n15268), .ZN(n15271) );
  AOI22_X1 U16845 ( .A1(P3_REG0_REG_4__SCAN_IN), .A2(keyinput232), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(keyinput155), .ZN(n15269) );
  OAI221_X1 U16846 ( .B1(P3_REG0_REG_4__SCAN_IN), .B2(keyinput232), .C1(
        P1_DATAO_REG_25__SCAN_IN), .C2(keyinput155), .A(n15269), .ZN(n15270)
         );
  NOR4_X1 U16847 ( .A1(n15273), .A2(n15272), .A3(n15271), .A4(n15270), .ZN(
        n15283) );
  AOI22_X1 U16848 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput170), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(keyinput161), .ZN(n15274) );
  OAI221_X1 U16849 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput170), .C1(
        P1_DATAO_REG_3__SCAN_IN), .C2(keyinput161), .A(n15274), .ZN(n15281) );
  AOI22_X1 U16850 ( .A1(P3_DATAO_REG_12__SCAN_IN), .A2(keyinput237), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(keyinput132), .ZN(n15275) );
  OAI221_X1 U16851 ( .B1(P3_DATAO_REG_12__SCAN_IN), .B2(keyinput237), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput132), .A(n15275), .ZN(n15280) );
  AOI22_X1 U16852 ( .A1(P2_REG0_REG_20__SCAN_IN), .A2(keyinput159), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput128), .ZN(n15276) );
  OAI221_X1 U16853 ( .B1(P2_REG0_REG_20__SCAN_IN), .B2(keyinput159), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput128), .A(n15276), .ZN(n15279) );
  AOI22_X1 U16854 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(keyinput213), .B1(
        P3_D_REG_22__SCAN_IN), .B2(keyinput210), .ZN(n15277) );
  OAI221_X1 U16855 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(keyinput213), .C1(
        P3_D_REG_22__SCAN_IN), .C2(keyinput210), .A(n15277), .ZN(n15278) );
  NOR4_X1 U16856 ( .A1(n15281), .A2(n15280), .A3(n15279), .A4(n15278), .ZN(
        n15282) );
  NAND4_X1 U16857 ( .A1(n15285), .A2(n15284), .A3(n15283), .A4(n15282), .ZN(
        n15432) );
  AOI22_X1 U16858 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(keyinput133), .B1(
        P3_D_REG_5__SCAN_IN), .B2(keyinput158), .ZN(n15286) );
  OAI221_X1 U16859 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(keyinput133), .C1(
        P3_D_REG_5__SCAN_IN), .C2(keyinput158), .A(n15286), .ZN(n15293) );
  AOI22_X1 U16860 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(keyinput226), .B1(
        P3_REG0_REG_31__SCAN_IN), .B2(keyinput244), .ZN(n15287) );
  OAI221_X1 U16861 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(keyinput226), .C1(
        P3_REG0_REG_31__SCAN_IN), .C2(keyinput244), .A(n15287), .ZN(n15292) );
  AOI22_X1 U16862 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(keyinput183), .B1(
        P2_REG0_REG_28__SCAN_IN), .B2(keyinput141), .ZN(n15288) );
  OAI221_X1 U16863 ( .B1(P2_REG0_REG_1__SCAN_IN), .B2(keyinput183), .C1(
        P2_REG0_REG_28__SCAN_IN), .C2(keyinput141), .A(n15288), .ZN(n15291) );
  AOI22_X1 U16864 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput150), .B1(
        P2_IR_REG_1__SCAN_IN), .B2(keyinput173), .ZN(n15289) );
  OAI221_X1 U16865 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput150), .C1(
        P2_IR_REG_1__SCAN_IN), .C2(keyinput173), .A(n15289), .ZN(n15290) );
  NOR4_X1 U16866 ( .A1(n15293), .A2(n15292), .A3(n15291), .A4(n15290), .ZN(
        n15321) );
  AOI22_X1 U16867 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(keyinput222), .B1(
        P3_IR_REG_22__SCAN_IN), .B2(keyinput234), .ZN(n15294) );
  OAI221_X1 U16868 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(keyinput222), .C1(
        P3_IR_REG_22__SCAN_IN), .C2(keyinput234), .A(n15294), .ZN(n15301) );
  AOI22_X1 U16869 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput253), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(keyinput129), .ZN(n15295) );
  OAI221_X1 U16870 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput253), .C1(
        P3_REG3_REG_2__SCAN_IN), .C2(keyinput129), .A(n15295), .ZN(n15300) );
  AOI22_X1 U16871 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(keyinput172), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(keyinput186), .ZN(n15296) );
  OAI221_X1 U16872 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(keyinput172), .C1(
        P1_DATAO_REG_13__SCAN_IN), .C2(keyinput186), .A(n15296), .ZN(n15299)
         );
  AOI22_X1 U16873 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput179), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput219), .ZN(n15297) );
  OAI221_X1 U16874 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput179), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput219), .A(n15297), .ZN(n15298)
         );
  NOR4_X1 U16875 ( .A1(n15301), .A2(n15300), .A3(n15299), .A4(n15298), .ZN(
        n15320) );
  AOI22_X1 U16876 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(keyinput151), .B1(SI_12_), 
        .B2(keyinput157), .ZN(n15302) );
  OAI221_X1 U16877 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(keyinput151), .C1(SI_12_), .C2(keyinput157), .A(n15302), .ZN(n15309) );
  AOI22_X1 U16878 ( .A1(P2_REG2_REG_30__SCAN_IN), .A2(keyinput255), .B1(
        P3_IR_REG_5__SCAN_IN), .B2(keyinput247), .ZN(n15303) );
  OAI221_X1 U16879 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(keyinput255), .C1(
        P3_IR_REG_5__SCAN_IN), .C2(keyinput247), .A(n15303), .ZN(n15308) );
  AOI22_X1 U16880 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput137), .B1(
        P3_REG2_REG_17__SCAN_IN), .B2(keyinput185), .ZN(n15304) );
  OAI221_X1 U16881 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput137), .C1(
        P3_REG2_REG_17__SCAN_IN), .C2(keyinput185), .A(n15304), .ZN(n15307) );
  AOI22_X1 U16882 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput175), .B1(
        P3_REG2_REG_15__SCAN_IN), .B2(keyinput142), .ZN(n15305) );
  OAI221_X1 U16883 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput175), .C1(
        P3_REG2_REG_15__SCAN_IN), .C2(keyinput142), .A(n15305), .ZN(n15306) );
  NOR4_X1 U16884 ( .A1(n15309), .A2(n15308), .A3(n15307), .A4(n15306), .ZN(
        n15319) );
  AOI22_X1 U16885 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput169), .B1(SI_26_), 
        .B2(keyinput229), .ZN(n15310) );
  OAI221_X1 U16886 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput169), .C1(SI_26_), 
        .C2(keyinput229), .A(n15310), .ZN(n15317) );
  AOI22_X1 U16887 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(keyinput214), .B1(
        P2_IR_REG_9__SCAN_IN), .B2(keyinput182), .ZN(n15311) );
  OAI221_X1 U16888 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(keyinput214), .C1(
        P2_IR_REG_9__SCAN_IN), .C2(keyinput182), .A(n15311), .ZN(n15316) );
  AOI22_X1 U16889 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput131), .B1(
        P2_REG2_REG_13__SCAN_IN), .B2(keyinput246), .ZN(n15312) );
  OAI221_X1 U16890 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput131), .C1(
        P2_REG2_REG_13__SCAN_IN), .C2(keyinput246), .A(n15312), .ZN(n15315) );
  AOI22_X1 U16891 ( .A1(P1_D_REG_17__SCAN_IN), .A2(keyinput168), .B1(
        P2_IR_REG_21__SCAN_IN), .B2(keyinput192), .ZN(n15313) );
  OAI221_X1 U16892 ( .B1(P1_D_REG_17__SCAN_IN), .B2(keyinput168), .C1(
        P2_IR_REG_21__SCAN_IN), .C2(keyinput192), .A(n15313), .ZN(n15314) );
  NOR4_X1 U16893 ( .A1(n15317), .A2(n15316), .A3(n15315), .A4(n15314), .ZN(
        n15318) );
  NAND4_X1 U16894 ( .A1(n15321), .A2(n15320), .A3(n15319), .A4(n15318), .ZN(
        n15431) );
  AOI22_X1 U16895 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput231), .B1(
        P3_D_REG_29__SCAN_IN), .B2(keyinput193), .ZN(n15322) );
  OAI221_X1 U16896 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput231), .C1(
        P3_D_REG_29__SCAN_IN), .C2(keyinput193), .A(n15322), .ZN(n15331) );
  AOI22_X1 U16897 ( .A1(P2_D_REG_6__SCAN_IN), .A2(keyinput249), .B1(SI_28_), 
        .B2(keyinput235), .ZN(n15323) );
  OAI221_X1 U16898 ( .B1(P2_D_REG_6__SCAN_IN), .B2(keyinput249), .C1(SI_28_), 
        .C2(keyinput235), .A(n15323), .ZN(n15330) );
  AOI22_X1 U16899 ( .A1(P1_D_REG_8__SCAN_IN), .A2(keyinput217), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput207), .ZN(n15324) );
  OAI221_X1 U16900 ( .B1(P1_D_REG_8__SCAN_IN), .B2(keyinput217), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput207), .A(n15324), .ZN(n15329) );
  AOI22_X1 U16901 ( .A1(n15327), .A2(keyinput164), .B1(keyinput156), .B2(
        n15326), .ZN(n15325) );
  OAI221_X1 U16902 ( .B1(n15327), .B2(keyinput164), .C1(n15326), .C2(
        keyinput156), .A(n15325), .ZN(n15328) );
  NOR4_X1 U16903 ( .A1(n15331), .A2(n15330), .A3(n15329), .A4(n15328), .ZN(
        n15373) );
  AOI22_X1 U16904 ( .A1(n15333), .A2(keyinput160), .B1(keyinput188), .B2(
        n15445), .ZN(n15332) );
  OAI221_X1 U16905 ( .B1(n15333), .B2(keyinput160), .C1(n15445), .C2(
        keyinput188), .A(n15332), .ZN(n15343) );
  INV_X1 U16906 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n15335) );
  AOI22_X1 U16907 ( .A1(n15335), .A2(keyinput212), .B1(n15502), .B2(
        keyinput152), .ZN(n15334) );
  OAI221_X1 U16908 ( .B1(n15335), .B2(keyinput212), .C1(n15502), .C2(
        keyinput152), .A(n15334), .ZN(n15342) );
  XNOR2_X1 U16909 ( .A(P3_REG1_REG_31__SCAN_IN), .B(keyinput251), .ZN(n15338)
         );
  XNOR2_X1 U16910 ( .A(P3_IR_REG_30__SCAN_IN), .B(keyinput202), .ZN(n15337) );
  XNOR2_X1 U16911 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput191), .ZN(n15336) );
  NAND3_X1 U16912 ( .A1(n15338), .A2(n15337), .A3(n15336), .ZN(n15341) );
  XNOR2_X1 U16913 ( .A(n15339), .B(keyinput181), .ZN(n15340) );
  NOR4_X1 U16914 ( .A1(n15343), .A2(n15342), .A3(n15341), .A4(n15340), .ZN(
        n15372) );
  INV_X1 U16915 ( .A(SI_0_), .ZN(n15508) );
  AOI22_X1 U16916 ( .A1(n15345), .A2(keyinput241), .B1(n15508), .B2(
        keyinput145), .ZN(n15344) );
  OAI221_X1 U16917 ( .B1(n15345), .B2(keyinput241), .C1(n15508), .C2(
        keyinput145), .A(n15344), .ZN(n15357) );
  INV_X1 U16918 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n15453) );
  AOI22_X1 U16919 ( .A1(n15347), .A2(keyinput250), .B1(n15453), .B2(
        keyinput221), .ZN(n15346) );
  OAI221_X1 U16920 ( .B1(n15347), .B2(keyinput250), .C1(n15453), .C2(
        keyinput221), .A(n15346), .ZN(n15356) );
  AOI22_X1 U16921 ( .A1(n15350), .A2(keyinput225), .B1(n15349), .B2(
        keyinput153), .ZN(n15348) );
  OAI221_X1 U16922 ( .B1(n15350), .B2(keyinput225), .C1(n15349), .C2(
        keyinput153), .A(n15348), .ZN(n15355) );
  XOR2_X1 U16923 ( .A(n15351), .B(keyinput227), .Z(n15353) );
  XNOR2_X1 U16924 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput208), .ZN(n15352)
         );
  NAND2_X1 U16925 ( .A1(n15353), .A2(n15352), .ZN(n15354) );
  NOR4_X1 U16926 ( .A1(n15357), .A2(n15356), .A3(n15355), .A4(n15354), .ZN(
        n15371) );
  AOI22_X1 U16927 ( .A1(n8459), .A2(keyinput230), .B1(n15359), .B2(keyinput184), .ZN(n15358) );
  OAI221_X1 U16928 ( .B1(n8459), .B2(keyinput230), .C1(n15359), .C2(
        keyinput184), .A(n15358), .ZN(n15369) );
  AOI22_X1 U16929 ( .A1(n15498), .A2(keyinput242), .B1(keyinput197), .B2(
        P2_U3088), .ZN(n15360) );
  OAI221_X1 U16930 ( .B1(n15498), .B2(keyinput242), .C1(P2_U3088), .C2(
        keyinput197), .A(n15360), .ZN(n15368) );
  AOI22_X1 U16931 ( .A1(n15363), .A2(keyinput187), .B1(n15362), .B2(
        keyinput162), .ZN(n15361) );
  OAI221_X1 U16932 ( .B1(n15363), .B2(keyinput187), .C1(n15362), .C2(
        keyinput162), .A(n15361), .ZN(n15367) );
  XNOR2_X1 U16933 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput174), .ZN(n15365)
         );
  XNOR2_X1 U16934 ( .A(P1_REG1_REG_29__SCAN_IN), .B(keyinput136), .ZN(n15364)
         );
  NAND2_X1 U16935 ( .A1(n15365), .A2(n15364), .ZN(n15366) );
  NOR4_X1 U16936 ( .A1(n15369), .A2(n15368), .A3(n15367), .A4(n15366), .ZN(
        n15370) );
  NAND4_X1 U16937 ( .A1(n15373), .A2(n15372), .A3(n15371), .A4(n15370), .ZN(
        n15430) );
  AOI22_X1 U16938 ( .A1(n15473), .A2(keyinput196), .B1(n15375), .B2(
        keyinput180), .ZN(n15374) );
  OAI221_X1 U16939 ( .B1(n15473), .B2(keyinput196), .C1(n15375), .C2(
        keyinput180), .A(n15374), .ZN(n15387) );
  AOI22_X1 U16940 ( .A1(n15378), .A2(keyinput224), .B1(keyinput233), .B2(
        n15377), .ZN(n15376) );
  OAI221_X1 U16941 ( .B1(n15378), .B2(keyinput224), .C1(n15377), .C2(
        keyinput233), .A(n15376), .ZN(n15386) );
  AOI22_X1 U16942 ( .A1(n8510), .A2(keyinput140), .B1(n15380), .B2(keyinput177), .ZN(n15379) );
  OAI221_X1 U16943 ( .B1(n8510), .B2(keyinput140), .C1(n15380), .C2(
        keyinput177), .A(n15379), .ZN(n15385) );
  AOI22_X1 U16944 ( .A1(n15383), .A2(keyinput203), .B1(n15382), .B2(
        keyinput178), .ZN(n15381) );
  OAI221_X1 U16945 ( .B1(n15383), .B2(keyinput203), .C1(n15382), .C2(
        keyinput178), .A(n15381), .ZN(n15384) );
  NOR4_X1 U16946 ( .A1(n15387), .A2(n15386), .A3(n15385), .A4(n15384), .ZN(
        n15428) );
  INV_X1 U16947 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U16948 ( .A1(n15389), .A2(keyinput198), .B1(keyinput190), .B2(
        n10759), .ZN(n15388) );
  OAI221_X1 U16949 ( .B1(n15389), .B2(keyinput198), .C1(n10759), .C2(
        keyinput190), .A(n15388), .ZN(n15399) );
  INV_X1 U16950 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n15537) );
  AOI22_X1 U16951 ( .A1(n15391), .A2(keyinput238), .B1(n15537), .B2(
        keyinput245), .ZN(n15390) );
  OAI221_X1 U16952 ( .B1(n15391), .B2(keyinput238), .C1(n15537), .C2(
        keyinput245), .A(n15390), .ZN(n15398) );
  AOI22_X1 U16953 ( .A1(n15521), .A2(keyinput223), .B1(n15393), .B2(
        keyinput163), .ZN(n15392) );
  OAI221_X1 U16954 ( .B1(n15521), .B2(keyinput223), .C1(n15393), .C2(
        keyinput163), .A(n15392), .ZN(n15397) );
  AOI22_X1 U16955 ( .A1(n15496), .A2(keyinput171), .B1(n15395), .B2(
        keyinput218), .ZN(n15394) );
  OAI221_X1 U16956 ( .B1(n15496), .B2(keyinput171), .C1(n15395), .C2(
        keyinput218), .A(n15394), .ZN(n15396) );
  NOR4_X1 U16957 ( .A1(n15399), .A2(n15398), .A3(n15397), .A4(n15396), .ZN(
        n15427) );
  AOI22_X1 U16958 ( .A1(n15459), .A2(keyinput138), .B1(keyinput205), .B2(
        n11498), .ZN(n15400) );
  OAI221_X1 U16959 ( .B1(n15459), .B2(keyinput138), .C1(n11498), .C2(
        keyinput205), .A(n15400), .ZN(n15409) );
  AOI22_X1 U16960 ( .A1(n15452), .A2(keyinput189), .B1(n15499), .B2(
        keyinput209), .ZN(n15401) );
  OAI221_X1 U16961 ( .B1(n15452), .B2(keyinput189), .C1(n15499), .C2(
        keyinput209), .A(n15401), .ZN(n15408) );
  AOI22_X1 U16962 ( .A1(n10146), .A2(keyinput236), .B1(n15531), .B2(
        keyinput154), .ZN(n15402) );
  OAI221_X1 U16963 ( .B1(n10146), .B2(keyinput236), .C1(n15531), .C2(
        keyinput154), .A(n15402), .ZN(n15407) );
  XOR2_X1 U16964 ( .A(n15403), .B(keyinput139), .Z(n15405) );
  XNOR2_X1 U16965 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput167), .ZN(n15404) );
  NAND2_X1 U16966 ( .A1(n15405), .A2(n15404), .ZN(n15406) );
  NOR4_X1 U16967 ( .A1(n15409), .A2(n15408), .A3(n15407), .A4(n15406), .ZN(
        n15426) );
  AOI22_X1 U16968 ( .A1(n11548), .A2(keyinput134), .B1(keyinput130), .B2(
        n15411), .ZN(n15410) );
  OAI221_X1 U16969 ( .B1(n11548), .B2(keyinput134), .C1(n15411), .C2(
        keyinput130), .A(n15410), .ZN(n15412) );
  INV_X1 U16970 ( .A(n15412), .ZN(n15424) );
  XNOR2_X1 U16971 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput146), .ZN(n15415) );
  XNOR2_X1 U16972 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput135), .ZN(n15414)
         );
  XNOR2_X1 U16973 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput228), .ZN(n15413) );
  AND3_X1 U16974 ( .A1(n15415), .A2(n15414), .A3(n15413), .ZN(n15423) );
  AOI22_X1 U16975 ( .A1(n15418), .A2(keyinput215), .B1(n15417), .B2(
        keyinput201), .ZN(n15416) );
  OAI221_X1 U16976 ( .B1(n15418), .B2(keyinput215), .C1(n15417), .C2(
        keyinput201), .A(n15416), .ZN(n15419) );
  INV_X1 U16977 ( .A(n15419), .ZN(n15422) );
  INV_X1 U16978 ( .A(keyinput199), .ZN(n15420) );
  XNOR2_X1 U16979 ( .A(n15450), .B(n15420), .ZN(n15421) );
  AND4_X1 U16980 ( .A1(n15424), .A2(n15423), .A3(n15422), .A4(n15421), .ZN(
        n15425) );
  NAND4_X1 U16981 ( .A1(n15428), .A2(n15427), .A3(n15426), .A4(n15425), .ZN(
        n15429) );
  NOR4_X1 U16982 ( .A1(n15432), .A2(n15431), .A3(n15430), .A4(n15429), .ZN(
        n15550) );
  AOI22_X1 U16983 ( .A1(P3_REG0_REG_17__SCAN_IN), .A2(keyinput70), .B1(n15434), 
        .B2(keyinput44), .ZN(n15433) );
  OAI221_X1 U16984 ( .B1(P3_REG0_REG_17__SCAN_IN), .B2(keyinput70), .C1(n15434), .C2(keyinput44), .A(n15433), .ZN(n15442) );
  AOI22_X1 U16985 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(keyinput78), .B1(
        P3_REG0_REG_5__SCAN_IN), .B2(keyinput37), .ZN(n15435) );
  OAI221_X1 U16986 ( .B1(P2_IR_REG_20__SCAN_IN), .B2(keyinput78), .C1(
        P3_REG0_REG_5__SCAN_IN), .C2(keyinput37), .A(n15435), .ZN(n15441) );
  AOI22_X1 U16987 ( .A1(P1_D_REG_17__SCAN_IN), .A2(keyinput40), .B1(
        P3_IR_REG_15__SCAN_IN), .B2(keyinput92), .ZN(n15436) );
  OAI221_X1 U16988 ( .B1(P1_D_REG_17__SCAN_IN), .B2(keyinput40), .C1(
        P3_IR_REG_15__SCAN_IN), .C2(keyinput92), .A(n15436), .ZN(n15440) );
  XNOR2_X1 U16989 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput80), .ZN(n15438) );
  XNOR2_X1 U16990 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(keyinput27), .ZN(n15437)
         );
  NAND2_X1 U16991 ( .A1(n15438), .A2(n15437), .ZN(n15439) );
  NOR4_X1 U16992 ( .A1(n15442), .A2(n15441), .A3(n15440), .A4(n15439), .ZN(
        n15490) );
  AOI22_X1 U16993 ( .A1(n15445), .A2(keyinput60), .B1(n15444), .B2(keyinput101), .ZN(n15443) );
  OAI221_X1 U16994 ( .B1(n15445), .B2(keyinput60), .C1(n15444), .C2(
        keyinput101), .A(n15443), .ZN(n15457) );
  INV_X1 U16995 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15447) );
  AOI22_X1 U16996 ( .A1(n15447), .A2(keyinput0), .B1(keyinput5), .B2(n10176), 
        .ZN(n15446) );
  OAI221_X1 U16997 ( .B1(n15447), .B2(keyinput0), .C1(n10176), .C2(keyinput5), 
        .A(n15446), .ZN(n15456) );
  AOI22_X1 U16998 ( .A1(n15450), .A2(keyinput71), .B1(n15449), .B2(keyinput116), .ZN(n15448) );
  OAI221_X1 U16999 ( .B1(n15450), .B2(keyinput71), .C1(n15449), .C2(
        keyinput116), .A(n15448), .ZN(n15455) );
  AOI22_X1 U17000 ( .A1(n15453), .A2(keyinput93), .B1(keyinput61), .B2(n15452), 
        .ZN(n15451) );
  OAI221_X1 U17001 ( .B1(n15453), .B2(keyinput93), .C1(n15452), .C2(keyinput61), .A(n15451), .ZN(n15454) );
  NOR4_X1 U17002 ( .A1(n15457), .A2(n15456), .A3(n15455), .A4(n15454), .ZN(
        n15489) );
  INV_X1 U17003 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n15460) );
  AOI22_X1 U17004 ( .A1(n15460), .A2(keyinput123), .B1(keyinput10), .B2(n15459), .ZN(n15458) );
  OAI221_X1 U17005 ( .B1(n15460), .B2(keyinput123), .C1(n15459), .C2(
        keyinput10), .A(n15458), .ZN(n15470) );
  AOI22_X1 U17006 ( .A1(n15463), .A2(keyinput89), .B1(keyinput126), .B2(n15462), .ZN(n15461) );
  OAI221_X1 U17007 ( .B1(n15463), .B2(keyinput89), .C1(n15462), .C2(
        keyinput126), .A(n15461), .ZN(n15469) );
  XOR2_X1 U17008 ( .A(n14139), .B(keyinput16), .Z(n15467) );
  XNOR2_X1 U17009 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput94), .ZN(n15466) );
  XNOR2_X1 U17010 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput79), .ZN(n15465) );
  XNOR2_X1 U17011 ( .A(P3_IR_REG_23__SCAN_IN), .B(keyinput15), .ZN(n15464) );
  NAND4_X1 U17012 ( .A1(n15467), .A2(n15466), .A3(n15465), .A4(n15464), .ZN(
        n15468) );
  NOR3_X1 U17013 ( .A1(n15470), .A2(n15469), .A3(n15468), .ZN(n15488) );
  XNOR2_X1 U17014 ( .A(n15471), .B(keyinput100), .ZN(n15476) );
  XNOR2_X1 U17015 ( .A(n15472), .B(keyinput21), .ZN(n15475) );
  XNOR2_X1 U17016 ( .A(n15473), .B(keyinput68), .ZN(n15474) );
  NOR3_X1 U17017 ( .A1(n15476), .A2(n15475), .A3(n15474), .ZN(n15479) );
  XNOR2_X1 U17018 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput7), .ZN(n15478) );
  XNOR2_X1 U17019 ( .A(SI_17_), .B(keyinput75), .ZN(n15477) );
  NAND3_X1 U17020 ( .A1(n15479), .A2(n15478), .A3(n15477), .ZN(n15486) );
  AOI22_X1 U17021 ( .A1(n15482), .A2(keyinput65), .B1(keyinput57), .B2(n15481), 
        .ZN(n15480) );
  OAI221_X1 U17022 ( .B1(n15482), .B2(keyinput65), .C1(n15481), .C2(keyinput57), .A(n15480), .ZN(n15485) );
  XNOR2_X1 U17023 ( .A(n15483), .B(keyinput66), .ZN(n15484) );
  NOR3_X1 U17024 ( .A1(n15486), .A2(n15485), .A3(n15484), .ZN(n15487) );
  NAND4_X1 U17025 ( .A1(n15490), .A2(n15489), .A3(n15488), .A4(n15487), .ZN(
        n15549) );
  AOI22_X1 U17026 ( .A1(n15493), .A2(keyinput120), .B1(keyinput38), .B2(n15492), .ZN(n15491) );
  OAI221_X1 U17027 ( .B1(n15493), .B2(keyinput120), .C1(n15492), .C2(
        keyinput38), .A(n15491), .ZN(n15506) );
  AOI22_X1 U17028 ( .A1(n15496), .A2(keyinput43), .B1(n15495), .B2(keyinput82), 
        .ZN(n15494) );
  OAI221_X1 U17029 ( .B1(n15496), .B2(keyinput43), .C1(n15495), .C2(keyinput82), .A(n15494), .ZN(n15505) );
  AOI22_X1 U17030 ( .A1(n15499), .A2(keyinput81), .B1(n15498), .B2(keyinput114), .ZN(n15497) );
  OAI221_X1 U17031 ( .B1(n15499), .B2(keyinput81), .C1(n15498), .C2(
        keyinput114), .A(n15497), .ZN(n15504) );
  AOI22_X1 U17032 ( .A1(n15502), .A2(keyinput24), .B1(keyinput115), .B2(n15501), .ZN(n15500) );
  OAI221_X1 U17033 ( .B1(n15502), .B2(keyinput24), .C1(n15501), .C2(
        keyinput115), .A(n15500), .ZN(n15503) );
  NOR4_X1 U17034 ( .A1(n15506), .A2(n15505), .A3(n15504), .A4(n15503), .ZN(
        n15547) );
  AOI22_X1 U17035 ( .A1(n13318), .A2(keyinput98), .B1(keyinput108), .B2(n10146), .ZN(n15507) );
  OAI221_X1 U17036 ( .B1(n13318), .B2(keyinput98), .C1(n10146), .C2(
        keyinput108), .A(n15507), .ZN(n15516) );
  XNOR2_X1 U17037 ( .A(keyinput17), .B(n15508), .ZN(n15515) );
  XNOR2_X1 U17038 ( .A(keyinput86), .B(n8649), .ZN(n15514) );
  XNOR2_X1 U17039 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput64), .ZN(n15512) );
  XNOR2_X1 U17040 ( .A(P1_REG1_REG_18__SCAN_IN), .B(keyinput113), .ZN(n15511)
         );
  XNOR2_X1 U17041 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput119), .ZN(n15510) );
  XNOR2_X1 U17042 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput19), .ZN(n15509) );
  NAND4_X1 U17043 ( .A1(n15512), .A2(n15511), .A3(n15510), .A4(n15509), .ZN(
        n15513) );
  NOR4_X1 U17044 ( .A1(n15516), .A2(n15515), .A3(n15514), .A4(n15513), .ZN(
        n15546) );
  AOI22_X1 U17045 ( .A1(n15519), .A2(keyinput85), .B1(keyinput67), .B2(n15518), 
        .ZN(n15517) );
  OAI221_X1 U17046 ( .B1(n15519), .B2(keyinput85), .C1(n15518), .C2(keyinput67), .A(n15517), .ZN(n15529) );
  AOI22_X1 U17047 ( .A1(n15522), .A2(keyinput31), .B1(n15521), .B2(keyinput95), 
        .ZN(n15520) );
  OAI221_X1 U17048 ( .B1(n15522), .B2(keyinput31), .C1(n15521), .C2(keyinput95), .A(n15520), .ZN(n15528) );
  XNOR2_X1 U17049 ( .A(SI_5_), .B(keyinput112), .ZN(n15526) );
  XNOR2_X1 U17050 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput25), .ZN(n15525)
         );
  XNOR2_X1 U17051 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput88), .ZN(n15524) );
  XNOR2_X1 U17052 ( .A(keyinput23), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n15523) );
  NAND4_X1 U17053 ( .A1(n15526), .A2(n15525), .A3(n15524), .A4(n15523), .ZN(
        n15527) );
  NOR3_X1 U17054 ( .A1(n15529), .A2(n15528), .A3(n15527), .ZN(n15545) );
  AOI22_X1 U17055 ( .A1(n15532), .A2(keyinput51), .B1(n15531), .B2(keyinput26), 
        .ZN(n15530) );
  OAI221_X1 U17056 ( .B1(n15532), .B2(keyinput51), .C1(n15531), .C2(keyinput26), .A(n15530), .ZN(n15543) );
  AOI22_X1 U17057 ( .A1(n15535), .A2(keyinput20), .B1(n15534), .B2(keyinput121), .ZN(n15533) );
  OAI221_X1 U17058 ( .B1(n15535), .B2(keyinput20), .C1(n15534), .C2(
        keyinput121), .A(n15533), .ZN(n15542) );
  AOI22_X1 U17059 ( .A1(n8459), .A2(keyinput102), .B1(n15537), .B2(keyinput117), .ZN(n15536) );
  OAI221_X1 U17060 ( .B1(n8459), .B2(keyinput102), .C1(n15537), .C2(
        keyinput117), .A(n15536), .ZN(n15541) );
  XNOR2_X1 U17061 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput33), .ZN(n15539)
         );
  XNOR2_X1 U17062 ( .A(SI_28_), .B(keyinput107), .ZN(n15538) );
  NAND2_X1 U17063 ( .A1(n15539), .A2(n15538), .ZN(n15540) );
  NOR4_X1 U17064 ( .A1(n15543), .A2(n15542), .A3(n15541), .A4(n15540), .ZN(
        n15544) );
  NAND4_X1 U17065 ( .A1(n15547), .A2(n15546), .A3(n15545), .A4(n15544), .ZN(
        n15548) );
  NOR3_X1 U17066 ( .A1(n15550), .A2(n15549), .A3(n15548), .ZN(n15588) );
  OAI22_X1 U17067 ( .A1(P3_D_REG_5__SCAN_IN), .A2(keyinput30), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput39), .ZN(n15551) );
  AOI221_X1 U17068 ( .B1(P3_D_REG_5__SCAN_IN), .B2(keyinput30), .C1(keyinput39), .C2(P1_IR_REG_8__SCAN_IN), .A(n15551), .ZN(n15558) );
  OAI22_X1 U17069 ( .A1(P3_IR_REG_30__SCAN_IN), .A2(keyinput74), .B1(
        keyinput76), .B2(P3_REG1_REG_3__SCAN_IN), .ZN(n15552) );
  AOI221_X1 U17070 ( .B1(P3_IR_REG_30__SCAN_IN), .B2(keyinput74), .C1(
        P3_REG1_REG_3__SCAN_IN), .C2(keyinput76), .A(n15552), .ZN(n15557) );
  OAI22_X1 U17071 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput1), .B1(
        keyinput105), .B2(P2_D_REG_13__SCAN_IN), .ZN(n15553) );
  AOI221_X1 U17072 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput1), .C1(
        P2_D_REG_13__SCAN_IN), .C2(keyinput105), .A(n15553), .ZN(n15556) );
  OAI22_X1 U17073 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(keyinput45), .B1(
        keyinput122), .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n15554) );
  AOI221_X1 U17074 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(keyinput45), .C1(
        P3_DATAO_REG_15__SCAN_IN), .C2(keyinput122), .A(n15554), .ZN(n15555)
         );
  NAND4_X1 U17075 ( .A1(n15558), .A2(n15557), .A3(n15556), .A4(n15555), .ZN(
        n15586) );
  OAI22_X1 U17076 ( .A1(P3_REG1_REG_25__SCAN_IN), .A2(keyinput73), .B1(
        keyinput54), .B2(P2_IR_REG_9__SCAN_IN), .ZN(n15559) );
  AOI221_X1 U17077 ( .B1(P3_REG1_REG_25__SCAN_IN), .B2(keyinput73), .C1(
        P2_IR_REG_9__SCAN_IN), .C2(keyinput54), .A(n15559), .ZN(n15566) );
  OAI22_X1 U17078 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(keyinput87), .B1(
        keyinput12), .B2(P1_REG1_REG_11__SCAN_IN), .ZN(n15560) );
  AOI221_X1 U17079 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(keyinput87), .C1(
        P1_REG1_REG_11__SCAN_IN), .C2(keyinput12), .A(n15560), .ZN(n15565) );
  OAI22_X1 U17080 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(keyinput46), .B1(SI_14_), 
        .B2(keyinput49), .ZN(n15561) );
  AOI221_X1 U17081 ( .B1(P1_DATAO_REG_4__SCAN_IN), .B2(keyinput46), .C1(
        keyinput49), .C2(SI_14_), .A(n15561), .ZN(n15564) );
  OAI22_X1 U17082 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput103), .B1(
        P2_REG0_REG_1__SCAN_IN), .B2(keyinput55), .ZN(n15562) );
  AOI221_X1 U17083 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput103), .C1(
        keyinput55), .C2(P2_REG0_REG_1__SCAN_IN), .A(n15562), .ZN(n15563) );
  NAND4_X1 U17084 ( .A1(n15566), .A2(n15565), .A3(n15564), .A4(n15563), .ZN(
        n15585) );
  OAI22_X1 U17085 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(keyinput97), .B1(
        keyinput127), .B2(P2_REG2_REG_30__SCAN_IN), .ZN(n15567) );
  AOI221_X1 U17086 ( .B1(P2_REG0_REG_26__SCAN_IN), .B2(keyinput97), .C1(
        P2_REG2_REG_30__SCAN_IN), .C2(keyinput127), .A(n15567), .ZN(n15574) );
  OAI22_X1 U17087 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput4), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput69), .ZN(n15568) );
  AOI221_X1 U17088 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput4), .C1(
        keyinput69), .C2(P2_STATE_REG_SCAN_IN), .A(n15568), .ZN(n15573) );
  OAI22_X1 U17089 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(keyinput58), .B1(
        keyinput62), .B2(P2_REG0_REG_13__SCAN_IN), .ZN(n15569) );
  AOI221_X1 U17090 ( .B1(P1_DATAO_REG_13__SCAN_IN), .B2(keyinput58), .C1(
        P2_REG0_REG_13__SCAN_IN), .C2(keyinput62), .A(n15569), .ZN(n15572) );
  OAI22_X1 U17091 ( .A1(P3_REG0_REG_4__SCAN_IN), .A2(keyinput104), .B1(
        keyinput42), .B2(P2_REG3_REG_13__SCAN_IN), .ZN(n15570) );
  AOI221_X1 U17092 ( .B1(P3_REG0_REG_4__SCAN_IN), .B2(keyinput104), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput42), .A(n15570), .ZN(n15571) );
  NAND4_X1 U17093 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        n15584) );
  OAI22_X1 U17094 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(keyinput106), .B1(
        keyinput18), .B2(P1_IR_REG_16__SCAN_IN), .ZN(n15575) );
  AOI221_X1 U17095 ( .B1(P3_IR_REG_22__SCAN_IN), .B2(keyinput106), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput18), .A(n15575), .ZN(n15582) );
  OAI22_X1 U17096 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(keyinput99), .B1(
        keyinput118), .B2(P2_REG2_REG_13__SCAN_IN), .ZN(n15576) );
  AOI221_X1 U17097 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(keyinput99), .C1(
        P2_REG2_REG_13__SCAN_IN), .C2(keyinput118), .A(n15576), .ZN(n15581) );
  OAI22_X1 U17098 ( .A1(P3_D_REG_7__SCAN_IN), .A2(keyinput53), .B1(
        P2_REG2_REG_19__SCAN_IN), .B2(keyinput77), .ZN(n15577) );
  AOI221_X1 U17099 ( .B1(P3_D_REG_7__SCAN_IN), .B2(keyinput53), .C1(keyinput77), .C2(P2_REG2_REG_19__SCAN_IN), .A(n15577), .ZN(n15580) );
  OAI22_X1 U17100 ( .A1(SI_24_), .A2(keyinput72), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(keyinput84), .ZN(n15578) );
  AOI221_X1 U17101 ( .B1(SI_24_), .B2(keyinput72), .C1(keyinput84), .C2(
        P2_REG2_REG_15__SCAN_IN), .A(n15578), .ZN(n15579) );
  NAND4_X1 U17102 ( .A1(n15582), .A2(n15581), .A3(n15580), .A4(n15579), .ZN(
        n15583) );
  NOR4_X1 U17103 ( .A1(n15586), .A2(n15585), .A3(n15584), .A4(n15583), .ZN(
        n15587) );
  NAND3_X1 U17104 ( .A1(n15589), .A2(n15588), .A3(n15587), .ZN(n15604) );
  AOI21_X1 U17105 ( .B1(n15591), .B2(n13441), .A(n15590), .ZN(n15602) );
  INV_X1 U17106 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n15593) );
  OAI22_X1 U17107 ( .A1(n15599), .A2(n15594), .B1(n15593), .B2(n15592), .ZN(
        n15598) );
  NOR2_X1 U17108 ( .A1(n15596), .A2(n15595), .ZN(n15597) );
  AOI211_X1 U17109 ( .C1(n15599), .C2(P2_REG2_REG_0__SCAN_IN), .A(n15598), .B(
        n15597), .ZN(n15600) );
  OAI21_X1 U17110 ( .B1(n15602), .B2(n15601), .A(n15600), .ZN(n15603) );
  XNOR2_X1 U17111 ( .A(n15604), .B(n15603), .ZN(P2_U3265) );
  XOR2_X1 U17112 ( .A(n15606), .B(n15605), .Z(SUB_1596_U59) );
  XNOR2_X1 U17113 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15607), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17114 ( .B1(n15609), .B2(n15608), .A(n15617), .ZN(SUB_1596_U53) );
  XOR2_X1 U17115 ( .A(n15611), .B(n15610), .Z(SUB_1596_U56) );
  AOI21_X1 U17116 ( .B1(n15614), .B2(n15613), .A(n15612), .ZN(n15615) );
  XOR2_X1 U17117 ( .A(n15615), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  XOR2_X1 U17118 ( .A(n15617), .B(n15616), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7508 ( .A(n13810), .Z(n6827) );
  CLKBUF_X1 U8443 ( .A(n9596), .Z(n13246) );
  CLKBUF_X1 U8823 ( .A(n11689), .Z(n11605) );
endmodule

