

module b22_C_AntiSAT_k_256_8 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6646, n6650, n6651, n6652, n6654, n6656, n6657, n6658, n6659, n6660,
         n6661, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6675, n6676, n6677, n6678, n6679, n6680, n6682, n6683,
         n6684, n6685, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15607;

  INV_X1 U7393 ( .A(n6665), .ZN(n13579) );
  OAI211_X1 U7395 ( .C1(n8463), .C2(n7518), .A(n6654), .B(n11835), .ZN(n7517)
         );
  AOI21_X1 U7396 ( .B1(n6999), .B2(n12806), .A(n6997), .ZN(n12813) );
  NOR2_X1 U7397 ( .A1(n6652), .A2(n6651), .ZN(n6650) );
  AOI222_X1 U7398 ( .A1(n14759), .A2(n14758), .B1(n14757), .B2(
        P1_STATE_REG_SCAN_IN), .C1(P2_DATAO_REG_20__SCAN_IN), .C2(n14756), 
        .ZN(n14760) );
  NOR2_X1 U7399 ( .A1(n15570), .A2(n13234), .ZN(n6651) );
  NOR2_X1 U7400 ( .A1(n13236), .A2(n13285), .ZN(n6652) );
  OAI21_X1 U7402 ( .B1(n9977), .B2(n15490), .A(n9976), .ZN(n12969) );
  AOI21_X1 U7403 ( .B1(n13741), .B2(n15297), .A(n13578), .ZN(n6666) );
  NAND2_X1 U7404 ( .A1(n12387), .A2(n12386), .ZN(n13886) );
  OAI21_X1 U7405 ( .B1(n12801), .B2(n12800), .A(n12799), .ZN(n12802) );
  NAND2_X1 U7406 ( .A1(n12379), .A2(n12378), .ZN(n13915) );
  XNOR2_X1 U7407 ( .A(n13521), .B(n13431), .ZN(n9294) );
  AND2_X1 U7408 ( .A1(n8451), .A2(n8440), .ZN(n8441) );
  NAND2_X1 U7409 ( .A1(n15018), .A2(n15016), .ZN(n15021) );
  NAND2_X1 U7410 ( .A1(n12451), .A2(n12450), .ZN(n12456) );
  INV_X1 U7411 ( .A(n12791), .ZN(n12795) );
  NAND2_X1 U7412 ( .A1(n6660), .A2(n6659), .ZN(n12791) );
  NAND2_X1 U7413 ( .A1(n12785), .A2(n12784), .ZN(n6660) );
  NAND2_X1 U7414 ( .A1(n13924), .A2(n13923), .ZN(n13922) );
  AND2_X1 U7415 ( .A1(n7376), .A2(n7380), .ZN(n15013) );
  NAND2_X1 U7416 ( .A1(n8397), .A2(n8396), .ZN(n8465) );
  NAND2_X1 U7417 ( .A1(n8426), .A2(n8425), .ZN(n13729) );
  CLKBUF_X1 U7418 ( .A(n14389), .Z(n6661) );
  CLKBUF_X1 U7419 ( .A(n10276), .Z(n6663) );
  NAND2_X1 U7420 ( .A1(n15007), .A2(n15008), .ZN(n15004) );
  NAND2_X1 U7421 ( .A1(n14950), .A2(n12325), .ZN(n13895) );
  NAND2_X1 U7422 ( .A1(n9417), .A2(n9416), .ZN(n15007) );
  NOR2_X1 U7423 ( .A1(n9416), .A2(n9417), .ZN(n15005) );
  XNOR2_X1 U7424 ( .A(n13752), .B(n13629), .ZN(n13602) );
  OAI21_X1 U7425 ( .B1(n8423), .B2(n8422), .A(n8372), .ZN(n8410) );
  AOI21_X1 U7426 ( .B1(n9917), .B2(n9522), .A(n9521), .ZN(n9934) );
  NAND2_X1 U7427 ( .A1(n14917), .A2(n12318), .ZN(n12322) );
  NAND2_X1 U7428 ( .A1(n12432), .A2(n12431), .ZN(n12583) );
  OR3_X1 U7429 ( .A1(n13046), .A2(n13079), .A3(n13065), .ZN(n12761) );
  NOR2_X1 U7430 ( .A1(n7388), .A2(n14788), .ZN(n15002) );
  NAND2_X1 U7431 ( .A1(n6839), .A2(n7221), .ZN(n7219) );
  AND2_X1 U7433 ( .A1(n12749), .A2(n12750), .ZN(n13052) );
  NAND2_X1 U7434 ( .A1(n9891), .A2(n9890), .ZN(n12453) );
  NAND2_X1 U7435 ( .A1(n9877), .A2(n9876), .ZN(n13258) );
  NAND2_X1 U7436 ( .A1(n7241), .A2(n11998), .ZN(n7243) );
  OAI21_X1 U7437 ( .B1(n11776), .B2(n7434), .A(n7432), .ZN(n7437) );
  OAI21_X2 U7438 ( .B1(n8281), .B2(n11415), .A(n8284), .ZN(n8301) );
  NAND2_X1 U7439 ( .A1(n8759), .A2(n9181), .ZN(n14973) );
  NAND2_X1 U7440 ( .A1(n8938), .A2(n8937), .ZN(n14235) );
  NAND2_X2 U7441 ( .A1(n8152), .A2(n8151), .ZN(n13787) );
  CLKBUF_X2 U7442 ( .A(n12404), .Z(n12409) );
  NAND2_X1 U7443 ( .A1(n10732), .A2(n10733), .ZN(n10731) );
  NAND2_X1 U7444 ( .A1(n7155), .A2(n9504), .ZN(n9829) );
  NAND2_X1 U7445 ( .A1(n10614), .A2(n10613), .ZN(n10612) );
  OAI21_X1 U7446 ( .B1(n10229), .B2(n10210), .A(n10209), .ZN(n10211) );
  NAND2_X1 U7447 ( .A1(n10250), .A2(n10251), .ZN(n10249) );
  NAND2_X1 U7449 ( .A1(n7040), .A2(n7039), .ZN(n10270) );
  OR2_X1 U7450 ( .A1(n12825), .A2(n11389), .ZN(n12669) );
  NAND2_X1 U7451 ( .A1(n6849), .A2(n9493), .ZN(n9752) );
  NAND2_X1 U7452 ( .A1(n7177), .A2(n9208), .ZN(n10276) );
  NAND2_X2 U7453 ( .A1(n6669), .A2(n10286), .ZN(n9591) );
  CLKBUF_X1 U7454 ( .A(n12609), .Z(n6668) );
  BUF_X1 U7455 ( .A(n9569), .Z(n6688) );
  INV_X1 U7456 ( .A(n10788), .ZN(n6848) );
  NAND3_X1 U7458 ( .A1(n9583), .A2(n9582), .A3(n9581), .ZN(n15503) );
  CLKBUF_X2 U7459 ( .A(n9867), .Z(n6684) );
  OAI21_X1 U7460 ( .B1(n9487), .B2(n7143), .A(n7141), .ZN(n9492) );
  XNOR2_X1 U7461 ( .A(n10004), .B(n10003), .ZN(n12268) );
  BUF_X1 U7462 ( .A(n12609), .Z(n6667) );
  NAND2_X2 U7464 ( .A1(n9461), .A2(n9460), .ZN(n9600) );
  BUF_X2 U7465 ( .A(n7802), .Z(n8424) );
  INV_X1 U7466 ( .A(n7917), .ZN(n8437) );
  INV_X1 U7467 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9328) );
  BUF_X2 U7468 ( .A(n9164), .Z(n9154) );
  NAND4_X2 U7469 ( .A1(n8612), .A2(n8611), .A3(n8610), .A4(n8609), .ZN(n13965)
         );
  OR2_X1 U7470 ( .A1(n9526), .A2(n9720), .ZN(n6657) );
  INV_X1 U7471 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n6656) );
  CLKBUF_X1 U7472 ( .A(n7810), .Z(n6670) );
  NAND4_X1 U7473 ( .A1(n7725), .A2(n7724), .A3(n7723), .A4(n7722), .ZN(n8478)
         );
  INV_X2 U7475 ( .A(n7810), .ZN(n7684) );
  INV_X1 U7476 ( .A(n8428), .ZN(n7929) );
  CLKBUF_X1 U7477 ( .A(n7680), .Z(n12273) );
  CLKBUF_X1 U7478 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n6664) );
  INV_X1 U7479 ( .A(n14206), .ZN(n11942) );
  CLKBUF_X1 U7481 ( .A(n8620), .Z(n6658) );
  XNOR2_X1 U7482 ( .A(n7167), .B(n8541), .ZN(n14389) );
  OR2_X1 U7483 ( .A1(n8542), .A2(n8787), .ZN(n7167) );
  INV_X1 U7484 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10809) );
  XNOR2_X1 U7485 ( .A(n7756), .B(n10294), .ZN(n7754) );
  NOR2_X1 U7486 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7663) );
  INV_X1 U7488 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13507) );
  INV_X1 U7489 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7520) );
  INV_X1 U7490 ( .A(n6646), .ZN(n8982) );
  NOR2_X2 U7491 ( .A1(n8963), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n6646) );
  AND2_X1 U7492 ( .A1(n7426), .A2(n6789), .ZN(n11506) );
  NAND4_X1 U7493 ( .A1(n8528), .A2(n8812), .A3(n7647), .A4(n8620), .ZN(n8901)
         );
  AND4_X2 U7494 ( .A1(n8523), .A2(n8524), .A3(n8522), .A4(n8525), .ZN(n8528)
         );
  OAI21_X1 U7495 ( .B1(n12208), .B2(n6933), .A(n6931), .ZN(n12244) );
  OAI21_X1 U7496 ( .B1(n11590), .B2(n11589), .A(n11588), .ZN(n11596) );
  INV_X4 U7497 ( .A(n12353), .ZN(n10208) );
  NAND2_X2 U7498 ( .A1(n10207), .A2(n10206), .ZN(n12353) );
  NAND2_X2 U7499 ( .A1(n15589), .A2(n9391), .ZN(n9393) );
  NOR2_X2 U7501 ( .A1(n15586), .A2(n9387), .ZN(n9389) );
  NOR2_X2 U7502 ( .A1(n9329), .A2(n6863), .ZN(n9331) );
  NOR2_X2 U7503 ( .A1(n15593), .A2(n9400), .ZN(n9403) );
  NOR2_X2 U7504 ( .A1(n9421), .A2(n9420), .ZN(n15017) );
  NAND2_X2 U7505 ( .A1(n6828), .A2(n8456), .ZN(n8463) );
  INV_X1 U7506 ( .A(n7730), .ZN(n7759) );
  NAND2_X1 U7507 ( .A1(n7504), .A2(n7503), .ZN(n8349) );
  NAND2_X1 U7509 ( .A1(n11843), .A2(n9689), .ZN(n11977) );
  NAND2_X1 U7510 ( .A1(n9812), .A2(n9811), .ZN(n13116) );
  OAI21_X1 U7511 ( .B1(n13243), .B2(n13013), .A(n12997), .ZN(n12984) );
  NAND2_X1 U7512 ( .A1(n7338), .A2(n6711), .ZN(n13155) );
  NAND2_X1 U7513 ( .A1(n13015), .A2(n9913), .ZN(n12999) );
  NAND2_X1 U7514 ( .A1(n7337), .A2(n9615), .ZN(n11555) );
  NAND2_X2 U7515 ( .A1(n9559), .A2(n15607), .ZN(n10788) );
  INV_X1 U7517 ( .A(n9730), .ZN(n12074) );
  OAI21_X1 U7518 ( .B1(n13233), .B2(n15568), .A(n6650), .ZN(P3_U3455) );
  XNOR2_X1 U7519 ( .A(n8495), .B(n13504), .ZN(n6654) );
  XNOR2_X2 U7520 ( .A(n6657), .B(n6656), .ZN(n9968) );
  XNOR2_X2 U7522 ( .A(n8301), .B(SI_24_), .ZN(n8299) );
  NAND2_X2 U7523 ( .A1(n7758), .A2(n7757), .ZN(n7776) );
  AND2_X2 U7524 ( .A1(n11232), .A2(n11231), .ZN(n11237) );
  AND2_X2 U7525 ( .A1(n9637), .A2(n7482), .ZN(n9746) );
  INV_X2 U7526 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U7527 ( .A1(n7450), .A2(n11006), .ZN(n11007) );
  NAND4_X1 U7528 ( .A1(n9571), .A2(n9574), .A3(n9572), .A4(n9573), .ZN(n10994)
         );
  OAI21_X1 U7529 ( .B1(n13573), .B2(n13574), .A(n13572), .ZN(n13576) );
  NAND2_X1 U7530 ( .A1(n13573), .A2(n13574), .ZN(n13572) );
  NAND2_X2 U7531 ( .A1(n8894), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8586) );
  NOR2_X1 U7532 ( .A1(n12974), .A2(n12783), .ZN(n6659) );
  NAND2_X2 U7533 ( .A1(n14377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8544) );
  OAI21_X2 U7534 ( .B1(n11905), .B2(n7182), .A(n7179), .ZN(n12116) );
  NAND2_X2 U7535 ( .A1(n7578), .A2(n9220), .ZN(n11905) );
  NAND2_X2 U7536 ( .A1(n9702), .A2(n9700), .ZN(n9487) );
  OAI21_X2 U7537 ( .B1(n9752), .B2(n10620), .A(n9493), .ZN(n9765) );
  OAI21_X1 U7538 ( .B1(n13744), .B2(n15301), .A(n6666), .ZN(n6665) );
  INV_X2 U7539 ( .A(n7685), .ZN(n7057) );
  INV_X2 U7540 ( .A(n7845), .ZN(n7917) );
  OR2_X1 U7541 ( .A1(n13887), .A2(n7431), .ZN(n7430) );
  INV_X1 U7542 ( .A(n12424), .ZN(n9461) );
  INV_X1 U7543 ( .A(n12780), .ZN(n12794) );
  INV_X1 U7544 ( .A(n13316), .ZN(n10161) );
  INV_X1 U7545 ( .A(n10362), .ZN(n8170) );
  AND2_X1 U7546 ( .A1(n13948), .A2(n7430), .ZN(n7429) );
  AOI21_X1 U7547 ( .B1(n7427), .B2(n6922), .A(n6921), .ZN(n6920) );
  INV_X1 U7548 ( .A(n13056), .ZN(n12554) );
  NAND2_X1 U7550 ( .A1(n12787), .A2(n12790), .ZN(n12974) );
  NAND2_X2 U7553 ( .A1(n8286), .A2(n8285), .ZN(n13752) );
  NOR2_X1 U7554 ( .A1(n7494), .A2(n7675), .ZN(n7696) );
  NAND2_X1 U7555 ( .A1(n7295), .A2(n8773), .ZN(n12097) );
  AOI21_X1 U7556 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(n9412), .A(n15000), .ZN(
        n9413) );
  NAND2_X1 U7558 ( .A1(n9530), .A2(n9529), .ZN(n9947) );
  NAND2_X1 U7559 ( .A1(n10005), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10004) );
  INV_X1 U7560 ( .A(n10302), .ZN(n10286) );
  NOR2_X1 U7561 ( .A1(n15002), .A2(n15001), .ZN(n15000) );
  INV_X1 U7562 ( .A(n11145), .ZN(n13964) );
  NAND2_X1 U7563 ( .A1(n12424), .A2(n9460), .ZN(n12609) );
  INV_X1 U7564 ( .A(n10861), .ZN(n10146) );
  AOI21_X2 U7565 ( .B1(n12281), .B2(n15495), .A(n12278), .ZN(n12279) );
  AND2_X2 U7566 ( .A1(n9299), .A2(n10911), .ZN(n9298) );
  OAI222_X1 U7567 ( .A1(P3_U3151), .A2(n12424), .B1(n12306), .B2(n12601), .C1(
        n12604), .C2(n12423), .ZN(P3_U3265) );
  NAND2_X1 U7568 ( .A1(n9968), .A2(n12936), .ZN(n6669) );
  OR2_X1 U7569 ( .A1(n9591), .A2(SI_3_), .ZN(n9595) );
  OAI21_X2 U7570 ( .B1(n7774), .B2(n7501), .A(n7777), .ZN(n7799) );
  XNOR2_X2 U7571 ( .A(n7776), .B(SI_2_), .ZN(n7774) );
  OR2_X2 U7572 ( .A1(n14786), .A2(n14787), .ZN(n7390) );
  AOI21_X2 U7573 ( .B1(n7429), .B2(n7431), .A(n6754), .ZN(n7427) );
  OAI21_X2 U7574 ( .B1(n9829), .B2(n9505), .A(n9506), .ZN(n9842) );
  NAND2_X2 U7575 ( .A1(n12168), .A2(n12167), .ZN(n12166) );
  XNOR2_X2 U7577 ( .A(n8367), .B(n8366), .ZN(n8365) );
  OAI21_X2 U7578 ( .B1(n8349), .B2(n8348), .A(n8347), .ZN(n8367) );
  XNOR2_X2 U7579 ( .A(n12456), .B(n12454), .ZN(n12555) );
  NAND2_X1 U7580 ( .A1(n12273), .A2(n7683), .ZN(n7810) );
  AOI21_X2 U7581 ( .B1(n12973), .B2(n12790), .A(n9994), .ZN(n12620) );
  NOR2_X2 U7582 ( .A1(n12274), .A2(n12788), .ZN(n12973) );
  NAND2_X2 U7583 ( .A1(n7733), .A2(n7062), .ZN(n7756) );
  NAND2_X2 U7584 ( .A1(n8802), .A2(n8801), .ZN(n14342) );
  NAND2_X1 U7586 ( .A1(n7683), .A2(n7682), .ZN(n8431) );
  OAI21_X2 U7587 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n9384), .A(n14770), .ZN(
        n15597) );
  NOR2_X2 U7588 ( .A1(n9332), .A2(n9333), .ZN(n9334) );
  NAND2_X1 U7589 ( .A1(n7269), .A2(n7272), .ZN(n14076) );
  XNOR2_X2 U7591 ( .A(n8283), .B(n8282), .ZN(n8281) );
  NOR2_X2 U7592 ( .A1(n14075), .A2(n7363), .ZN(n7362) );
  XNOR2_X2 U7593 ( .A(n9328), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n9378) );
  NAND2_X2 U7594 ( .A1(n9100), .A2(n9101), .ZN(n14217) );
  NAND2_X1 U7595 ( .A1(n8261), .A2(n8260), .ZN(n13759) );
  AND2_X1 U7596 ( .A1(n10843), .A2(n11100), .ZN(n11439) );
  NAND2_X2 U7597 ( .A1(n12669), .A2(n12668), .ZN(n12626) );
  INV_X1 U7598 ( .A(n8473), .ZN(n7176) );
  INV_X2 U7599 ( .A(n10067), .ZN(n8476) );
  INV_X2 U7600 ( .A(n9167), .ZN(n9142) );
  CLKBUF_X2 U7601 ( .A(n11511), .Z(n12404) );
  NAND2_X2 U7602 ( .A1(n10362), .A2(n10302), .ZN(n8030) );
  OAI21_X1 U7604 ( .B1(n8982), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8965) );
  AND3_X1 U7605 ( .A1(n14098), .A2(n14097), .A3(n14096), .ZN(n14291) );
  NOR2_X1 U7606 ( .A1(n12284), .A2(n6748), .ZN(n13172) );
  AOI21_X1 U7607 ( .B1(n7002), .B2(n7001), .A(n6766), .ZN(n7000) );
  NOR2_X1 U7608 ( .A1(n7654), .A2(n14282), .ZN(n14283) );
  MUX2_X1 U7609 ( .A(n13238), .B(n13237), .S(n15570), .Z(n13239) );
  AND2_X1 U7610 ( .A1(n13537), .A2(n13536), .ZN(n13731) );
  MUX2_X1 U7611 ( .A(n13177), .B(n13237), .S(n15585), .Z(n13178) );
  NAND2_X1 U7612 ( .A1(n7486), .A2(n10146), .ZN(n13723) );
  OR2_X1 U7613 ( .A1(n8298), .A2(n6897), .ZN(n6895) );
  AOI21_X1 U7614 ( .B1(n7211), .B2(n13586), .A(n13554), .ZN(n13740) );
  OR2_X1 U7615 ( .A1(n14122), .A2(n14123), .ZN(n14120) );
  NAND2_X1 U7616 ( .A1(n10168), .A2(n7565), .ZN(n7563) );
  CLKBUF_X2 U7617 ( .A(n14274), .Z(n6685) );
  OR2_X1 U7618 ( .A1(n13593), .A2(n13594), .ZN(n13591) );
  AOI21_X1 U7620 ( .B1(n12272), .B2(n9154), .A(n6826), .ZN(n14277) );
  NAND2_X1 U7621 ( .A1(n6961), .A2(n6840), .ZN(n10164) );
  AND2_X1 U7622 ( .A1(n12786), .A2(n9993), .ZN(n12645) );
  NOR2_X1 U7623 ( .A1(n12931), .A2(n12930), .ZN(n12932) );
  AOI211_X1 U7624 ( .C1(n12954), .C2(n12953), .A(n12952), .B(n12951), .ZN(
        n12955) );
  AOI21_X1 U7625 ( .B1(n7204), .B2(n7208), .A(n7203), .ZN(n7202) );
  NAND2_X1 U7626 ( .A1(n7017), .A2(n7016), .ZN(n12931) );
  OAI21_X1 U7627 ( .B1(n8395), .B2(n8393), .A(n8379), .ZN(n8382) );
  XNOR2_X1 U7628 ( .A(n8395), .B(n8394), .ZN(n12272) );
  NAND2_X1 U7629 ( .A1(n8377), .A2(n8376), .ZN(n8395) );
  OAI21_X1 U7630 ( .B1(n12547), .B2(n12446), .A(n12448), .ZN(n12499) );
  OAI21_X1 U7631 ( .B1(n10153), .B2(n6962), .A(n10160), .ZN(n6841) );
  NAND2_X1 U7632 ( .A1(n9936), .A2(n9935), .ZN(n12470) );
  OR2_X1 U7633 ( .A1(n10152), .A2(n6962), .ZN(n6961) );
  OR2_X1 U7634 ( .A1(n14833), .A2(n7018), .ZN(n7017) );
  NAND2_X1 U7635 ( .A1(n8824), .A2(n7308), .ZN(n14208) );
  AOI21_X1 U7636 ( .B1(n13373), .B2(n13302), .A(n13377), .ZN(n10152) );
  NAND2_X2 U7637 ( .A1(n7061), .A2(n8567), .ZN(n14285) );
  NAND2_X1 U7638 ( .A1(n8324), .A2(n8323), .ZN(n13742) );
  OR2_X1 U7639 ( .A1(n7207), .A2(n13580), .ZN(n7206) );
  NAND2_X1 U7640 ( .A1(n8888), .A2(n8887), .ZN(n14112) );
  XNOR2_X1 U7641 ( .A(n8423), .B(n8422), .ZN(n14387) );
  OAI21_X1 U7642 ( .B1(n15021), .B2(n15022), .A(n7375), .ZN(n7374) );
  OR2_X1 U7643 ( .A1(n12324), .A2(n12323), .ZN(n12325) );
  NAND2_X1 U7644 ( .A1(n14914), .A2(n12314), .ZN(n14917) );
  OR2_X1 U7645 ( .A1(n9517), .A2(n12190), .ZN(n9519) );
  NAND2_X1 U7646 ( .A1(n8861), .A2(n8860), .ZN(n14313) );
  AOI21_X1 U7647 ( .B1(n8302), .B2(n7506), .A(n7505), .ZN(n7503) );
  NAND2_X1 U7648 ( .A1(n11937), .A2(n9069), .ZN(n12086) );
  OR2_X1 U7649 ( .A1(n14229), .A2(n14199), .ZN(n9100) );
  AND2_X1 U7650 ( .A1(n14912), .A2(n14913), .ZN(n12314) );
  NAND2_X1 U7651 ( .A1(n11938), .A2(n11944), .ZN(n11937) );
  NAND2_X1 U7652 ( .A1(n8172), .A2(n8171), .ZN(n13782) );
  NAND2_X1 U7653 ( .A1(n12244), .A2(n12243), .ZN(n14914) );
  OAI21_X1 U7654 ( .B1(n11725), .B2(n7551), .A(n7549), .ZN(n6976) );
  INV_X1 U7655 ( .A(n14212), .ZN(n14329) );
  NAND2_X1 U7656 ( .A1(n8837), .A2(n8836), .ZN(n14324) );
  NAND2_X1 U7657 ( .A1(n7542), .A2(n9271), .ZN(n12113) );
  AND2_X1 U7658 ( .A1(n12843), .A2(n7418), .ZN(n12846) );
  CLKBUF_X1 U7659 ( .A(n8258), .Z(n8846) );
  NAND2_X1 U7660 ( .A1(n12050), .A2(n12049), .ZN(n12141) );
  OR2_X1 U7661 ( .A1(n12036), .A2(n9270), .ZN(n7542) );
  XNOR2_X1 U7662 ( .A(n8169), .B(n8168), .ZN(n8811) );
  NAND3_X1 U7663 ( .A1(n7417), .A2(P3_REG2_REG_13__SCAN_IN), .A3(n12843), .ZN(
        n7418) );
  OAI21_X1 U7664 ( .B1(n8166), .B2(n8165), .A(n8167), .ZN(n8169) );
  NAND4_X1 U7665 ( .A1(n7243), .A2(n7244), .A3(n7242), .A4(n12049), .ZN(n12050) );
  NAND2_X1 U7666 ( .A1(n8750), .A2(n8749), .ZN(n14971) );
  XNOR2_X1 U7667 ( .A(n8189), .B(n10654), .ZN(n8166) );
  NAND2_X1 U7668 ( .A1(n11995), .A2(n7245), .ZN(n12049) );
  OAI21_X1 U7669 ( .B1(n8147), .B2(n7084), .A(n6699), .ZN(n8232) );
  NAND2_X1 U7670 ( .A1(n8038), .A2(n8037), .ZN(n12039) );
  NAND2_X1 U7671 ( .A1(n8098), .A2(n8097), .ZN(n8118) );
  OR3_X1 U7672 ( .A1(n7898), .A2(n7897), .A3(n6909), .ZN(n6904) );
  NAND2_X1 U7673 ( .A1(n11357), .A2(n9215), .ZN(n11423) );
  NAND2_X1 U7674 ( .A1(n14782), .A2(n9405), .ZN(n9407) );
  NAND2_X1 U7675 ( .A1(n11444), .A2(n9214), .ZN(n11357) );
  AOI22_X1 U7676 ( .A1(n11510), .A2(n11509), .B1(n11508), .B2(n11507), .ZN(
        n11590) );
  XNOR2_X1 U7677 ( .A(n15177), .B(n8921), .ZN(n11371) );
  NAND2_X1 U7678 ( .A1(n7928), .A2(n7927), .ZN(n15355) );
  NAND2_X1 U7679 ( .A1(n7909), .A2(n7908), .ZN(n11484) );
  NAND2_X1 U7680 ( .A1(n8670), .A2(n8669), .ZN(n15177) );
  NAND2_X1 U7681 ( .A1(n11439), .A2(n15343), .ZN(n11438) );
  INV_X2 U7682 ( .A(n15501), .ZN(n13166) );
  NAND2_X2 U7683 ( .A1(n11008), .A2(n15506), .ZN(n15505) );
  NAND2_X2 U7684 ( .A1(n10801), .A2(n15479), .ZN(n15501) );
  OR2_X1 U7685 ( .A1(n9864), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U7686 ( .A1(n7901), .A2(n7900), .ZN(n7904) );
  NAND2_X1 U7687 ( .A1(n9492), .A2(n10618), .ZN(n9493) );
  OR2_X1 U7688 ( .A1(n9492), .A2(n10618), .ZN(n6849) );
  OR2_X1 U7689 ( .A1(n10192), .A2(n10186), .ZN(n13417) );
  AND2_X1 U7690 ( .A1(n12678), .A2(n12682), .ZN(n12676) );
  NOR2_X1 U7691 ( .A1(n10860), .A2(n10780), .ZN(n10843) );
  INV_X1 U7692 ( .A(n15470), .ZN(n6673) );
  AND2_X1 U7693 ( .A1(n9210), .A2(n8481), .ZN(n10762) );
  NAND2_X1 U7694 ( .A1(n9579), .A2(n9580), .ZN(n10802) );
  NAND2_X1 U7695 ( .A1(n9485), .A2(n9484), .ZN(n9702) );
  AND2_X1 U7696 ( .A1(n8623), .A2(n8622), .ZN(n15149) );
  NAND2_X1 U7697 ( .A1(n7809), .A2(n7808), .ZN(n10780) );
  NAND4_X2 U7698 ( .A1(n9588), .A2(n9587), .A3(n9586), .A4(n9585), .ZN(n12825)
         );
  NAND4_X1 U7699 ( .A1(n9553), .A2(n9552), .A3(n9551), .A4(n9550), .ZN(n12826)
         );
  INV_X1 U7700 ( .A(n6946), .ZN(n11150) );
  AOI21_X1 U7701 ( .B1(n7075), .B2(n7079), .A(n7073), .ZN(n7072) );
  OR2_X1 U7702 ( .A1(n9591), .A2(n10294), .ZN(n9583) );
  AND2_X1 U7703 ( .A1(n8607), .A2(n8608), .ZN(n6946) );
  CLKBUF_X2 U7704 ( .A(n8478), .Z(n10062) );
  BUF_X2 U7705 ( .A(n9591), .Z(n6687) );
  NAND4_X2 U7706 ( .A1(n7840), .A2(n7839), .A3(n7838), .A4(n7837), .ZN(n13449)
         );
  OR2_X1 U7707 ( .A1(n9805), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9820) );
  AND4_X1 U7708 ( .A1(n8618), .A2(n8617), .A3(n8616), .A4(n8615), .ZN(n11145)
         );
  INV_X1 U7709 ( .A(n14262), .ZN(n6857) );
  OAI21_X1 U7710 ( .B1(n10979), .B2(n11388), .A(n10966), .ZN(n10967) );
  NAND2_X1 U7711 ( .A1(n10980), .A2(n7034), .ZN(n10959) );
  AND3_X1 U7712 ( .A1(n8584), .A2(n8583), .A3(n8582), .ZN(n15124) );
  INV_X1 U7713 ( .A(n9459), .ZN(n9460) );
  AOI21_X1 U7714 ( .B1(n7069), .B2(n7071), .A(n7941), .ZN(n7068) );
  CLKBUF_X1 U7715 ( .A(n8973), .Z(n15111) );
  AOI21_X1 U7716 ( .B1(n7923), .B2(n7070), .A(n6772), .ZN(n7069) );
  INV_X1 U7717 ( .A(n8320), .ZN(n7505) );
  AND2_X1 U7718 ( .A1(n7708), .A2(n10262), .ZN(n10911) );
  NAND2_X1 U7719 ( .A1(n8496), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7688) );
  AND2_X1 U7720 ( .A1(n6677), .A2(n10286), .ZN(n8600) );
  AND2_X1 U7721 ( .A1(n6677), .A2(n10302), .ZN(n9164) );
  NAND2_X1 U7722 ( .A1(n7703), .A2(n7702), .ZN(n12270) );
  XNOR2_X1 U7723 ( .A(n7677), .B(n13835), .ZN(n7680) );
  NAND2_X1 U7724 ( .A1(n8904), .A2(n8963), .ZN(n11079) );
  NAND2_X1 U7725 ( .A1(n13834), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7677) );
  XNOR2_X1 U7726 ( .A(n8907), .B(n8906), .ZN(n11834) );
  AND2_X2 U7727 ( .A1(n8813), .A2(n6728), .ZN(n8542) );
  INV_X1 U7728 ( .A(n7336), .ZN(n7333) );
  XOR2_X1 U7729 ( .A(n9378), .B(n9379), .Z(n9381) );
  AND3_X2 U7730 ( .A1(n8528), .A2(n8620), .A3(n7647), .ZN(n8813) );
  NAND2_X1 U7731 ( .A1(n9380), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9379) );
  AND2_X1 U7732 ( .A1(n9330), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6863) );
  AND2_X1 U7733 ( .A1(n9465), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U7734 ( .A1(n10316), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9469) );
  NAND4_X1 U7735 ( .A1(n7466), .A2(n9564), .A3(n9443), .A4(n10809), .ZN(n9606)
         );
  AND2_X1 U7736 ( .A1(n8533), .A2(n8532), .ZN(n8812) );
  AND3_X1 U7737 ( .A1(n8531), .A2(n8530), .A3(n8529), .ZN(n8968) );
  INV_X1 U7738 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9380) );
  NOR2_X1 U7739 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8522) );
  NOR2_X1 U7740 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8523) );
  NOR2_X1 U7741 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8524) );
  NOR2_X1 U7742 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n8532) );
  NOR2_X1 U7743 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n8533) );
  INV_X4 U7744 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7745 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7746 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8527) );
  INV_X1 U7747 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8127) );
  INV_X1 U7748 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8639) );
  INV_X1 U7749 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8643) );
  NOR2_X1 U7750 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n9450) );
  INV_X4 U7751 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7752 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8543) );
  NOR2_X1 U7753 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n9451) );
  INV_X1 U7754 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9698) );
  INV_X1 U7755 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9744) );
  NOR2_X1 U7756 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n7015) );
  NOR2_X2 U7757 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7466) );
  INV_X1 U7758 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9443) );
  INV_X1 U7759 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8964) );
  INV_X1 U7760 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U7761 ( .A1(n9461), .A2(n9459), .ZN(n9867) );
  NOR2_X1 U7762 ( .A1(n14776), .A2(n14775), .ZN(n14774) );
  XNOR2_X1 U7763 ( .A(n9393), .B(n9392), .ZN(n14776) );
  OAI21_X1 U7764 ( .B1(n10011), .B2(n7333), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9458) );
  OAI21_X1 U7765 ( .B1(n9636), .B2(n9477), .A(n9478), .ZN(n6675) );
  XNOR2_X1 U7766 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n6676) );
  OAI21_X1 U7767 ( .B1(n9636), .B2(n9477), .A(n9478), .ZN(n9655) );
  XNOR2_X1 U7768 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n9562) );
  AND2_X2 U7769 ( .A1(n8549), .A2(n8548), .ZN(n8851) );
  AOI21_X1 U7770 ( .B1(n12262), .B2(n15198), .A(n7358), .ZN(n7357) );
  NAND2_X1 U7771 ( .A1(n9706), .A2(n9705), .ZN(n14850) );
  OAI22_X1 U7772 ( .A1(n10229), .A2(n14261), .B1(n15124), .B2(n12363), .ZN(
        n10218) );
  NAND2_X1 U7773 ( .A1(n14071), .A2(n8951), .ZN(n7172) );
  NAND4_X2 U7774 ( .A1(n8597), .A2(n8595), .A3(n8594), .A4(n8596), .ZN(n14267)
         );
  NAND2_X2 U7775 ( .A1(n9297), .A2(n13504), .ZN(n10061) );
  OAI21_X2 U7776 ( .B1(n15080), .B2(n8919), .A(n8920), .ZN(n11367) );
  NAND2_X1 U7777 ( .A1(n8918), .A2(n8917), .ZN(n15080) );
  NAND2_X1 U7778 ( .A1(n9568), .A2(n10788), .ZN(n12657) );
  NAND2_X1 U7779 ( .A1(n9009), .A2(n9010), .ZN(n14264) );
  NAND2_X1 U7780 ( .A1(n14389), .A2(n15026), .ZN(n6677) );
  INV_X1 U7781 ( .A(n8754), .ZN(n6678) );
  INV_X1 U7782 ( .A(n8796), .ZN(n6679) );
  NAND2_X1 U7783 ( .A1(n8549), .A2(n14386), .ZN(n8754) );
  OAI222_X1 U7784 ( .A1(P1_U3086), .A2(n14386), .B1(n14398), .B2(n14385), .C1(
        n14597), .C2(n14395), .ZN(P1_U3326) );
  NAND2_X1 U7785 ( .A1(n9968), .A2(n12936), .ZN(n6680) );
  NAND2_X2 U7786 ( .A1(n9968), .A2(n12936), .ZN(n10807) );
  NAND2_X4 U7787 ( .A1(n7448), .A2(n7447), .ZN(n13966) );
  BUF_X1 U7788 ( .A(n13749), .Z(n6682) );
  CLKBUF_X2 U7789 ( .A(n7917), .Z(n7843) );
  NAND4_X4 U7790 ( .A1(n8585), .A2(n8587), .A3(n8588), .A4(n8586), .ZN(n14262)
         );
  NAND2_X1 U7791 ( .A1(n13155), .A2(n13156), .ZN(n13139) );
  XNOR2_X1 U7792 ( .A(n10848), .B(n13449), .ZN(n10836) );
  AND2_X1 U7793 ( .A1(n7709), .A2(n11719), .ZN(n9296) );
  XNOR2_X2 U7794 ( .A(n7691), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7709) );
  AOI21_X2 U7795 ( .B1(n11367), .B2(n8923), .A(n8922), .ZN(n15066) );
  OAI21_X2 U7796 ( .B1(n15471), .B2(n7350), .A(n6755), .ZN(n11843) );
  NAND2_X2 U7797 ( .A1(n11529), .A2(n9643), .ZN(n15471) );
  AOI21_X2 U7798 ( .B1(n13139), .B2(n9798), .A(n6722), .ZN(n13127) );
  OAI21_X2 U7799 ( .B1(n9008), .B2(n9175), .A(n9010), .ZN(n11190) );
  NAND2_X2 U7800 ( .A1(n6857), .A2(n6858), .ZN(n9175) );
  OAI21_X2 U7801 ( .B1(n8933), .B2(n7163), .A(n7161), .ZN(n14236) );
  OAI222_X1 U7802 ( .A1(P1_U3086), .A2(n14384), .B1(n14383), .B2(n14382), .C1(
        n14381), .C2(n14395), .ZN(P1_U3325) );
  NAND2_X2 U7803 ( .A1(n12086), .A2(n7298), .ZN(n8933) );
  NAND2_X4 U7804 ( .A1(n10208), .A2(n15125), .ZN(n10229) );
  INV_X2 U7805 ( .A(n9152), .ZN(n8593) );
  NAND2_X2 U7806 ( .A1(n14384), .A2(n8548), .ZN(n9152) );
  AND2_X1 U7807 ( .A1(n9459), .A2(n12424), .ZN(n9569) );
  NOR2_X1 U7808 ( .A1(n12645), .A2(n7345), .ZN(n7344) );
  INV_X1 U7809 ( .A(n9930), .ZN(n7345) );
  AND2_X1 U7810 ( .A1(n10802), .A2(n9978), .ZN(n15504) );
  NOR2_X1 U7811 ( .A1(n9234), .A2(n7194), .ZN(n7191) );
  INV_X1 U7812 ( .A(n7051), .ZN(n7050) );
  OAI21_X1 U7813 ( .B1(n7053), .B2(n7052), .A(n13657), .ZN(n7051) );
  INV_X1 U7814 ( .A(n7760), .ZN(n7802) );
  NAND2_X1 U7815 ( .A1(n9247), .A2(n10489), .ZN(n9208) );
  AND3_X1 U7816 ( .A1(n7673), .A2(n7672), .A3(n7671), .ZN(n8505) );
  INV_X1 U7817 ( .A(n12394), .ZN(n7431) );
  NOR2_X1 U7818 ( .A1(n7305), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n7302) );
  OR2_X1 U7819 ( .A1(n11381), .A2(n11061), .ZN(n12650) );
  NAND2_X1 U7820 ( .A1(n13109), .A2(n6739), .ZN(n7474) );
  OR2_X1 U7821 ( .A1(n13267), .A2(n13118), .ZN(n12740) );
  NOR2_X1 U7822 ( .A1(n9964), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n9962) );
  AOI21_X1 U7823 ( .B1(n10848), .B2(n8437), .A(n7844), .ZN(n7848) );
  NAND2_X1 U7824 ( .A1(n7631), .A2(n7633), .ZN(n7629) );
  INV_X1 U7825 ( .A(n7634), .ZN(n7631) );
  AND2_X1 U7826 ( .A1(n8093), .A2(n8094), .ZN(n7638) );
  AND2_X1 U7827 ( .A1(n9102), .A2(n7287), .ZN(n7286) );
  OR2_X1 U7828 ( .A1(n7614), .A2(n8163), .ZN(n6702) );
  INV_X1 U7829 ( .A(n8162), .ZN(n7614) );
  NAND2_X1 U7830 ( .A1(n6898), .A2(n6743), .ZN(n6896) );
  AOI21_X1 U7831 ( .B1(n6699), .B2(n7084), .A(n8231), .ZN(n7080) );
  NOR2_X1 U7832 ( .A1(n8318), .A2(n6770), .ZN(n7619) );
  NOR2_X1 U7833 ( .A1(n14925), .A2(n12029), .ZN(n6959) );
  NAND2_X1 U7834 ( .A1(n8121), .A2(n10579), .ZN(n8148) );
  NAND2_X1 U7835 ( .A1(n12618), .A2(n12616), .ZN(n12623) );
  OR2_X1 U7836 ( .A1(n12968), .A2(n12977), .ZN(n12792) );
  NOR2_X1 U7837 ( .A1(n12470), .A2(n9945), .ZN(n9946) );
  NAND2_X1 U7838 ( .A1(n9928), .A2(n9927), .ZN(n9929) );
  NAND2_X1 U7839 ( .A1(n13008), .A2(n13009), .ZN(n12773) );
  OR2_X1 U7840 ( .A1(n12767), .A2(n13043), .ZN(n13009) );
  OR2_X1 U7841 ( .A1(n12453), .A2(n12554), .ZN(n12756) );
  NAND2_X1 U7842 ( .A1(n13116), .A2(n13115), .ZN(n9827) );
  OR2_X1 U7843 ( .A1(n12821), .A2(n11824), .ZN(n12694) );
  OR2_X1 U7844 ( .A1(n12823), .A2(n15546), .ZN(n12686) );
  OR2_X1 U7845 ( .A1(n10792), .A2(n11001), .ZN(n10046) );
  OR2_X1 U7846 ( .A1(n10472), .A2(n10028), .ZN(n10049) );
  INV_X1 U7847 ( .A(n12810), .ZN(n10032) );
  NOR2_X1 U7848 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), .ZN(
        n7215) );
  INV_X1 U7849 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n10029) );
  INV_X1 U7850 ( .A(n13365), .ZN(n7565) );
  INV_X1 U7851 ( .A(n12293), .ZN(n7683) );
  NAND2_X1 U7852 ( .A1(n13549), .A2(n7603), .ZN(n7601) );
  INV_X1 U7853 ( .A(n7605), .ZN(n7603) );
  NAND2_X1 U7854 ( .A1(n9249), .A2(n9248), .ZN(n7525) );
  XNOR2_X1 U7855 ( .A(n7698), .B(n7697), .ZN(n8516) );
  NAND2_X1 U7856 ( .A1(n7699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7698) );
  NAND2_X1 U7857 ( .A1(n13966), .A2(n15124), .ZN(n9009) );
  NAND2_X1 U7858 ( .A1(n8953), .A2(n11079), .ZN(n9170) );
  NOR2_X1 U7859 ( .A1(n9170), .A2(n8961), .ZN(n8973) );
  AND2_X1 U7860 ( .A1(n8119), .A2(n8101), .ZN(n8117) );
  OAI22_X1 U7861 ( .A1(n9351), .A2(P1_ADDR_REG_11__SCAN_IN), .B1(n9410), .B2(
        n9350), .ZN(n9415) );
  AOI21_X1 U7862 ( .B1(n7248), .B2(n7247), .A(n6773), .ZN(n7246) );
  INV_X1 U7863 ( .A(n7251), .ZN(n7247) );
  NAND2_X1 U7864 ( .A1(n6698), .A2(n7231), .ZN(n7230) );
  OR2_X1 U7865 ( .A1(n7238), .A2(n6727), .ZN(n7231) );
  NAND2_X1 U7866 ( .A1(n12465), .A2(n13013), .ZN(n7240) );
  INV_X1 U7867 ( .A(n12936), .ZN(n10825) );
  NAND2_X1 U7868 ( .A1(n12620), .A2(n12792), .ZN(n7002) );
  INV_X1 U7869 ( .A(n9600), .ZN(n9954) );
  OR3_X1 U7870 ( .A1(n11883), .A2(n12268), .A3(n11976), .ZN(n10922) );
  INV_X1 U7871 ( .A(n6688), .ZN(n9908) );
  NAND2_X1 U7872 ( .A1(n10981), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10980) );
  XNOR2_X1 U7873 ( .A(n7037), .B(n7036), .ZN(n14826) );
  NAND2_X1 U7874 ( .A1(n7348), .A2(n7346), .ZN(n12976) );
  AND2_X1 U7875 ( .A1(n12974), .A2(n7347), .ZN(n7346) );
  INV_X1 U7876 ( .A(n9946), .ZN(n7347) );
  OR2_X1 U7877 ( .A1(n7005), .A2(n12624), .ZN(n6861) );
  OR2_X1 U7878 ( .A1(n13264), .A2(n13100), .ZN(n12758) );
  AND2_X1 U7879 ( .A1(n13095), .A2(n12736), .ZN(n7481) );
  NAND2_X1 U7880 ( .A1(n14857), .A2(n12703), .ZN(n12077) );
  INV_X1 U7881 ( .A(n12711), .ZN(n9987) );
  NAND2_X1 U7882 ( .A1(n11838), .A2(n9984), .ZN(n7009) );
  OR2_X1 U7883 ( .A1(n10995), .A2(n12794), .ZN(n15509) );
  NAND2_X2 U7884 ( .A1(n6680), .A2(n10302), .ZN(n9742) );
  INV_X1 U7885 ( .A(n9742), .ZN(n12602) );
  AND2_X1 U7886 ( .A1(n10922), .A2(n10471), .ZN(n10932) );
  NAND2_X1 U7887 ( .A1(n10032), .A2(n12651), .ZN(n15545) );
  NAND2_X1 U7888 ( .A1(n10013), .A2(n10014), .ZN(n10472) );
  AND2_X1 U7889 ( .A1(n13845), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U7890 ( .A(n9963), .B(P3_IR_REG_21__SCAN_IN), .ZN(n11381) );
  NAND2_X1 U7891 ( .A1(n9847), .A2(n9846), .ZN(n9964) );
  INV_X1 U7892 ( .A(n7570), .ZN(n6982) );
  INV_X1 U7893 ( .A(n10090), .ZN(n6980) );
  NAND2_X1 U7894 ( .A1(n7558), .A2(n7557), .ZN(n7556) );
  NAND2_X1 U7895 ( .A1(n13312), .A2(n13318), .ZN(n7557) );
  NAND2_X1 U7896 ( .A1(n7560), .A2(n7559), .ZN(n7558) );
  INV_X1 U7897 ( .A(n13318), .ZN(n7559) );
  INV_X1 U7898 ( .A(n6975), .ZN(n6970) );
  AOI21_X1 U7899 ( .B1(n6969), .B2(n13331), .A(n6970), .ZN(n6968) );
  INV_X1 U7900 ( .A(n6974), .ZN(n6969) );
  NAND2_X2 U7901 ( .A1(n8516), .A2(n12270), .ZN(n10362) );
  AND2_X1 U7902 ( .A1(n11829), .A2(n7709), .ZN(n10360) );
  OR3_X1 U7903 ( .A1(n10196), .A2(n10195), .A3(n15311), .ZN(n10192) );
  AND2_X1 U7904 ( .A1(n15246), .A2(n15245), .ZN(n15248) );
  NAND2_X1 U7905 ( .A1(n12292), .A2(n8424), .ZN(n7502) );
  NAND2_X1 U7906 ( .A1(n6866), .A2(n6865), .ZN(n13565) );
  NOR2_X1 U7907 ( .A1(n13742), .A2(n7488), .ZN(n6865) );
  INV_X1 U7908 ( .A(n13642), .ZN(n6866) );
  AOI21_X1 U7909 ( .B1(n7187), .B2(n7186), .A(n7594), .ZN(n7185) );
  AND2_X1 U7910 ( .A1(n13765), .A2(n13662), .ZN(n7594) );
  INV_X1 U7911 ( .A(n7191), .ZN(n7186) );
  NOR2_X1 U7912 ( .A1(n7054), .A2(n9282), .ZN(n7053) );
  INV_X1 U7913 ( .A(n9281), .ZN(n7054) );
  AOI21_X1 U7914 ( .B1(n9277), .B2(n7537), .A(n6723), .ZN(n7536) );
  INV_X1 U7915 ( .A(n9276), .ZN(n7537) );
  NAND2_X1 U7916 ( .A1(n12162), .A2(n7058), .ZN(n7535) );
  AND2_X1 U7917 ( .A1(n9277), .A2(n12161), .ZN(n7058) );
  AOI21_X1 U7918 ( .B1(n7181), .B2(n7180), .A(n6762), .ZN(n7179) );
  INV_X1 U7919 ( .A(n9221), .ZN(n7180) );
  INV_X2 U7920 ( .A(n8030), .ZN(n8259) );
  INV_X1 U7921 ( .A(n13661), .ZN(n13607) );
  NOR2_X1 U7922 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n7674) );
  OR2_X1 U7923 ( .A1(n7830), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7881) );
  INV_X1 U7924 ( .A(n7422), .ZN(n7421) );
  INV_X1 U7925 ( .A(n7429), .ZN(n6922) );
  INV_X1 U7926 ( .A(n13855), .ZN(n6921) );
  NAND2_X1 U7927 ( .A1(n13966), .A2(n11511), .ZN(n7446) );
  NAND2_X1 U7928 ( .A1(n14254), .A2(n10208), .ZN(n7445) );
  AOI21_X1 U7929 ( .B1(n12404), .B2(n6858), .A(n10211), .ZN(n10614) );
  NAND2_X1 U7930 ( .A1(n10212), .A2(n6664), .ZN(n10209) );
  NOR2_X1 U7931 ( .A1(n14099), .A2(n14279), .ZN(n14079) );
  AND2_X1 U7932 ( .A1(n8951), .A2(n8900), .ZN(n14077) );
  NAND2_X1 U7933 ( .A1(n7367), .A2(n7366), .ZN(n14099) );
  INV_X1 U7934 ( .A(n14285), .ZN(n7366) );
  NAND2_X1 U7935 ( .A1(n14208), .A2(n7306), .ZN(n14191) );
  NOR2_X1 U7936 ( .A1(n14194), .A2(n7307), .ZN(n7306) );
  INV_X1 U7937 ( .A(n8835), .ZN(n7307) );
  INV_X1 U7938 ( .A(n8973), .ZN(n15125) );
  NAND2_X1 U7939 ( .A1(n11079), .A2(n8954), .ZN(n15185) );
  AOI21_X1 U7940 ( .B1(n10398), .B2(n10404), .A(n10402), .ZN(n11064) );
  AND2_X1 U7941 ( .A1(n10207), .A2(n10403), .ZN(n11067) );
  NAND2_X1 U7942 ( .A1(n8813), .A2(n7449), .ZN(n8536) );
  AND3_X1 U7943 ( .A1(n8968), .A2(n8812), .A3(n8534), .ZN(n7449) );
  AND2_X1 U7944 ( .A1(n9373), .A2(n9372), .ZN(n9347) );
  AND2_X1 U7945 ( .A1(n15506), .A2(n11004), .ZN(n7252) );
  INV_X1 U7946 ( .A(n7092), .ZN(n13497) );
  AND2_X1 U7947 ( .A1(n10371), .A2(n10370), .ZN(n15277) );
  NAND2_X1 U7948 ( .A1(n9017), .A2(n7643), .ZN(n9021) );
  INV_X1 U7949 ( .A(n9028), .ZN(n7320) );
  OR2_X1 U7950 ( .A1(n7323), .A2(n9038), .ZN(n7322) );
  INV_X1 U7951 ( .A(n9037), .ZN(n7323) );
  INV_X1 U7952 ( .A(n7921), .ZN(n6908) );
  AOI21_X1 U7953 ( .B1(n6909), .B2(n6907), .A(n6709), .ZN(n6906) );
  NOR2_X1 U7954 ( .A1(n8094), .A2(n8093), .ZN(n7636) );
  AND2_X1 U7955 ( .A1(n8022), .A2(n6785), .ZN(n6901) );
  NAND2_X1 U7956 ( .A1(n7628), .A2(n7625), .ZN(n8144) );
  AND2_X1 U7957 ( .A1(n7627), .A2(n7626), .ZN(n7625) );
  NAND2_X1 U7958 ( .A1(n7634), .A2(n7637), .ZN(n7626) );
  NOR2_X1 U7959 ( .A1(n7292), .A2(n7290), .ZN(n7289) );
  INV_X1 U7960 ( .A(n7292), .ZN(n7288) );
  INV_X1 U7961 ( .A(n6888), .ZN(n6887) );
  OAI21_X1 U7962 ( .B1(n6889), .B2(n6702), .A(n6890), .ZN(n6888) );
  NAND2_X1 U7963 ( .A1(n7064), .A2(n9137), .ZN(n7063) );
  OR2_X1 U7964 ( .A1(n9133), .A2(n9134), .ZN(n9135) );
  NAND2_X1 U7965 ( .A1(n9136), .A2(n7294), .ZN(n7293) );
  INV_X1 U7966 ( .A(n9137), .ZN(n7294) );
  INV_X1 U7967 ( .A(n8146), .ZN(n7083) );
  NOR2_X1 U7968 ( .A1(n8188), .A2(n7086), .ZN(n7085) );
  INV_X1 U7969 ( .A(n8148), .ZN(n7086) );
  OR2_X1 U7970 ( .A1(n8187), .A2(n8186), .ZN(n8188) );
  NAND2_X1 U7971 ( .A1(n8238), .A2(n8237), .ZN(n8255) );
  NAND2_X1 U7972 ( .A1(n7081), .A2(n7080), .ZN(n8238) );
  INV_X1 U7973 ( .A(n15014), .ZN(n7383) );
  XNOR2_X1 U7974 ( .A(n12466), .B(n11242), .ZN(n11233) );
  AND2_X1 U7975 ( .A1(n12526), .A2(n12438), .ZN(n7251) );
  INV_X1 U7976 ( .A(n12178), .ZN(n7222) );
  NAND2_X1 U7977 ( .A1(n7154), .A2(n7153), .ZN(n7152) );
  NOR2_X1 U7978 ( .A1(n12646), .A2(n12974), .ZN(n7153) );
  NAND2_X1 U7979 ( .A1(n15401), .A2(n7032), .ZN(n11276) );
  OR2_X1 U7980 ( .A1(n11297), .A2(n11295), .ZN(n7032) );
  NAND2_X1 U7981 ( .A1(n7026), .A2(n6819), .ZN(n11269) );
  NAND2_X1 U7982 ( .A1(n7022), .A2(n6812), .ZN(n11464) );
  INV_X1 U7983 ( .A(n11463), .ZN(n7022) );
  OR2_X1 U7984 ( .A1(n11952), .A2(n11951), .ZN(n11953) );
  INV_X1 U7985 ( .A(n9953), .ZN(n12960) );
  OR2_X1 U7986 ( .A1(n12470), .A2(n12986), .ZN(n12786) );
  OR2_X1 U7987 ( .A1(n12467), .A2(n9927), .ZN(n12782) );
  INV_X1 U7988 ( .A(n12771), .ZN(n7476) );
  OAI21_X1 U7989 ( .B1(n7330), .B2(n7329), .A(n9898), .ZN(n7328) );
  NAND2_X1 U7990 ( .A1(n13255), .A2(n12554), .ZN(n7332) );
  NAND2_X1 U7991 ( .A1(n9992), .A2(n12756), .ZN(n13027) );
  AND2_X1 U7992 ( .A1(n13027), .A2(n13026), .ZN(n13029) );
  NOR2_X1 U7993 ( .A1(n13052), .A2(n7331), .ZN(n7330) );
  INV_X1 U7994 ( .A(n9872), .ZN(n7331) );
  NOR2_X1 U7995 ( .A1(n13128), .A2(n9988), .ZN(n7468) );
  NOR2_X1 U7996 ( .A1(n14846), .A2(n12818), .ZN(n7341) );
  INV_X1 U7997 ( .A(n9751), .ZN(n7343) );
  NOR2_X1 U7998 ( .A1(n7341), .A2(n7340), .ZN(n7339) );
  NOR2_X1 U7999 ( .A1(n12690), .A2(n7352), .ZN(n7351) );
  INV_X1 U8000 ( .A(n9658), .ZN(n7352) );
  NAND2_X1 U8001 ( .A1(n7351), .A2(n6673), .ZN(n7349) );
  NAND2_X1 U8002 ( .A1(n15471), .A2(n15470), .ZN(n7353) );
  NAND2_X1 U8003 ( .A1(n7353), .A2(n7351), .ZN(n11841) );
  INV_X1 U8004 ( .A(n9981), .ZN(n6996) );
  OR2_X1 U8005 ( .A1(n11859), .A2(n11558), .ZN(n12678) );
  INV_X1 U8006 ( .A(n9512), .ZN(n7140) );
  INV_X1 U8007 ( .A(n7139), .ZN(n7138) );
  OAI21_X1 U8008 ( .B1(n9874), .B2(n7140), .A(n9887), .ZN(n7139) );
  INV_X1 U8009 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9846) );
  NOR2_X1 U8010 ( .A1(n9489), .A2(n7148), .ZN(n7147) );
  INV_X1 U8011 ( .A(n9486), .ZN(n7148) );
  NAND2_X1 U8012 ( .A1(n9466), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U8013 ( .A1(n7575), .A2(n10145), .ZN(n7574) );
  INV_X1 U8014 ( .A(n13355), .ZN(n7575) );
  INV_X1 U8015 ( .A(n10139), .ZN(n6989) );
  OR2_X1 U8016 ( .A1(n13395), .A2(n7577), .ZN(n7576) );
  INV_X1 U8017 ( .A(n10145), .ZN(n7577) );
  INV_X1 U8018 ( .A(n13345), .ZN(n7545) );
  AND2_X1 U8019 ( .A1(n7617), .A2(n8341), .ZN(n7616) );
  NAND2_X1 U8020 ( .A1(n7619), .A2(n7618), .ZN(n7617) );
  AOI21_X1 U8021 ( .B1(n6696), .B2(n6897), .A(n6893), .ZN(n6892) );
  INV_X1 U8022 ( .A(n13602), .ZN(n7207) );
  AND2_X1 U8023 ( .A1(n13759), .A2(n13640), .ZN(n7592) );
  INV_X1 U8024 ( .A(n9229), .ZN(n7199) );
  INV_X1 U8025 ( .A(n7200), .ZN(n7196) );
  AND2_X1 U8026 ( .A1(n12154), .A2(n9227), .ZN(n7200) );
  INV_X1 U8027 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U8028 ( .A1(n7057), .A2(n7686), .ZN(n7692) );
  NOR2_X1 U8029 ( .A1(n8125), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8006) );
  NOR2_X1 U8030 ( .A1(n8899), .A2(n7279), .ZN(n7278) );
  INV_X1 U8031 ( .A(n8886), .ZN(n7279) );
  NAND2_X1 U8032 ( .A1(n14109), .A2(n8949), .ZN(n7159) );
  NOR2_X1 U8033 ( .A1(n14142), .A2(n7175), .ZN(n7174) );
  INV_X1 U8034 ( .A(n8944), .ZN(n7175) );
  OR2_X1 U8035 ( .A1(n8936), .A2(n7164), .ZN(n7163) );
  INV_X1 U8036 ( .A(n8934), .ZN(n7164) );
  NAND2_X1 U8037 ( .A1(n14342), .A2(n14222), .ZN(n8937) );
  OR2_X1 U8038 ( .A1(n14342), .A2(n14222), .ZN(n8938) );
  INV_X1 U8039 ( .A(n9089), .ZN(n9183) );
  NOR2_X1 U8040 ( .A1(n12098), .A2(n7166), .ZN(n7165) );
  INV_X1 U8041 ( .A(n9077), .ZN(n7166) );
  INV_X1 U8042 ( .A(n8760), .ZN(n7297) );
  INV_X1 U8043 ( .A(n14815), .ZN(n7371) );
  NOR2_X1 U8044 ( .A1(n9178), .A2(n7261), .ZN(n7260) );
  NOR2_X1 U8045 ( .A1(n11371), .A2(n7262), .ZN(n7261) );
  INV_X1 U8046 ( .A(n8677), .ZN(n7262) );
  NAND2_X1 U8047 ( .A1(n8961), .A2(n8953), .ZN(n10206) );
  INV_X1 U8048 ( .A(n11834), .ZN(n8961) );
  INV_X1 U8049 ( .A(n12259), .ZN(n9143) );
  AOI21_X1 U8050 ( .B1(n14811), .B2(n7266), .A(n6760), .ZN(n7265) );
  INV_X1 U8051 ( .A(n8732), .ZN(n7266) );
  NOR2_X1 U8052 ( .A1(n12227), .A2(n6958), .ZN(n6957) );
  INV_X1 U8053 ( .A(n6959), .ZN(n6958) );
  AND2_X1 U8054 ( .A1(n8812), .A2(n8814), .ZN(n6942) );
  NAND2_X1 U8055 ( .A1(n7087), .A2(n8148), .ZN(n8189) );
  NAND2_X1 U8056 ( .A1(n8050), .A2(n8049), .ZN(n8052) );
  INV_X1 U8057 ( .A(n7903), .ZN(n7070) );
  INV_X1 U8058 ( .A(n7923), .ZN(n7071) );
  NAND2_X1 U8059 ( .A1(n7880), .A2(n7879), .ZN(n7901) );
  INV_X1 U8060 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9337) );
  XNOR2_X1 U8061 ( .A(n9336), .B(n9337), .ZN(n9388) );
  OAI22_X1 U8062 ( .A1(n9394), .A2(n9341), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n9340), .ZN(n9342) );
  AND2_X1 U8063 ( .A1(n9340), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9341) );
  INV_X1 U8064 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U8065 ( .A1(n7378), .A2(n7383), .ZN(n7377) );
  INV_X1 U8066 ( .A(n7380), .ZN(n7378) );
  AOI21_X1 U8067 ( .B1(n7221), .B2(n7218), .A(n7217), .ZN(n7216) );
  INV_X1 U8068 ( .A(n7224), .ZN(n7218) );
  INV_X1 U8069 ( .A(n12180), .ZN(n7217) );
  AND2_X1 U8070 ( .A1(n6727), .A2(n7238), .ZN(n7228) );
  NOR2_X1 U8071 ( .A1(n6725), .A2(n7235), .ZN(n7234) );
  INV_X1 U8072 ( .A(n12490), .ZN(n7235) );
  AND3_X1 U8073 ( .A1(n9750), .A2(n9749), .A3(n9748), .ZN(n12079) );
  NAND2_X1 U8074 ( .A1(n9437), .A2(n9436), .ZN(n9905) );
  NAND2_X1 U8075 ( .A1(n12445), .A2(n12444), .ZN(n12547) );
  NAND2_X1 U8076 ( .A1(n9853), .A2(n9434), .ZN(n9864) );
  AND3_X1 U8077 ( .A1(n9727), .A2(n9726), .A3(n9725), .ZN(n11996) );
  NAND2_X1 U8078 ( .A1(n12518), .A2(n7251), .ZN(n12524) );
  INV_X1 U8079 ( .A(n12141), .ZN(n6839) );
  NAND2_X1 U8080 ( .A1(n9570), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9571) );
  NAND2_X1 U8081 ( .A1(n10967), .A2(n10968), .ZN(n11263) );
  NAND2_X1 U8082 ( .A1(n10955), .A2(n10964), .ZN(n7034) );
  NAND2_X1 U8083 ( .A1(n11263), .A2(n7030), .ZN(n7029) );
  NAND2_X1 U8084 ( .A1(n11264), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7030) );
  NAND2_X1 U8085 ( .A1(n15403), .A2(n15402), .ZN(n15401) );
  AND2_X1 U8086 ( .A1(n7029), .A2(n7028), .ZN(n11265) );
  XNOR2_X1 U8087 ( .A(n11276), .B(n11304), .ZN(n15421) );
  OR2_X1 U8088 ( .A1(n15428), .A2(n15427), .ZN(n7026) );
  NAND2_X1 U8089 ( .A1(n7409), .A2(n11317), .ZN(n7407) );
  INV_X1 U8090 ( .A(n11269), .ZN(n7409) );
  NOR2_X1 U8091 ( .A1(n11657), .A2(n9708), .ZN(n7413) );
  OR2_X1 U8092 ( .A1(n11953), .A2(n12836), .ZN(n7417) );
  INV_X1 U8093 ( .A(n12910), .ZN(n7021) );
  XNOR2_X1 U8094 ( .A(n12909), .B(n7036), .ZN(n14833) );
  NOR2_X1 U8095 ( .A1(n12909), .A2(n7036), .ZN(n7419) );
  OR2_X1 U8096 ( .A1(n14833), .A2(n14834), .ZN(n7019) );
  NAND2_X1 U8097 ( .A1(n12605), .A2(n7652), .ZN(n12618) );
  NAND2_X1 U8098 ( .A1(n12603), .A2(n12602), .ZN(n12605) );
  INV_X1 U8099 ( .A(n12974), .ZN(n6871) );
  NAND2_X1 U8100 ( .A1(n9931), .A2(n9930), .ZN(n12277) );
  NOR2_X1 U8101 ( .A1(n12773), .A2(n7480), .ZN(n7479) );
  INV_X1 U8102 ( .A(n12756), .ZN(n7480) );
  NAND2_X1 U8103 ( .A1(n9873), .A2(n7330), .ZN(n7326) );
  NOR2_X1 U8104 ( .A1(n13095), .A2(n7355), .ZN(n7354) );
  INV_X1 U8105 ( .A(n9826), .ZN(n7355) );
  OR2_X1 U8106 ( .A1(n13271), .A2(n13101), .ZN(n12736) );
  NAND2_X1 U8107 ( .A1(n13150), .A2(n13149), .ZN(n13152) );
  AND4_X1 U8108 ( .A1(n9795), .A2(n9794), .A3(n9793), .A4(n9792), .ZN(n13159)
         );
  AND2_X1 U8109 ( .A1(n12718), .A2(n12719), .ZN(n14844) );
  OR2_X1 U8110 ( .A1(n14854), .A2(n12079), .ZN(n12717) );
  NAND2_X1 U8111 ( .A1(n12074), .A2(n12073), .ZN(n12072) );
  NAND2_X1 U8112 ( .A1(n11978), .A2(n6744), .ZN(n14857) );
  AOI21_X1 U8113 ( .B1(n7455), .B2(n7457), .A(n7452), .ZN(n7451) );
  INV_X1 U8114 ( .A(n12694), .ZN(n7452) );
  AND2_X1 U8115 ( .A1(n12694), .A2(n12693), .ZN(n12690) );
  NAND2_X1 U8116 ( .A1(n11854), .A2(n12671), .ZN(n11856) );
  INV_X1 U8117 ( .A(n15509), .ZN(n14851) );
  OR2_X1 U8118 ( .A1(n9742), .A2(n10322), .ZN(n9556) );
  NAND2_X1 U8119 ( .A1(n10000), .A2(n10036), .ZN(n15495) );
  NAND2_X1 U8120 ( .A1(n10995), .A2(n12780), .ZN(n15507) );
  INV_X1 U8121 ( .A(n15490), .ZN(n15511) );
  NAND2_X1 U8122 ( .A1(n9534), .A2(n9533), .ZN(n9914) );
  INV_X1 U8123 ( .A(n15507), .ZN(n14853) );
  OAI21_X1 U8124 ( .B1(P1_DATAO_REG_25__SCAN_IN), .B2(n14396), .A(n9520), .ZN(
        n9917) );
  NAND2_X1 U8125 ( .A1(n9518), .A2(n7157), .ZN(n7156) );
  AND2_X1 U8126 ( .A1(n7215), .A2(n10029), .ZN(n7214) );
  XNOR2_X1 U8127 ( .A(n9509), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n9861) );
  AND2_X1 U8128 ( .A1(n11549), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9505) );
  AND2_X1 U8129 ( .A1(n9746), .A2(n6778), .ZN(n9847) );
  NOR2_X1 U8130 ( .A1(n9738), .A2(n7145), .ZN(n7144) );
  INV_X1 U8131 ( .A(n9488), .ZN(n7145) );
  NAND2_X1 U8132 ( .A1(n9487), .A2(n7147), .ZN(n7146) );
  XNOR2_X1 U8133 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9667) );
  XNOR2_X1 U8134 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9592) );
  NAND2_X1 U8135 ( .A1(n9468), .A2(n9467), .ZN(n9555) );
  OR2_X1 U8136 ( .A1(n13640), .A2(n10146), .ZN(n7566) );
  NAND2_X1 U8137 ( .A1(n10362), .A2(n10286), .ZN(n7760) );
  AND2_X1 U8138 ( .A1(n6750), .A2(n10170), .ZN(n6974) );
  NAND2_X1 U8139 ( .A1(n11259), .A2(n7569), .ZN(n11784) );
  AND2_X1 U8140 ( .A1(n10108), .A2(n10103), .ZN(n7569) );
  AND2_X1 U8141 ( .A1(n10089), .A2(n10084), .ZN(n7570) );
  OR2_X1 U8142 ( .A1(n7836), .A2(n10372), .ZN(n7746) );
  NOR2_X1 U8143 ( .A1(n15248), .A2(n6734), .ZN(n10407) );
  OR2_X1 U8144 ( .A1(n10407), .A2(n10406), .ZN(n7100) );
  OR2_X1 U8145 ( .A1(n10870), .A2(n10871), .ZN(n7098) );
  AND2_X1 U8146 ( .A1(n7098), .A2(n7097), .ZN(n11221) );
  NAND2_X1 U8147 ( .A1(n11219), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7097) );
  OR2_X1 U8148 ( .A1(n11221), .A2(n11220), .ZN(n7096) );
  NAND2_X1 U8149 ( .A1(n9162), .A2(n8424), .ZN(n8384) );
  NAND2_X1 U8150 ( .A1(n13515), .A2(n13726), .ZN(n13514) );
  INV_X1 U8151 ( .A(n9236), .ZN(n13594) );
  OR2_X1 U8152 ( .A1(n13580), .A2(n7592), .ZN(n7208) );
  NOR2_X1 U8153 ( .A1(n13625), .A2(n7592), .ZN(n13603) );
  NOR2_X1 U8154 ( .A1(n13603), .A2(n13602), .ZN(n13601) );
  INV_X1 U8155 ( .A(n13584), .ZN(n13629) );
  INV_X1 U8156 ( .A(n7044), .ZN(n13624) );
  NAND2_X1 U8157 ( .A1(n7538), .A2(n7046), .ZN(n7045) );
  INV_X1 U8158 ( .A(n7539), .ZN(n7538) );
  NAND2_X1 U8159 ( .A1(n13673), .A2(n7191), .ZN(n7189) );
  AOI21_X1 U8160 ( .B1(n7191), .B2(n13674), .A(n6707), .ZN(n7190) );
  NAND2_X1 U8161 ( .A1(n7047), .A2(n7050), .ZN(n9285) );
  NAND2_X1 U8162 ( .A1(n7048), .A2(n9283), .ZN(n7047) );
  OR2_X1 U8163 ( .A1(n13673), .A2(n13674), .ZN(n7192) );
  NOR2_X1 U8164 ( .A1(n13719), .A2(n7534), .ZN(n7533) );
  INV_X1 U8165 ( .A(n7536), .ZN(n7534) );
  INV_X1 U8166 ( .A(n9278), .ZN(n13719) );
  NAND2_X1 U8167 ( .A1(n12166), .A2(n7200), .ZN(n12153) );
  OAI21_X1 U8168 ( .B1(n12113), .B2(n9272), .A(n9273), .ZN(n12165) );
  NAND2_X1 U8169 ( .A1(n7043), .A2(n7530), .ZN(n11636) );
  AOI21_X1 U8170 ( .B1(n7528), .B2(n9264), .A(n7527), .ZN(n7530) );
  NOR2_X1 U8171 ( .A1(n7531), .A2(n7042), .ZN(n7041) );
  NAND2_X1 U8172 ( .A1(n11352), .A2(n11355), .ZN(n9263) );
  NAND2_X1 U8173 ( .A1(n9263), .A2(n7532), .ZN(n11418) );
  INV_X1 U8174 ( .A(n7528), .ZN(n7532) );
  NAND2_X1 U8175 ( .A1(n7861), .A2(n7860), .ZN(n11442) );
  NAND2_X1 U8176 ( .A1(n7526), .A2(n9256), .ZN(n10835) );
  NAND2_X1 U8177 ( .A1(n10360), .A2(n8518), .ZN(n13661) );
  NAND2_X1 U8178 ( .A1(n10062), .A2(n15316), .ZN(n7177) );
  AND2_X1 U8179 ( .A1(n10360), .A2(n8517), .ZN(n13604) );
  AOI21_X1 U8180 ( .B1(n15356), .B2(n13521), .A(n13527), .ZN(n9300) );
  INV_X1 U8181 ( .A(n15342), .ZN(n15356) );
  NOR2_X1 U8182 ( .A1(n7667), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7496) );
  NAND2_X1 U8183 ( .A1(n7057), .A2(n6911), .ZN(n8508) );
  INV_X1 U8184 ( .A(n7675), .ZN(n6911) );
  AND2_X1 U8185 ( .A1(n7057), .A2(n8505), .ZN(n8510) );
  INV_X1 U8186 ( .A(n8496), .ZN(n8498) );
  OR2_X1 U8187 ( .A1(n8008), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8033) );
  OR2_X1 U8188 ( .A1(n8689), .A2(n8688), .ZN(n8698) );
  AND2_X1 U8189 ( .A1(n6729), .A2(n13896), .ZN(n6940) );
  AOI21_X1 U8190 ( .B1(n6920), .B2(n6923), .A(n6756), .ZN(n6918) );
  INV_X1 U8191 ( .A(n7427), .ZN(n6923) );
  NAND2_X1 U8192 ( .A1(n12228), .A2(n7442), .ZN(n7441) );
  INV_X1 U8193 ( .A(n7649), .ZN(n7442) );
  OR2_X1 U8194 ( .A1(n12207), .A2(n12206), .ZN(n7648) );
  NOR2_X1 U8195 ( .A1(n7441), .A2(n6935), .ZN(n6934) );
  INV_X1 U8196 ( .A(n14930), .ZN(n6935) );
  AND2_X1 U8197 ( .A1(n12359), .A2(n12357), .ZN(n7444) );
  AOI21_X1 U8198 ( .B1(n13904), .B2(n7423), .A(n6777), .ZN(n7422) );
  INV_X1 U8199 ( .A(n12334), .ZN(n7423) );
  NAND2_X1 U8200 ( .A1(n13895), .A2(n13896), .ZN(n13894) );
  INV_X1 U8201 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10645) );
  NAND2_X1 U8202 ( .A1(n14079), .A2(n12259), .ZN(n14060) );
  AOI21_X1 U8203 ( .B1(n7273), .B2(n14090), .A(n6768), .ZN(n7272) );
  NAND2_X1 U8204 ( .A1(n14120), .A2(n7278), .ZN(n7277) );
  NAND2_X1 U8205 ( .A1(n7276), .A2(n7280), .ZN(n7275) );
  AOI21_X1 U8206 ( .B1(n7284), .B2(n6695), .A(n6758), .ZN(n7283) );
  AND2_X1 U8207 ( .A1(n14209), .A2(n8823), .ZN(n7308) );
  OR2_X1 U8208 ( .A1(n14354), .A2(n14908), .ZN(n9077) );
  NAND2_X1 U8209 ( .A1(n8933), .A2(n7165), .ZN(n12101) );
  OR2_X1 U8210 ( .A1(n8698), .A2(n10645), .ZN(n8725) );
  NAND2_X1 U8211 ( .A1(n9143), .A2(n14980), .ZN(n7360) );
  NAND2_X1 U8212 ( .A1(n8740), .A2(n8739), .ZN(n14981) );
  OR2_X1 U8213 ( .A1(n8848), .A2(n10594), .ZN(n8582) );
  AND2_X1 U8214 ( .A1(n8972), .A2(n8977), .ZN(n10398) );
  XNOR2_X1 U8215 ( .A(n8410), .B(n8409), .ZN(n12292) );
  INV_X1 U8216 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8535) );
  XNOR2_X1 U8217 ( .A(n8365), .B(SI_27_), .ZN(n12269) );
  MUX2_X1 U8218 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8903), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8904) );
  XNOR2_X1 U8219 ( .A(n9388), .B(n7385), .ZN(n9390) );
  INV_X1 U8220 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7385) );
  AOI22_X1 U8221 ( .A1(n15048), .A2(P3_ADDR_REG_12__SCAN_IN), .B1(n9352), .B2(
        n9415), .ZN(n9370) );
  OR2_X1 U8222 ( .A1(n15010), .A2(n7384), .ZN(n7380) );
  NAND2_X1 U8223 ( .A1(n15010), .A2(n7384), .ZN(n7381) );
  INV_X1 U8224 ( .A(n13101), .ZN(n13130) );
  AND4_X1 U8225 ( .A1(n9838), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(n13118)
         );
  AND3_X1 U8226 ( .A1(n9544), .A2(n9543), .A3(n9542), .ZN(n13043) );
  AND2_X1 U8227 ( .A1(n9540), .A2(n9539), .ZN(n13013) );
  NAND2_X1 U8228 ( .A1(n10928), .A2(n10927), .ZN(n12578) );
  NAND2_X1 U8229 ( .A1(n10934), .A2(n10933), .ZN(n12572) );
  XNOR2_X1 U8230 ( .A(n7000), .B(n12942), .ZN(n6999) );
  NOR2_X1 U8231 ( .A1(n12619), .A2(n12796), .ZN(n7001) );
  NAND2_X1 U8232 ( .A1(n6781), .A2(n6998), .ZN(n6997) );
  INV_X1 U8233 ( .A(n12805), .ZN(n6998) );
  INV_X1 U8234 ( .A(n13042), .ZN(n13070) );
  AND2_X1 U8235 ( .A1(n10819), .A2(n10818), .ZN(n14832) );
  AND3_X1 U8236 ( .A1(n7407), .A2(n11268), .A3(P3_REG2_REG_9__SCAN_IN), .ZN(
        n15446) );
  AOI21_X1 U8237 ( .B1(n14826), .B2(P3_REG1_REG_17__SCAN_IN), .A(n6726), .ZN(
        n12946) );
  INV_X1 U8238 ( .A(n12618), .ZN(n14867) );
  NOR2_X1 U8239 ( .A1(n9975), .A2(n9974), .ZN(n9976) );
  NOR2_X1 U8240 ( .A1(n12473), .A2(n15509), .ZN(n9975) );
  NAND2_X1 U8241 ( .A1(n9952), .A2(n9951), .ZN(n12968) );
  NOR2_X1 U8242 ( .A1(n13079), .A2(n7473), .ZN(n7472) );
  INV_X1 U8243 ( .A(n12758), .ZN(n7473) );
  OR2_X1 U8244 ( .A1(n9742), .A2(n10288), .ZN(n9580) );
  NAND2_X1 U8245 ( .A1(n10016), .A2(n10015), .ZN(n10792) );
  XNOR2_X1 U8246 ( .A(n9961), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12810) );
  NAND2_X1 U8247 ( .A1(n9962), .A2(n9446), .ZN(n9960) );
  NAND2_X1 U8248 ( .A1(n7952), .A2(n7951), .ZN(n11803) );
  NOR2_X1 U8249 ( .A1(n6708), .A2(n13417), .ZN(n7553) );
  NAND2_X1 U8250 ( .A1(n7556), .A2(n7561), .ZN(n7555) );
  NAND2_X1 U8251 ( .A1(n7562), .A2(n13318), .ZN(n7561) );
  INV_X1 U8252 ( .A(n10183), .ZN(n7562) );
  AOI21_X1 U8253 ( .B1(n7563), .B2(n6968), .A(n6965), .ZN(n6963) );
  NOR2_X1 U8254 ( .A1(n6970), .A2(n10175), .ZN(n6967) );
  NAND2_X1 U8255 ( .A1(n8106), .A2(n8105), .ZN(n13798) );
  INV_X1 U8256 ( .A(n13450), .ZN(n10838) );
  NAND2_X1 U8257 ( .A1(n10080), .A2(n10701), .ZN(n10706) );
  NAND2_X1 U8258 ( .A1(n8240), .A2(n8239), .ZN(n13765) );
  NAND2_X1 U8259 ( .A1(n10486), .A2(n10066), .ZN(n7548) );
  NAND2_X1 U8260 ( .A1(n10190), .A2(n13683), .ZN(n13425) );
  OR2_X1 U8261 ( .A1(n6672), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7785) );
  AND3_X1 U8262 ( .A1(n7783), .A2(n7782), .A3(n7781), .ZN(n7784) );
  OAI21_X1 U8263 ( .B1(n13502), .B2(n15271), .A(n7091), .ZN(n7090) );
  AOI21_X1 U8264 ( .B1(n13501), .B2(n15277), .A(n15281), .ZN(n7091) );
  NAND2_X1 U8265 ( .A1(n9292), .A2(n6716), .ZN(n13736) );
  NAND2_X1 U8266 ( .A1(n9292), .A2(n9291), .ZN(n13561) );
  NAND2_X1 U8267 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  XNOR2_X1 U8268 ( .A(n13550), .B(n13549), .ZN(n7211) );
  NAND2_X1 U8269 ( .A1(n8196), .A2(n8195), .ZN(n13777) );
  INV_X1 U8270 ( .A(n13519), .ZN(n15297) );
  INV_X1 U8271 ( .A(n15293), .ZN(n13652) );
  NAND2_X1 U8272 ( .A1(n7833), .A2(n7832), .ZN(n10848) );
  OR2_X1 U8273 ( .A1(n15311), .A2(n10194), .ZN(n13683) );
  INV_X1 U8274 ( .A(n9294), .ZN(n9240) );
  NOR2_X1 U8275 ( .A1(n15371), .A2(n13676), .ZN(n7587) );
  INV_X1 U8276 ( .A(n9300), .ZN(n7585) );
  OR2_X1 U8277 ( .A1(n7591), .A2(n15371), .ZN(n7583) );
  INV_X1 U8278 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7590) );
  NOR2_X1 U8279 ( .A1(n15371), .A2(n15360), .ZN(n7581) );
  NAND2_X1 U8280 ( .A1(n9322), .A2(n9321), .ZN(n15310) );
  AND2_X1 U8281 ( .A1(n8978), .A2(n8977), .ZN(n8979) );
  INV_X1 U8282 ( .A(n8976), .ZN(n8980) );
  INV_X1 U8283 ( .A(n13958), .ZN(n14911) );
  INV_X1 U8284 ( .A(n7437), .ZN(n12031) );
  INV_X1 U8285 ( .A(n7435), .ZN(n7434) );
  AOI21_X1 U8286 ( .B1(n7435), .B2(n7433), .A(n6780), .ZN(n7432) );
  INV_X1 U8287 ( .A(n13966), .ZN(n14261) );
  NOR2_X1 U8288 ( .A1(n11338), .A2(n11339), .ZN(n11921) );
  NAND2_X1 U8289 ( .A1(n14060), .A2(n6953), .ZN(n12252) );
  OR2_X1 U8290 ( .A1(n14079), .A2(n12259), .ZN(n6953) );
  XNOR2_X1 U8291 ( .A(n7362), .B(n7361), .ZN(n12262) );
  AND2_X1 U8292 ( .A1(n14279), .A2(n14095), .ZN(n7363) );
  OR3_X1 U8293 ( .A1(n14079), .A2(n14078), .A3(n15125), .ZN(n14281) );
  INV_X1 U8294 ( .A(n14074), .ZN(n6870) );
  NAND2_X1 U8295 ( .A1(n7285), .A2(n7284), .ZN(n14135) );
  AND2_X1 U8296 ( .A1(n7285), .A2(n6730), .ZN(n14136) );
  OR2_X1 U8297 ( .A1(n14152), .A2(n6695), .ZN(n7285) );
  NAND2_X1 U8298 ( .A1(n8811), .A2(n9154), .ZN(n8817) );
  AND2_X1 U8299 ( .A1(n10479), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10403) );
  NAND2_X1 U8300 ( .A1(n7387), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7386) );
  OAI21_X1 U8301 ( .B1(n14765), .B2(n14766), .A(n7396), .ZN(n7395) );
  INV_X1 U8302 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7396) );
  OAI21_X1 U8303 ( .B1(n9013), .B2(n9012), .A(n7644), .ZN(n9017) );
  AND2_X1 U8304 ( .A1(n7695), .A2(n9296), .ZN(n7715) );
  NAND2_X1 U8305 ( .A1(n7320), .A2(n9027), .ZN(n7319) );
  AND2_X1 U8306 ( .A1(n6874), .A2(n7846), .ZN(n6875) );
  NAND2_X1 U8307 ( .A1(n9046), .A2(n7311), .ZN(n7310) );
  NAND2_X1 U8308 ( .A1(n6905), .A2(n6906), .ZN(n7938) );
  NAND2_X1 U8309 ( .A1(n9056), .A2(n9058), .ZN(n7315) );
  NAND2_X1 U8310 ( .A1(n9104), .A2(n9105), .ZN(n7287) );
  AND2_X1 U8311 ( .A1(n8115), .A2(n7635), .ZN(n7634) );
  NAND2_X1 U8312 ( .A1(n7630), .A2(n8116), .ZN(n7637) );
  INV_X1 U8313 ( .A(n7638), .ZN(n7630) );
  NAND2_X1 U8314 ( .A1(n7624), .A2(n6741), .ZN(n7623) );
  NOR2_X1 U8315 ( .A1(n6759), .A2(n6901), .ZN(n6900) );
  AND2_X1 U8316 ( .A1(n7629), .A2(n6878), .ZN(n6877) );
  NOR2_X1 U8317 ( .A1(n6880), .A2(n8068), .ZN(n6878) );
  INV_X1 U8318 ( .A(n8067), .ZN(n6880) );
  AND2_X1 U8319 ( .A1(n7629), .A2(n6784), .ZN(n6879) );
  NAND2_X1 U8320 ( .A1(n7632), .A2(n7638), .ZN(n7627) );
  INV_X1 U8321 ( .A(n9109), .ZN(n7290) );
  NAND2_X1 U8322 ( .A1(n9111), .A2(n9113), .ZN(n7313) );
  OAI211_X1 U8323 ( .C1(n9108), .C2(n9109), .A(n9110), .B(n6769), .ZN(n7312)
         );
  NOR2_X1 U8324 ( .A1(n8207), .A2(n6742), .ZN(n7612) );
  INV_X1 U8325 ( .A(n8226), .ZN(n7610) );
  INV_X1 U8326 ( .A(n8224), .ZN(n7609) );
  INV_X1 U8327 ( .A(n7612), .ZN(n6882) );
  NAND2_X1 U8328 ( .A1(n6887), .A2(n6889), .ZN(n6883) );
  NAND2_X1 U8329 ( .A1(n8207), .A2(n6742), .ZN(n7611) );
  NOR2_X1 U8330 ( .A1(n6886), .A2(n8185), .ZN(n6885) );
  NAND2_X1 U8331 ( .A1(n9129), .A2(n7317), .ZN(n7316) );
  AND2_X1 U8332 ( .A1(n12458), .A2(n12511), .ZN(n12771) );
  INV_X1 U8333 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7014) );
  NAND2_X1 U8334 ( .A1(n6895), .A2(n6896), .ZN(n8319) );
  NAND2_X1 U8335 ( .A1(n6770), .A2(n8318), .ZN(n7618) );
  INV_X1 U8336 ( .A(n6896), .ZN(n6894) );
  INV_X1 U8337 ( .A(n7618), .ZN(n6893) );
  NAND2_X1 U8338 ( .A1(n13511), .A2(n6690), .ZN(n8391) );
  INV_X1 U8339 ( .A(n9238), .ZN(n7604) );
  NAND2_X1 U8340 ( .A1(n9138), .A2(n9141), .ZN(n7065) );
  NOR2_X1 U8341 ( .A1(n9141), .A2(n9138), .ZN(n7066) );
  OAI21_X1 U8342 ( .B1(n6721), .B2(n6859), .A(n7293), .ZN(n9139) );
  AND2_X1 U8343 ( .A1(n14349), .A2(n13943), .ZN(n9089) );
  NOR2_X1 U8344 ( .A1(n7267), .A2(n11751), .ZN(n7264) );
  INV_X1 U8345 ( .A(n8321), .ZN(n7507) );
  NOR2_X1 U8346 ( .A1(n8321), .A2(n8300), .ZN(n7506) );
  NAND2_X1 U8347 ( .A1(n7085), .A2(n7083), .ZN(n7082) );
  INV_X1 U8348 ( .A(n7085), .ZN(n7084) );
  INV_X1 U8349 ( .A(n8095), .ZN(n7073) );
  NAND2_X1 U8350 ( .A1(n8099), .A2(n10494), .ZN(n8119) );
  NAND2_X1 U8351 ( .A1(n8072), .A2(n10474), .ZN(n8097) );
  INV_X1 U8352 ( .A(n8025), .ZN(n7077) );
  OR2_X1 U8353 ( .A1(n6701), .A2(n8070), .ZN(n7512) );
  NAND4_X1 U8354 ( .A1(n13507), .A2(n7524), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n7523), .ZN(n7522) );
  INV_X1 U8355 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7524) );
  INV_X1 U8356 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7523) );
  NAND4_X1 U8357 ( .A1(n7521), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(n7520), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7519) );
  INV_X1 U8358 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7521) );
  INV_X1 U8359 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9335) );
  INV_X1 U8360 ( .A(n12441), .ZN(n7250) );
  NAND2_X1 U8361 ( .A1(n12499), .A2(n12500), .ZN(n12451) );
  NAND2_X1 U8362 ( .A1(n15439), .A2(n7031), .ZN(n11278) );
  OR2_X1 U8363 ( .A1(n11311), .A2(n11309), .ZN(n7031) );
  OR2_X1 U8364 ( .A1(n9947), .A2(n12473), .ZN(n12787) );
  INV_X1 U8365 ( .A(n12782), .ZN(n7006) );
  AND2_X1 U8366 ( .A1(n7007), .A2(n12781), .ZN(n7004) );
  OR2_X1 U8367 ( .A1(n13258), .A2(n13042), .ZN(n12749) );
  NAND2_X1 U8368 ( .A1(n9873), .A2(n9872), .ZN(n13053) );
  INV_X1 U8369 ( .A(n12717), .ZN(n7463) );
  INV_X1 U8370 ( .A(n7456), .ZN(n7455) );
  OAI21_X1 U8371 ( .B1(n6673), .B2(n7457), .A(n12690), .ZN(n7456) );
  INV_X1 U8372 ( .A(n12688), .ZN(n7457) );
  NAND2_X1 U8373 ( .A1(n14597), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7127) );
  NOR2_X1 U8374 ( .A1(n9949), .A2(n7124), .ZN(n7123) );
  INV_X1 U8375 ( .A(n9523), .ZN(n7124) );
  NAND2_X1 U8376 ( .A1(n7128), .A2(n7127), .ZN(n7126) );
  NAND2_X1 U8377 ( .A1(n7122), .A2(n6825), .ZN(n7121) );
  INV_X1 U8378 ( .A(n9949), .ZN(n7122) );
  NAND2_X1 U8379 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n7129), .ZN(n7128) );
  INV_X1 U8380 ( .A(n7142), .ZN(n7141) );
  OAI21_X1 U8381 ( .B1(n7147), .B2(n7143), .A(n9491), .ZN(n7142) );
  INV_X1 U8382 ( .A(n7144), .ZN(n7143) );
  INV_X1 U8383 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U8384 ( .A1(n9650), .A2(n9651), .ZN(n9669) );
  INV_X1 U8385 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9444) );
  INV_X1 U8386 ( .A(n11723), .ZN(n7550) );
  NAND2_X1 U8387 ( .A1(n13312), .A2(n10183), .ZN(n7560) );
  INV_X1 U8388 ( .A(n8288), .ZN(n8289) );
  OR2_X1 U8389 ( .A1(n7490), .A2(n13752), .ZN(n7488) );
  NAND2_X1 U8390 ( .A1(n7492), .A2(n7491), .ZN(n7490) );
  OAI21_X1 U8391 ( .B1(n6719), .B2(n7540), .A(n13626), .ZN(n7539) );
  NAND2_X1 U8392 ( .A1(n6703), .A2(n7052), .ZN(n7046) );
  AND2_X1 U8393 ( .A1(n8133), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8153) );
  INV_X1 U8394 ( .A(n9222), .ZN(n7183) );
  NAND2_X1 U8395 ( .A1(n6868), .A2(n6867), .ZN(n11810) );
  OR2_X1 U8396 ( .A1(n11421), .A2(n7529), .ZN(n7528) );
  INV_X1 U8397 ( .A(n9262), .ZN(n7529) );
  NOR2_X1 U8398 ( .A1(n9212), .A2(n7598), .ZN(n7597) );
  INV_X1 U8399 ( .A(n9211), .ZN(n7598) );
  INV_X1 U8400 ( .A(n10268), .ZN(n7039) );
  INV_X1 U8401 ( .A(n10276), .ZN(n7040) );
  NOR2_X2 U8402 ( .A1(n13696), .A2(n13777), .ZN(n13680) );
  INV_X1 U8403 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7666) );
  INV_X1 U8404 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7665) );
  NOR2_X1 U8405 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n7670) );
  NOR2_X1 U8406 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7668) );
  INV_X1 U8407 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8499) );
  INV_X1 U8408 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7687) );
  INV_X1 U8409 ( .A(n7497), .ZN(n7906) );
  AOI21_X1 U8410 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14027), .A(n14026), .ZN(
        n14036) );
  NOR2_X1 U8411 ( .A1(n7274), .A2(n7271), .ZN(n7270) );
  INV_X1 U8412 ( .A(n7278), .ZN(n7271) );
  INV_X1 U8413 ( .A(n7275), .ZN(n7273) );
  NOR2_X1 U8414 ( .A1(n6691), .A2(n14313), .ZN(n7368) );
  NAND2_X1 U8415 ( .A1(n6951), .A2(n6950), .ZN(n6949) );
  INV_X1 U8416 ( .A(n6952), .ZN(n6951) );
  NAND2_X1 U8417 ( .A1(n14335), .A2(n14212), .ZN(n6952) );
  NAND2_X1 U8418 ( .A1(n7365), .A2(n6959), .ZN(n6960) );
  INV_X1 U8419 ( .A(n7368), .ZN(n14163) );
  NAND2_X1 U8420 ( .A1(n7365), .A2(n7364), .ZN(n15075) );
  AND2_X1 U8421 ( .A1(n6946), .A2(n15135), .ZN(n6944) );
  AND2_X1 U8422 ( .A1(n6946), .A2(n6945), .ZN(n11171) );
  AND2_X1 U8423 ( .A1(n14258), .A2(n15135), .ZN(n6945) );
  NAND2_X1 U8424 ( .A1(n14258), .A2(n15135), .ZN(n11185) );
  AND2_X1 U8425 ( .A1(n15124), .A2(n14256), .ZN(n14258) );
  AND2_X1 U8426 ( .A1(n8376), .A2(n8375), .ZN(n8409) );
  XNOR2_X1 U8427 ( .A(n8255), .B(SI_22_), .ZN(n8258) );
  AND2_X1 U8428 ( .A1(n8148), .A2(n8123), .ZN(n8146) );
  AND2_X1 U8429 ( .A1(n7510), .A2(n7076), .ZN(n7075) );
  AND2_X1 U8430 ( .A1(n7512), .A2(n7511), .ZN(n7510) );
  NAND2_X1 U8431 ( .A1(n7078), .A2(n7077), .ZN(n7076) );
  OR2_X1 U8432 ( .A1(n8051), .A2(SI_14_), .ZN(n7511) );
  NAND2_X1 U8433 ( .A1(n8052), .A2(n8051), .ZN(n7509) );
  AND2_X1 U8434 ( .A1(n8051), .A2(n8029), .ZN(n8049) );
  NAND2_X1 U8435 ( .A1(n8026), .A2(n8025), .ZN(n8050) );
  OR2_X1 U8436 ( .A1(n8627), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8638) );
  INV_X1 U8437 ( .A(n7775), .ZN(n7501) );
  INV_X1 U8438 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9330) );
  XNOR2_X1 U8439 ( .A(n9334), .B(n9335), .ZN(n9374) );
  NOR2_X1 U8440 ( .A1(n9344), .A2(n9343), .ZN(n9401) );
  AND2_X1 U8441 ( .A1(n9397), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n9343) );
  AOI21_X1 U8442 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n9346), .A(n9345), .ZN(
        n9372) );
  NOR2_X1 U8443 ( .A1(n9401), .A2(n9402), .ZN(n9345) );
  INV_X1 U8444 ( .A(n12507), .ZN(n7236) );
  NAND2_X1 U8445 ( .A1(n12468), .A2(n9927), .ZN(n7239) );
  OR2_X1 U8446 ( .A1(n12570), .A2(n7240), .ZN(n7237) );
  OR2_X1 U8447 ( .A1(n9939), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U8448 ( .A1(n15504), .A2(n12657), .ZN(n7450) );
  NAND2_X1 U8449 ( .A1(n7253), .A2(n7255), .ZN(n7254) );
  INV_X1 U8450 ( .A(n12650), .ZN(n7255) );
  AND2_X1 U8451 ( .A1(n11453), .A2(n11235), .ZN(n11236) );
  NAND2_X1 U8452 ( .A1(n7225), .A2(n14854), .ZN(n7224) );
  INV_X1 U8453 ( .A(n12139), .ZN(n7225) );
  AND2_X1 U8454 ( .A1(n11994), .A2(n11997), .ZN(n7245) );
  OR2_X1 U8455 ( .A1(n11994), .A2(n11997), .ZN(n7244) );
  XNOR2_X1 U8456 ( .A(n11046), .B(n11040), .ZN(n11045) );
  NAND2_X1 U8457 ( .A1(n9439), .A2(n9438), .ZN(n9920) );
  OR2_X1 U8458 ( .A1(n9920), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9937) );
  NOR2_X1 U8459 ( .A1(n12800), .A2(n7150), .ZN(n7149) );
  NAND2_X1 U8460 ( .A1(n7151), .A2(n12799), .ZN(n7150) );
  NOR2_X1 U8461 ( .A1(n12647), .A2(n7152), .ZN(n7151) );
  OAI21_X1 U8462 ( .B1(n10828), .B2(n11093), .A(n7645), .ZN(n10901) );
  NAND2_X1 U8463 ( .A1(n7023), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10903) );
  INV_X1 U8464 ( .A(n10901), .ZN(n7023) );
  NAND2_X1 U8465 ( .A1(n10903), .A2(n7645), .ZN(n10820) );
  XNOR2_X1 U8466 ( .A(n10965), .B(n10964), .ZN(n10979) );
  INV_X1 U8467 ( .A(n9566), .ZN(n7212) );
  NAND2_X1 U8468 ( .A1(n15382), .A2(n11275), .ZN(n15403) );
  NAND2_X1 U8469 ( .A1(n15420), .A2(n11277), .ZN(n15441) );
  NAND2_X1 U8470 ( .A1(n15441), .A2(n15440), .ZN(n15439) );
  XNOR2_X1 U8471 ( .A(n11278), .B(n11317), .ZN(n15462) );
  INV_X1 U8472 ( .A(n11272), .ZN(n7408) );
  NAND2_X1 U8473 ( .A1(n12871), .A2(n12898), .ZN(n7402) );
  OR2_X1 U8474 ( .A1(n12872), .A2(n13146), .ZN(n7025) );
  NAND2_X1 U8475 ( .A1(n12911), .A2(n7038), .ZN(n7037) );
  OR2_X1 U8476 ( .A1(n12912), .A2(n13220), .ZN(n7038) );
  NAND2_X1 U8477 ( .A1(n9947), .A2(n6831), .ZN(n6830) );
  INV_X1 U8478 ( .A(n12473), .ZN(n6831) );
  INV_X1 U8479 ( .A(n12645), .ZN(n12783) );
  AND2_X1 U8480 ( .A1(n12781), .A2(n12782), .ZN(n12987) );
  AND2_X1 U8481 ( .A1(n7477), .A2(n7475), .ZN(n12995) );
  NAND2_X1 U8482 ( .A1(n7478), .A2(n7477), .ZN(n13011) );
  INV_X1 U8483 ( .A(n7332), .ZN(n7324) );
  NAND2_X1 U8484 ( .A1(n7332), .A2(n9886), .ZN(n7325) );
  INV_X1 U8485 ( .A(n7328), .ZN(n7327) );
  OR2_X1 U8486 ( .A1(n13029), .A2(n13028), .ZN(n13035) );
  INV_X1 U8487 ( .A(n9881), .ZN(n9435) );
  NAND2_X1 U8488 ( .A1(n9827), .A2(n9826), .ZN(n13096) );
  NAND2_X1 U8489 ( .A1(n9432), .A2(n12528), .ZN(n9834) );
  INV_X1 U8490 ( .A(n9820), .ZN(n9432) );
  AOI21_X1 U8491 ( .B1(n13125), .B2(n7471), .A(n7470), .ZN(n7469) );
  INV_X1 U8492 ( .A(n12731), .ZN(n7471) );
  AND4_X1 U8493 ( .A1(n9810), .A2(n9809), .A3(n9808), .A4(n9807), .ZN(n13142)
         );
  INV_X1 U8494 ( .A(n9790), .ZN(n9431) );
  INV_X1 U8495 ( .A(n12818), .ZN(n13158) );
  AOI21_X1 U8496 ( .B1(n14846), .B2(n12818), .A(n7343), .ZN(n7342) );
  AOI21_X1 U8497 ( .B1(n7462), .B2(n12073), .A(n7461), .ZN(n7460) );
  INV_X1 U8498 ( .A(n12719), .ZN(n7461) );
  NAND2_X1 U8499 ( .A1(n14857), .A2(n7011), .ZN(n7459) );
  NOR2_X1 U8500 ( .A1(n7013), .A2(n7012), .ZN(n7011) );
  INV_X1 U8501 ( .A(n12703), .ZN(n7012) );
  INV_X1 U8502 ( .A(n7462), .ZN(n7013) );
  NAND2_X1 U8503 ( .A1(n7459), .A2(n7458), .ZN(n13160) );
  AND2_X1 U8504 ( .A1(n7465), .A2(n7460), .ZN(n7458) );
  NOR2_X1 U8505 ( .A1(n9732), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9756) );
  OR2_X1 U8506 ( .A1(n9690), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9709) );
  OR2_X1 U8507 ( .A1(n9709), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9732) );
  AND3_X1 U8508 ( .A1(n9686), .A2(n9685), .A3(n9684), .ZN(n12698) );
  INV_X1 U8509 ( .A(n7351), .ZN(n7350) );
  NAND2_X1 U8510 ( .A1(n7353), .A2(n9658), .ZN(n11708) );
  NOR2_X1 U8511 ( .A1(n9644), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9660) );
  AOI21_X1 U8512 ( .B1(n6995), .B2(n6996), .A(n6993), .ZN(n6992) );
  INV_X1 U8513 ( .A(n11854), .ZN(n6994) );
  INV_X1 U8514 ( .A(n12678), .ZN(n6993) );
  NAND2_X1 U8515 ( .A1(n9615), .A2(n9614), .ZN(n11553) );
  NAND2_X1 U8516 ( .A1(n7450), .A2(n12663), .ZN(n15487) );
  NAND2_X1 U8517 ( .A1(n9919), .A2(n9918), .ZN(n12467) );
  OR2_X1 U8518 ( .A1(n6687), .A2(n11975), .ZN(n9918) );
  NAND2_X1 U8519 ( .A1(n9548), .A2(n9547), .ZN(n12767) );
  AND3_X1 U8520 ( .A1(n9641), .A2(n9640), .A3(n9639), .ZN(n15546) );
  OR2_X1 U8521 ( .A1(n12650), .A2(n10047), .ZN(n10930) );
  NOR2_X1 U8522 ( .A1(n10046), .A2(n10045), .ZN(n10917) );
  AND2_X1 U8523 ( .A1(n10032), .A2(n12804), .ZN(n15566) );
  AOI21_X1 U8524 ( .B1(n7114), .B2(n7117), .A(n7112), .ZN(n7111) );
  INV_X1 U8525 ( .A(n12594), .ZN(n7112) );
  AOI21_X1 U8526 ( .B1(n7116), .B2(n7121), .A(n7115), .ZN(n7114) );
  NOR2_X1 U8527 ( .A1(n7125), .A2(n12421), .ZN(n7115) );
  NOR2_X1 U8528 ( .A1(n7123), .A2(n7126), .ZN(n7116) );
  INV_X1 U8529 ( .A(n7127), .ZN(n7125) );
  NAND2_X1 U8530 ( .A1(n7121), .A2(n7118), .ZN(n7117) );
  INV_X1 U8531 ( .A(n7126), .ZN(n7118) );
  NAND2_X1 U8532 ( .A1(n7336), .A2(n9457), .ZN(n7335) );
  AND2_X1 U8533 ( .A1(n6656), .A2(n9528), .ZN(n7336) );
  INV_X1 U8534 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9457) );
  INV_X1 U8535 ( .A(n7120), .ZN(n7119) );
  OAI21_X1 U8536 ( .B1(n6825), .B2(n9523), .A(n7122), .ZN(n7120) );
  INV_X1 U8537 ( .A(n7128), .ZN(n7108) );
  AND2_X1 U8539 ( .A1(n10012), .A2(n10011), .ZN(n10014) );
  AOI21_X1 U8540 ( .B1(n7138), .B2(n7140), .A(n6823), .ZN(n7136) );
  XNOR2_X1 U8541 ( .A(n10030), .B(n10029), .ZN(n10918) );
  AND2_X1 U8542 ( .A1(n9498), .A2(n9497), .ZN(n9776) );
  INV_X1 U8543 ( .A(n9746), .ZN(n9843) );
  AND2_X1 U8544 ( .A1(n9495), .A2(n9494), .ZN(n9764) );
  OR2_X1 U8545 ( .A1(n9697), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9718) );
  AND2_X1 U8546 ( .A1(n10342), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9477) );
  XNOR2_X1 U8547 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9653) );
  AND2_X1 U8548 ( .A1(n9637), .A2(n9444), .ZN(n9650) );
  XNOR2_X1 U8549 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9623) );
  XNOR2_X1 U8550 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9610) );
  XNOR2_X1 U8551 ( .A(n7033), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U8552 ( .A1(n9566), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8553 ( .A1(n10809), .A2(n9564), .ZN(n9566) );
  NOR2_X1 U8554 ( .A1(n8039), .A2(n11630), .ZN(n8056) );
  AOI21_X1 U8555 ( .B1(n6984), .B2(n6988), .A(n7573), .ZN(n6987) );
  NAND2_X1 U8556 ( .A1(n6988), .A2(n6985), .ZN(n6986) );
  NAND2_X1 U8557 ( .A1(n6966), .A2(n10180), .ZN(n6965) );
  NAND2_X1 U8558 ( .A1(n6968), .A2(n6973), .ZN(n6966) );
  NOR2_X1 U8559 ( .A1(n8108), .A2(n8107), .ZN(n8133) );
  NAND2_X1 U8560 ( .A1(n13418), .A2(n13416), .ZN(n7546) );
  NAND2_X1 U8561 ( .A1(n13342), .A2(n10139), .ZN(n13354) );
  INV_X1 U8562 ( .A(n7566), .ZN(n7564) );
  INV_X1 U8563 ( .A(n6841), .ZN(n6840) );
  NAND2_X1 U8564 ( .A1(n13354), .A2(n13355), .ZN(n13353) );
  AND3_X1 U8565 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n7863) );
  AND2_X1 U8566 ( .A1(n13410), .A2(n10176), .ZN(n6975) );
  CLKBUF_X1 U8567 ( .A(n8030), .Z(n8031) );
  INV_X1 U8568 ( .A(n9296), .ZN(n10060) );
  NAND2_X1 U8569 ( .A1(n8441), .A2(n6844), .ZN(n6843) );
  NOR2_X1 U8570 ( .A1(n6746), .A2(n6845), .ZN(n6844) );
  NAND2_X1 U8571 ( .A1(n8343), .A2(n6753), .ZN(n6845) );
  NAND2_X1 U8572 ( .A1(n8441), .A2(n6745), .ZN(n6902) );
  AOI21_X1 U8573 ( .B1(n8451), .B2(n8452), .A(n7646), .ZN(n8453) );
  OR2_X1 U8574 ( .A1(n6671), .A2(n7780), .ZN(n7782) );
  OR2_X1 U8575 ( .A1(n7810), .A2(n10356), .ZN(n7725) );
  NAND2_X1 U8576 ( .A1(n7684), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7713) );
  OR2_X1 U8577 ( .A1(n8428), .A2(n7681), .ZN(n7716) );
  OR2_X1 U8578 ( .A1(n6672), .A2(n10660), .ZN(n7717) );
  OR2_X1 U8579 ( .A1(n10353), .A2(n10352), .ZN(n10365) );
  NAND2_X1 U8580 ( .A1(n10415), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7099) );
  NOR2_X1 U8581 ( .A1(n10666), .A2(n7101), .ZN(n10670) );
  NOR2_X1 U8582 ( .A1(n7103), .A2(n7102), .ZN(n7101) );
  NAND2_X1 U8583 ( .A1(n10670), .A2(n10669), .ZN(n10868) );
  AND2_X1 U8584 ( .A1(n7096), .A2(n7095), .ZN(n11399) );
  NAND2_X1 U8585 ( .A1(n11396), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7095) );
  OR2_X1 U8586 ( .A1(n11626), .A2(n11625), .ZN(n11894) );
  NOR2_X1 U8587 ( .A1(n11896), .A2(n7106), .ZN(n11899) );
  NOR2_X1 U8588 ( .A1(n11629), .A2(n11616), .ZN(n7106) );
  NOR2_X1 U8589 ( .A1(n11899), .A2(n11898), .ZN(n13466) );
  XNOR2_X1 U8590 ( .A(n13469), .B(n13468), .ZN(n15260) );
  NOR2_X1 U8591 ( .A1(n13466), .A2(n7105), .ZN(n13469) );
  AND2_X1 U8592 ( .A1(n13467), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7105) );
  NOR2_X1 U8593 ( .A1(n13482), .A2(n7094), .ZN(n15273) );
  AND2_X1 U8594 ( .A1(n13483), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7094) );
  NOR2_X1 U8595 ( .A1(n15273), .A2(n15272), .ZN(n15270) );
  XNOR2_X1 U8596 ( .A(n7092), .B(n13492), .ZN(n13485) );
  OR2_X1 U8597 ( .A1(n15270), .A2(n7093), .ZN(n7092) );
  AND2_X1 U8598 ( .A1(n15280), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7093) );
  OAI211_X1 U8599 ( .C1(n9292), .C2(n6705), .A(n13531), .B(n6779), .ZN(n13532)
         );
  INV_X1 U8600 ( .A(n9237), .ZN(n7203) );
  NOR2_X1 U8601 ( .A1(n13642), .A2(n7488), .ZN(n13587) );
  INV_X1 U8602 ( .A(n7198), .ZN(n7197) );
  AOI21_X1 U8603 ( .B1(n7198), .B2(n7196), .A(n6733), .ZN(n7195) );
  NOR2_X1 U8604 ( .A1(n12191), .A2(n7199), .ZN(n7198) );
  NAND2_X1 U8605 ( .A1(n7500), .A2(n7499), .ZN(n12171) );
  OR2_X1 U8606 ( .A1(n8013), .A2(n8012), .ZN(n8039) );
  NOR2_X1 U8607 ( .A1(n11644), .A2(n11803), .ZN(n6868) );
  NAND2_X1 U8608 ( .A1(n11643), .A2(n11648), .ZN(n11644) );
  AOI21_X1 U8609 ( .B1(n11423), .B2(n11421), .A(n6761), .ZN(n11640) );
  AND2_X1 U8610 ( .A1(n7911), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U8611 ( .A1(n7485), .A2(n7484), .ZN(n11428) );
  INV_X1 U8612 ( .A(n11438), .ZN(n7485) );
  INV_X1 U8613 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7886) );
  NOR2_X1 U8614 ( .A1(n7887), .A2(n7886), .ZN(n7911) );
  NAND2_X1 U8615 ( .A1(n10854), .A2(n9211), .ZN(n10837) );
  NAND2_X1 U8616 ( .A1(n9254), .A2(n9253), .ZN(n10853) );
  NAND2_X1 U8617 ( .A1(n10761), .A2(n10762), .ZN(n10760) );
  AND2_X1 U8618 ( .A1(n9299), .A2(n11835), .ZN(n10696) );
  NAND2_X1 U8619 ( .A1(n13535), .A2(n13534), .ZN(n13533) );
  NAND2_X1 U8620 ( .A1(n8055), .A2(n8054), .ZN(n13811) );
  CLKBUF_X1 U8621 ( .A(n8516), .Z(n8517) );
  INV_X1 U8622 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8506) );
  INV_X1 U8623 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7693) );
  OR2_X1 U8624 ( .A1(n7772), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7804) );
  AOI21_X1 U8626 ( .B1(n13931), .B2(n6929), .A(n6776), .ZN(n6928) );
  INV_X1 U8627 ( .A(n12362), .ZN(n6929) );
  INV_X1 U8628 ( .A(n13931), .ZN(n6930) );
  INV_X1 U8629 ( .A(n14156), .ZN(n13881) );
  NAND2_X1 U8630 ( .A1(n12208), .A2(n7648), .ZN(n14931) );
  NAND3_X1 U8631 ( .A1(n7425), .A2(n10227), .A3(n10731), .ZN(n7426) );
  OR2_X1 U8632 ( .A1(n10226), .A2(n10225), .ZN(n10227) );
  INV_X1 U8633 ( .A(n8871), .ZN(n8880) );
  NOR2_X1 U8634 ( .A1(n14660), .A2(n8862), .ZN(n8872) );
  AOI21_X1 U8635 ( .B1(n6928), .B2(n6930), .A(n6927), .ZN(n6926) );
  INV_X1 U8636 ( .A(n13863), .ZN(n6927) );
  INV_X1 U8637 ( .A(n11775), .ZN(n7433) );
  NOR2_X1 U8638 ( .A1(n11874), .A2(n7436), .ZN(n7435) );
  INV_X1 U8639 ( .A(n11871), .ZN(n7436) );
  NOR2_X1 U8640 ( .A1(n8818), .A2(n13872), .ZN(n8827) );
  AND2_X1 U8641 ( .A1(n8838), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8849) );
  NAND2_X1 U8642 ( .A1(n8849), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U8643 ( .A1(n14931), .A2(n14930), .ZN(n14940) );
  AND2_X1 U8644 ( .A1(n14940), .A2(n12219), .ZN(n14942) );
  OR2_X1 U8645 ( .A1(n8752), .A2(n8751), .ZN(n8767) );
  NOR2_X1 U8646 ( .A1(n8767), .A2(n8766), .ZN(n8780) );
  INV_X1 U8647 ( .A(n8894), .ZN(n8873) );
  AND4_X1 U8648 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n12310)
         );
  NAND2_X1 U8649 ( .A1(n8894), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8595) );
  AOI21_X1 U8650 ( .B1(n13991), .B2(P1_REG1_REG_4__SCAN_IN), .A(n13992), .ZN(
        n10507) );
  AOI21_X1 U8651 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10535), .A(n10595), .ZN(
        n14002) );
  AOI21_X1 U8652 ( .B1(n10745), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10744), .ZN(
        n10747) );
  INV_X1 U8653 ( .A(n7159), .ZN(n14089) );
  AND2_X1 U8654 ( .A1(n14123), .A2(n8946), .ZN(n7173) );
  AND2_X1 U8655 ( .A1(n7368), .A2(n6943), .ZN(n14145) );
  NAND2_X1 U8656 ( .A1(n14145), .A2(n14301), .ZN(n14124) );
  AND2_X1 U8657 ( .A1(n14142), .A2(n6730), .ZN(n7284) );
  NAND2_X1 U8658 ( .A1(n14191), .A2(n8845), .ZN(n14171) );
  NOR2_X1 U8659 ( .A1(n7300), .A2(n9087), .ZN(n7299) );
  INV_X1 U8660 ( .A(n8937), .ZN(n7300) );
  NAND2_X1 U8661 ( .A1(n8794), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8803) );
  INV_X1 U8662 ( .A(n7162), .ZN(n7161) );
  OAI21_X1 U8663 ( .B1(n7165), .B2(n7163), .A(n8935), .ZN(n7162) );
  AND2_X1 U8664 ( .A1(n7371), .A2(n14349), .ZN(n6954) );
  NAND2_X1 U8665 ( .A1(n6704), .A2(n7371), .ZN(n12131) );
  NOR2_X1 U8666 ( .A1(n7298), .A2(n7297), .ZN(n7296) );
  NAND2_X1 U8667 ( .A1(n7373), .A2(n7372), .ZN(n14815) );
  NAND2_X1 U8668 ( .A1(n7371), .A2(n7370), .ZN(n12088) );
  NOR2_X1 U8669 ( .A1(n8725), .A2(n8550), .ZN(n8741) );
  OR2_X1 U8670 ( .A1(n6960), .A2(n12216), .ZN(n11759) );
  NAND2_X1 U8671 ( .A1(n8697), .A2(n8696), .ZN(n14925) );
  INV_X1 U8672 ( .A(n11496), .ZN(n6872) );
  AOI21_X1 U8673 ( .B1(n7260), .B2(n7262), .A(n6757), .ZN(n7258) );
  NAND2_X1 U8674 ( .A1(n15090), .A2(n15171), .ZN(n15089) );
  NAND2_X1 U8675 ( .A1(n6948), .A2(n6947), .ZN(n15110) );
  NOR2_X1 U8676 ( .A1(n15110), .A2(n11594), .ZN(n15090) );
  NAND2_X1 U8677 ( .A1(n11140), .A2(n8613), .ZN(n11170) );
  INV_X1 U8678 ( .A(n14220), .ZN(n14812) );
  INV_X1 U8679 ( .A(n15185), .ZN(n14980) );
  INV_X1 U8680 ( .A(n14265), .ZN(n14979) );
  XNOR2_X1 U8681 ( .A(n8382), .B(n8381), .ZN(n9162) );
  AND2_X1 U8682 ( .A1(n8971), .A2(n8536), .ZN(n8977) );
  OAI21_X1 U8683 ( .B1(n8299), .B2(n7508), .A(n8302), .ZN(n8322) );
  AND2_X1 U8684 ( .A1(n8983), .A2(n8982), .ZN(n9196) );
  XNOR2_X1 U8685 ( .A(n8908), .B(n8902), .ZN(n8953) );
  XNOR2_X1 U8686 ( .A(n8071), .B(n8070), .ZN(n10754) );
  NAND2_X1 U8687 ( .A1(n7514), .A2(n7515), .ZN(n8071) );
  NAND2_X1 U8688 ( .A1(n8052), .A2(n6701), .ZN(n7515) );
  NAND2_X1 U8689 ( .A1(n7509), .A2(n14777), .ZN(n7514) );
  AND2_X1 U8690 ( .A1(n8747), .A2(n8738), .ZN(n11024) );
  XNOR2_X1 U8691 ( .A(n8050), .B(n8049), .ZN(n10617) );
  OR2_X1 U8692 ( .A1(n8678), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8680) );
  OAI21_X1 U8693 ( .B1(n7904), .B2(n7071), .A(n7069), .ZN(n7942) );
  OR2_X1 U8694 ( .A1(n8667), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8678) );
  XNOR2_X1 U8695 ( .A(n7825), .B(n7823), .ZN(n10311) );
  OAI21_X1 U8696 ( .B1(n9378), .B2(n9379), .A(n7398), .ZN(n7397) );
  NAND2_X1 U8697 ( .A1(n9328), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7398) );
  NOR2_X1 U8698 ( .A1(n9339), .A2(n9338), .ZN(n9394) );
  OAI21_X1 U8699 ( .B1(n14572), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n9349), .ZN(
        n9410) );
  OAI22_X1 U8700 ( .A1(n9354), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(n9370), .B2(
        n9353), .ZN(n9419) );
  AND2_X1 U8701 ( .A1(n15012), .A2(n6852), .ZN(n9421) );
  INV_X1 U8702 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U8703 ( .A1(n7219), .A2(n7216), .ZN(n12427) );
  AND4_X1 U8704 ( .A1(n9871), .A2(n9870), .A3(n9869), .A4(n9868), .ZN(n13058)
         );
  NAND2_X1 U8705 ( .A1(n6698), .A2(n12492), .ZN(n7232) );
  OAI21_X1 U8706 ( .B1(n6698), .B2(n7238), .A(n7230), .ZN(n7229) );
  AND3_X1 U8707 ( .A1(n9673), .A2(n9672), .A3(n9671), .ZN(n11824) );
  AND2_X1 U8708 ( .A1(n12518), .A2(n12438), .ZN(n12525) );
  NAND2_X1 U8709 ( .A1(n11695), .A2(n11694), .ZN(n11697) );
  NAND2_X1 U8710 ( .A1(n7220), .A2(n7224), .ZN(n12179) );
  OR2_X1 U8711 ( .A1(n12141), .A2(n12140), .ZN(n7220) );
  INV_X1 U8712 ( .A(n11996), .ZN(n14859) );
  NAND2_X1 U8713 ( .A1(n12524), .A2(n12441), .ZN(n12563) );
  NAND2_X1 U8714 ( .A1(n10998), .A2(n10937), .ZN(n12584) );
  INV_X1 U8715 ( .A(n7240), .ZN(n7227) );
  NAND2_X1 U8716 ( .A1(n7219), .A2(n6737), .ZN(n12432) );
  AND2_X1 U8717 ( .A1(n12612), .A2(n9972), .ZN(n12616) );
  AND2_X1 U8718 ( .A1(n12612), .A2(n9958), .ZN(n12977) );
  INV_X1 U8719 ( .A(n13058), .ZN(n13085) );
  OR2_X1 U8720 ( .A1(n6668), .A2(n15572), .ZN(n9552) );
  OR2_X1 U8721 ( .A1(n6684), .A2(n10827), .ZN(n9573) );
  OR2_X1 U8722 ( .A1(n9600), .A2(n10941), .ZN(n9572) );
  INV_X1 U8723 ( .A(n10959), .ZN(n10956) );
  NOR2_X1 U8724 ( .A1(n7029), .A2(n7028), .ZN(n7027) );
  NOR2_X1 U8725 ( .A1(n15408), .A2(n11267), .ZN(n15428) );
  INV_X1 U8726 ( .A(n7026), .ZN(n15426) );
  NAND2_X1 U8727 ( .A1(n7407), .A2(n11268), .ZN(n15447) );
  INV_X1 U8728 ( .A(n15446), .ZN(n7405) );
  AND2_X1 U8729 ( .A1(n6694), .A2(n7414), .ZN(n11653) );
  INV_X1 U8730 ( .A(n11653), .ZN(n7411) );
  NAND2_X1 U8731 ( .A1(n11654), .A2(n7415), .ZN(n7410) );
  NAND2_X1 U8732 ( .A1(n7417), .A2(n12843), .ZN(n11954) );
  OAI22_X1 U8733 ( .A1(n12872), .A2(n7024), .B1(n12880), .B2(n12882), .ZN(
        n12908) );
  OR2_X1 U8734 ( .A1(n12882), .A2(n13146), .ZN(n7024) );
  INV_X1 U8735 ( .A(n7019), .ZN(n14835) );
  NAND2_X1 U8736 ( .A1(n7021), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7018) );
  INV_X1 U8737 ( .A(n7419), .ZN(n7020) );
  INV_X1 U8738 ( .A(n12949), .ZN(n15463) );
  OAI21_X1 U8739 ( .B1(n12946), .B2(n12945), .A(n7035), .ZN(n12948) );
  OR2_X1 U8740 ( .A1(n12944), .A2(n12943), .ZN(n7035) );
  OAI21_X1 U8741 ( .B1(n12280), .B2(n15490), .A(n12279), .ZN(n12284) );
  OR2_X1 U8742 ( .A1(n9591), .A2(n12304), .ZN(n9935) );
  NAND2_X1 U8743 ( .A1(n7326), .A2(n9886), .ZN(n13041) );
  NAND2_X1 U8744 ( .A1(n9863), .A2(n9862), .ZN(n13076) );
  NAND2_X1 U8745 ( .A1(n13109), .A2(n12740), .ZN(n13082) );
  NAND2_X1 U8746 ( .A1(n15501), .A2(n12078), .ZN(n13137) );
  NAND2_X1 U8747 ( .A1(n13152), .A2(n12731), .ZN(n13126) );
  NAND2_X1 U8748 ( .A1(n12072), .A2(n9751), .ZN(n14840) );
  NAND2_X1 U8749 ( .A1(n7464), .A2(n12717), .ZN(n14845) );
  NAND2_X1 U8750 ( .A1(n12077), .A2(n7340), .ZN(n7464) );
  AND2_X1 U8751 ( .A1(n11978), .A2(n12710), .ZN(n14858) );
  NAND2_X1 U8752 ( .A1(n7009), .A2(n9985), .ZN(n11980) );
  NAND2_X1 U8753 ( .A1(n15469), .A2(n6673), .ZN(n7454) );
  NAND2_X1 U8754 ( .A1(n11856), .A2(n9981), .ZN(n11551) );
  INV_X1 U8755 ( .A(n13148), .ZN(n13163) );
  AND2_X1 U8756 ( .A1(n10932), .A2(n10800), .ZN(n15517) );
  NOR2_X1 U8757 ( .A1(n15482), .A2(n15545), .ZN(n13148) );
  AND2_X1 U8758 ( .A1(n14865), .A2(n14868), .ZN(n14885) );
  AND2_X1 U8759 ( .A1(n14869), .A2(n14868), .ZN(n14886) );
  INV_X1 U8760 ( .A(n12467), .ZN(n9928) );
  INV_X1 U8761 ( .A(n9914), .ZN(n13243) );
  INV_X1 U8762 ( .A(n12767), .ZN(n13251) );
  INV_X1 U8763 ( .A(n12453), .ZN(n13255) );
  NAND2_X1 U8764 ( .A1(n9852), .A2(n9851), .ZN(n13264) );
  NAND2_X1 U8765 ( .A1(n9833), .A2(n9832), .ZN(n13267) );
  NAND2_X1 U8766 ( .A1(n9819), .A2(n9818), .ZN(n13271) );
  INV_X1 U8767 ( .A(n10802), .ZN(n10790) );
  OR2_X1 U8768 ( .A1(n15568), .A2(n15545), .ZN(n13285) );
  INV_X1 U8769 ( .A(n10471), .ZN(n10436) );
  INV_X1 U8770 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13287) );
  NAND2_X1 U8771 ( .A1(n7110), .A2(n7114), .ZN(n12595) );
  OR2_X1 U8772 ( .A1(n9934), .A2(n7117), .ZN(n7110) );
  NAND2_X1 U8773 ( .A1(n7109), .A2(n7107), .ZN(n12420) );
  AOI21_X1 U8774 ( .B1(n7119), .B2(n6825), .A(n7108), .ZN(n7107) );
  NAND2_X1 U8775 ( .A1(n10011), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7010) );
  AND2_X1 U8776 ( .A1(n7156), .A2(n9519), .ZN(n9532) );
  XNOR2_X1 U8777 ( .A(n10007), .B(n10006), .ZN(n11883) );
  OAI21_X1 U8778 ( .B1(n10005), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n10007) );
  INV_X1 U8779 ( .A(SI_25_), .ZN(n14664) );
  NAND2_X1 U8780 ( .A1(n7137), .A2(n9512), .ZN(n9888) );
  NAND2_X1 U8781 ( .A1(n9875), .A2(n9874), .ZN(n7137) );
  INV_X1 U8782 ( .A(n11381), .ZN(n12651) );
  INV_X1 U8783 ( .A(SI_20_), .ZN(n11059) );
  NAND2_X1 U8784 ( .A1(n9967), .A2(n9966), .ZN(n11061) );
  INV_X1 U8785 ( .A(SI_19_), .ZN(n10711) );
  INV_X1 U8786 ( .A(SI_18_), .ZN(n10654) );
  INV_X1 U8787 ( .A(SI_16_), .ZN(n10494) );
  INV_X1 U8788 ( .A(SI_15_), .ZN(n10474) );
  INV_X1 U8789 ( .A(SI_13_), .ZN(n10434) );
  INV_X1 U8790 ( .A(n11665), .ZN(n11958) );
  INV_X1 U8791 ( .A(SI_12_), .ZN(n10339) );
  NAND2_X1 U8792 ( .A1(n7146), .A2(n7144), .ZN(n9741) );
  NAND2_X1 U8793 ( .A1(n7146), .A2(n9488), .ZN(n9739) );
  INV_X1 U8794 ( .A(SI_11_), .ZN(n10321) );
  INV_X1 U8795 ( .A(SI_10_), .ZN(n10308) );
  NAND2_X1 U8796 ( .A1(n7134), .A2(n9469), .ZN(n9593) );
  NAND2_X1 U8797 ( .A1(n9555), .A2(n9554), .ZN(n7134) );
  NAND2_X1 U8798 ( .A1(n6978), .A2(n6717), .ZN(n11159) );
  NOR2_X1 U8799 ( .A1(n13294), .A2(n7566), .ZN(n13301) );
  NAND2_X1 U8800 ( .A1(n11259), .A2(n10103), .ZN(n11799) );
  OR2_X1 U8801 ( .A1(n10362), .A2(n10374), .ZN(n7599) );
  OR2_X1 U8802 ( .A1(n7760), .A2(n10304), .ZN(n7600) );
  NAND2_X1 U8803 ( .A1(n13384), .A2(n7571), .ZN(n13325) );
  AND2_X1 U8804 ( .A1(n13384), .A2(n10156), .ZN(n7572) );
  NAND2_X1 U8805 ( .A1(n11793), .A2(n10114), .ZN(n11725) );
  NAND2_X1 U8806 ( .A1(n7546), .A2(n10133), .ZN(n13344) );
  INV_X1 U8807 ( .A(n8474), .ZN(n10655) );
  OAI21_X1 U8808 ( .B1(n11725), .B2(n11722), .A(n11723), .ZN(n11885) );
  XNOR2_X1 U8809 ( .A(n10164), .B(n10162), .ZN(n13386) );
  OR2_X1 U8810 ( .A1(n10486), .A2(n10485), .ZN(n10681) );
  OR2_X1 U8811 ( .A1(n10192), .A2(n10191), .ZN(n13397) );
  NAND2_X1 U8812 ( .A1(n13353), .A2(n10145), .ZN(n13396) );
  NAND2_X1 U8813 ( .A1(n10487), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13406) );
  NAND2_X1 U8814 ( .A1(n10706), .A2(n7570), .ZN(n11126) );
  NAND2_X1 U8815 ( .A1(n10706), .A2(n10084), .ZN(n10889) );
  NOR2_X1 U8816 ( .A1(n13397), .A2(n13661), .ZN(n13421) );
  NOR3_X1 U8817 ( .A1(n8494), .A2(n8493), .A3(n8492), .ZN(n8495) );
  INV_X1 U8818 ( .A(n10911), .ZN(n7518) );
  OR3_X1 U8819 ( .A1(n8390), .A2(n8389), .A3(n8388), .ZN(n13510) );
  OR2_X1 U8820 ( .A1(n6672), .A2(n10676), .ZN(n7747) );
  OR2_X1 U8821 ( .A1(n6670), .A2(n10357), .ZN(n7745) );
  OR2_X2 U8822 ( .A1(n10365), .A2(P2_U3088), .ZN(n13451) );
  INV_X1 U8823 ( .A(n7100), .ZN(n10405) );
  NOR2_X1 U8824 ( .A1(n10564), .A2(n10563), .ZN(n10666) );
  NOR2_X1 U8825 ( .A1(n10562), .A2(n7104), .ZN(n10564) );
  AND2_X1 U8826 ( .A1(n10565), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7104) );
  INV_X1 U8827 ( .A(n7098), .ZN(n11218) );
  INV_X1 U8828 ( .A(n7096), .ZN(n11395) );
  XNOR2_X1 U8829 ( .A(n13514), .B(n7487), .ZN(n7486) );
  INV_X1 U8830 ( .A(n8465), .ZN(n13726) );
  NAND2_X1 U8831 ( .A1(n13532), .A2(n7059), .ZN(n13732) );
  NAND2_X1 U8832 ( .A1(n13736), .A2(n7060), .ZN(n7059) );
  NOR2_X1 U8833 ( .A1(n13531), .A2(n6705), .ZN(n7060) );
  OAI21_X1 U8834 ( .B1(n13625), .B2(n7208), .A(n7204), .ZN(n13582) );
  INV_X1 U8835 ( .A(n13617), .ZN(n13755) );
  INV_X1 U8836 ( .A(n7593), .ZN(n13627) );
  NAND2_X1 U8837 ( .A1(n13767), .A2(n9286), .ZN(n13622) );
  NAND2_X1 U8838 ( .A1(n9285), .A2(n6719), .ZN(n13767) );
  NAND2_X1 U8839 ( .A1(n7189), .A2(n7190), .ZN(n13638) );
  AND2_X1 U8840 ( .A1(n7189), .A2(n7187), .ZN(n13637) );
  NAND2_X1 U8841 ( .A1(n9285), .A2(n9284), .ZN(n13651) );
  NAND2_X1 U8842 ( .A1(n7192), .A2(n7193), .ZN(n13658) );
  NAND2_X1 U8843 ( .A1(n7049), .A2(n9283), .ZN(n13656) );
  NAND2_X1 U8844 ( .A1(n7543), .A2(n7053), .ZN(n7049) );
  NAND2_X1 U8845 ( .A1(n7543), .A2(n9281), .ZN(n13672) );
  NAND2_X1 U8846 ( .A1(n7535), .A2(n7536), .ZN(n13718) );
  NAND2_X1 U8847 ( .A1(n13799), .A2(n9276), .ZN(n12197) );
  NAND2_X1 U8848 ( .A1(n12153), .A2(n9229), .ZN(n12192) );
  NAND2_X1 U8849 ( .A1(n12162), .A2(n12161), .ZN(n13799) );
  AND2_X1 U8850 ( .A1(n12166), .A2(n9227), .ZN(n12155) );
  NAND2_X1 U8851 ( .A1(n7184), .A2(n9222), .ZN(n12042) );
  NAND2_X1 U8852 ( .A1(n11905), .A2(n9221), .ZN(n7184) );
  NAND2_X1 U8853 ( .A1(n8011), .A2(n8010), .ZN(n11917) );
  NAND2_X1 U8854 ( .A1(n11418), .A2(n9264), .ZN(n11637) );
  NAND2_X1 U8855 ( .A1(n9263), .A2(n9262), .ZN(n11416) );
  OR2_X1 U8856 ( .A1(n15301), .A2(n10262), .ZN(n13519) );
  AND2_X1 U8857 ( .A1(n9300), .A2(n7591), .ZN(n7579) );
  NAND2_X1 U8858 ( .A1(n13528), .A2(n15339), .ZN(n7544) );
  NAND2_X1 U8859 ( .A1(n13740), .A2(n13739), .ZN(n13820) );
  AND2_X1 U8860 ( .A1(n13738), .A2(n13737), .ZN(n13739) );
  OR2_X1 U8861 ( .A1(n9315), .A2(P2_U3088), .ZN(n15311) );
  INV_X1 U8862 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13835) );
  NOR2_X1 U8863 ( .A1(n7675), .A2(n7210), .ZN(n7209) );
  NAND2_X1 U8864 ( .A1(n7606), .A2(n7679), .ZN(n7210) );
  AOI21_X1 U8865 ( .B1(n7057), .B2(n7056), .A(n7678), .ZN(n7055) );
  NOR2_X1 U8866 ( .A1(n7675), .A2(n7607), .ZN(n7056) );
  NAND2_X1 U8867 ( .A1(n8508), .A2(n7701), .ZN(n7702) );
  NOR2_X1 U8868 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7700) );
  OAI21_X1 U8869 ( .B1(n8503), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8504) );
  INV_X1 U8870 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n14521) );
  INV_X1 U8871 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11548) );
  INV_X1 U8872 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11227) );
  INV_X1 U8873 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n14648) );
  INV_X1 U8874 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10993) );
  INV_X1 U8875 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10620) );
  INV_X1 U8876 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10559) );
  INV_X1 U8877 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10469) );
  AND2_X1 U8878 ( .A1(n7950), .A2(n7976), .ZN(n11219) );
  INV_X1 U8879 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10342) );
  AND2_X1 U8880 ( .A1(n7831), .A2(n7881), .ZN(n10429) );
  INV_X1 U8881 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10318) );
  NAND2_X1 U8882 ( .A1(n11776), .A2(n11775), .ZN(n11872) );
  NAND2_X1 U8883 ( .A1(n6919), .A2(n7427), .ZN(n13854) );
  OAI21_X1 U8884 ( .B1(n13877), .B2(n6930), .A(n6928), .ZN(n13862) );
  NAND2_X1 U8885 ( .A1(n10731), .A2(n10227), .ZN(n11111) );
  NAND2_X1 U8886 ( .A1(n6938), .A2(n6936), .ZN(n13869) );
  NOR2_X1 U8887 ( .A1(n6937), .A2(n6939), .ZN(n6936) );
  INV_X1 U8888 ( .A(n13870), .ZN(n6937) );
  AND2_X1 U8889 ( .A1(n6938), .A2(n7420), .ZN(n13871) );
  NAND2_X1 U8890 ( .A1(n6916), .A2(n12413), .ZN(n6915) );
  INV_X1 U8891 ( .A(n6920), .ZN(n6916) );
  NAND2_X1 U8892 ( .A1(n6918), .A2(n12413), .ZN(n6917) );
  NAND2_X1 U8893 ( .A1(n11872), .A2(n11871), .ZN(n11873) );
  NAND2_X1 U8894 ( .A1(n10215), .A2(n10223), .ZN(n10216) );
  AND2_X1 U8895 ( .A1(n10219), .A2(n10218), .ZN(n10220) );
  NAND2_X1 U8896 ( .A1(n13922), .A2(n12357), .ZN(n13879) );
  NAND2_X1 U8897 ( .A1(n7440), .A2(n7439), .ZN(n12240) );
  INV_X1 U8898 ( .A(n7441), .ZN(n7439) );
  INV_X1 U8899 ( .A(n14942), .ZN(n7440) );
  NOR2_X1 U8900 ( .A1(n14942), .A2(n7649), .ZN(n12229) );
  AND2_X1 U8901 ( .A1(n8779), .A2(n8778), .ZN(n14967) );
  NAND2_X1 U8902 ( .A1(n13894), .A2(n12334), .ZN(n13905) );
  AOI21_X1 U8903 ( .B1(n6934), .B2(n6932), .A(n7438), .ZN(n6931) );
  INV_X1 U8904 ( .A(n6934), .ZN(n6933) );
  INV_X1 U8905 ( .A(n7648), .ZN(n6932) );
  NAND2_X1 U8906 ( .A1(n13930), .A2(n13931), .ZN(n13929) );
  NAND2_X1 U8907 ( .A1(n13877), .A2(n12362), .ZN(n13930) );
  INV_X1 U8908 ( .A(n14909), .ZN(n14954) );
  OAI21_X1 U8909 ( .B1(n13894), .B2(n7424), .A(n7422), .ZN(n13937) );
  OR2_X1 U8910 ( .A1(n10243), .A2(n10237), .ZN(n14916) );
  NAND2_X1 U8911 ( .A1(n7428), .A2(n12394), .ZN(n13947) );
  NAND2_X1 U8912 ( .A1(n13886), .A2(n13887), .ZN(n7428) );
  AND2_X1 U8913 ( .A1(n14926), .A2(n14980), .ZN(n14921) );
  INV_X1 U8914 ( .A(n14916), .ZN(n14960) );
  AND2_X1 U8915 ( .A1(n10242), .A2(n12011), .ZN(n14964) );
  NAND2_X1 U8916 ( .A1(n6834), .A2(n6763), .ZN(n6833) );
  INV_X1 U8917 ( .A(n9173), .ZN(n6834) );
  NAND2_X1 U8918 ( .A1(n8894), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7447) );
  AOI21_X1 U8919 ( .B1(n10533), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10545), .ZN(
        n10597) );
  NAND2_X1 U8920 ( .A1(n15049), .A2(n6718), .ZN(n11924) );
  INV_X1 U8921 ( .A(n15056), .ZN(n15044) );
  AOI22_X1 U8922 ( .A1(n14376), .A2(n9154), .B1(P2_DATAO_REG_31__SCAN_IN), 
        .B2(n9163), .ZN(n14274) );
  AND2_X1 U8923 ( .A1(n8540), .A2(n8539), .ZN(n12259) );
  NAND2_X1 U8924 ( .A1(n14086), .A2(n14090), .ZN(n14088) );
  NAND2_X1 U8925 ( .A1(n7277), .A2(n7275), .ZN(n14086) );
  NAND2_X1 U8926 ( .A1(n12269), .A2(n9154), .ZN(n7061) );
  NAND2_X1 U8927 ( .A1(n14120), .A2(n8886), .ZN(n14108) );
  NAND2_X1 U8928 ( .A1(n6854), .A2(n8946), .ZN(n14119) );
  NAND2_X1 U8929 ( .A1(n14153), .A2(n8944), .ZN(n14141) );
  NAND2_X1 U8930 ( .A1(n14208), .A2(n8835), .ZN(n14193) );
  NAND2_X1 U8931 ( .A1(n7301), .A2(n9182), .ZN(n14234) );
  NAND2_X1 U8932 ( .A1(n12101), .A2(n8934), .ZN(n12130) );
  INV_X1 U8933 ( .A(n14967), .ZN(n12106) );
  NAND2_X1 U8934 ( .A1(n8933), .A2(n9077), .ZN(n12099) );
  NAND2_X1 U8935 ( .A1(n14973), .A2(n8760), .ZN(n12093) );
  NAND2_X1 U8936 ( .A1(n7268), .A2(n8732), .ZN(n14800) );
  NAND2_X1 U8937 ( .A1(n11752), .A2(n11754), .ZN(n7268) );
  NAND2_X1 U8938 ( .A1(n8724), .A2(n8723), .ZN(n12227) );
  NAND2_X1 U8939 ( .A1(n11370), .A2(n11371), .ZN(n7259) );
  NAND2_X1 U8940 ( .A1(n12255), .A2(n14801), .ZN(n14804) );
  INV_X1 U8941 ( .A(n11758), .ZN(n15102) );
  OR2_X1 U8942 ( .A1(n15118), .A2(n11120), .ZN(n14210) );
  INV_X1 U8943 ( .A(n11765), .ZN(n15114) );
  NAND2_X1 U8944 ( .A1(n11067), .A2(n11066), .ZN(n14801) );
  INV_X1 U8945 ( .A(n14210), .ZN(n14809) );
  AND2_X2 U8946 ( .A1(n9206), .A2(n9205), .ZN(n15215) );
  OAI21_X1 U8947 ( .B1(n12252), .B2(n15125), .A(n6775), .ZN(n7358) );
  INV_X1 U8948 ( .A(n8962), .ZN(n7359) );
  NAND2_X1 U8949 ( .A1(n15199), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U8950 ( .A1(n14281), .A2(n14280), .ZN(n14282) );
  NOR2_X1 U8951 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n7443) );
  INV_X1 U8953 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14597) );
  INV_X1 U8954 ( .A(n8542), .ZN(n7256) );
  INV_X1 U8955 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14396) );
  NAND2_X1 U8956 ( .A1(n8982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8966) );
  INV_X1 U8957 ( .A(n11079), .ZN(n14400) );
  NAND2_X1 U8958 ( .A1(n7303), .A2(n7304), .ZN(n8905) );
  AND2_X1 U8959 ( .A1(n8902), .A2(n8814), .ZN(n7304) );
  INV_X1 U8960 ( .A(n8953), .ZN(n14757) );
  XNOR2_X1 U8961 ( .A(n8815), .B(n8814), .ZN(n14206) );
  INV_X1 U8962 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n14610) );
  INV_X1 U8963 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n14636) );
  INV_X1 U8964 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10991) );
  INV_X1 U8965 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10755) );
  INV_X1 U8966 ( .A(n11024), .ZN(n11342) );
  INV_X1 U8967 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10560) );
  INV_X1 U8968 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10467) );
  INV_X1 U8969 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10438) );
  INV_X1 U8970 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10395) );
  INV_X1 U8971 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10348) );
  INV_X1 U8972 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10343) );
  CLKBUF_X1 U8973 ( .A(P1_RD_REG_SCAN_IN), .Z(n6829) );
  NOR2_X1 U8974 ( .A1(n9383), .A2(n15601), .ZN(n14771) );
  AOI21_X1 U8975 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n9385), .A(n15596), .ZN(
        n15588) );
  XNOR2_X1 U8976 ( .A(n9389), .B(n6864), .ZN(n15591) );
  NAND2_X1 U8977 ( .A1(n15591), .A2(n15590), .ZN(n15589) );
  XNOR2_X1 U8978 ( .A(n9403), .B(n7392), .ZN(n14784) );
  INV_X1 U8979 ( .A(n9404), .ZN(n7392) );
  NAND2_X1 U8980 ( .A1(n14784), .A2(n14783), .ZN(n14782) );
  AND2_X1 U8981 ( .A1(n12476), .A2(n6809), .ZN(n6837) );
  NOR2_X1 U8982 ( .A1(n10040), .A2(n10042), .ZN(n10043) );
  NAND2_X1 U8983 ( .A1(n9947), .A2(n13226), .ZN(n6847) );
  NOR2_X1 U8984 ( .A1(n10055), .A2(n10057), .ZN(n10058) );
  NAND2_X1 U8985 ( .A1(n10188), .A2(n10187), .ZN(n10203) );
  AND2_X1 U8986 ( .A1(n10686), .A2(n10071), .ZN(n10629) );
  NAND2_X1 U8987 ( .A1(n7555), .A2(n10187), .ZN(n7554) );
  OAI21_X1 U8988 ( .B1(n13505), .B2(n10262), .A(n7088), .ZN(P2_U3233) );
  AOI21_X1 U8989 ( .B1(n7090), .B2(n10262), .A(n7089), .ZN(n7088) );
  OAI21_X1 U8990 ( .B1(n15269), .B2(n13507), .A(n13506), .ZN(n7089) );
  AND2_X1 U8991 ( .A1(n7589), .A2(n7591), .ZN(n13520) );
  AND2_X1 U8992 ( .A1(n7583), .A2(n6824), .ZN(n7582) );
  NAND2_X1 U8993 ( .A1(n7585), .A2(n13815), .ZN(n7584) );
  NAND2_X1 U8994 ( .A1(n7588), .A2(n7587), .ZN(n7586) );
  INV_X1 U8995 ( .A(n10403), .ZN(n10204) );
  OAI21_X1 U8996 ( .B1(n12264), .B2(n7170), .A(n7168), .ZN(P1_U3525) );
  NAND2_X1 U8997 ( .A1(n15201), .A2(n15098), .ZN(n7170) );
  INV_X1 U8998 ( .A(n7169), .ZN(n7168) );
  OAI21_X1 U8999 ( .B1(n7357), .B2(n15199), .A(n7171), .ZN(n7169) );
  CLKBUF_X1 U9000 ( .A(P2_RD_REG_SCAN_IN), .Z(n6842) );
  AND2_X1 U9001 ( .A1(n7390), .A2(n6697), .ZN(n14790) );
  NAND2_X1 U9002 ( .A1(n15006), .A2(n15004), .ZN(n15009) );
  XNOR2_X1 U9003 ( .A(n9429), .B(n9423), .ZN(n7393) );
  OR3_X1 U9004 ( .A1(n14242), .A2(n6949), .A3(n12364), .ZN(n6691) );
  AND2_X1 U9005 ( .A1(n6884), .A2(n6883), .ZN(n6692) );
  AND2_X1 U9006 ( .A1(n7370), .A2(n6955), .ZN(n6693) );
  AND2_X1 U9007 ( .A1(n11652), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6694) );
  INV_X1 U9008 ( .A(n8262), .ZN(n7990) );
  CLKBUF_X3 U9009 ( .A(n7917), .Z(n8262) );
  NAND2_X2 U9010 ( .A1(n8817), .A2(n8816), .ZN(n14229) );
  INV_X1 U9011 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8787) );
  INV_X1 U9012 ( .A(n14811), .ZN(n7267) );
  NOR2_X1 U9013 ( .A1(n14313), .A2(n14174), .ZN(n6695) );
  NOR2_X1 U9014 ( .A1(n7619), .A2(n6894), .ZN(n6696) );
  OR2_X1 U9015 ( .A1(n9407), .A2(n9406), .ZN(n6697) );
  NOR2_X1 U9016 ( .A1(n7234), .A2(n6782), .ZN(n6698) );
  OAI21_X1 U9017 ( .B1(n10362), .B2(n7707), .A(n7706), .ZN(n8474) );
  AND2_X1 U9018 ( .A1(n7082), .A2(n8194), .ZN(n6699) );
  INV_X1 U9019 ( .A(n11519), .ZN(n6947) );
  AND2_X1 U9020 ( .A1(n8051), .A2(SI_14_), .ZN(n6701) );
  INV_X1 U9021 ( .A(n12073), .ZN(n7340) );
  AND2_X1 U9022 ( .A1(n7050), .A2(n9286), .ZN(n6703) );
  INV_X1 U9023 ( .A(n12092), .ZN(n7298) );
  AND2_X1 U9024 ( .A1(n6693), .A2(n14967), .ZN(n6704) );
  AND2_X1 U9025 ( .A1(n13734), .A2(n13575), .ZN(n6705) );
  NAND2_X1 U9026 ( .A1(n8213), .A2(n8212), .ZN(n13772) );
  INV_X1 U9027 ( .A(n11638), .ZN(n7527) );
  XOR2_X1 U9028 ( .A(n7149), .B(n12942), .Z(n6706) );
  NAND2_X1 U9029 ( .A1(n7493), .A2(n7497), .ZN(n7685) );
  NAND2_X1 U9030 ( .A1(n7522), .A2(n7519), .ZN(n7732) );
  AND2_X1 U9031 ( .A1(n13669), .A2(n13433), .ZN(n6707) );
  AND2_X1 U9032 ( .A1(n7556), .A2(n6765), .ZN(n6708) );
  INV_X1 U9033 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8541) );
  AND2_X1 U9034 ( .A1(n7935), .A2(n7934), .ZN(n6709) );
  NOR2_X1 U9035 ( .A1(n7612), .A2(n7610), .ZN(n6710) );
  OR2_X1 U9036 ( .A1(n7341), .A2(n7342), .ZN(n6711) );
  AND2_X1 U9037 ( .A1(n7356), .A2(n9839), .ZN(n6712) );
  NAND2_X2 U9038 ( .A1(n10696), .A2(n11719), .ZN(n10861) );
  INV_X1 U9039 ( .A(n13650), .ZN(n7541) );
  INV_X1 U9040 ( .A(n13156), .ZN(n7465) );
  NOR2_X1 U9041 ( .A1(n14242), .A2(n6949), .ZN(n6713) );
  INV_X1 U9042 ( .A(n13759), .ZN(n7491) );
  INV_X1 U9043 ( .A(n11657), .ZN(n7415) );
  INV_X1 U9044 ( .A(n9947), .ZN(n13236) );
  AND2_X1 U9045 ( .A1(n7408), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6714) );
  INV_X1 U9046 ( .A(n12216), .ZN(n6956) );
  INV_X1 U9047 ( .A(n14981), .ZN(n7372) );
  NAND2_X1 U9048 ( .A1(n8765), .A2(n8764), .ZN(n14354) );
  INV_X1 U9049 ( .A(n14354), .ZN(n6955) );
  NAND2_X1 U9050 ( .A1(n8687), .A2(n8686), .ZN(n12029) );
  NAND2_X2 U9051 ( .A1(n9001), .A2(n10206), .ZN(n10223) );
  INV_X1 U9052 ( .A(n8600), .ZN(n8684) );
  OR2_X1 U9053 ( .A1(n12871), .A2(n12898), .ZN(n12880) );
  INV_X1 U9054 ( .A(n13752), .ZN(n13616) );
  XNOR2_X1 U9055 ( .A(n9458), .B(n9457), .ZN(n9459) );
  NAND4_X2 U9056 ( .A1(n7748), .A2(n7747), .A3(n7746), .A4(n7745), .ZN(n8475)
         );
  INV_X1 U9057 ( .A(n14107), .ZN(n7276) );
  INV_X1 U9058 ( .A(n9189), .ZN(n7361) );
  OR2_X1 U9059 ( .A1(n11265), .A2(n7027), .ZN(n6715) );
  NAND2_X1 U9060 ( .A1(n7785), .A2(n7784), .ZN(n8479) );
  NAND2_X1 U9061 ( .A1(n10207), .A2(n10205), .ZN(n12363) );
  INV_X1 U9062 ( .A(n12413), .ZN(n6924) );
  NAND2_X1 U9063 ( .A1(n7779), .A2(n7778), .ZN(n8480) );
  AND2_X1 U9064 ( .A1(n13549), .A2(n9291), .ZN(n6716) );
  AND2_X1 U9065 ( .A1(n6977), .A2(n11124), .ZN(n6717) );
  OR2_X1 U9066 ( .A1(n11923), .A2(n11928), .ZN(n6718) );
  AND2_X1 U9067 ( .A1(n7541), .A2(n9284), .ZN(n6719) );
  NAND2_X1 U9068 ( .A1(n9298), .A2(n7709), .ZN(n7845) );
  AND2_X1 U9069 ( .A1(n7622), .A2(n7623), .ZN(n6720) );
  AND2_X1 U9070 ( .A1(n9132), .A2(n9131), .ZN(n6721) );
  NOR2_X1 U9071 ( .A1(n9797), .A2(n9988), .ZN(n6722) );
  INV_X1 U9072 ( .A(n14090), .ZN(n7274) );
  NAND2_X1 U9073 ( .A1(n7303), .A2(n7302), .ZN(n8963) );
  NAND2_X1 U9074 ( .A1(n8980), .A2(n8979), .ZN(n10207) );
  AND2_X1 U9075 ( .A1(n12201), .A2(n13437), .ZN(n6723) );
  NOR2_X1 U9076 ( .A1(n12570), .A2(n7236), .ZN(n6724) );
  NAND2_X1 U9077 ( .A1(n11953), .A2(n12836), .ZN(n12843) );
  INV_X1 U9078 ( .A(n14256), .ZN(n6858) );
  NAND2_X1 U9079 ( .A1(n8712), .A2(n8711), .ZN(n12216) );
  AND2_X1 U9080 ( .A1(n7237), .A2(n7239), .ZN(n6725) );
  INV_X1 U9081 ( .A(n7079), .ZN(n7078) );
  NAND2_X1 U9082 ( .A1(n8049), .A2(n6736), .ZN(n7079) );
  AND2_X1 U9083 ( .A1(n7037), .A2(n14824), .ZN(n6726) );
  AND2_X1 U9084 ( .A1(n12490), .A2(n6724), .ZN(n6727) );
  AND4_X1 U9085 ( .A1(n8968), .A2(n8812), .A3(n8535), .A4(n8534), .ZN(n6728)
         );
  INV_X1 U9086 ( .A(n13511), .ZN(n7487) );
  INV_X1 U9087 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7679) );
  INV_X1 U9088 ( .A(n13904), .ZN(n7424) );
  AND2_X1 U9089 ( .A1(n13938), .A2(n13904), .ZN(n6729) );
  INV_X1 U9090 ( .A(n9178), .ZN(n15067) );
  NAND2_X1 U9091 ( .A1(n12293), .A2(n7682), .ZN(n7836) );
  BUF_X1 U9092 ( .A(n7836), .Z(n8387) );
  NAND2_X1 U9093 ( .A1(n14313), .A2(n14174), .ZN(n6730) );
  INV_X1 U9094 ( .A(n9047), .ZN(n7311) );
  INV_X1 U9095 ( .A(n9130), .ZN(n7317) );
  AND2_X1 U9096 ( .A1(n7100), .A2(n7099), .ZN(n6731) );
  AND2_X1 U9097 ( .A1(n6697), .A2(n14789), .ZN(n6732) );
  NOR2_X1 U9098 ( .A1(n13792), .A2(n13437), .ZN(n6733) );
  AND2_X1 U9099 ( .A1(n15251), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6734) );
  AND2_X1 U9100 ( .A1(n12467), .A2(n9927), .ZN(n12624) );
  AND2_X1 U9101 ( .A1(n10133), .A2(n7545), .ZN(n6735) );
  NAND2_X1 U9102 ( .A1(n8132), .A2(n8131), .ZN(n12201) );
  OR2_X1 U9103 ( .A1(n7513), .A2(n14777), .ZN(n6736) );
  INV_X1 U9104 ( .A(n9264), .ZN(n7531) );
  AND2_X1 U9105 ( .A1(n7216), .A2(n7223), .ZN(n6737) );
  NOR2_X1 U9106 ( .A1(n13301), .A2(n10168), .ZN(n6738) );
  AND2_X1 U9107 ( .A1(n12759), .A2(n12740), .ZN(n6739) );
  AND2_X1 U9108 ( .A1(n8363), .A2(n8362), .ZN(n6740) );
  INV_X1 U9109 ( .A(n8252), .ZN(n7640) );
  INV_X1 U9110 ( .A(n7489), .ZN(n13612) );
  NOR3_X1 U9111 ( .A1(n13642), .A2(n13752), .A3(n13759), .ZN(n7489) );
  AND2_X1 U9112 ( .A1(n8047), .A2(n8046), .ZN(n6741) );
  AND2_X1 U9113 ( .A1(n8205), .A2(n8204), .ZN(n6742) );
  AND2_X1 U9114 ( .A1(n8296), .A2(n8295), .ZN(n6743) );
  NOR2_X1 U9115 ( .A1(n6898), .A2(n6743), .ZN(n6897) );
  INV_X1 U9116 ( .A(n7367), .ZN(n14111) );
  NOR2_X1 U9117 ( .A1(n14124), .A2(n14112), .ZN(n7367) );
  INV_X1 U9118 ( .A(n13095), .ZN(n13107) );
  AND2_X1 U9119 ( .A1(n12740), .A2(n12743), .ZN(n13095) );
  AOI21_X1 U9120 ( .B1(n12140), .B2(n7224), .A(n7222), .ZN(n7221) );
  INV_X1 U9121 ( .A(n13331), .ZN(n6973) );
  AND2_X1 U9122 ( .A1(n9987), .A2(n12710), .ZN(n6744) );
  INV_X1 U9123 ( .A(n12648), .ZN(n7154) );
  AND2_X1 U9124 ( .A1(n6903), .A2(n6740), .ZN(n6745) );
  AND2_X1 U9125 ( .A1(n8340), .A2(n8339), .ZN(n6746) );
  INV_X1 U9126 ( .A(n9286), .ZN(n7540) );
  NOR2_X1 U9127 ( .A1(n12908), .A2(n12907), .ZN(n12909) );
  AND2_X1 U9128 ( .A1(n9123), .A2(n9122), .ZN(n6747) );
  AND2_X1 U9129 ( .A1(n12281), .A2(n15566), .ZN(n6748) );
  INV_X1 U9130 ( .A(n15010), .ZN(n7382) );
  INV_X1 U9131 ( .A(n9886), .ZN(n7329) );
  AND2_X1 U9132 ( .A1(n10628), .A2(n10071), .ZN(n6749) );
  NAND2_X1 U9133 ( .A1(n7565), .A2(n7564), .ZN(n6750) );
  AND2_X1 U9134 ( .A1(n9986), .A2(n9985), .ZN(n6751) );
  INV_X1 U9135 ( .A(n12029), .ZN(n7364) );
  OR2_X1 U9136 ( .A1(n8901), .A2(n7305), .ZN(n6752) );
  OR2_X1 U9137 ( .A1(n6903), .A2(n6740), .ZN(n6753) );
  INV_X1 U9138 ( .A(n9988), .ZN(n13149) );
  AND2_X1 U9139 ( .A1(n12400), .A2(n12399), .ZN(n6754) );
  AND2_X1 U9140 ( .A1(n14399), .A2(n8848), .ZN(n12364) );
  INV_X1 U9141 ( .A(n12364), .ZN(n7369) );
  AND2_X1 U9142 ( .A1(n9688), .A2(n7349), .ZN(n6755) );
  AND2_X1 U9143 ( .A1(n12407), .A2(n12406), .ZN(n6756) );
  NAND2_X1 U9144 ( .A1(n8793), .A2(n8792), .ZN(n13912) );
  INV_X1 U9145 ( .A(n13912), .ZN(n14349) );
  INV_X1 U9146 ( .A(n9283), .ZN(n7052) );
  NOR2_X1 U9147 ( .A1(n12029), .A2(n14927), .ZN(n6757) );
  NOR2_X1 U9148 ( .A1(n14308), .A2(n14157), .ZN(n6758) );
  NOR2_X1 U9149 ( .A1(n7624), .A2(n6741), .ZN(n6759) );
  NOR2_X1 U9150 ( .A1(n14981), .A2(n13958), .ZN(n6760) );
  NOR2_X1 U9151 ( .A1(n11484), .A2(n11248), .ZN(n6761) );
  NOR2_X1 U9152 ( .A1(n12039), .A2(n12119), .ZN(n6762) );
  INV_X1 U9153 ( .A(n9185), .ZN(n12098) );
  AND2_X1 U9154 ( .A1(n8934), .A2(n8784), .ZN(n9185) );
  AND2_X1 U9155 ( .A1(n9195), .A2(n9171), .ZN(n6763) );
  INV_X1 U9156 ( .A(n7633), .ZN(n7632) );
  OR2_X1 U9157 ( .A1(n7636), .A2(n8116), .ZN(n7633) );
  INV_X1 U9158 ( .A(n7194), .ZN(n7193) );
  NOR2_X1 U9159 ( .A1(n9233), .A2(n13434), .ZN(n7194) );
  AND2_X1 U9160 ( .A1(n6891), .A2(n6892), .ZN(n6764) );
  OR2_X1 U9161 ( .A1(n13318), .A2(n13313), .ZN(n6765) );
  AND2_X1 U9162 ( .A1(n12800), .A2(n12621), .ZN(n6766) );
  AND2_X1 U9163 ( .A1(n6835), .A2(n9198), .ZN(n6767) );
  NOR2_X1 U9164 ( .A1(n14285), .A2(n14069), .ZN(n6768) );
  NOR2_X1 U9165 ( .A1(n12636), .A2(n7463), .ZN(n7462) );
  OR2_X1 U9166 ( .A1(n9113), .A2(n9111), .ZN(n6769) );
  AND2_X1 U9167 ( .A1(n8315), .A2(n8314), .ZN(n6770) );
  AND2_X1 U9168 ( .A1(n6904), .A2(n6907), .ZN(n6771) );
  INV_X1 U9169 ( .A(n7607), .ZN(n7606) );
  NAND2_X1 U9170 ( .A1(n7676), .A2(n7697), .ZN(n7607) );
  AND2_X1 U9171 ( .A1(n7925), .A2(SI_8_), .ZN(n6772) );
  NOR2_X1 U9172 ( .A1(n12561), .A2(n13118), .ZN(n6773) );
  OAI21_X1 U9173 ( .B1(n12671), .B2(n6996), .A(n12676), .ZN(n6991) );
  INV_X1 U9174 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n10002) );
  AND2_X1 U9175 ( .A1(n7818), .A2(n7817), .ZN(n6774) );
  AND2_X1 U9176 ( .A1(n7360), .A2(n7359), .ZN(n6775) );
  AND2_X1 U9177 ( .A1(n12371), .A2(n12370), .ZN(n6776) );
  AND2_X1 U9178 ( .A1(n12341), .A2(n12340), .ZN(n6777) );
  INV_X1 U9179 ( .A(n7188), .ZN(n7187) );
  NAND2_X1 U9180 ( .A1(n13650), .A2(n7190), .ZN(n7188) );
  AND4_X1 U9181 ( .A1(n9451), .A2(n9450), .A3(n9780), .A4(n9816), .ZN(n6778)
         );
  OR2_X1 U9182 ( .A1(n6716), .A2(n6705), .ZN(n6779) );
  INV_X1 U9183 ( .A(n7249), .ZN(n7248) );
  OR2_X1 U9184 ( .A1(n12442), .A2(n7250), .ZN(n7249) );
  INV_X1 U9185 ( .A(n7182), .ZN(n7181) );
  OR2_X1 U9186 ( .A1(n9223), .A2(n7183), .ZN(n7182) );
  OAI21_X1 U9187 ( .B1(n12219), .B2(n7441), .A(n12239), .ZN(n7438) );
  OAI21_X1 U9188 ( .B1(n13395), .B2(n7574), .A(n10151), .ZN(n7573) );
  NOR2_X1 U9189 ( .A1(n7576), .A2(n6989), .ZN(n6988) );
  AND3_X1 U9190 ( .A1(n9583), .A2(n9582), .A3(n9581), .ZN(n9568) );
  INV_X1 U9191 ( .A(n9136), .ZN(n7064) );
  AND2_X1 U9192 ( .A1(n12023), .A2(n12022), .ZN(n6780) );
  OR2_X1 U9193 ( .A1(n6706), .A2(n12650), .ZN(n6781) );
  AND2_X1 U9194 ( .A1(n12489), .A2(n12986), .ZN(n6782) );
  AND2_X1 U9195 ( .A1(n6920), .A2(n6924), .ZN(n6783) );
  INV_X1 U9196 ( .A(n9235), .ZN(n13626) );
  OR2_X1 U9197 ( .A1(n8067), .A2(n8069), .ZN(n6784) );
  AND2_X1 U9198 ( .A1(n8020), .A2(n8019), .ZN(n6785) );
  OR2_X1 U9199 ( .A1(n13251), .A2(n13043), .ZN(n6786) );
  NOR2_X1 U9200 ( .A1(n7605), .A2(n7604), .ZN(n6787) );
  OR2_X1 U9201 ( .A1(n9334), .A2(n9335), .ZN(n6788) );
  INV_X1 U9202 ( .A(n8070), .ZN(n7513) );
  AND2_X1 U9203 ( .A1(n13326), .A2(n10156), .ZN(n7571) );
  INV_X1 U9204 ( .A(n7571), .ZN(n6962) );
  NAND2_X1 U9205 ( .A1(n10233), .A2(n10232), .ZN(n6789) );
  AND2_X1 U9206 ( .A1(n10014), .A2(n7213), .ZN(n6790) );
  OR2_X1 U9207 ( .A1(n7320), .A2(n9027), .ZN(n6791) );
  OR2_X1 U9208 ( .A1(n7311), .A2(n9046), .ZN(n6792) );
  AND2_X1 U9209 ( .A1(n7379), .A2(n7377), .ZN(n6793) );
  OR2_X1 U9210 ( .A1(n7317), .A2(n9129), .ZN(n6794) );
  OR2_X1 U9211 ( .A1(n8162), .A2(n8164), .ZN(n6795) );
  OR2_X1 U9212 ( .A1(n9056), .A2(n9058), .ZN(n6796) );
  OR2_X1 U9213 ( .A1(n9037), .A2(n9039), .ZN(n6797) );
  AND2_X1 U9214 ( .A1(n7025), .A2(n12880), .ZN(n6798) );
  OR2_X1 U9215 ( .A1(n7965), .A2(n7966), .ZN(n6799) );
  OR2_X1 U9216 ( .A1(n8252), .A2(n8253), .ZN(n6800) );
  OR2_X1 U9217 ( .A1(n6887), .A2(n6885), .ZN(n6801) );
  AND2_X1 U9218 ( .A1(n6883), .A2(n6882), .ZN(n6802) );
  AOI21_X1 U9219 ( .B1(n11884), .B2(n7550), .A(n10123), .ZN(n7549) );
  AND2_X1 U9220 ( .A1(n7381), .A2(n7383), .ZN(n6803) );
  OAI21_X1 U9221 ( .B1(n7611), .B2(n7610), .A(n7609), .ZN(n7608) );
  AND2_X1 U9222 ( .A1(n7020), .A2(n7019), .ZN(n6804) );
  INV_X1 U9223 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8814) );
  INV_X1 U9224 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9528) );
  OR2_X1 U9225 ( .A1(n8022), .A2(n6785), .ZN(n6805) );
  OR2_X1 U9226 ( .A1(n7640), .A2(n7641), .ZN(n6806) );
  INV_X1 U9227 ( .A(n7205), .ZN(n7204) );
  NAND2_X1 U9228 ( .A1(n13594), .A2(n7206), .ZN(n7205) );
  INV_X1 U9229 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6862) );
  INV_X1 U9230 ( .A(n11293), .ZN(n7028) );
  INV_X1 U9231 ( .A(n13302), .ZN(n6990) );
  INV_X1 U9232 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9720) );
  OR2_X1 U9233 ( .A1(n14242), .A2(n14229), .ZN(n6807) );
  AND2_X1 U9234 ( .A1(n7371), .A2(n6693), .ZN(n6808) );
  NAND2_X1 U9235 ( .A1(n7467), .A2(n7469), .ZN(n13113) );
  INV_X1 U9236 ( .A(n14324), .ZN(n6950) );
  INV_X1 U9237 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U9238 ( .A1(n8870), .A2(n8869), .ZN(n14308) );
  INV_X1 U9239 ( .A(n14308), .ZN(n6943) );
  INV_X1 U9240 ( .A(n12732), .ZN(n7470) );
  INV_X1 U9241 ( .A(n11317), .ZN(n15455) );
  OR2_X1 U9242 ( .A1(n13174), .A2(n12581), .ZN(n6809) );
  NAND2_X1 U9243 ( .A1(n7474), .A2(n12758), .ZN(n13078) );
  INV_X1 U9244 ( .A(n11667), .ZN(n11658) );
  NOR2_X1 U9245 ( .A1(n9724), .A2(n9723), .ZN(n11667) );
  NAND2_X1 U9246 ( .A1(n8307), .A2(n8306), .ZN(n13747) );
  INV_X1 U9247 ( .A(n13747), .ZN(n7492) );
  NAND2_X1 U9248 ( .A1(n9989), .A2(n12736), .ZN(n13106) );
  AND2_X1 U9249 ( .A1(n7459), .A2(n7460), .ZN(n6810) );
  INV_X1 U9250 ( .A(n7500), .ZN(n12170) );
  INV_X1 U9251 ( .A(n7498), .ZN(n12198) );
  OR2_X1 U9252 ( .A1(n13174), .A2(n13232), .ZN(n6811) );
  NAND2_X1 U9253 ( .A1(n11470), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6812) );
  OR2_X1 U9254 ( .A1(n14242), .A2(n6952), .ZN(n6813) );
  AND2_X1 U9255 ( .A1(n7411), .A2(n11652), .ZN(n6814) );
  NAND2_X1 U9256 ( .A1(n7009), .A2(n6751), .ZN(n11978) );
  AND2_X1 U9257 ( .A1(n13098), .A2(n9839), .ZN(n6815) );
  AND2_X1 U9258 ( .A1(n12758), .A2(n12759), .ZN(n13083) );
  INV_X1 U9259 ( .A(n13083), .ZN(n7356) );
  AND3_X1 U9260 ( .A1(n15006), .A2(n15004), .A3(n7382), .ZN(n6816) );
  OR2_X1 U9261 ( .A1(n13174), .A2(n13285), .ZN(n6817) );
  INV_X1 U9262 ( .A(n7420), .ZN(n6939) );
  AOI21_X1 U9263 ( .B1(n13938), .B2(n7421), .A(n12348), .ZN(n7420) );
  AND2_X1 U9264 ( .A1(n8824), .A2(n8823), .ZN(n6818) );
  INV_X1 U9265 ( .A(n15348), .ZN(n7484) );
  XNOR2_X1 U9266 ( .A(n8965), .B(n8964), .ZN(n8976) );
  INV_X1 U9267 ( .A(n11355), .ZN(n7042) );
  NAND2_X1 U9268 ( .A1(n7259), .A2(n8677), .ZN(n15065) );
  OAI21_X1 U9269 ( .B1(n6991), .B2(n6994), .A(n6992), .ZN(n11527) );
  NAND2_X1 U9270 ( .A1(n7453), .A2(n7451), .ZN(n11838) );
  NAND2_X1 U9271 ( .A1(n7454), .A2(n12688), .ZN(n11707) );
  NAND2_X1 U9272 ( .A1(n8082), .A2(n8081), .ZN(n13805) );
  INV_X1 U9273 ( .A(n13805), .ZN(n7499) );
  OR2_X1 U9274 ( .A1(n11311), .A2(n11310), .ZN(n6819) );
  XNOR2_X1 U9275 ( .A(n8966), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8978) );
  INV_X1 U9276 ( .A(n14971), .ZN(n7370) );
  INV_X1 U9277 ( .A(n6868), .ZN(n11811) );
  AND2_X1 U9278 ( .A1(n11464), .A2(n11658), .ZN(n11654) );
  INV_X1 U9279 ( .A(n11654), .ZN(n11652) );
  NAND2_X1 U9280 ( .A1(n11269), .A2(n15455), .ZN(n11268) );
  AND2_X1 U9281 ( .A1(n11872), .A2(n7435), .ZN(n6820) );
  AND2_X1 U9282 ( .A1(n7405), .A2(n11268), .ZN(n6821) );
  INV_X1 U9283 ( .A(n8300), .ZN(n7508) );
  OR2_X1 U9284 ( .A1(n15089), .A2(n15177), .ZN(n15074) );
  INV_X1 U9285 ( .A(n15074), .ZN(n7365) );
  NAND2_X1 U9286 ( .A1(n9962), .A2(n7215), .ZN(n6822) );
  AND2_X1 U9287 ( .A1(n9513), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6823) );
  INV_X1 U9288 ( .A(n7373), .ZN(n14814) );
  AND3_X1 U9289 ( .A1(n6956), .A2(n6957), .A3(n7365), .ZN(n7373) );
  INV_X1 U9290 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7102) );
  OR2_X1 U9291 ( .A1(n13815), .A2(n7590), .ZN(n6824) );
  INV_X1 U9292 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7129) );
  AND2_X1 U9293 ( .A1(n14390), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6825) );
  INV_X1 U9294 ( .A(n12819), .ZN(n7242) );
  INV_X1 U9295 ( .A(n10701), .ZN(n6981) );
  INV_X1 U9296 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14552) );
  NAND2_X1 U9297 ( .A1(n7979), .A2(n7978), .ZN(n15286) );
  INV_X1 U9298 ( .A(n15286), .ZN(n6867) );
  NOR2_X1 U9299 ( .A1(n9786), .A2(n9785), .ZN(n12898) );
  NAND3_X1 U9300 ( .A1(n15149), .A2(n14258), .A3(n6944), .ZN(n15109) );
  INV_X1 U9301 ( .A(n15109), .ZN(n6948) );
  AND2_X1 U9302 ( .A1(n9163), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6826) );
  OR2_X1 U9303 ( .A1(n15215), .A2(n8547), .ZN(n6827) );
  INV_X1 U9304 ( .A(n14824), .ZN(n7036) );
  INV_X1 U9305 ( .A(n10262), .ZN(n13504) );
  XNOR2_X1 U9306 ( .A(n7689), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10262) );
  INV_X1 U9307 ( .A(n10667), .ZN(n7103) );
  INV_X1 U9308 ( .A(n12942), .ZN(n12649) );
  AND2_X1 U9309 ( .A1(n8952), .A2(n9153), .ZN(n15083) );
  INV_X1 U9310 ( .A(n15083), .ZN(n15098) );
  INV_X1 U9311 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7375) );
  NAND3_X1 U9312 ( .A1(n6843), .A2(n6902), .A3(n8453), .ZN(n6828) );
  NAND2_X1 U9313 ( .A1(n11446), .A2(n11445), .ZN(n11444) );
  NAND2_X1 U9314 ( .A1(n7588), .A2(n13705), .ZN(n7589) );
  NAND2_X1 U9315 ( .A1(n11640), .A2(n7527), .ZN(n11639) );
  NAND2_X1 U9316 ( .A1(n7602), .A2(n7601), .ZN(n13535) );
  NAND2_X1 U9317 ( .A1(n9225), .A2(n9224), .ZN(n12114) );
  AOI21_X1 U9318 ( .B1(n13375), .B2(n13782), .A(n9232), .ZN(n13673) );
  OAI211_X1 U9319 ( .C1(n10856), .C2(n7596), .A(n7595), .B(n9213), .ZN(n7178)
         );
  XNOR2_X1 U9320 ( .A(n9374), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U9321 ( .A1(n15021), .A2(n15022), .ZN(n15020) );
  INV_X1 U9322 ( .A(n7397), .ZN(n9377) );
  OAI21_X2 U9323 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n9422), .A(n14820), .ZN(
        n14765) );
  NAND2_X1 U9324 ( .A1(n6793), .A2(n6853), .ZN(n6852) );
  NAND2_X1 U9325 ( .A1(n15013), .A2(n15014), .ZN(n15012) );
  XNOR2_X1 U9326 ( .A(n9331), .B(n6862), .ZN(n9375) );
  NAND2_X1 U9327 ( .A1(n7374), .A2(n15020), .ZN(n14822) );
  OAI21_X1 U9328 ( .B1(n9374), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6788), .ZN(
        n7391) );
  XNOR2_X1 U9329 ( .A(n9398), .B(n9399), .ZN(n15594) );
  NAND2_X2 U9330 ( .A1(n13084), .A2(n9860), .ZN(n13069) );
  AND2_X1 U9331 ( .A1(n9627), .A2(n9614), .ZN(n7337) );
  NAND2_X1 U9332 ( .A1(n12976), .A2(n6830), .ZN(n9959) );
  NAND2_X1 U9333 ( .A1(n9979), .A2(n9584), .ZN(n15492) );
  NAND2_X1 U9334 ( .A1(n6846), .A2(n7650), .ZN(n13168) );
  NAND2_X1 U9335 ( .A1(n13098), .A2(n6712), .ZN(n13084) );
  NAND2_X1 U9336 ( .A1(n11858), .A2(n12630), .ZN(n9615) );
  NAND2_X1 U9337 ( .A1(n13032), .A2(n13031), .ZN(n13030) );
  NAND2_X1 U9338 ( .A1(n6832), .A2(n9201), .ZN(P1_U3242) );
  NAND3_X1 U9339 ( .A1(n6767), .A2(n7281), .A3(n6833), .ZN(n6832) );
  OAI21_X2 U9340 ( .B1(n13673), .B2(n7188), .A(n7185), .ZN(n7593) );
  NAND2_X1 U9341 ( .A1(n6836), .A2(n11080), .ZN(n6835) );
  XNOR2_X1 U9342 ( .A(n9194), .B(n11942), .ZN(n6836) );
  INV_X1 U9343 ( .A(n7178), .ZN(n11446) );
  NAND2_X2 U9344 ( .A1(n15503), .A2(n6848), .ZN(n12663) );
  NAND2_X1 U9345 ( .A1(n6838), .A2(n6837), .ZN(P3_U3154) );
  NAND2_X1 U9346 ( .A1(n12471), .A2(n12572), .ZN(n6838) );
  NAND2_X1 U9347 ( .A1(n11237), .A2(n11236), .ZN(n11454) );
  MUX2_X1 U9348 ( .A(n11005), .B(n12663), .S(n11046), .Z(n11010) );
  NAND2_X1 U9349 ( .A1(n11010), .A2(n11007), .ZN(n11035) );
  NAND2_X1 U9351 ( .A1(n7233), .A2(n6725), .ZN(n12491) );
  XNOR2_X2 U9352 ( .A(n9456), .B(n13287), .ZN(n12424) );
  INV_X1 U9353 ( .A(n7334), .ZN(n13286) );
  OAI21_X1 U9354 ( .B1(n7475), .B2(n12998), .A(n12777), .ZN(n7008) );
  NOR2_X1 U9355 ( .A1(n12275), .A2(n12783), .ZN(n12274) );
  NAND2_X1 U9356 ( .A1(n9562), .A2(n9577), .ZN(n9468) );
  NAND2_X1 U9357 ( .A1(n6851), .A2(n13031), .ZN(n7478) );
  INV_X1 U9358 ( .A(n7008), .ZN(n7007) );
  INV_X1 U9359 ( .A(n7546), .ZN(n6984) );
  NAND2_X1 U9360 ( .A1(n13403), .A2(n6975), .ZN(n13402) );
  INV_X1 U9361 ( .A(n10167), .ZN(n7568) );
  NAND2_X1 U9362 ( .A1(n14072), .A2(n14077), .ZN(n14071) );
  NAND2_X1 U9363 ( .A1(n8930), .A2(n8929), .ZN(n14810) );
  OAI21_X2 U9364 ( .B1(n14216), .B2(n14217), .A(n9101), .ZN(n14198) );
  OAI21_X2 U9365 ( .B1(n14173), .B2(n14172), .A(n8943), .ZN(n14155) );
  NAND2_X1 U9366 ( .A1(n6869), .A2(n6872), .ZN(n11493) );
  NAND2_X1 U9367 ( .A1(n11191), .A2(n11190), .ZN(n11189) );
  NAND2_X1 U9368 ( .A1(n14153), .A2(n7174), .ZN(n14139) );
  NAND2_X1 U9369 ( .A1(n11555), .A2(n9642), .ZN(n11529) );
  NAND3_X1 U9370 ( .A1(n12975), .A2(n12976), .A3(n15511), .ZN(n6846) );
  NAND2_X1 U9371 ( .A1(n13171), .A2(n6847), .ZN(P3_U3487) );
  NAND2_X1 U9372 ( .A1(n12283), .A2(n6817), .ZN(P3_U3454) );
  NAND2_X1 U9373 ( .A1(n13173), .A2(n6811), .ZN(P3_U3486) );
  XNOR2_X2 U9374 ( .A(n11150), .B(n13965), .ZN(n11142) );
  NAND2_X1 U9375 ( .A1(n13030), .A2(n6786), .ZN(n13017) );
  NAND2_X1 U9376 ( .A1(n9931), .A2(n7344), .ZN(n7348) );
  NAND2_X1 U9377 ( .A1(n11382), .A2(n9597), .ZN(n11858) );
  AND2_X1 U9378 ( .A1(n12964), .A2(n14883), .ZN(n10001) );
  NAND2_X2 U9379 ( .A1(n9511), .A2(n9510), .ZN(n9875) );
  INV_X1 U9380 ( .A(n12773), .ZN(n6851) );
  NAND2_X1 U9381 ( .A1(n6850), .A2(n9471), .ZN(n9611) );
  NAND2_X1 U9382 ( .A1(n9499), .A2(n9498), .ZN(n9801) );
  NAND2_X1 U9383 ( .A1(n9682), .A2(n9680), .ZN(n9485) );
  NAND2_X1 U9384 ( .A1(n9473), .A2(n9472), .ZN(n9624) );
  NAND3_X1 U9385 ( .A1(n7133), .A2(n9592), .A3(n7132), .ZN(n6850) );
  NAND2_X1 U9386 ( .A1(n9508), .A2(n9507), .ZN(n9509) );
  NAND2_X1 U9387 ( .A1(n9516), .A2(n9515), .ZN(n9517) );
  NAND2_X1 U9388 ( .A1(n14155), .A2(n14154), .ZN(n14153) );
  NAND2_X1 U9389 ( .A1(n14765), .A2(n14766), .ZN(n14764) );
  XNOR2_X2 U9390 ( .A(n12458), .B(n12511), .ZN(n13016) );
  NAND2_X2 U9391 ( .A1(n9902), .A2(n9901), .ZN(n12458) );
  NAND3_X1 U9392 ( .A1(n15006), .A2(n7381), .A3(n15004), .ZN(n7376) );
  NOR2_X1 U9393 ( .A1(n14822), .A2(n14821), .ZN(n9422) );
  NOR2_X2 U9394 ( .A1(n14774), .A2(n9396), .ZN(n9398) );
  AOI21_X1 U9395 ( .B1(n7007), .B2(n12998), .A(n7006), .ZN(n7005) );
  AOI21_X1 U9396 ( .B1(n6732), .B2(n7390), .A(n7389), .ZN(n7388) );
  INV_X1 U9397 ( .A(n9009), .ZN(n9008) );
  NAND2_X1 U9399 ( .A1(n7159), .A2(n7274), .ZN(n14092) );
  OR2_X1 U9400 ( .A1(n8893), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U9401 ( .A1(n7160), .A2(n8834), .ZN(n14202) );
  NAND2_X1 U9402 ( .A1(n6855), .A2(n7801), .ZN(n7825) );
  NAND2_X1 U9403 ( .A1(n7799), .A2(n7798), .ZN(n6855) );
  AOI21_X2 U9404 ( .B1(n9166), .B2(n9165), .A(n9193), .ZN(n9173) );
  NAND2_X1 U9405 ( .A1(n6856), .A2(n6827), .ZN(P1_U3557) );
  NAND2_X1 U9406 ( .A1(n9207), .A2(n15215), .ZN(n6856) );
  NAND2_X1 U9407 ( .A1(n14092), .A2(n8950), .ZN(n14072) );
  OAI211_X1 U9408 ( .C1(n13511), .C2(n13510), .A(n8392), .B(n8391), .ZN(n8421)
         );
  OAI21_X1 U9409 ( .B1(n12264), .B2(n15083), .A(n7357), .ZN(n9207) );
  NAND2_X1 U9410 ( .A1(n6861), .A2(n7003), .ZN(n12275) );
  NAND2_X1 U9411 ( .A1(n9519), .A2(n9518), .ZN(n9900) );
  NAND2_X1 U9412 ( .A1(n14110), .A2(n7276), .ZN(n14109) );
  NOR2_X1 U9413 ( .A1(n11924), .A2(n11925), .ZN(n12063) );
  NOR2_X2 U9414 ( .A1(n8599), .A2(n6658), .ZN(n10724) );
  NAND2_X1 U9415 ( .A1(n9135), .A2(n7063), .ZN(n6859) );
  OAI21_X1 U9416 ( .B1(n6747), .B2(n6860), .A(n7316), .ZN(n9133) );
  NAND2_X1 U9417 ( .A1(n9128), .A2(n6794), .ZN(n6860) );
  NAND2_X1 U9418 ( .A1(n9476), .A2(n9475), .ZN(n9636) );
  NAND2_X1 U9419 ( .A1(n9814), .A2(n9503), .ZN(n7155) );
  NAND2_X1 U9420 ( .A1(n9655), .A2(n9653), .ZN(n9480) );
  AND2_X2 U9421 ( .A1(n7478), .A2(n7476), .ZN(n7475) );
  INV_X1 U9422 ( .A(n7391), .ZN(n9336) );
  INV_X1 U9423 ( .A(n9390), .ZN(n6864) );
  NAND2_X1 U9424 ( .A1(n7395), .A2(n14764), .ZN(n7394) );
  XNOR2_X1 U9425 ( .A(n7394), .B(n7393), .ZN(SUB_1596_U4) );
  NAND3_X1 U9426 ( .A1(n7495), .A2(n7496), .A3(n7497), .ZN(n7494) );
  AND4_X2 U9427 ( .A1(n7669), .A2(n7727), .A3(n7670), .A4(n7668), .ZN(n7497)
         );
  NAND2_X1 U9428 ( .A1(n7498), .A2(n13792), .ZN(n13707) );
  INV_X1 U9429 ( .A(n11495), .ZN(n6869) );
  NAND2_X1 U9430 ( .A1(n8925), .A2(n8924), .ZN(n11495) );
  AOI21_X2 U9431 ( .B1(n14073), .B2(n15098), .A(n6870), .ZN(n14284) );
  NAND2_X2 U9432 ( .A1(n13069), .A2(n13079), .ZN(n9873) );
  OAI21_X2 U9433 ( .B1(n12276), .B2(n9946), .A(n6871), .ZN(n12975) );
  NAND2_X1 U9434 ( .A1(n7158), .A2(n8942), .ZN(n14173) );
  NAND2_X1 U9435 ( .A1(n7904), .A2(n7903), .ZN(n7924) );
  OR2_X2 U9436 ( .A1(n14267), .A2(n15135), .ZN(n9014) );
  AND3_X2 U9437 ( .A1(n8574), .A2(n8575), .A3(n8576), .ZN(n7448) );
  NAND2_X1 U9438 ( .A1(n8940), .A2(n8939), .ZN(n14216) );
  INV_X1 U9439 ( .A(n14198), .ZN(n7160) );
  NAND2_X1 U9440 ( .A1(n7742), .A2(n6873), .ZN(n7741) );
  NAND2_X1 U9441 ( .A1(n7736), .A2(n7737), .ZN(n6873) );
  INV_X1 U9442 ( .A(n6873), .ZN(n7743) );
  NAND2_X1 U9443 ( .A1(n7820), .A2(n6774), .ZN(n6874) );
  NAND2_X1 U9444 ( .A1(n6876), .A2(n6875), .ZN(n7852) );
  OAI211_X1 U9445 ( .C1(n7820), .C2(n6774), .A(n7821), .B(n7822), .ZN(n6876)
         );
  AOI21_X1 U9446 ( .B1(n6720), .B2(n6879), .A(n6877), .ZN(n7628) );
  NAND2_X1 U9447 ( .A1(n7613), .A2(n6801), .ZN(n6884) );
  NAND2_X1 U9448 ( .A1(n6881), .A2(n7611), .ZN(n8227) );
  NAND2_X1 U9449 ( .A1(n6884), .A2(n6802), .ZN(n6881) );
  INV_X1 U9450 ( .A(n6702), .ZN(n6886) );
  INV_X1 U9451 ( .A(n8185), .ZN(n6889) );
  INV_X1 U9452 ( .A(n8184), .ZN(n6890) );
  NAND2_X1 U9453 ( .A1(n8298), .A2(n6696), .ZN(n6891) );
  INV_X1 U9454 ( .A(n8297), .ZN(n6898) );
  NAND2_X1 U9455 ( .A1(n6899), .A2(n6900), .ZN(n7622) );
  NAND3_X1 U9456 ( .A1(n7998), .A2(n6805), .A3(n7997), .ZN(n6899) );
  INV_X1 U9457 ( .A(n8364), .ZN(n6903) );
  OAI21_X1 U9458 ( .B1(n7898), .B2(n7897), .A(n6907), .ZN(n6905) );
  NAND2_X1 U9459 ( .A1(n6908), .A2(n6910), .ZN(n6907) );
  AND2_X1 U9460 ( .A1(n7920), .A2(n7921), .ZN(n6909) );
  INV_X1 U9461 ( .A(n7920), .ZN(n6910) );
  NAND2_X1 U9462 ( .A1(n13886), .A2(n7429), .ZN(n6919) );
  OAI211_X1 U9463 ( .C1(n13886), .C2(n6917), .A(n6913), .B(n6912), .ZN(n12419)
         );
  NAND2_X1 U9464 ( .A1(n13886), .A2(n6783), .ZN(n6912) );
  OAI21_X1 U9465 ( .B1(n6918), .B2(n6924), .A(n6914), .ZN(n6913) );
  NAND2_X1 U9466 ( .A1(n6918), .A2(n6915), .ZN(n6914) );
  NAND2_X1 U9467 ( .A1(n13877), .A2(n6928), .ZN(n6925) );
  NAND2_X1 U9468 ( .A1(n6925), .A2(n6926), .ZN(n12379) );
  NAND2_X1 U9469 ( .A1(n13895), .A2(n6940), .ZN(n6938) );
  NAND4_X1 U9470 ( .A1(n7647), .A2(n8528), .A3(n6942), .A4(n6658), .ZN(n6941)
         );
  INV_X1 U9471 ( .A(n8813), .ZN(n8761) );
  NAND2_X1 U9472 ( .A1(n6954), .A2(n6704), .ZN(n14244) );
  INV_X1 U9473 ( .A(n6960), .ZN(n11541) );
  NAND2_X1 U9474 ( .A1(n10153), .A2(n10152), .ZN(n13384) );
  NAND2_X1 U9475 ( .A1(n6964), .A2(n6963), .ZN(n10184) );
  NAND3_X1 U9476 ( .A1(n7563), .A2(n6967), .A3(n13294), .ZN(n6964) );
  AOI21_X1 U9477 ( .B1(n7563), .B2(n6974), .A(n6973), .ZN(n6971) );
  OAI21_X1 U9478 ( .B1(n13294), .B2(n6750), .A(n7563), .ZN(n13364) );
  NAND3_X1 U9479 ( .A1(n7563), .A2(n13294), .A3(n10170), .ZN(n6972) );
  NAND2_X1 U9480 ( .A1(n6971), .A2(n6972), .ZN(n13403) );
  NAND2_X1 U9481 ( .A1(n11784), .A2(n10110), .ZN(n11793) );
  INV_X1 U9482 ( .A(n6976), .ZN(n12015) );
  NAND2_X1 U9483 ( .A1(n6979), .A2(n6982), .ZN(n6977) );
  NAND2_X1 U9484 ( .A1(n10080), .A2(n6979), .ZN(n6978) );
  AOI21_X1 U9485 ( .B1(n7570), .B2(n6981), .A(n6980), .ZN(n6979) );
  NOR2_X2 U9486 ( .A1(n7692), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7690) );
  NAND2_X1 U9487 ( .A1(n10686), .A2(n6749), .ZN(n10774) );
  NAND2_X1 U9488 ( .A1(n6983), .A2(n7548), .ZN(n10686) );
  AND2_X1 U9489 ( .A1(n7547), .A2(n10680), .ZN(n6983) );
  INV_X1 U9490 ( .A(n6735), .ZN(n6985) );
  NAND2_X1 U9491 ( .A1(n6986), .A2(n6987), .ZN(n13373) );
  NAND3_X1 U9492 ( .A1(n6987), .A2(n6990), .A3(n6986), .ZN(n13372) );
  NAND2_X1 U9493 ( .A1(n6735), .A2(n7546), .ZN(n13342) );
  INV_X1 U9494 ( .A(n6991), .ZN(n6995) );
  NAND2_X1 U9495 ( .A1(n7477), .A2(n7004), .ZN(n7003) );
  OAI21_X1 U9496 ( .B1(n7477), .B2(n12998), .A(n7007), .ZN(n12988) );
  XNOR2_X2 U9497 ( .A(n7010), .B(n9528), .ZN(n12936) );
  NAND2_X2 U9498 ( .A1(n9455), .A2(n9454), .ZN(n10011) );
  NAND2_X1 U9499 ( .A1(n7474), .A2(n7472), .ZN(n13077) );
  NAND4_X1 U9500 ( .A1(n7015), .A2(n9698), .A3(n7014), .A4(n9744), .ZN(n9445)
         );
  NAND2_X1 U9501 ( .A1(n7419), .A2(n7021), .ZN(n7016) );
  NAND2_X1 U9502 ( .A1(n9567), .A2(n9566), .ZN(n10828) );
  INV_X1 U9503 ( .A(n7025), .ZN(n12881) );
  NAND2_X1 U9504 ( .A1(n11352), .A2(n7041), .ZN(n7043) );
  NAND2_X1 U9505 ( .A1(n9261), .A2(n9260), .ZN(n11352) );
  NAND2_X1 U9506 ( .A1(n11636), .A2(n9265), .ZN(n11567) );
  AOI21_X1 U9507 ( .B1(n7543), .B2(n6703), .A(n7045), .ZN(n7044) );
  INV_X1 U9508 ( .A(n7543), .ZN(n7048) );
  XNOR2_X2 U9509 ( .A(n7055), .B(P2_IR_REG_29__SCAN_IN), .ZN(n12293) );
  NAND2_X1 U9510 ( .A1(n7535), .A2(n7533), .ZN(n13716) );
  NAND3_X1 U9511 ( .A1(n7522), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(n7519), .ZN(
        n7062) );
  OAI21_X2 U9512 ( .B1(n9139), .B2(n7066), .A(n7065), .ZN(n9148) );
  INV_X1 U9513 ( .A(n9148), .ZN(n9146) );
  NAND2_X1 U9514 ( .A1(n7904), .A2(n7069), .ZN(n7067) );
  NAND2_X1 U9515 ( .A1(n7067), .A2(n7068), .ZN(n7945) );
  OAI21_X1 U9516 ( .B1(n8026), .B2(n7079), .A(n7075), .ZN(n8096) );
  NAND2_X1 U9517 ( .A1(n7074), .A2(n7072), .ZN(n8098) );
  NAND2_X1 U9518 ( .A1(n8026), .A2(n7075), .ZN(n7074) );
  NAND2_X1 U9519 ( .A1(n8147), .A2(n6699), .ZN(n7081) );
  NAND2_X1 U9520 ( .A1(n8147), .A2(n8146), .ZN(n7087) );
  NAND2_X1 U9521 ( .A1(n9934), .A2(n7114), .ZN(n7113) );
  AOI21_X1 U9522 ( .B1(n9934), .B2(n9523), .A(n6825), .ZN(n9948) );
  NAND2_X1 U9523 ( .A1(n9934), .A2(n7119), .ZN(n7109) );
  NAND2_X1 U9524 ( .A1(n7113), .A2(n7111), .ZN(n12596) );
  NAND2_X1 U9525 ( .A1(n9468), .A2(n7130), .ZN(n7133) );
  AND2_X1 U9526 ( .A1(n9469), .A2(n9467), .ZN(n7130) );
  NAND2_X1 U9527 ( .A1(n7131), .A2(n9469), .ZN(n7132) );
  INV_X1 U9528 ( .A(n9554), .ZN(n7131) );
  NAND2_X1 U9529 ( .A1(n9875), .A2(n7138), .ZN(n7135) );
  NAND2_X1 U9530 ( .A1(n7135), .A2(n7136), .ZN(n9546) );
  NAND2_X1 U9531 ( .A1(n9487), .A2(n9486), .ZN(n9717) );
  NAND3_X1 U9532 ( .A1(n7156), .A2(n9531), .A3(n9519), .ZN(n9520) );
  INV_X1 U9533 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7157) );
  NAND2_X1 U9534 ( .A1(n14185), .A2(n14194), .ZN(n7158) );
  INV_X4 U9535 ( .A(n8848), .ZN(n10477) );
  XNOR2_X2 U9537 ( .A(n7172), .B(n7361), .ZN(n12264) );
  NAND2_X1 U9538 ( .A1(n14139), .A2(n7173), .ZN(n8948) );
  NAND2_X1 U9539 ( .A1(n7176), .A2(n8474), .ZN(n10268) );
  NAND2_X1 U9540 ( .A1(n10760), .A2(n9210), .ZN(n10856) );
  INV_X1 U9541 ( .A(n12116), .ZN(n9225) );
  OAI21_X1 U9542 ( .B1(n12166), .B2(n7197), .A(n7195), .ZN(n13704) );
  INV_X1 U9543 ( .A(n13625), .ZN(n7201) );
  OAI21_X1 U9544 ( .B1(n7201), .B2(n7205), .A(n7202), .ZN(n13573) );
  NAND2_X1 U9545 ( .A1(n7209), .A2(n7057), .ZN(n13834) );
  NAND2_X1 U9546 ( .A1(n7212), .A2(n7466), .ZN(n9607) );
  NAND2_X1 U9547 ( .A1(n10013), .A2(n6790), .ZN(n10018) );
  INV_X1 U9548 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7213) );
  NAND2_X1 U9549 ( .A1(n9962), .A2(n7214), .ZN(n10005) );
  INV_X1 U9550 ( .A(n12426), .ZN(n7223) );
  NAND2_X1 U9551 ( .A1(n12508), .A2(n7228), .ZN(n7226) );
  OAI211_X1 U9552 ( .C1(n12508), .C2(n7232), .A(n7229), .B(n7226), .ZN(n12493)
         );
  NAND2_X1 U9553 ( .A1(n12508), .A2(n6724), .ZN(n7233) );
  AOI21_X1 U9554 ( .B1(n12508), .B2(n12507), .A(n7227), .ZN(n12571) );
  INV_X1 U9555 ( .A(n12492), .ZN(n7238) );
  INV_X1 U9556 ( .A(n11995), .ZN(n7241) );
  NAND3_X1 U9557 ( .A1(n7243), .A2(n7244), .A3(n12049), .ZN(n12000) );
  INV_X1 U9558 ( .A(n11001), .ZN(n7253) );
  NAND2_X1 U9559 ( .A1(n7254), .A2(n7252), .ZN(n11006) );
  INV_X2 U9560 ( .A(n11046), .ZN(n12452) );
  NAND2_X2 U9561 ( .A1(n7254), .A2(n11004), .ZN(n11046) );
  AND2_X1 U9562 ( .A1(n7483), .A2(n9444), .ZN(n7482) );
  INV_X4 U9563 ( .A(n12452), .ZN(n12466) );
  NAND2_X2 U9564 ( .A1(n8538), .A2(n7256), .ZN(n15026) );
  NAND2_X1 U9565 ( .A1(n7257), .A2(n7258), .ZN(n11492) );
  NAND2_X1 U9566 ( .A1(n11370), .A2(n7260), .ZN(n7257) );
  NAND2_X1 U9567 ( .A1(n7263), .A2(n7265), .ZN(n11943) );
  NAND2_X1 U9568 ( .A1(n11752), .A2(n7264), .ZN(n7263) );
  NAND2_X1 U9569 ( .A1(n14120), .A2(n7270), .ZN(n7269) );
  INV_X1 U9570 ( .A(n8899), .ZN(n7280) );
  NAND2_X1 U9571 ( .A1(n9173), .A2(n7642), .ZN(n7281) );
  NAND2_X1 U9572 ( .A1(n14152), .A2(n7284), .ZN(n7282) );
  NAND2_X1 U9573 ( .A1(n7282), .A2(n7283), .ZN(n14122) );
  NAND2_X1 U9574 ( .A1(n9103), .A2(n7286), .ZN(n7291) );
  NAND2_X1 U9575 ( .A1(n7291), .A2(n7289), .ZN(n9107) );
  AND2_X1 U9576 ( .A1(n7291), .A2(n7288), .ZN(n9108) );
  NOR2_X1 U9577 ( .A1(n9104), .A2(n9105), .ZN(n7292) );
  NAND2_X1 U9578 ( .A1(n14973), .A2(n7296), .ZN(n7295) );
  NAND2_X1 U9579 ( .A1(n12128), .A2(n9183), .ZN(n7301) );
  NAND2_X1 U9580 ( .A1(n7301), .A2(n7299), .ZN(n8810) );
  INV_X1 U9581 ( .A(n8901), .ZN(n7303) );
  NAND3_X1 U9582 ( .A1(n8902), .A2(n8814), .A3(n8906), .ZN(n7305) );
  NAND3_X1 U9583 ( .A1(n9045), .A2(n9044), .A3(n6792), .ZN(n7309) );
  NAND2_X1 U9584 ( .A1(n7309), .A2(n7310), .ZN(n9050) );
  NAND2_X1 U9585 ( .A1(n7312), .A2(n7313), .ZN(n9116) );
  NAND3_X1 U9586 ( .A1(n9055), .A2(n9054), .A3(n6796), .ZN(n7314) );
  NAND2_X1 U9587 ( .A1(n7314), .A2(n7315), .ZN(n9063) );
  AND2_X4 U9588 ( .A1(n14384), .A2(n14386), .ZN(n8894) );
  XNOR2_X2 U9589 ( .A(n8544), .B(n8543), .ZN(n14384) );
  INV_X2 U9590 ( .A(n8548), .ZN(n14386) );
  NAND3_X1 U9591 ( .A1(n9026), .A2(n9025), .A3(n6791), .ZN(n7318) );
  NAND2_X1 U9592 ( .A1(n7318), .A2(n7319), .ZN(n9031) );
  NAND3_X1 U9593 ( .A1(n9036), .A2(n9035), .A3(n6797), .ZN(n7321) );
  NAND2_X1 U9594 ( .A1(n7321), .A2(n7322), .ZN(n9043) );
  OAI22_X2 U9595 ( .A1(n9873), .A2(n7325), .B1(n7324), .B2(n7327), .ZN(n13032)
         );
  NOR2_X1 U9596 ( .A1(n10011), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n9526) );
  NOR2_X2 U9597 ( .A1(n10011), .A2(n7335), .ZN(n7334) );
  NAND2_X1 U9598 ( .A1(n12074), .A2(n7339), .ZN(n7338) );
  INV_X1 U9599 ( .A(n7348), .ZN(n12276) );
  NAND2_X2 U9600 ( .A1(n9827), .A2(n7354), .ZN(n13098) );
  NAND3_X1 U9601 ( .A1(n15006), .A2(n15004), .A3(n6803), .ZN(n7379) );
  INV_X1 U9602 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7384) );
  OAI22_X1 U9603 ( .A1(n14786), .A2(n7386), .B1(n6697), .B2(n14789), .ZN(
        n14788) );
  INV_X1 U9604 ( .A(n14789), .ZN(n7387) );
  INV_X1 U9605 ( .A(n7390), .ZN(n14785) );
  INV_X1 U9606 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7389) );
  NAND2_X1 U9607 ( .A1(n10963), .A2(n7399), .ZN(n10821) );
  OR2_X1 U9608 ( .A1(n10820), .A2(n7400), .ZN(n7399) );
  NAND2_X1 U9609 ( .A1(n10820), .A2(n7400), .ZN(n10963) );
  OAI21_X1 U9610 ( .B1(n10945), .B2(P3_REG2_REG_2__SCAN_IN), .A(n7401), .ZN(
        n7400) );
  NAND2_X1 U9611 ( .A1(n10945), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7401) );
  INV_X1 U9612 ( .A(n12847), .ZN(n12869) );
  NAND2_X1 U9613 ( .A1(n12880), .A2(n7402), .ZN(n12872) );
  NOR2_X1 U9614 ( .A1(n12847), .A2(n7403), .ZN(n12871) );
  INV_X1 U9615 ( .A(n12870), .ZN(n7403) );
  NAND2_X1 U9616 ( .A1(n11270), .A2(n7408), .ZN(n7404) );
  NAND2_X1 U9617 ( .A1(n7406), .A2(n7404), .ZN(n11463) );
  NAND3_X1 U9618 ( .A1(n7407), .A2(n11268), .A3(n6714), .ZN(n7406) );
  NAND2_X1 U9619 ( .A1(n7410), .A2(n7412), .ZN(n11952) );
  NAND3_X1 U9620 ( .A1(n7414), .A2(n11652), .A3(n7413), .ZN(n7412) );
  INV_X1 U9621 ( .A(n11464), .ZN(n7416) );
  NAND2_X1 U9622 ( .A1(n7414), .A2(n11652), .ZN(n11465) );
  NAND2_X1 U9623 ( .A1(n7416), .A2(n11667), .ZN(n7414) );
  INV_X1 U9624 ( .A(n7418), .ZN(n12844) );
  INV_X1 U9625 ( .A(n11112), .ZN(n7425) );
  INV_X1 U9626 ( .A(n7426), .ZN(n11110) );
  NAND2_X1 U9627 ( .A1(n8542), .A2(n8541), .ZN(n8545) );
  NAND2_X1 U9628 ( .A1(n8542), .A2(n7443), .ZN(n14377) );
  NAND2_X1 U9629 ( .A1(n13922), .A2(n7444), .ZN(n13877) );
  NAND2_X1 U9630 ( .A1(n7446), .A2(n7445), .ZN(n10217) );
  NAND2_X1 U9631 ( .A1(n15469), .A2(n7455), .ZN(n7453) );
  NAND2_X1 U9632 ( .A1(n13150), .A2(n7468), .ZN(n7467) );
  NAND2_X1 U9633 ( .A1(n9992), .A2(n7479), .ZN(n7477) );
  NAND2_X1 U9634 ( .A1(n9989), .A2(n7481), .ZN(n13109) );
  NOR2_X1 U9635 ( .A1(n9445), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U9636 ( .A1(n9746), .A2(n9453), .ZN(n10009) );
  NOR2_X2 U9637 ( .A1(n13541), .A2(n13521), .ZN(n13515) );
  NOR2_X1 U9638 ( .A1(n13642), .A2(n13759), .ZN(n13630) );
  NOR2_X1 U9639 ( .A1(n8124), .A2(n7667), .ZN(n7493) );
  INV_X1 U9640 ( .A(n8124), .ZN(n7495) );
  NOR2_X2 U9641 ( .A1(n11810), .A2(n11917), .ZN(n12037) );
  NOR2_X2 U9642 ( .A1(n12171), .A2(n13798), .ZN(n7498) );
  NOR2_X2 U9643 ( .A1(n12120), .A2(n13811), .ZN(n7500) );
  NAND2_X2 U9644 ( .A1(n7502), .A2(n8411), .ZN(n13521) );
  NAND3_X1 U9645 ( .A1(n8299), .A2(n8302), .A3(n7507), .ZN(n7504) );
  NAND2_X1 U9646 ( .A1(n8502), .A2(n8501), .ZN(n7516) );
  OAI211_X1 U9647 ( .C1(n7517), .C2(n12009), .A(n7516), .B(n8521), .ZN(
        P2_U3328) );
  OAI21_X2 U9648 ( .B1(n8365), .B2(n12304), .A(n8368), .ZN(n8423) );
  NAND2_X1 U9649 ( .A1(n7525), .A2(n10253), .ZN(n9251) );
  XNOR2_X1 U9650 ( .A(n7525), .B(n10253), .ZN(n15324) );
  NAND2_X1 U9651 ( .A1(n10835), .A2(n9257), .ZN(n9259) );
  NAND2_X1 U9652 ( .A1(n10853), .A2(n9255), .ZN(n7526) );
  OR2_X2 U9653 ( .A1(n13691), .A2(n9280), .ZN(n7543) );
  NAND3_X1 U9654 ( .A1(n7579), .A2(n7589), .A3(n7544), .ZN(n13727) );
  XNOR2_X2 U9655 ( .A(n9295), .B(n9294), .ZN(n13528) );
  XNOR2_X1 U9657 ( .A(n10132), .B(n10130), .ZN(n13418) );
  NAND2_X1 U9658 ( .A1(n10485), .A2(n10066), .ZN(n7547) );
  NAND2_X1 U9659 ( .A1(n10063), .A2(n10656), .ZN(n10485) );
  XNOR2_X1 U9660 ( .A(n10064), .B(n10065), .ZN(n10486) );
  NAND2_X1 U9661 ( .A1(n10115), .A2(n11884), .ZN(n7551) );
  NAND2_X1 U9662 ( .A1(n10184), .A2(n7553), .ZN(n7552) );
  NOR2_X1 U9663 ( .A1(n10184), .A2(n10183), .ZN(n13314) );
  OAI211_X1 U9664 ( .C1(n10184), .C2(n7554), .A(n13324), .B(n7552), .ZN(
        P2_U3192) );
  XNOR2_X2 U9665 ( .A(n7568), .B(n7567), .ZN(n13294) );
  INV_X1 U9666 ( .A(n10166), .ZN(n7567) );
  NAND2_X1 U9667 ( .A1(n10099), .A2(n11245), .ZN(n11259) );
  OAI211_X1 U9668 ( .C1(n7572), .C2(n13326), .A(n13325), .B(n10187), .ZN(
        n13330) );
  NAND2_X1 U9669 ( .A1(n7685), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U9670 ( .A1(n11806), .A2(n11807), .ZN(n7578) );
  NAND4_X1 U9671 ( .A1(n7586), .A2(n7584), .A3(n7582), .A4(n7580), .ZN(
        P2_U3528) );
  NAND2_X1 U9672 ( .A1(n13528), .A2(n7581), .ZN(n7580) );
  XNOR2_X2 U9673 ( .A(n9241), .B(n9240), .ZN(n7588) );
  INV_X1 U9674 ( .A(n9245), .ZN(n7591) );
  AND2_X2 U9675 ( .A1(n7593), .A2(n9235), .ZN(n13625) );
  NAND2_X1 U9676 ( .A1(n10856), .A2(n10855), .ZN(n10854) );
  NAND2_X1 U9677 ( .A1(n7597), .A2(n9255), .ZN(n7595) );
  INV_X1 U9678 ( .A(n7597), .ZN(n7596) );
  OAI211_X2 U9679 ( .C1(n8030), .C2(n9466), .A(n7600), .B(n7599), .ZN(n10489)
         );
  AND2_X1 U9680 ( .A1(n13572), .A2(n9238), .ZN(n13550) );
  NAND2_X1 U9681 ( .A1(n13572), .A2(n6787), .ZN(n7602) );
  AND2_X1 U9682 ( .A1(n13734), .A2(n9239), .ZN(n7605) );
  OAI21_X1 U9683 ( .B1(n8459), .B2(n8463), .A(n8462), .ZN(n8502) );
  AOI21_X1 U9684 ( .B1(n6692), .B2(n6710), .A(n7608), .ZN(n8225) );
  NAND3_X1 U9685 ( .A1(n7657), .A2(n8145), .A3(n6795), .ZN(n7613) );
  NAND2_X1 U9686 ( .A1(n7615), .A2(n7616), .ZN(n8340) );
  NAND2_X1 U9687 ( .A1(n8319), .A2(n7618), .ZN(n7615) );
  NAND3_X1 U9688 ( .A1(n7940), .A2(n7939), .A3(n7620), .ZN(n7621) );
  NAND2_X1 U9689 ( .A1(n7966), .A2(n7965), .ZN(n7620) );
  NAND2_X1 U9690 ( .A1(n7621), .A2(n6799), .ZN(n7993) );
  INV_X1 U9691 ( .A(n8048), .ZN(n7624) );
  NAND2_X1 U9692 ( .A1(n7636), .A2(n8116), .ZN(n7635) );
  NAND3_X1 U9693 ( .A1(n7658), .A2(n8228), .A3(n6806), .ZN(n7639) );
  NAND2_X1 U9694 ( .A1(n7639), .A2(n6800), .ZN(n8275) );
  INV_X1 U9695 ( .A(n8253), .ZN(n7641) );
  OAI211_X2 U9696 ( .C1(n12535), .C2(n12463), .A(n12462), .B(n12461), .ZN(
        n12508) );
  NOR2_X1 U9697 ( .A1(n12969), .A2(n10001), .ZN(n10053) );
  AND2_X1 U9698 ( .A1(n8473), .A2(n8474), .ZN(n10275) );
  NAND2_X1 U9699 ( .A1(n13077), .A2(n9990), .ZN(n13066) );
  XNOR2_X1 U9700 ( .A(n10217), .B(n10223), .ZN(n10219) );
  OAI21_X1 U9701 ( .B1(n9299), .B2(n13504), .A(n9242), .ZN(n13586) );
  INV_X1 U9702 ( .A(n9299), .ZN(n11829) );
  INV_X1 U9703 ( .A(n14384), .ZN(n8549) );
  NAND2_X1 U9704 ( .A1(n10184), .A2(n10183), .ZN(n10188) );
  XNOR2_X1 U9705 ( .A(n12620), .B(n7154), .ZN(n12964) );
  OR2_X1 U9706 ( .A1(n7690), .A2(n7678), .ZN(n7691) );
  NOR2_X2 U9707 ( .A1(n11484), .A2(n11428), .ZN(n11643) );
  AOI22_X1 U9708 ( .A1(n8475), .A2(n8437), .B1(n7917), .B2(n10067), .ZN(n7769)
         );
  XNOR2_X1 U9709 ( .A(n7799), .B(n7797), .ZN(n8605) );
  OR2_X1 U9710 ( .A1(n7874), .A2(n7873), .ZN(n7660) );
  NAND2_X1 U9711 ( .A1(n8463), .A2(n8461), .ZN(n8462) );
  NOR2_X1 U9712 ( .A1(n10054), .A2(n13285), .ZN(n10055) );
  INV_X2 U9713 ( .A(n15568), .ZN(n15570) );
  AND2_X1 U9714 ( .A1(n10052), .A2(n10051), .ZN(n15568) );
  NOR2_X1 U9715 ( .A1(n10054), .A2(n13232), .ZN(n10040) );
  AND2_X2 U9716 ( .A1(n10799), .A2(n10039), .ZN(n15585) );
  AND2_X1 U9717 ( .A1(n9172), .A2(n11078), .ZN(n7642) );
  CLKBUF_X3 U9718 ( .A(n9070), .Z(n9167) );
  AND2_X1 U9719 ( .A1(n11142), .A2(n9016), .ZN(n7643) );
  AND2_X1 U9720 ( .A1(n11191), .A2(n9011), .ZN(n7644) );
  INV_X1 U9721 ( .A(n12458), .ZN(n13247) );
  OR3_X1 U9722 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n10827), .ZN(n7645) );
  AND2_X1 U9723 ( .A1(n8450), .A2(n8449), .ZN(n7646) );
  AND4_X1 U9724 ( .A1(n8619), .A2(n8639), .A3(n8643), .A4(n8526), .ZN(n7647)
         );
  XNOR2_X1 U9725 ( .A(n15316), .B(n13316), .ZN(n10064) );
  AND2_X1 U9726 ( .A1(n12222), .A2(n12221), .ZN(n7649) );
  AND2_X1 U9727 ( .A1(n12978), .A2(n7653), .ZN(n7650) );
  OR2_X1 U9728 ( .A1(n10807), .A2(n10809), .ZN(n7651) );
  OR2_X1 U9729 ( .A1(n9591), .A2(n12604), .ZN(n7652) );
  OR2_X1 U9730 ( .A1(n12977), .A2(n15507), .ZN(n7653) );
  AND2_X1 U9731 ( .A1(n14278), .A2(n15198), .ZN(n7654) );
  INV_X1 U9732 ( .A(n12996), .ZN(n9927) );
  INV_X1 U9733 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9659) );
  OR2_X1 U9734 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11091), .ZN(n7655) );
  AND2_X1 U9735 ( .A1(n9944), .A2(n9943), .ZN(n12986) );
  INV_X1 U9736 ( .A(n12363), .ZN(n11511) );
  AND2_X1 U9737 ( .A1(n9911), .A2(n9910), .ZN(n12511) );
  INV_X1 U9738 ( .A(n12511), .ZN(n9912) );
  NAND3_X1 U9739 ( .A1(n9094), .A2(n9093), .A3(n14235), .ZN(n7656) );
  OR2_X1 U9740 ( .A1(n8144), .A2(n8143), .ZN(n7657) );
  OR2_X1 U9741 ( .A1(n8227), .A2(n8226), .ZN(n7658) );
  NAND2_X1 U9742 ( .A1(n12659), .A2(n12664), .ZN(n9979) );
  INV_X1 U9743 ( .A(n13417), .ZN(n10187) );
  AND2_X1 U9744 ( .A1(n9732), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7659) );
  INV_X1 U9745 ( .A(n14262), .ZN(n10210) );
  AND3_X1 U9746 ( .A1(n7714), .A2(n10655), .A3(n7713), .ZN(n7719) );
  OR2_X1 U9747 ( .A1(n7770), .A2(n7769), .ZN(n7791) );
  AOI21_X1 U9748 ( .B1(n7660), .B2(n7896), .A(n7895), .ZN(n7898) );
  NAND2_X1 U9749 ( .A1(n8113), .A2(n8112), .ZN(n8116) );
  NAND2_X1 U9750 ( .A1(n8280), .A2(n8279), .ZN(n8298) );
  INV_X1 U9751 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9446) );
  INV_X1 U9752 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8526) );
  INV_X1 U9753 ( .A(n12986), .ZN(n9945) );
  INV_X1 U9754 ( .A(n9834), .ZN(n9433) );
  AND2_X1 U9755 ( .A1(n9452), .A2(n6778), .ZN(n9453) );
  INV_X1 U9756 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7676) );
  OAI21_X1 U9757 ( .B1(n9146), .B2(n9145), .A(n9144), .ZN(n9147) );
  INV_X1 U9758 ( .A(n15504), .ZN(n10789) );
  NAND2_X1 U9759 ( .A1(n12458), .A2(n9912), .ZN(n9913) );
  AND2_X1 U9760 ( .A1(n9433), .A2(n12564), .ZN(n9853) );
  INV_X1 U9761 ( .A(n12676), .ZN(n9627) );
  INV_X1 U9762 ( .A(n12701), .ZN(n9986) );
  INV_X1 U9763 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9780) );
  INV_X1 U9764 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9481) );
  AND2_X1 U9765 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n7956) );
  INV_X1 U9766 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11215) );
  INV_X1 U9767 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8012) );
  INV_X1 U9768 ( .A(n10253), .ZN(n10251) );
  INV_X1 U9769 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8497) );
  NOR2_X1 U9770 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7669) );
  INV_X1 U9771 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8658) );
  INV_X1 U9772 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8619) );
  INV_X1 U9773 ( .A(n9903), .ZN(n9437) );
  OR2_X1 U9774 ( .A1(n9769), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9790) );
  NOR2_X1 U9775 ( .A1(n12616), .A2(n12957), .ZN(n9974) );
  INV_X1 U9776 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n12564) );
  NAND2_X1 U9777 ( .A1(n9431), .A2(n9430), .ZN(n9805) );
  INV_X1 U9778 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U9779 ( .A1(n10018), .A2(n10017), .ZN(n11001) );
  INV_X1 U9780 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9454) );
  AND2_X1 U9781 ( .A1(n9501), .A2(n9500), .ZN(n9799) );
  AND2_X1 U9782 ( .A1(n10467), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9489) );
  INV_X1 U9783 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U9784 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8289), .ZN(n8327) );
  OR2_X1 U9785 ( .A1(n8174), .A2(n8173), .ZN(n8197) );
  OR2_X1 U9786 ( .A1(n7981), .A2(n11215), .ZN(n8013) );
  INV_X1 U9787 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11630) );
  INV_X1 U9788 ( .A(n15221), .ZN(n10389) );
  NOR2_X1 U9789 ( .A1(n14574), .A2(n8241), .ZN(n8264) );
  NAND2_X1 U9790 ( .A1(n8498), .A2(n8497), .ZN(n8503) );
  INV_X1 U9791 ( .A(n11767), .ZN(n11768) );
  INV_X1 U9792 ( .A(n13880), .ZN(n12359) );
  INV_X1 U9793 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8688) );
  OAI21_X1 U9794 ( .B1(n9161), .B2(n9160), .A(n9159), .ZN(n9166) );
  OR2_X1 U9795 ( .A1(n8803), .A2(n13940), .ZN(n8818) );
  OR2_X1 U9796 ( .A1(n9894), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9903) );
  NAND2_X1 U9797 ( .A1(n9674), .A2(n11700), .ZN(n9690) );
  AND2_X1 U9798 ( .A1(n9660), .A2(n9659), .ZN(n9674) );
  NAND2_X1 U9799 ( .A1(n9435), .A2(n12501), .ZN(n9892) );
  INV_X1 U9800 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12528) );
  INV_X1 U9801 ( .A(n12698), .ZN(n11703) );
  OR2_X1 U9802 ( .A1(n9892), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U9803 ( .A1(n10998), .A2(n10997), .ZN(n12576) );
  INV_X1 U9804 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n14661) );
  INV_X1 U9805 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11700) );
  AND2_X1 U9806 ( .A1(n10815), .A2(n10813), .ZN(n10819) );
  AND3_X1 U9807 ( .A1(n10797), .A2(n10796), .A3(n10795), .ZN(n10798) );
  OR3_X1 U9808 ( .A1(n10792), .A2(n10793), .A3(n10920), .ZN(n10037) );
  INV_X1 U9809 ( .A(n9591), .ZN(n9850) );
  AND2_X1 U9810 ( .A1(n10047), .A2(n12622), .ZN(n15490) );
  AND3_X1 U9811 ( .A1(n10792), .A2(n11001), .A3(n10049), .ZN(n10998) );
  INV_X1 U9812 ( .A(SI_14_), .ZN(n14777) );
  OR2_X1 U9813 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  NAND2_X1 U9814 ( .A1(n8214), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8241) );
  INV_X1 U9815 ( .A(n11800), .ZN(n10108) );
  INV_X1 U9816 ( .A(n13422), .ZN(n13390) );
  INV_X1 U9817 ( .A(n13421), .ZN(n13389) );
  OR2_X1 U9818 ( .A1(n8083), .A2(n15257), .ZN(n8108) );
  INV_X1 U9819 ( .A(n8387), .ZN(n8352) );
  NOR2_X1 U9820 ( .A1(n8197), .A2(n13379), .ZN(n8214) );
  NAND2_X1 U9821 ( .A1(n8153), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8174) );
  OR2_X1 U9822 ( .A1(n11212), .A2(n11211), .ZN(n11405) );
  INV_X1 U9823 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n15257) );
  OR2_X1 U9824 ( .A1(n8429), .A2(n13321), .ZN(n13523) );
  INV_X1 U9825 ( .A(n13441), .ZN(n12119) );
  INV_X1 U9826 ( .A(n13586), .ZN(n13676) );
  OR3_X1 U9827 ( .A1(n10195), .A2(P2_U3088), .A3(n9316), .ZN(n10257) );
  NOR2_X1 U9828 ( .A1(n7676), .A2(n7678), .ZN(n7701) );
  NOR2_X1 U9829 ( .A1(n8033), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U9830 ( .A1(n11870), .A2(n11869), .ZN(n11871) );
  AND3_X1 U9831 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8648) );
  AND2_X1 U9832 ( .A1(n8827), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8838) );
  OR2_X1 U9833 ( .A1(n13949), .A2(n14265), .ZN(n14910) );
  INV_X1 U9834 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8766) );
  AND2_X1 U9835 ( .A1(n8780), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8794) );
  INV_X1 U9836 ( .A(n10236), .ZN(n10478) );
  INV_X1 U9837 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n13940) );
  OR2_X1 U9838 ( .A1(n11120), .A2(n11942), .ZN(n11758) );
  AND2_X1 U9839 ( .A1(n8097), .A2(n8074), .ZN(n8095) );
  AND2_X1 U9840 ( .A1(n8025), .A2(n8004), .ZN(n8023) );
  XNOR2_X1 U9841 ( .A(n7855), .B(n7853), .ZN(n8626) );
  NOR2_X1 U9842 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9388), .ZN(n9338) );
  AOI21_X1 U9843 ( .B1(n14696), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n9347), .ZN(
        n9409) );
  AOI22_X1 U9844 ( .A1(n9357), .A2(n9356), .B1(P1_ADDR_REG_14__SCAN_IN), .B2(
        n9355), .ZN(n9368) );
  OR2_X1 U9845 ( .A1(n9629), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9644) );
  INV_X1 U9846 ( .A(n12581), .ZN(n12590) );
  AND3_X1 U9847 ( .A1(n9885), .A2(n9884), .A3(n9883), .ZN(n13042) );
  INV_X1 U9848 ( .A(n15454), .ZN(n14825) );
  AND2_X1 U9849 ( .A1(P3_U3897), .A2(n9968), .ZN(n12954) );
  INV_X1 U9850 ( .A(n13035), .ZN(n13188) );
  INV_X1 U9851 ( .A(n13137), .ZN(n14861) );
  INV_X1 U9852 ( .A(n15517), .ZN(n15479) );
  NOR2_X1 U9853 ( .A1(n15585), .A2(n10041), .ZN(n10042) );
  AND2_X1 U9854 ( .A1(n10046), .A2(n10031), .ZN(n10799) );
  OR2_X1 U9855 ( .A1(n15495), .A2(n15566), .ZN(n14883) );
  OR2_X1 U9856 ( .A1(n10935), .A2(n10930), .ZN(n10052) );
  INV_X1 U9857 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n10006) );
  INV_X1 U9858 ( .A(n9962), .ZN(n9966) );
  INV_X1 U9859 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9816) );
  INV_X1 U9860 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9651) );
  INV_X1 U9861 ( .A(n12009), .ZN(n8501) );
  OR2_X1 U9862 ( .A1(n6672), .A2(n13568), .ZN(n8333) );
  OR2_X1 U9863 ( .A1(n6670), .A2(n7811), .ZN(n7816) );
  OR2_X1 U9864 ( .A1(n10369), .A2(n10370), .ZN(n15271) );
  INV_X1 U9865 ( .A(n15236), .ZN(n15281) );
  INV_X1 U9866 ( .A(n9290), .ZN(n13574) );
  INV_X1 U9867 ( .A(n13676), .ZN(n13705) );
  NAND2_X1 U9868 ( .A1(n10696), .A2(n10191), .ZN(n15342) );
  INV_X1 U9869 ( .A(n15339), .ZN(n15360) );
  NAND2_X1 U9870 ( .A1(n10061), .A2(n13756), .ZN(n15339) );
  OR2_X1 U9871 ( .A1(n10257), .A2(n9319), .ZN(n11104) );
  AND2_X1 U9872 ( .A1(n9303), .A2(n9320), .ZN(n15302) );
  XNOR2_X1 U9873 ( .A(n8504), .B(P2_IR_REG_24__SCAN_IN), .ZN(n12187) );
  AND2_X1 U9874 ( .A1(n8080), .A2(n8102), .ZN(n15263) );
  INV_X1 U9875 ( .A(n13852), .ZN(n12008) );
  OR2_X1 U9876 ( .A1(n10243), .A2(n10610), .ZN(n13949) );
  AND2_X1 U9877 ( .A1(n8833), .A2(n8832), .ZN(n14221) );
  OR2_X1 U9878 ( .A1(n15029), .A2(n10509), .ZN(n15056) );
  OR3_X1 U9879 ( .A1(n11931), .A2(n15052), .A3(n11930), .ZN(n12059) );
  AOI22_X1 U9880 ( .A1(n14070), .A2(n14812), .B1(n14069), .B2(n14979), .ZN(
        n14074) );
  NAND2_X1 U9881 ( .A1(n8859), .A2(n8858), .ZN(n14152) );
  OR2_X1 U9882 ( .A1(n15118), .A2(n11081), .ZN(n15107) );
  INV_X1 U9883 ( .A(n14816), .ZN(n15113) );
  INV_X1 U9884 ( .A(n15107), .ZN(n14255) );
  INV_X1 U9885 ( .A(n15198), .ZN(n14359) );
  NAND2_X1 U9886 ( .A1(n11758), .A2(n14345), .ZN(n15198) );
  AND3_X1 U9887 ( .A1(n8998), .A2(n8997), .A3(n8996), .ZN(n11065) );
  INV_X1 U9888 ( .A(n9196), .ZN(n10479) );
  INV_X1 U9889 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8906) );
  AND2_X1 U9890 ( .A1(n8763), .A2(n8775), .ZN(n11928) );
  AND2_X1 U9891 ( .A1(n10815), .A2(n10814), .ZN(n15460) );
  INV_X1 U9892 ( .A(n12578), .ZN(n12588) );
  AND2_X1 U9893 ( .A1(n10936), .A2(n15479), .ZN(n12581) );
  NAND2_X1 U9894 ( .A1(n9926), .A2(n9925), .ZN(n12996) );
  OR2_X1 U9895 ( .A1(n10922), .A2(n10436), .ZN(n12816) );
  INV_X1 U9896 ( .A(n12954), .ZN(n15456) );
  INV_X1 U9897 ( .A(n14832), .ZN(n15467) );
  AND2_X1 U9898 ( .A1(n13103), .A2(n13102), .ZN(n13210) );
  INV_X1 U9899 ( .A(n15585), .ZN(n15583) );
  INV_X1 U9900 ( .A(n12470), .ZN(n13174) );
  AND2_X1 U9901 ( .A1(n15557), .A2(n15556), .ZN(n15581) );
  NAND2_X1 U9902 ( .A1(n10472), .A2(n10471), .ZN(n10481) );
  AND2_X1 U9903 ( .A1(n10918), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10471) );
  INV_X1 U9904 ( .A(n10014), .ZN(n11976) );
  INV_X1 U9905 ( .A(SI_21_), .ZN(n11206) );
  INV_X1 U9906 ( .A(SI_17_), .ZN(n10579) );
  INV_X1 U9907 ( .A(n11297), .ZN(n15397) );
  INV_X1 U9908 ( .A(n10201), .ZN(n10202) );
  INV_X1 U9909 ( .A(n13425), .ZN(n13369) );
  OR2_X1 U9910 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  NAND2_X1 U9911 ( .A1(n8249), .A2(n8248), .ZN(n13432) );
  INV_X1 U9912 ( .A(n15275), .ZN(n15269) );
  AND2_X1 U9913 ( .A1(n10260), .A2(n13683), .ZN(n15301) );
  INV_X1 U9914 ( .A(n13689), .ZN(n15290) );
  OR2_X1 U9915 ( .A1(n15301), .A2(n10852), .ZN(n15293) );
  OR2_X1 U9916 ( .A1(n15301), .A2(n10851), .ZN(n13618) );
  OR2_X1 U9917 ( .A1(n11104), .A2(n15310), .ZN(n15371) );
  OR2_X1 U9918 ( .A1(n15364), .A2(n9324), .ZN(n9325) );
  OR2_X1 U9919 ( .A1(n11104), .A2(n9323), .ZN(n15362) );
  INV_X2 U9920 ( .A(n15362), .ZN(n15364) );
  NOR2_X1 U9921 ( .A1(n15311), .A2(n15302), .ZN(n15307) );
  INV_X1 U9922 ( .A(n15307), .ZN(n15308) );
  INV_X1 U9923 ( .A(n7709), .ZN(n11835) );
  INV_X1 U9924 ( .A(n15263), .ZN(n13468) );
  INV_X1 U9925 ( .A(n12008), .ZN(n13844) );
  INV_X1 U9926 ( .A(n14229), .ZN(n14335) );
  OR2_X1 U9927 ( .A1(n13949), .A2(n14220), .ZN(n14909) );
  INV_X1 U9928 ( .A(n14921), .ZN(n14958) );
  INV_X1 U9929 ( .A(n9003), .ZN(n14070) );
  OAI21_X1 U9930 ( .B1(n14188), .B2(n8893), .A(n8844), .ZN(n14175) );
  INV_X1 U9931 ( .A(n12310), .ZN(n14955) );
  OR2_X1 U9932 ( .A1(n15029), .A2(n10715), .ZN(n15054) );
  OR2_X1 U9933 ( .A1(n15029), .A2(n10508), .ZN(n12065) );
  OR2_X1 U9934 ( .A1(n12255), .A2(n11942), .ZN(n14816) );
  INV_X1 U9935 ( .A(n14804), .ZN(n15105) );
  INV_X1 U9936 ( .A(n14804), .ZN(n14251) );
  INV_X1 U9937 ( .A(n14804), .ZN(n15118) );
  OR2_X1 U9938 ( .A1(n15118), .A2(n11069), .ZN(n11765) );
  INV_X1 U9939 ( .A(n15215), .ZN(n15213) );
  NAND2_X1 U9940 ( .A1(n14284), .A2(n14283), .ZN(n14363) );
  INV_X1 U9941 ( .A(n15201), .ZN(n15199) );
  AND2_X2 U9942 ( .A1(n8999), .A2(n11065), .ZN(n15201) );
  AND2_X1 U9943 ( .A1(n8976), .A2(n14394), .ZN(n10402) );
  INV_X1 U9944 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10618) );
  INV_X1 U9945 ( .A(n14758), .ZN(n14383) );
  INV_X2 U9946 ( .A(n12816), .ZN(P3_U3897) );
  NAND2_X1 U9947 ( .A1(n9326), .A2(n9325), .ZN(P2_U3496) );
  NOR2_X1 U9948 ( .A1(n10207), .A2(n10204), .ZN(P1_U4016) );
  NOR2_X1 U9949 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7664) );
  NOR2_X2 U9950 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7662) );
  NOR2_X2 U9951 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7661) );
  NAND4_X1 U9952 ( .A1(n7664), .A2(n7663), .A3(n7662), .A4(n7661), .ZN(n8124)
         );
  NAND3_X1 U9953 ( .A1(n7666), .A2(n8127), .A3(n7665), .ZN(n7667) );
  NOR2_X2 U9954 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7727) );
  NOR2_X1 U9955 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n7673) );
  NOR2_X1 U9956 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n7672) );
  NOR2_X1 U9957 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n7671) );
  NAND2_X1 U9958 ( .A1(n8505), .A2(n7674), .ZN(n7675) );
  INV_X1 U9959 ( .A(n7680), .ZN(n7682) );
  INV_X1 U9960 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7678) );
  INV_X1 U9961 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10660) );
  NAND2_X2 U9962 ( .A1(n12293), .A2(n12273), .ZN(n8428) );
  INV_X1 U9963 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7681) );
  INV_X1 U9964 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10442) );
  OR2_X1 U9965 ( .A1(n7836), .A2(n10442), .ZN(n7714) );
  NAND4_X1 U9966 ( .A1(n7717), .A2(n7716), .A3(n7714), .A4(n7713), .ZN(n8473)
         );
  INV_X1 U9967 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U9968 ( .A1(n7690), .A2(n7687), .ZN(n8496) );
  NAND2_X1 U9969 ( .A1(n9299), .A2(n10262), .ZN(n7695) );
  NAND2_X1 U9970 ( .A1(n7692), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7694) );
  XNOR2_X1 U9971 ( .A(n7694), .B(n7693), .ZN(n7708) );
  INV_X1 U9972 ( .A(n7696), .ZN(n7699) );
  NOR2_X1 U9973 ( .A1(n7696), .A2(n7700), .ZN(n7703) );
  INV_X1 U9974 ( .A(SI_0_), .ZN(n10287) );
  INV_X1 U9975 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9465) );
  OAI21_X1 U9976 ( .B1(n10302), .B2(n10287), .A(n9465), .ZN(n7705) );
  INV_X1 U9977 ( .A(n7732), .ZN(n7730) );
  AND2_X1 U9978 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U9979 ( .A1(n7730), .A2(n7704), .ZN(n7735) );
  AND2_X1 U9980 ( .A1(n7705), .A2(n7735), .ZN(n13853) );
  NAND2_X1 U9981 ( .A1(n10362), .A2(n13853), .ZN(n7706) );
  NAND2_X1 U9982 ( .A1(n7715), .A2(n8474), .ZN(n7710) );
  AND2_X1 U9983 ( .A1(n7710), .A2(n7845), .ZN(n7712) );
  NOR2_X1 U9984 ( .A1(n10655), .A2(n7845), .ZN(n7711) );
  AOI21_X1 U9985 ( .B1(n8473), .B2(n7712), .A(n7711), .ZN(n7721) );
  INV_X1 U9986 ( .A(n7715), .ZN(n7718) );
  NAND4_X1 U9987 ( .A1(n7719), .A2(n7718), .A3(n7717), .A4(n7716), .ZN(n7720)
         );
  NAND2_X1 U9988 ( .A1(n7721), .A2(n7720), .ZN(n7742) );
  INV_X1 U9989 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10356) );
  INV_X1 U9990 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10279) );
  OR2_X1 U9991 ( .A1(n8431), .A2(n10279), .ZN(n7724) );
  NAND2_X1 U9992 ( .A1(n7929), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7723) );
  INV_X1 U9993 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10373) );
  OR2_X1 U9994 ( .A1(n7836), .A2(n10373), .ZN(n7722) );
  NAND2_X1 U9995 ( .A1(n10062), .A2(n8437), .ZN(n7737) );
  NAND2_X1 U9996 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7726) );
  MUX2_X1 U9997 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7726), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7729) );
  INV_X1 U9998 ( .A(n7752), .ZN(n7728) );
  NAND2_X1 U9999 ( .A1(n7729), .A2(n7728), .ZN(n10374) );
  INV_X1 U10000 ( .A(n7730), .ZN(n7731) );
  NAND2_X1 U10001 ( .A1(n7732), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7733) );
  INV_X1 U10002 ( .A(SI_1_), .ZN(n10294) );
  AND2_X1 U10003 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7734) );
  NAND2_X1 U10004 ( .A1(n7759), .A2(n7734), .ZN(n8590) );
  NAND2_X1 U10005 ( .A1(n7735), .A2(n8590), .ZN(n7755) );
  XNOR2_X1 U10006 ( .A(n7755), .B(n7754), .ZN(n10304) );
  CLKBUF_X3 U10007 ( .A(n7759), .Z(n10302) );
  INV_X1 U10008 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U10009 ( .A1(n10489), .A2(n7843), .ZN(n7736) );
  NAND2_X1 U10010 ( .A1(n8478), .A2(n7917), .ZN(n7739) );
  NAND2_X1 U10011 ( .A1(n10489), .A2(n8437), .ZN(n7738) );
  NAND2_X1 U10012 ( .A1(n7739), .A2(n7738), .ZN(n7740) );
  NAND2_X1 U10013 ( .A1(n7741), .A2(n7740), .ZN(n7768) );
  INV_X1 U10014 ( .A(n7742), .ZN(n7744) );
  NAND2_X1 U10015 ( .A1(n7744), .A2(n7743), .ZN(n7767) );
  NAND2_X1 U10016 ( .A1(n7929), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7748) );
  INV_X1 U10017 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10676) );
  INV_X1 U10018 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10372) );
  INV_X1 U10019 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10357) );
  NOR2_X1 U10020 ( .A1(n7752), .A2(n7678), .ZN(n7749) );
  MUX2_X1 U10021 ( .A(n7678), .B(n7749), .S(P2_IR_REG_2__SCAN_IN), .Z(n7750)
         );
  INV_X1 U10022 ( .A(n7750), .ZN(n7753) );
  INV_X1 U10023 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7751) );
  NAND2_X1 U10024 ( .A1(n7752), .A2(n7751), .ZN(n7772) );
  NAND2_X1 U10025 ( .A1(n7753), .A2(n7772), .ZN(n15235) );
  NAND2_X1 U10026 ( .A1(n7755), .A2(n7754), .ZN(n7758) );
  NAND2_X1 U10027 ( .A1(n7756), .A2(SI_1_), .ZN(n7757) );
  MUX2_X1 U10028 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n7731), .Z(n7775) );
  XNOR2_X1 U10029 ( .A(n7774), .B(n7775), .ZN(n8601) );
  NAND2_X1 U10030 ( .A1(n8601), .A2(n7802), .ZN(n7763) );
  INV_X1 U10031 ( .A(n8030), .ZN(n7761) );
  NAND2_X1 U10032 ( .A1(n7761), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7762) );
  OAI211_X1 U10033 ( .C1(n10362), .C2(n15235), .A(n7763), .B(n7762), .ZN(
        n10067) );
  NAND2_X1 U10034 ( .A1(n8475), .A2(n7843), .ZN(n7765) );
  NAND2_X1 U10035 ( .A1(n10067), .A2(n8437), .ZN(n7764) );
  NAND2_X1 U10036 ( .A1(n7765), .A2(n7764), .ZN(n7770) );
  NAND2_X1 U10037 ( .A1(n7769), .A2(n7770), .ZN(n7766) );
  NAND3_X1 U10038 ( .A1(n7768), .A2(n7767), .A3(n7766), .ZN(n7792) );
  NAND2_X1 U10039 ( .A1(n7772), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7771) );
  MUX2_X1 U10040 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7771), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7773) );
  AND2_X1 U10041 ( .A1(n7773), .A2(n7804), .ZN(n15251) );
  AOI22_X1 U10042 ( .A1(n8259), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8170), .B2(
        n15251), .ZN(n7779) );
  NAND2_X1 U10043 ( .A1(n7776), .A2(SI_2_), .ZN(n7777) );
  MUX2_X1 U10044 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7731), .Z(n7800) );
  XNOR2_X1 U10045 ( .A(n7800), .B(SI_3_), .ZN(n7797) );
  NAND2_X1 U10046 ( .A1(n8605), .A2(n7802), .ZN(n7778) );
  NAND2_X1 U10047 ( .A1(n8480), .A2(n8437), .ZN(n7787) );
  INV_X1 U10048 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10376) );
  OR2_X1 U10049 ( .A1(n7836), .A2(n10376), .ZN(n7783) );
  INV_X1 U10050 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U10051 ( .A1(n7929), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7781) );
  NAND2_X1 U10052 ( .A1(n7843), .A2(n8479), .ZN(n7786) );
  AND2_X1 U10053 ( .A1(n7787), .A2(n7786), .ZN(n7794) );
  NAND2_X1 U10054 ( .A1(n8479), .A2(n8437), .ZN(n7789) );
  NAND2_X1 U10055 ( .A1(n8480), .A2(n7917), .ZN(n7788) );
  NAND2_X1 U10056 ( .A1(n7789), .A2(n7788), .ZN(n7793) );
  NAND2_X1 U10057 ( .A1(n7794), .A2(n7793), .ZN(n7790) );
  NAND3_X1 U10058 ( .A1(n7792), .A2(n7791), .A3(n7790), .ZN(n7822) );
  INV_X1 U10059 ( .A(n7793), .ZN(n7796) );
  INV_X1 U10060 ( .A(n7794), .ZN(n7795) );
  NAND2_X1 U10061 ( .A1(n7796), .A2(n7795), .ZN(n7821) );
  INV_X1 U10062 ( .A(n7797), .ZN(n7798) );
  NAND2_X1 U10063 ( .A1(n7800), .A2(SI_3_), .ZN(n7801) );
  MUX2_X1 U10064 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7759), .Z(n7826) );
  XNOR2_X1 U10065 ( .A(n7826), .B(SI_4_), .ZN(n7823) );
  NAND2_X1 U10066 ( .A1(n10311), .A2(n8424), .ZN(n7809) );
  NAND2_X1 U10067 ( .A1(n7804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7803) );
  MUX2_X1 U10068 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7803), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7807) );
  INV_X1 U10069 ( .A(n7804), .ZN(n7806) );
  INV_X1 U10070 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U10071 ( .A1(n7806), .A2(n7805), .ZN(n7830) );
  NAND2_X1 U10072 ( .A1(n7807), .A2(n7830), .ZN(n10408) );
  INV_X1 U10073 ( .A(n10408), .ZN(n10415) );
  AOI22_X1 U10074 ( .A1(n8259), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8170), .B2(
        n10415), .ZN(n7808) );
  NAND2_X1 U10075 ( .A1(n10780), .A2(n7845), .ZN(n7818) );
  INV_X1 U10076 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7811) );
  INV_X1 U10077 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7812) );
  OR2_X1 U10078 ( .A1(n8428), .A2(n7812), .ZN(n7815) );
  XNOR2_X1 U10079 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10859) );
  OR2_X1 U10080 ( .A1(n6672), .A2(n10859), .ZN(n7814) );
  INV_X1 U10081 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10858) );
  OR2_X1 U10082 ( .A1(n7836), .A2(n10858), .ZN(n7813) );
  NAND4_X1 U10083 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n13450) );
  NAND2_X1 U10084 ( .A1(n13450), .A2(n7843), .ZN(n7817) );
  NAND2_X1 U10085 ( .A1(n10780), .A2(n7843), .ZN(n7819) );
  OAI21_X1 U10086 ( .B1(n7843), .B2(n10838), .A(n7819), .ZN(n7820) );
  INV_X1 U10087 ( .A(n7823), .ZN(n7824) );
  NAND2_X1 U10088 ( .A1(n7825), .A2(n7824), .ZN(n7828) );
  NAND2_X1 U10089 ( .A1(n7826), .A2(SI_4_), .ZN(n7827) );
  NAND2_X1 U10090 ( .A1(n7828), .A2(n7827), .ZN(n7855) );
  MUX2_X1 U10091 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7731), .Z(n7856) );
  XNOR2_X1 U10092 ( .A(n7856), .B(SI_5_), .ZN(n7853) );
  NAND2_X1 U10093 ( .A1(n8626), .A2(n8424), .ZN(n7833) );
  NAND2_X1 U10094 ( .A1(n7830), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7829) );
  MUX2_X1 U10095 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7829), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n7831) );
  AOI22_X1 U10096 ( .A1(n8259), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8170), .B2(
        n10429), .ZN(n7832) );
  NAND2_X1 U10097 ( .A1(n10848), .A2(n7843), .ZN(n7842) );
  INV_X1 U10098 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7834) );
  OR2_X1 U10099 ( .A1(n8428), .A2(n7834), .ZN(n7840) );
  INV_X1 U10100 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10358) );
  OR2_X1 U10101 ( .A1(n6671), .A2(n10358), .ZN(n7839) );
  INV_X1 U10102 ( .A(n6672), .ZN(n8216) );
  AOI21_X1 U10103 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7835) );
  NOR2_X1 U10104 ( .A1(n7835), .A2(n7863), .ZN(n10844) );
  NAND2_X1 U10105 ( .A1(n8216), .A2(n10844), .ZN(n7838) );
  INV_X1 U10106 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10379) );
  OR2_X1 U10107 ( .A1(n8387), .A2(n10379), .ZN(n7837) );
  NAND2_X1 U10108 ( .A1(n13449), .A2(n7845), .ZN(n7841) );
  NAND2_X1 U10109 ( .A1(n7842), .A2(n7841), .ZN(n7847) );
  AND2_X1 U10110 ( .A1(n13449), .A2(n7843), .ZN(n7844) );
  NAND2_X1 U10111 ( .A1(n7847), .A2(n7848), .ZN(n7846) );
  INV_X1 U10112 ( .A(n7847), .ZN(n7850) );
  INV_X1 U10113 ( .A(n7848), .ZN(n7849) );
  NAND2_X1 U10114 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  NAND2_X1 U10115 ( .A1(n7852), .A2(n7851), .ZN(n7872) );
  INV_X1 U10116 ( .A(n7853), .ZN(n7854) );
  NAND2_X1 U10117 ( .A1(n7855), .A2(n7854), .ZN(n7858) );
  NAND2_X1 U10118 ( .A1(n7856), .A2(SI_5_), .ZN(n7857) );
  NAND2_X1 U10119 ( .A1(n7858), .A2(n7857), .ZN(n7877) );
  MUX2_X1 U10120 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n10302), .Z(n7878) );
  XNOR2_X1 U10121 ( .A(n7878), .B(SI_6_), .ZN(n7875) );
  XNOR2_X1 U10122 ( .A(n7877), .B(n7875), .ZN(n10340) );
  NAND2_X1 U10123 ( .A1(n10340), .A2(n8424), .ZN(n7861) );
  NAND2_X1 U10124 ( .A1(n7881), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7859) );
  XNOR2_X1 U10125 ( .A(n7859), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U10126 ( .A1(n8259), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8170), .B2(
        n10454), .ZN(n7860) );
  NAND2_X1 U10127 ( .A1(n11442), .A2(n7990), .ZN(n7869) );
  NAND2_X1 U10128 ( .A1(n7684), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7867) );
  INV_X1 U10129 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7862) );
  OR2_X1 U10130 ( .A1(n8428), .A2(n7862), .ZN(n7866) );
  NAND2_X1 U10131 ( .A1(n7863), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7887) );
  OAI21_X1 U10132 ( .B1(n7863), .B2(P2_REG3_REG_6__SCAN_IN), .A(n7887), .ZN(
        n11440) );
  OR2_X1 U10133 ( .A1(n6672), .A2(n11440), .ZN(n7865) );
  INV_X1 U10134 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10382) );
  OR2_X1 U10135 ( .A1(n8387), .A2(n10382), .ZN(n7864) );
  NAND4_X1 U10136 ( .A1(n7867), .A2(n7866), .A3(n7865), .A4(n7864), .ZN(n13448) );
  NAND2_X1 U10137 ( .A1(n13448), .A2(n8262), .ZN(n7868) );
  NAND2_X1 U10138 ( .A1(n7869), .A2(n7868), .ZN(n7871) );
  AOI22_X1 U10139 ( .A1(n11442), .A2(n8262), .B1(n7990), .B2(n13448), .ZN(
        n7870) );
  AOI21_X1 U10140 ( .B1(n7872), .B2(n7871), .A(n7870), .ZN(n7874) );
  NOR2_X1 U10141 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  INV_X1 U10142 ( .A(n7875), .ZN(n7876) );
  NAND2_X1 U10143 ( .A1(n7877), .A2(n7876), .ZN(n7880) );
  NAND2_X1 U10144 ( .A1(n7878), .A2(SI_6_), .ZN(n7879) );
  MUX2_X1 U10145 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n10302), .Z(n7902) );
  XNOR2_X1 U10146 ( .A(n7902), .B(SI_7_), .ZN(n7899) );
  XNOR2_X1 U10147 ( .A(n7901), .B(n7899), .ZN(n10345) );
  NAND2_X1 U10148 ( .A1(n10345), .A2(n8424), .ZN(n7884) );
  OAI21_X1 U10149 ( .B1(n7881), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7882) );
  XNOR2_X1 U10150 ( .A(n7882), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U10151 ( .A1(n8259), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8170), .B2(
        n10565), .ZN(n7883) );
  NAND2_X1 U10152 ( .A1(n7884), .A2(n7883), .ZN(n15348) );
  NAND2_X1 U10153 ( .A1(n15348), .A2(n8262), .ZN(n7894) );
  NAND2_X1 U10154 ( .A1(n7684), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7892) );
  INV_X1 U10155 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7885) );
  OR2_X1 U10156 ( .A1(n8428), .A2(n7885), .ZN(n7891) );
  AND2_X1 U10157 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  OR2_X1 U10158 ( .A1(n7888), .A2(n7911), .ZN(n11363) );
  OR2_X1 U10159 ( .A1(n6672), .A2(n11363), .ZN(n7890) );
  INV_X1 U10160 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10455) );
  OR2_X1 U10161 ( .A1(n7836), .A2(n10455), .ZN(n7889) );
  NAND4_X1 U10162 ( .A1(n7892), .A2(n7891), .A3(n7890), .A4(n7889), .ZN(n13447) );
  NAND2_X1 U10163 ( .A1(n13447), .A2(n8437), .ZN(n7893) );
  NAND2_X1 U10164 ( .A1(n7894), .A2(n7893), .ZN(n7896) );
  AOI22_X1 U10165 ( .A1(n15348), .A2(n6690), .B1(n8262), .B2(n13447), .ZN(
        n7895) );
  NOR2_X1 U10166 ( .A1(n7660), .A2(n7896), .ZN(n7897) );
  INV_X1 U10167 ( .A(n7899), .ZN(n7900) );
  NAND2_X1 U10168 ( .A1(n7902), .A2(SI_7_), .ZN(n7903) );
  MUX2_X1 U10169 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n10302), .Z(n7925) );
  XNOR2_X1 U10170 ( .A(n7925), .B(SI_8_), .ZN(n7922) );
  XNOR2_X1 U10171 ( .A(n7924), .B(n7922), .ZN(n10350) );
  NAND2_X1 U10172 ( .A1(n10350), .A2(n8424), .ZN(n7909) );
  NAND2_X1 U10173 ( .A1(n7906), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7905) );
  MUX2_X1 U10174 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7905), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n7907) );
  OR2_X1 U10175 ( .A1(n7906), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8125) );
  AND2_X1 U10176 ( .A1(n7907), .A2(n8125), .ZN(n10667) );
  AOI22_X1 U10177 ( .A1(n8259), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8170), .B2(
        n10667), .ZN(n7908) );
  NAND2_X1 U10178 ( .A1(n11484), .A2(n7990), .ZN(n7919) );
  NAND2_X1 U10179 ( .A1(n7684), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7916) );
  INV_X1 U10180 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7910) );
  OR2_X1 U10181 ( .A1(n8428), .A2(n7910), .ZN(n7915) );
  NOR2_X1 U10182 ( .A1(n7911), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7912) );
  OR2_X1 U10183 ( .A1(n7957), .A2(n7912), .ZN(n11431) );
  OR2_X1 U10184 ( .A1(n6672), .A2(n11431), .ZN(n7914) );
  INV_X1 U10185 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10566) );
  OR2_X1 U10186 ( .A1(n7836), .A2(n10566), .ZN(n7913) );
  NAND4_X1 U10187 ( .A1(n7916), .A2(n7915), .A3(n7914), .A4(n7913), .ZN(n13446) );
  NAND2_X1 U10188 ( .A1(n13446), .A2(n8262), .ZN(n7918) );
  NAND2_X1 U10189 ( .A1(n7919), .A2(n7918), .ZN(n7921) );
  AOI22_X1 U10190 ( .A1(n11484), .A2(n8262), .B1(n6690), .B2(n13446), .ZN(
        n7920) );
  INV_X1 U10191 ( .A(n7922), .ZN(n7923) );
  MUX2_X1 U10192 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n10302), .Z(n7943) );
  XNOR2_X1 U10193 ( .A(n7943), .B(SI_9_), .ZN(n7941) );
  XNOR2_X1 U10194 ( .A(n7942), .B(n7941), .ZN(n10394) );
  NAND2_X1 U10195 ( .A1(n10394), .A2(n8424), .ZN(n7928) );
  NAND2_X1 U10196 ( .A1(n8125), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7926) );
  XNOR2_X1 U10197 ( .A(n7926), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U10198 ( .A1(n8259), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8170), .B2(
        n10869), .ZN(n7927) );
  NAND2_X1 U10199 ( .A1(n15355), .A2(n8262), .ZN(n7935) );
  NAND2_X1 U10200 ( .A1(n8412), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7933) );
  INV_X1 U10201 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10668) );
  OR2_X1 U10202 ( .A1(n6670), .A2(n10668), .ZN(n7932) );
  XNOR2_X1 U10203 ( .A(n7957), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n11647) );
  OR2_X1 U10204 ( .A1(n6672), .A2(n11647), .ZN(n7931) );
  INV_X1 U10205 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11642) );
  OR2_X1 U10206 ( .A1(n8387), .A2(n11642), .ZN(n7930) );
  NAND4_X1 U10207 ( .A1(n7933), .A2(n7932), .A3(n7931), .A4(n7930), .ZN(n13445) );
  NAND2_X1 U10208 ( .A1(n13445), .A2(n6690), .ZN(n7934) );
  INV_X1 U10209 ( .A(n13445), .ZN(n11165) );
  NAND2_X1 U10210 ( .A1(n15355), .A2(n6690), .ZN(n7936) );
  OAI21_X1 U10211 ( .B1(n11165), .B2(n6690), .A(n7936), .ZN(n7937) );
  NAND2_X1 U10212 ( .A1(n7938), .A2(n7937), .ZN(n7940) );
  NAND2_X1 U10213 ( .A1(n6771), .A2(n6709), .ZN(n7939) );
  NAND2_X1 U10214 ( .A1(n7943), .A2(SI_9_), .ZN(n7944) );
  NAND2_X1 U10215 ( .A1(n7945), .A2(n7944), .ZN(n7969) );
  MUX2_X1 U10216 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n10302), .Z(n7970) );
  XNOR2_X1 U10217 ( .A(n7970), .B(SI_10_), .ZN(n7946) );
  XNOR2_X1 U10218 ( .A(n7969), .B(n7946), .ZN(n10437) );
  NAND2_X1 U10219 ( .A1(n10437), .A2(n8424), .ZN(n7952) );
  NOR2_X1 U10220 ( .A1(n8006), .A2(n7678), .ZN(n7947) );
  NAND2_X1 U10221 ( .A1(n7947), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n7950) );
  INV_X1 U10222 ( .A(n7947), .ZN(n7949) );
  INV_X1 U10223 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U10224 ( .A1(n7949), .A2(n7948), .ZN(n7976) );
  AOI22_X1 U10225 ( .A1(n8259), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8170), 
        .B2(n11219), .ZN(n7951) );
  NAND2_X1 U10226 ( .A1(n11803), .A2(n6690), .ZN(n7964) );
  NAND2_X1 U10227 ( .A1(n7684), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7962) );
  INV_X1 U10228 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7953) );
  OR2_X1 U10229 ( .A1(n8428), .A2(n7953), .ZN(n7961) );
  NAND2_X1 U10230 ( .A1(n7957), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7955) );
  INV_X1 U10231 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7954) );
  NAND2_X1 U10232 ( .A1(n7955), .A2(n7954), .ZN(n7958) );
  NAND2_X1 U10233 ( .A1(n7957), .A2(n7956), .ZN(n7981) );
  NAND2_X1 U10234 ( .A1(n7958), .A2(n7981), .ZN(n11797) );
  OR2_X1 U10235 ( .A1(n6672), .A2(n11797), .ZN(n7960) );
  INV_X1 U10236 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10875) );
  OR2_X1 U10237 ( .A1(n8387), .A2(n10875), .ZN(n7959) );
  NAND4_X1 U10238 ( .A1(n7962), .A2(n7961), .A3(n7960), .A4(n7959), .ZN(n13444) );
  NAND2_X1 U10239 ( .A1(n13444), .A2(n8262), .ZN(n7963) );
  NAND2_X1 U10240 ( .A1(n7964), .A2(n7963), .ZN(n7966) );
  AOI22_X1 U10241 ( .A1(n11803), .A2(n8262), .B1(n6690), .B2(n13444), .ZN(
        n7965) );
  INV_X1 U10242 ( .A(n7970), .ZN(n7967) );
  NAND2_X1 U10243 ( .A1(n7967), .A2(n10308), .ZN(n7968) );
  NAND2_X1 U10244 ( .A1(n7969), .A2(n7968), .ZN(n7972) );
  NAND2_X1 U10245 ( .A1(n7970), .A2(SI_10_), .ZN(n7971) );
  NAND2_X1 U10246 ( .A1(n7972), .A2(n7971), .ZN(n8001) );
  MUX2_X1 U10247 ( .A(n10469), .B(n10467), .S(n10302), .Z(n7973) );
  NAND2_X1 U10248 ( .A1(n7973), .A2(n10321), .ZN(n7999) );
  INV_X1 U10249 ( .A(n7973), .ZN(n7974) );
  NAND2_X1 U10250 ( .A1(n7974), .A2(SI_11_), .ZN(n7975) );
  NAND2_X1 U10251 ( .A1(n7999), .A2(n7975), .ZN(n8000) );
  XNOR2_X1 U10252 ( .A(n8001), .B(n8000), .ZN(n10466) );
  NAND2_X1 U10253 ( .A1(n10466), .A2(n8424), .ZN(n7979) );
  NAND2_X1 U10254 ( .A1(n7976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7977) );
  XNOR2_X1 U10255 ( .A(n7977), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U10256 ( .A1(n8259), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8170), 
        .B2(n11396), .ZN(n7978) );
  NAND2_X1 U10257 ( .A1(n15286), .A2(n8262), .ZN(n7988) );
  NAND2_X1 U10258 ( .A1(n7684), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7986) );
  INV_X1 U10259 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7980) );
  OR2_X1 U10260 ( .A1(n8428), .A2(n7980), .ZN(n7985) );
  NAND2_X1 U10261 ( .A1(n7981), .A2(n11215), .ZN(n7982) );
  NAND2_X1 U10262 ( .A1(n8013), .A2(n7982), .ZN(n15287) );
  OR2_X1 U10263 ( .A1(n6672), .A2(n15287), .ZN(n7984) );
  INV_X1 U10264 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11210) );
  OR2_X1 U10265 ( .A1(n8387), .A2(n11210), .ZN(n7983) );
  NAND4_X1 U10266 ( .A1(n7986), .A2(n7985), .A3(n7984), .A4(n7983), .ZN(n13443) );
  NAND2_X1 U10267 ( .A1(n13443), .A2(n7990), .ZN(n7987) );
  NAND2_X1 U10268 ( .A1(n7988), .A2(n7987), .ZN(n7994) );
  NAND2_X1 U10269 ( .A1(n7993), .A2(n7994), .ZN(n7992) );
  INV_X1 U10270 ( .A(n13443), .ZN(n11907) );
  NAND2_X1 U10271 ( .A1(n15286), .A2(n6690), .ZN(n7989) );
  OAI21_X1 U10272 ( .B1(n11907), .B2(n6690), .A(n7989), .ZN(n7991) );
  NAND2_X1 U10273 ( .A1(n7992), .A2(n7991), .ZN(n7998) );
  INV_X1 U10274 ( .A(n7993), .ZN(n7996) );
  INV_X1 U10275 ( .A(n7994), .ZN(n7995) );
  NAND2_X1 U10276 ( .A1(n7996), .A2(n7995), .ZN(n7997) );
  OAI21_X2 U10277 ( .B1(n8001), .B2(n8000), .A(n7999), .ZN(n8024) );
  MUX2_X1 U10278 ( .A(n10559), .B(n10560), .S(n10302), .Z(n8002) );
  NAND2_X1 U10279 ( .A1(n8002), .A2(n10339), .ZN(n8025) );
  INV_X1 U10280 ( .A(n8002), .ZN(n8003) );
  NAND2_X1 U10281 ( .A1(n8003), .A2(SI_12_), .ZN(n8004) );
  XNOR2_X1 U10282 ( .A(n8024), .B(n8023), .ZN(n10558) );
  NAND2_X1 U10283 ( .A1(n10558), .A2(n8424), .ZN(n8011) );
  NOR2_X1 U10284 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .ZN(n8005) );
  NAND2_X1 U10285 ( .A1(n8006), .A2(n8005), .ZN(n8008) );
  NAND2_X1 U10286 ( .A1(n8008), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8007) );
  MUX2_X1 U10287 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8007), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8009) );
  AND2_X1 U10288 ( .A1(n8009), .A2(n8033), .ZN(n11618) );
  AOI22_X1 U10289 ( .A1(n8259), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8170), 
        .B2(n11618), .ZN(n8010) );
  NAND2_X1 U10290 ( .A1(n11917), .A2(n6690), .ZN(n8020) );
  NAND2_X1 U10291 ( .A1(n8412), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8018) );
  INV_X1 U10292 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11397) );
  OR2_X1 U10293 ( .A1(n6671), .A2(n11397), .ZN(n8017) );
  NAND2_X1 U10294 ( .A1(n8013), .A2(n8012), .ZN(n8014) );
  NAND2_X1 U10295 ( .A1(n8039), .A2(n8014), .ZN(n11911) );
  OR2_X1 U10296 ( .A1(n6672), .A2(n11911), .ZN(n8016) );
  INV_X1 U10297 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11912) );
  OR2_X1 U10298 ( .A1(n7836), .A2(n11912), .ZN(n8015) );
  NAND4_X1 U10299 ( .A1(n8018), .A2(n8017), .A3(n8016), .A4(n8015), .ZN(n13442) );
  NAND2_X1 U10300 ( .A1(n13442), .A2(n8262), .ZN(n8019) );
  AOI22_X1 U10301 ( .A1(n11917), .A2(n8262), .B1(n8437), .B2(n13442), .ZN(
        n8021) );
  INV_X1 U10302 ( .A(n8021), .ZN(n8022) );
  NAND2_X1 U10303 ( .A1(n8024), .A2(n8023), .ZN(n8026) );
  MUX2_X1 U10304 ( .A(n10620), .B(n10618), .S(n10302), .Z(n8027) );
  NAND2_X1 U10305 ( .A1(n8027), .A2(n10434), .ZN(n8051) );
  INV_X1 U10306 ( .A(n8027), .ZN(n8028) );
  NAND2_X1 U10307 ( .A1(n8028), .A2(SI_13_), .ZN(n8029) );
  NAND2_X1 U10308 ( .A1(n10617), .A2(n8424), .ZN(n8038) );
  NAND2_X1 U10309 ( .A1(n8033), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8032) );
  MUX2_X1 U10310 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8032), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8035) );
  INV_X1 U10311 ( .A(n8076), .ZN(n8034) );
  NAND2_X1 U10312 ( .A1(n8035), .A2(n8034), .ZN(n11629) );
  OAI22_X1 U10313 ( .A1(n8031), .A2(n10620), .B1(n11629), .B2(n10362), .ZN(
        n8036) );
  INV_X1 U10314 ( .A(n8036), .ZN(n8037) );
  NAND2_X1 U10315 ( .A1(n12039), .A2(n8262), .ZN(n8047) );
  AND2_X1 U10316 ( .A1(n8039), .A2(n11630), .ZN(n8040) );
  NOR2_X1 U10317 ( .A1(n8056), .A2(n8040), .ZN(n12038) );
  NAND2_X1 U10318 ( .A1(n8216), .A2(n12038), .ZN(n8045) );
  INV_X1 U10319 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8041) );
  OR2_X1 U10320 ( .A1(n8428), .A2(n8041), .ZN(n8044) );
  INV_X1 U10321 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11624) );
  OR2_X1 U10322 ( .A1(n8387), .A2(n11624), .ZN(n8043) );
  INV_X1 U10323 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11616) );
  OR2_X1 U10324 ( .A1(n6670), .A2(n11616), .ZN(n8042) );
  NAND4_X1 U10325 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8042), .ZN(n13441) );
  NAND2_X1 U10326 ( .A1(n13441), .A2(n6690), .ZN(n8046) );
  AOI22_X1 U10327 ( .A1(n12039), .A2(n6690), .B1(n8262), .B2(n13441), .ZN(
        n8048) );
  MUX2_X1 U10328 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n10302), .Z(n8070) );
  NAND2_X1 U10329 ( .A1(n10754), .A2(n8424), .ZN(n8055) );
  OR2_X1 U10330 ( .A1(n8076), .A2(n7678), .ZN(n8053) );
  XNOR2_X1 U10331 ( .A(n8053), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U10332 ( .A1(n8259), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n13467), 
        .B2(n8170), .ZN(n8054) );
  NAND2_X1 U10333 ( .A1(n13811), .A2(n6690), .ZN(n8065) );
  NAND2_X1 U10334 ( .A1(n8056), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8083) );
  OR2_X1 U10335 ( .A1(n8056), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10336 ( .A1(n8083), .A2(n8057), .ZN(n12121) );
  OR2_X1 U10337 ( .A1(n12121), .A2(n6672), .ZN(n8063) );
  INV_X1 U10338 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8058) );
  OR2_X1 U10339 ( .A1(n6670), .A2(n8058), .ZN(n8062) );
  INV_X1 U10340 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8059) );
  OR2_X1 U10341 ( .A1(n8428), .A2(n8059), .ZN(n8061) );
  INV_X1 U10342 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n13453) );
  OR2_X1 U10343 ( .A1(n8387), .A2(n13453), .ZN(n8060) );
  NAND4_X1 U10344 ( .A1(n8063), .A2(n8062), .A3(n8061), .A4(n8060), .ZN(n13440) );
  NAND2_X1 U10345 ( .A1(n13440), .A2(n8262), .ZN(n8064) );
  NAND2_X1 U10346 ( .A1(n8065), .A2(n8064), .ZN(n8068) );
  INV_X1 U10347 ( .A(n13440), .ZN(n8469) );
  NAND2_X1 U10348 ( .A1(n13811), .A2(n8262), .ZN(n8066) );
  OAI21_X1 U10349 ( .B1(n7843), .B2(n8469), .A(n8066), .ZN(n8067) );
  INV_X1 U10350 ( .A(n8068), .ZN(n8069) );
  MUX2_X1 U10351 ( .A(n10993), .B(n10991), .S(n10302), .Z(n8072) );
  INV_X1 U10352 ( .A(n8072), .ZN(n8073) );
  NAND2_X1 U10353 ( .A1(n8073), .A2(SI_15_), .ZN(n8074) );
  XNOR2_X1 U10354 ( .A(n8096), .B(n8095), .ZN(n10990) );
  NAND2_X1 U10355 ( .A1(n10990), .A2(n8424), .ZN(n8082) );
  INV_X1 U10356 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8075) );
  AOI21_X1 U10357 ( .B1(n8076), .B2(n8075), .A(n7678), .ZN(n8077) );
  NAND2_X1 U10358 ( .A1(n8077), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8080) );
  INV_X1 U10359 ( .A(n8077), .ZN(n8079) );
  INV_X1 U10360 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U10361 ( .A1(n8079), .A2(n8078), .ZN(n8102) );
  AOI22_X1 U10362 ( .A1(n15263), .A2(n8170), .B1(n8259), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10363 ( .A1(n13805), .A2(n8262), .ZN(n8092) );
  NAND2_X1 U10364 ( .A1(n8083), .A2(n15257), .ZN(n8084) );
  AND2_X1 U10365 ( .A1(n8108), .A2(n8084), .ZN(n13423) );
  NAND2_X1 U10366 ( .A1(n8216), .A2(n13423), .ZN(n8090) );
  INV_X1 U10367 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15259) );
  OR2_X1 U10368 ( .A1(n6671), .A2(n15259), .ZN(n8089) );
  INV_X1 U10369 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8085) );
  OR2_X1 U10370 ( .A1(n8428), .A2(n8085), .ZN(n8088) );
  INV_X1 U10371 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8086) );
  OR2_X1 U10372 ( .A1(n7836), .A2(n8086), .ZN(n8087) );
  NAND4_X1 U10373 ( .A1(n8090), .A2(n8089), .A3(n8088), .A4(n8087), .ZN(n13439) );
  NAND2_X1 U10374 ( .A1(n13439), .A2(n6690), .ZN(n8091) );
  NAND2_X1 U10375 ( .A1(n8092), .A2(n8091), .ZN(n8094) );
  AOI22_X1 U10376 ( .A1(n13805), .A2(n8437), .B1(n8262), .B2(n13439), .ZN(
        n8093) );
  MUX2_X1 U10377 ( .A(n14648), .B(n14636), .S(n10302), .Z(n8099) );
  INV_X1 U10378 ( .A(n8099), .ZN(n8100) );
  NAND2_X1 U10379 ( .A1(n8100), .A2(SI_16_), .ZN(n8101) );
  XNOR2_X1 U10380 ( .A(n8118), .B(n8117), .ZN(n11135) );
  NAND2_X1 U10381 ( .A1(n11135), .A2(n8424), .ZN(n8106) );
  NAND2_X1 U10382 ( .A1(n8102), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8103) );
  XNOR2_X1 U10383 ( .A(n8103), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13483) );
  NOR2_X1 U10384 ( .A1(n8031), .A2(n14648), .ZN(n8104) );
  AOI21_X1 U10385 ( .B1(n13483), .B2(n8170), .A(n8104), .ZN(n8105) );
  NAND2_X1 U10386 ( .A1(n13798), .A2(n6690), .ZN(n8113) );
  INV_X1 U10387 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8107) );
  AND2_X1 U10388 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  OR2_X1 U10389 ( .A1(n8109), .A2(n8133), .ZN(n13347) );
  AOI22_X1 U10390 ( .A1(n7684), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8412), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n8111) );
  INV_X1 U10391 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13459) );
  OR2_X1 U10392 ( .A1(n7836), .A2(n13459), .ZN(n8110) );
  OAI211_X1 U10393 ( .C1(n13347), .C2(n6672), .A(n8111), .B(n8110), .ZN(n13438) );
  NAND2_X1 U10394 ( .A1(n13438), .A2(n8262), .ZN(n8112) );
  INV_X1 U10395 ( .A(n13438), .ZN(n9228) );
  NAND2_X1 U10396 ( .A1(n13798), .A2(n8262), .ZN(n8114) );
  OAI21_X1 U10397 ( .B1(n7843), .B2(n9228), .A(n8114), .ZN(n8115) );
  INV_X1 U10398 ( .A(n8144), .ZN(n8142) );
  NAND2_X1 U10399 ( .A1(n8118), .A2(n8117), .ZN(n8120) );
  NAND2_X2 U10400 ( .A1(n8120), .A2(n8119), .ZN(n8147) );
  MUX2_X1 U10401 ( .A(n11227), .B(n14610), .S(n10302), .Z(n8121) );
  INV_X1 U10402 ( .A(n8121), .ZN(n8122) );
  NAND2_X1 U10403 ( .A1(n8122), .A2(SI_17_), .ZN(n8123) );
  XNOR2_X1 U10404 ( .A(n8147), .B(n8146), .ZN(n11226) );
  NAND2_X1 U10405 ( .A1(n11226), .A2(n8424), .ZN(n8132) );
  NOR2_X1 U10406 ( .A1(n8125), .A2(n8124), .ZN(n8128) );
  NOR2_X1 U10407 ( .A1(n8128), .A2(n7678), .ZN(n8126) );
  MUX2_X1 U10408 ( .A(n7678), .B(n8126), .S(P2_IR_REG_17__SCAN_IN), .Z(n8130)
         );
  NAND2_X1 U10409 ( .A1(n8128), .A2(n8127), .ZN(n8149) );
  INV_X1 U10410 ( .A(n8149), .ZN(n8129) );
  NOR2_X1 U10411 ( .A1(n8130), .A2(n8129), .ZN(n15280) );
  AOI22_X1 U10412 ( .A1(n8259), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8170), 
        .B2(n15280), .ZN(n8131) );
  NAND2_X1 U10413 ( .A1(n12201), .A2(n8262), .ZN(n8138) );
  NOR2_X1 U10414 ( .A1(n8133), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8134) );
  OR2_X1 U10415 ( .A1(n8153), .A2(n8134), .ZN(n13357) );
  AOI22_X1 U10416 ( .A1(n7684), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8412), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n8136) );
  INV_X1 U10417 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13477) );
  OR2_X1 U10418 ( .A1(n8387), .A2(n13477), .ZN(n8135) );
  OAI211_X1 U10419 ( .C1(n13357), .C2(n6672), .A(n8136), .B(n8135), .ZN(n13437) );
  NAND2_X1 U10420 ( .A1(n13437), .A2(n8437), .ZN(n8137) );
  NAND2_X1 U10421 ( .A1(n8138), .A2(n8137), .ZN(n8143) );
  INV_X1 U10422 ( .A(n8143), .ZN(n8141) );
  AOI22_X1 U10423 ( .A1(n12201), .A2(n6690), .B1(n8262), .B2(n13437), .ZN(
        n8139) );
  INV_X1 U10424 ( .A(n8139), .ZN(n8140) );
  OAI21_X1 U10425 ( .B1(n8142), .B2(n8141), .A(n8140), .ZN(n8145) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n10302), .Z(n8191) );
  XNOR2_X1 U10427 ( .A(n8166), .B(n8191), .ZN(n11547) );
  NAND2_X1 U10428 ( .A1(n11547), .A2(n8424), .ZN(n8152) );
  NAND2_X1 U10429 ( .A1(n8149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8150) );
  XNOR2_X1 U10430 ( .A(n8150), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13492) );
  AOI22_X1 U10431 ( .A1(n8259), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8170), 
        .B2(n13492), .ZN(n8151) );
  NAND2_X1 U10432 ( .A1(n13787), .A2(n8437), .ZN(n8159) );
  OR2_X1 U10433 ( .A1(n8153), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U10434 ( .A1(n8174), .A2(n8154), .ZN(n13712) );
  AOI22_X1 U10435 ( .A1(n7684), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8412), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n8157) );
  INV_X1 U10436 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8155) );
  OR2_X1 U10437 ( .A1(n7836), .A2(n8155), .ZN(n8156) );
  OAI211_X1 U10438 ( .C1(n13712), .C2(n6672), .A(n8157), .B(n8156), .ZN(n13436) );
  NAND2_X1 U10439 ( .A1(n13436), .A2(n8262), .ZN(n8158) );
  NAND2_X1 U10440 ( .A1(n8159), .A2(n8158), .ZN(n8163) );
  NAND2_X1 U10441 ( .A1(n13787), .A2(n8262), .ZN(n8161) );
  NAND2_X1 U10442 ( .A1(n13436), .A2(n6690), .ZN(n8160) );
  NAND2_X1 U10443 ( .A1(n8161), .A2(n8160), .ZN(n8162) );
  INV_X1 U10444 ( .A(n8163), .ZN(n8164) );
  INV_X1 U10445 ( .A(n8191), .ZN(n8165) );
  OR2_X1 U10446 ( .A1(n8189), .A2(n10654), .ZN(n8167) );
  MUX2_X1 U10447 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n10302), .Z(n8192) );
  XNOR2_X1 U10448 ( .A(n8192), .B(SI_19_), .ZN(n8168) );
  NAND2_X1 U10449 ( .A1(n8811), .A2(n8424), .ZN(n8172) );
  AOI22_X1 U10450 ( .A1(n8259), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10262), 
        .B2(n8170), .ZN(n8171) );
  NAND2_X1 U10451 ( .A1(n13782), .A2(n8262), .ZN(n8183) );
  INV_X1 U10452 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8173) );
  NAND2_X1 U10453 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  AND2_X1 U10454 ( .A1(n8197), .A2(n8175), .ZN(n13698) );
  NAND2_X1 U10455 ( .A1(n13698), .A2(n8216), .ZN(n8181) );
  INV_X1 U10456 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U10457 ( .A1(n8352), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8177) );
  NAND2_X1 U10458 ( .A1(n8412), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8176) );
  OAI211_X1 U10459 ( .C1(n6670), .C2(n8178), .A(n8177), .B(n8176), .ZN(n8179)
         );
  INV_X1 U10460 ( .A(n8179), .ZN(n8180) );
  NAND2_X1 U10461 ( .A1(n8181), .A2(n8180), .ZN(n13435) );
  NAND2_X1 U10462 ( .A1(n13435), .A2(n8437), .ZN(n8182) );
  NAND2_X1 U10463 ( .A1(n8183), .A2(n8182), .ZN(n8185) );
  AOI22_X1 U10464 ( .A1(n13782), .A2(n6690), .B1(n8262), .B2(n13435), .ZN(
        n8184) );
  NOR2_X1 U10465 ( .A1(n8191), .A2(SI_18_), .ZN(n8187) );
  NOR2_X1 U10466 ( .A1(n8192), .A2(SI_19_), .ZN(n8186) );
  OAI21_X1 U10467 ( .B1(n8165), .B2(n10654), .A(n10711), .ZN(n8193) );
  AND2_X1 U10468 ( .A1(SI_18_), .A2(SI_19_), .ZN(n8190) );
  AOI22_X1 U10469 ( .A1(n8193), .A2(n8192), .B1(n8191), .B2(n8190), .ZN(n8194)
         );
  XNOR2_X1 U10470 ( .A(n8232), .B(SI_20_), .ZN(n8209) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n10302), .Z(n8230) );
  XNOR2_X1 U10472 ( .A(n8209), .B(n8230), .ZN(n14759) );
  NAND2_X1 U10473 ( .A1(n14759), .A2(n8424), .ZN(n8196) );
  NAND2_X1 U10474 ( .A1(n8259), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10475 ( .A1(n13777), .A2(n7990), .ZN(n8205) );
  INV_X1 U10476 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13379) );
  AND2_X1 U10477 ( .A1(n8197), .A2(n13379), .ZN(n8198) );
  OR2_X1 U10478 ( .A1(n8198), .A2(n8214), .ZN(n13682) );
  INV_X1 U10479 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8201) );
  NAND2_X1 U10480 ( .A1(n8352), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10481 ( .A1(n8412), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8199) );
  OAI211_X1 U10482 ( .C1(n6671), .C2(n8201), .A(n8200), .B(n8199), .ZN(n8202)
         );
  INV_X1 U10483 ( .A(n8202), .ZN(n8203) );
  OAI21_X1 U10484 ( .B1(n13682), .B2(n6672), .A(n8203), .ZN(n13434) );
  NAND2_X1 U10485 ( .A1(n13434), .A2(n8262), .ZN(n8204) );
  INV_X1 U10486 ( .A(n13434), .ZN(n13660) );
  NAND2_X1 U10487 ( .A1(n13777), .A2(n8262), .ZN(n8206) );
  OAI21_X1 U10488 ( .B1(n7843), .B2(n13660), .A(n8206), .ZN(n8207) );
  INV_X1 U10489 ( .A(n8230), .ZN(n8233) );
  INV_X1 U10490 ( .A(n8232), .ZN(n8208) );
  OAI22_X1 U10491 ( .A1(n8209), .A2(n8233), .B1(n8208), .B2(n11059), .ZN(n8211) );
  MUX2_X1 U10492 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n10302), .Z(n8234) );
  XNOR2_X1 U10493 ( .A(n8234), .B(SI_21_), .ZN(n8210) );
  XNOR2_X1 U10494 ( .A(n8211), .B(n8210), .ZN(n11832) );
  NAND2_X1 U10495 ( .A1(n11832), .A2(n8424), .ZN(n8213) );
  NAND2_X1 U10496 ( .A1(n8259), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U10497 ( .A1(n13772), .A2(n8262), .ZN(n8223) );
  OR2_X1 U10498 ( .A1(n8214), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8215) );
  AND2_X1 U10499 ( .A1(n8241), .A2(n8215), .ZN(n13666) );
  NAND2_X1 U10500 ( .A1(n13666), .A2(n8216), .ZN(n8221) );
  INV_X1 U10501 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14541) );
  NAND2_X1 U10502 ( .A1(n8352), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8218) );
  NAND2_X1 U10503 ( .A1(n8412), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8217) );
  OAI211_X1 U10504 ( .C1(n6671), .C2(n14541), .A(n8218), .B(n8217), .ZN(n8219)
         );
  INV_X1 U10505 ( .A(n8219), .ZN(n8220) );
  NAND2_X1 U10506 ( .A1(n8221), .A2(n8220), .ZN(n13433) );
  NAND2_X1 U10507 ( .A1(n13433), .A2(n8437), .ZN(n8222) );
  NAND2_X1 U10508 ( .A1(n8223), .A2(n8222), .ZN(n8226) );
  AOI22_X1 U10509 ( .A1(n13772), .A2(n7990), .B1(n8262), .B2(n13433), .ZN(
        n8224) );
  INV_X1 U10510 ( .A(n8225), .ZN(n8228) );
  INV_X1 U10511 ( .A(n8234), .ZN(n8229) );
  NAND2_X1 U10512 ( .A1(n8229), .A2(n11206), .ZN(n8235) );
  OAI21_X1 U10513 ( .B1(n8230), .B2(SI_20_), .A(n8235), .ZN(n8231) );
  NOR2_X1 U10514 ( .A1(n8233), .A2(n11059), .ZN(n8236) );
  AOI22_X1 U10515 ( .A1(n8236), .A2(n8235), .B1(n8234), .B2(SI_21_), .ZN(n8237) );
  MUX2_X1 U10516 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n10302), .Z(n8254) );
  XNOR2_X1 U10517 ( .A(n8846), .B(n8254), .ZN(n11830) );
  NAND2_X1 U10518 ( .A1(n11830), .A2(n8424), .ZN(n8240) );
  NAND2_X1 U10519 ( .A1(n8259), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10520 ( .A1(n13765), .A2(n6690), .ZN(n8251) );
  INV_X1 U10521 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14574) );
  NAND2_X1 U10522 ( .A1(n8241), .A2(n14574), .ZN(n8243) );
  INV_X1 U10523 ( .A(n8264), .ZN(n8242) );
  NAND2_X1 U10524 ( .A1(n8243), .A2(n8242), .ZN(n13644) );
  OR2_X1 U10525 ( .A1(n13644), .A2(n6672), .ZN(n8249) );
  INV_X1 U10526 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U10527 ( .A1(n7684), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8245) );
  INV_X1 U10528 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14500) );
  OR2_X1 U10529 ( .A1(n8428), .A2(n14500), .ZN(n8244) );
  OAI211_X1 U10530 ( .C1(n8246), .C2(n8387), .A(n8245), .B(n8244), .ZN(n8247)
         );
  INV_X1 U10531 ( .A(n8247), .ZN(n8248) );
  NAND2_X1 U10532 ( .A1(n13432), .A2(n8262), .ZN(n8250) );
  NAND2_X1 U10533 ( .A1(n8251), .A2(n8250), .ZN(n8253) );
  AOI22_X1 U10534 ( .A1(n13765), .A2(n8262), .B1(n8437), .B2(n13432), .ZN(
        n8252) );
  INV_X1 U10535 ( .A(n8254), .ZN(n8257) );
  NAND2_X1 U10536 ( .A1(n8255), .A2(SI_22_), .ZN(n8256) );
  OAI21_X2 U10537 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8283) );
  MUX2_X1 U10538 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n7731), .Z(n8282) );
  XNOR2_X1 U10539 ( .A(n8281), .B(SI_23_), .ZN(n12007) );
  NAND2_X1 U10540 ( .A1(n12007), .A2(n8424), .ZN(n8261) );
  NAND2_X1 U10541 ( .A1(n8259), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U10542 ( .A1(n13759), .A2(n8262), .ZN(n8270) );
  NAND2_X1 U10543 ( .A1(n7684), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8268) );
  INV_X1 U10544 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8263) );
  OR2_X1 U10545 ( .A1(n8428), .A2(n8263), .ZN(n8267) );
  NAND2_X1 U10546 ( .A1(n8264), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8288) );
  OAI21_X1 U10547 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n8264), .A(n8288), .ZN(
        n13631) );
  OR2_X1 U10548 ( .A1(n6672), .A2(n13631), .ZN(n8266) );
  INV_X1 U10549 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13632) );
  OR2_X1 U10550 ( .A1(n8387), .A2(n13632), .ZN(n8265) );
  NAND4_X1 U10551 ( .A1(n8268), .A2(n8267), .A3(n8266), .A4(n8265), .ZN(n13606) );
  NAND2_X1 U10552 ( .A1(n13606), .A2(n6690), .ZN(n8269) );
  NAND2_X1 U10553 ( .A1(n8270), .A2(n8269), .ZN(n8276) );
  NAND2_X1 U10554 ( .A1(n8275), .A2(n8276), .ZN(n8274) );
  NAND2_X1 U10555 ( .A1(n13759), .A2(n6690), .ZN(n8272) );
  NAND2_X1 U10556 ( .A1(n13606), .A2(n8262), .ZN(n8271) );
  NAND2_X1 U10557 ( .A1(n8272), .A2(n8271), .ZN(n8273) );
  NAND2_X1 U10558 ( .A1(n8274), .A2(n8273), .ZN(n8280) );
  INV_X1 U10559 ( .A(n8275), .ZN(n8278) );
  INV_X1 U10560 ( .A(n8276), .ZN(n8277) );
  NAND2_X1 U10561 ( .A1(n8278), .A2(n8277), .ZN(n8279) );
  NAND2_X1 U10562 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  MUX2_X1 U10563 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n10302), .Z(n8300) );
  XNOR2_X1 U10564 ( .A(n8299), .B(n8300), .ZN(n12151) );
  NAND2_X1 U10565 ( .A1(n12151), .A2(n8424), .ZN(n8286) );
  INV_X1 U10566 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12190) );
  OR2_X1 U10567 ( .A1(n8031), .A2(n12190), .ZN(n8285) );
  NAND2_X1 U10568 ( .A1(n13752), .A2(n8437), .ZN(n8296) );
  NAND2_X1 U10569 ( .A1(n7684), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8294) );
  INV_X1 U10570 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8287) );
  OR2_X1 U10571 ( .A1(n8428), .A2(n8287), .ZN(n8293) );
  OAI21_X1 U10572 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8289), .A(n8327), .ZN(
        n13366) );
  OR2_X1 U10573 ( .A1(n6672), .A2(n13366), .ZN(n8292) );
  INV_X1 U10574 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8290) );
  OR2_X1 U10575 ( .A1(n8387), .A2(n8290), .ZN(n8291) );
  NAND4_X1 U10576 ( .A1(n8294), .A2(n8293), .A3(n8292), .A4(n8291), .ZN(n13584) );
  NAND2_X1 U10577 ( .A1(n13584), .A2(n7843), .ZN(n8295) );
  AOI22_X1 U10578 ( .A1(n13752), .A2(n8262), .B1(n8437), .B2(n13584), .ZN(
        n8297) );
  NAND2_X1 U10579 ( .A1(n8301), .A2(SI_24_), .ZN(n8302) );
  INV_X1 U10580 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13851) );
  MUX2_X1 U10581 ( .A(n13851), .B(n14396), .S(n10302), .Z(n8303) );
  NAND2_X1 U10582 ( .A1(n8303), .A2(n14664), .ZN(n8320) );
  INV_X1 U10583 ( .A(n8303), .ZN(n8304) );
  NAND2_X1 U10584 ( .A1(n8304), .A2(SI_25_), .ZN(n8305) );
  NAND2_X1 U10585 ( .A1(n8320), .A2(n8305), .ZN(n8321) );
  XNOR2_X1 U10586 ( .A(n8322), .B(n8321), .ZN(n13847) );
  NAND2_X1 U10587 ( .A1(n13847), .A2(n8424), .ZN(n8307) );
  OR2_X1 U10588 ( .A1(n8031), .A2(n13851), .ZN(n8306) );
  NAND2_X1 U10589 ( .A1(n13747), .A2(n7843), .ZN(n8315) );
  NAND2_X1 U10590 ( .A1(n7684), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8313) );
  INV_X1 U10591 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8308) );
  OR2_X1 U10592 ( .A1(n8428), .A2(n8308), .ZN(n8312) );
  INV_X1 U10593 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13335) );
  XNOR2_X1 U10594 ( .A(n8327), .B(n13335), .ZN(n13588) );
  OR2_X1 U10595 ( .A1(n6672), .A2(n13588), .ZN(n8311) );
  INV_X1 U10596 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8309) );
  OR2_X1 U10597 ( .A1(n7836), .A2(n8309), .ZN(n8310) );
  NAND4_X1 U10598 ( .A1(n8313), .A2(n8312), .A3(n8311), .A4(n8310), .ZN(n13605) );
  NAND2_X1 U10599 ( .A1(n13605), .A2(n7990), .ZN(n8314) );
  NAND2_X1 U10600 ( .A1(n13747), .A2(n7990), .ZN(n8317) );
  NAND2_X1 U10601 ( .A1(n13605), .A2(n8262), .ZN(n8316) );
  NAND2_X1 U10602 ( .A1(n8317), .A2(n8316), .ZN(n8318) );
  INV_X1 U10603 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13845) );
  INV_X1 U10604 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14392) );
  MUX2_X1 U10605 ( .A(n13845), .B(n14392), .S(n10302), .Z(n8345) );
  XNOR2_X1 U10606 ( .A(n8345), .B(SI_26_), .ZN(n8344) );
  XNOR2_X1 U10607 ( .A(n8349), .B(n8344), .ZN(n13843) );
  NAND2_X1 U10608 ( .A1(n13843), .A2(n8424), .ZN(n8324) );
  OR2_X1 U10609 ( .A1(n8031), .A2(n13845), .ZN(n8323) );
  NAND2_X1 U10610 ( .A1(n13742), .A2(n7990), .ZN(n8337) );
  NAND2_X1 U10611 ( .A1(n7684), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8335) );
  INV_X1 U10612 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8325) );
  OR2_X1 U10613 ( .A1(n8428), .A2(n8325), .ZN(n8334) );
  INV_X1 U10614 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8326) );
  OAI21_X1 U10615 ( .B1(n8327), .B2(n13335), .A(n8326), .ZN(n8330) );
  INV_X1 U10616 ( .A(n8327), .ZN(n8329) );
  AND2_X1 U10617 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8328) );
  NAND2_X1 U10618 ( .A1(n8329), .A2(n8328), .ZN(n8356) );
  NAND2_X1 U10619 ( .A1(n8330), .A2(n8356), .ZN(n13568) );
  INV_X1 U10620 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8331) );
  OR2_X1 U10621 ( .A1(n8387), .A2(n8331), .ZN(n8332) );
  NAND4_X1 U10622 ( .A1(n8335), .A2(n8334), .A3(n8333), .A4(n8332), .ZN(n13583) );
  NAND2_X1 U10623 ( .A1(n13583), .A2(n8262), .ZN(n8336) );
  NAND2_X1 U10624 ( .A1(n8337), .A2(n8336), .ZN(n8341) );
  INV_X1 U10625 ( .A(n13583), .ZN(n13336) );
  NAND2_X1 U10626 ( .A1(n13742), .A2(n7843), .ZN(n8338) );
  OAI21_X1 U10627 ( .B1(n7843), .B2(n13336), .A(n8338), .ZN(n8339) );
  INV_X1 U10628 ( .A(n8341), .ZN(n8342) );
  NAND2_X1 U10629 ( .A1(n6764), .A2(n8342), .ZN(n8343) );
  INV_X1 U10630 ( .A(n8344), .ZN(n8348) );
  INV_X1 U10631 ( .A(n8345), .ZN(n8346) );
  NAND2_X1 U10632 ( .A1(n8346), .A2(SI_26_), .ZN(n8347) );
  MUX2_X1 U10633 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n10302), .Z(n8366) );
  NAND2_X1 U10634 ( .A1(n12269), .A2(n8424), .ZN(n8351) );
  INV_X1 U10635 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12271) );
  OR2_X1 U10636 ( .A1(n8031), .A2(n12271), .ZN(n8350) );
  NAND2_X2 U10637 ( .A1(n8351), .A2(n8350), .ZN(n13734) );
  NAND2_X1 U10638 ( .A1(n13734), .A2(n8262), .ZN(n8363) );
  NAND2_X1 U10639 ( .A1(n8352), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8361) );
  INV_X1 U10640 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8353) );
  OR2_X1 U10641 ( .A1(n6670), .A2(n8353), .ZN(n8360) );
  INV_X1 U10642 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14581) );
  OR2_X1 U10643 ( .A1(n8428), .A2(n14581), .ZN(n8359) );
  INV_X1 U10644 ( .A(n8356), .ZN(n8354) );
  NAND2_X1 U10645 ( .A1(n8354), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8429) );
  INV_X1 U10646 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U10647 ( .A1(n8356), .A2(n8355), .ZN(n8357) );
  NAND2_X1 U10648 ( .A1(n8429), .A2(n8357), .ZN(n10193) );
  OR2_X1 U10649 ( .A1(n6672), .A2(n10193), .ZN(n8358) );
  NAND4_X1 U10650 ( .A1(n8361), .A2(n8360), .A3(n8359), .A4(n8358), .ZN(n13575) );
  NAND2_X1 U10651 ( .A1(n13575), .A2(n7990), .ZN(n8362) );
  AOI22_X1 U10652 ( .A1(n13734), .A2(n8437), .B1(n8262), .B2(n13575), .ZN(
        n8364) );
  NAND2_X1 U10653 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  MUX2_X1 U10654 ( .A(n14552), .B(n7129), .S(n10302), .Z(n8369) );
  INV_X1 U10655 ( .A(SI_28_), .ZN(n12111) );
  NAND2_X1 U10656 ( .A1(n8369), .A2(n12111), .ZN(n8372) );
  INV_X1 U10657 ( .A(n8369), .ZN(n8370) );
  NAND2_X1 U10658 ( .A1(n8370), .A2(SI_28_), .ZN(n8371) );
  NAND2_X1 U10659 ( .A1(n8372), .A2(n8371), .ZN(n8422) );
  INV_X1 U10660 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12294) );
  MUX2_X1 U10661 ( .A(n12294), .B(n14597), .S(n7731), .Z(n8373) );
  INV_X1 U10662 ( .A(SI_29_), .ZN(n12297) );
  NAND2_X1 U10663 ( .A1(n8373), .A2(n12297), .ZN(n8376) );
  INV_X1 U10664 ( .A(n8373), .ZN(n8374) );
  NAND2_X1 U10665 ( .A1(n8374), .A2(SI_29_), .ZN(n8375) );
  NAND2_X1 U10666 ( .A1(n8410), .A2(n8409), .ZN(n8377) );
  MUX2_X1 U10667 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n10302), .Z(n8378) );
  XNOR2_X1 U10668 ( .A(n8378), .B(SI_30_), .ZN(n8393) );
  NAND2_X1 U10669 ( .A1(n8378), .A2(SI_30_), .ZN(n8379) );
  MUX2_X1 U10670 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n10302), .Z(n8380) );
  XNOR2_X1 U10671 ( .A(n8380), .B(SI_31_), .ZN(n8381) );
  INV_X1 U10672 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13836) );
  OR2_X1 U10673 ( .A1(n8031), .A2(n13836), .ZN(n8383) );
  INV_X1 U10674 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8385) );
  NOR2_X1 U10675 ( .A1(n6671), .A2(n8385), .ZN(n8390) );
  INV_X1 U10676 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8386) );
  NOR2_X1 U10677 ( .A1(n8387), .A2(n8386), .ZN(n8389) );
  INV_X1 U10678 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14657) );
  NOR2_X1 U10679 ( .A1(n8428), .A2(n14657), .ZN(n8388) );
  NAND2_X1 U10680 ( .A1(n13510), .A2(n7917), .ZN(n8392) );
  INV_X1 U10681 ( .A(n8393), .ZN(n8394) );
  NAND2_X1 U10682 ( .A1(n12272), .A2(n8424), .ZN(n8397) );
  INV_X1 U10683 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12422) );
  OR2_X1 U10684 ( .A1(n8031), .A2(n12422), .ZN(n8396) );
  NAND2_X1 U10685 ( .A1(n11829), .A2(n10911), .ZN(n8460) );
  NAND2_X1 U10686 ( .A1(n11719), .A2(n13504), .ZN(n10191) );
  AND2_X1 U10687 ( .A1(n7709), .A2(n10191), .ZN(n8398) );
  AND2_X1 U10688 ( .A1(n8460), .A2(n8398), .ZN(n8405) );
  NAND2_X1 U10689 ( .A1(n13510), .A2(n7990), .ZN(n8454) );
  INV_X1 U10690 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8399) );
  OR2_X1 U10691 ( .A1(n6670), .A2(n8399), .ZN(n8404) );
  INV_X1 U10692 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8400) );
  OR2_X1 U10693 ( .A1(n7836), .A2(n8400), .ZN(n8403) );
  INV_X1 U10694 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8401) );
  OR2_X1 U10695 ( .A1(n8428), .A2(n8401), .ZN(n8402) );
  AND3_X1 U10696 ( .A1(n8404), .A2(n8403), .A3(n8402), .ZN(n9243) );
  AOI21_X1 U10697 ( .B1(n8405), .B2(n8454), .A(n9243), .ZN(n8406) );
  AOI21_X1 U10698 ( .B1(n8465), .B2(n8262), .A(n8406), .ZN(n8450) );
  NAND2_X1 U10699 ( .A1(n8465), .A2(n6690), .ZN(n8408) );
  INV_X1 U10700 ( .A(n9243), .ZN(n13430) );
  NAND2_X1 U10701 ( .A1(n13430), .A2(n8262), .ZN(n8407) );
  NAND2_X1 U10702 ( .A1(n8408), .A2(n8407), .ZN(n8449) );
  OR2_X1 U10703 ( .A1(n8031), .A2(n12294), .ZN(n8411) );
  NAND2_X1 U10704 ( .A1(n7684), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U10705 ( .A1(n8412), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8415) );
  INV_X1 U10706 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13321) );
  OR2_X1 U10707 ( .A1(n6672), .A2(n13523), .ZN(n8414) );
  INV_X1 U10708 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13524) );
  OR2_X1 U10709 ( .A1(n7836), .A2(n13524), .ZN(n8413) );
  NAND4_X1 U10710 ( .A1(n8416), .A2(n8415), .A3(n8414), .A4(n8413), .ZN(n13431) );
  AND2_X1 U10711 ( .A1(n13431), .A2(n6690), .ZN(n8417) );
  AOI21_X1 U10712 ( .B1(n13521), .B2(n8262), .A(n8417), .ZN(n8447) );
  NAND2_X1 U10713 ( .A1(n13521), .A2(n6690), .ZN(n8419) );
  NAND2_X1 U10714 ( .A1(n13431), .A2(n8262), .ZN(n8418) );
  NAND2_X1 U10715 ( .A1(n8419), .A2(n8418), .ZN(n8446) );
  OAI22_X1 U10716 ( .A1(n8450), .A2(n8449), .B1(n8447), .B2(n8446), .ZN(n8420)
         );
  NAND2_X1 U10717 ( .A1(n8421), .A2(n8420), .ZN(n8451) );
  NAND2_X1 U10718 ( .A1(n14387), .A2(n8424), .ZN(n8426) );
  OR2_X1 U10719 ( .A1(n8031), .A2(n14552), .ZN(n8425) );
  NAND2_X1 U10720 ( .A1(n7684), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8435) );
  INV_X1 U10721 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8427) );
  OR2_X1 U10722 ( .A1(n8428), .A2(n8427), .ZN(n8434) );
  NAND2_X1 U10723 ( .A1(n8429), .A2(n13321), .ZN(n8430) );
  NAND2_X1 U10724 ( .A1(n13523), .A2(n8430), .ZN(n13538) );
  OR2_X1 U10725 ( .A1(n6672), .A2(n13538), .ZN(n8433) );
  INV_X1 U10726 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13544) );
  OR2_X1 U10727 ( .A1(n7836), .A2(n13544), .ZN(n8432) );
  NAND4_X1 U10728 ( .A1(n8435), .A2(n8434), .A3(n8433), .A4(n8432), .ZN(n13551) );
  AND2_X1 U10729 ( .A1(n13551), .A2(n8262), .ZN(n8436) );
  AOI21_X1 U10730 ( .B1(n13729), .B2(n7990), .A(n8436), .ZN(n8443) );
  NAND2_X1 U10731 ( .A1(n13729), .A2(n7917), .ZN(n8439) );
  NAND2_X1 U10732 ( .A1(n13551), .A2(n8437), .ZN(n8438) );
  NAND2_X1 U10733 ( .A1(n8439), .A2(n8438), .ZN(n8442) );
  NAND2_X1 U10734 ( .A1(n8443), .A2(n8442), .ZN(n8440) );
  XNOR2_X1 U10735 ( .A(n13511), .B(n13510), .ZN(n8464) );
  INV_X1 U10736 ( .A(n8442), .ZN(n8445) );
  INV_X1 U10737 ( .A(n8443), .ZN(n8444) );
  AOI22_X1 U10738 ( .A1(n8447), .A2(n8446), .B1(n8445), .B2(n8444), .ZN(n8448)
         );
  NAND2_X1 U10739 ( .A1(n8464), .A2(n8448), .ZN(n8452) );
  NAND2_X1 U10740 ( .A1(n13511), .A2(n7917), .ZN(n8455) );
  OAI211_X1 U10741 ( .C1(n13511), .C2(n13510), .A(n8455), .B(n8454), .ZN(n8456) );
  NAND2_X1 U10742 ( .A1(n7709), .A2(n13504), .ZN(n8457) );
  OAI211_X1 U10743 ( .C1(n11829), .C2(n10060), .A(n10191), .B(n8457), .ZN(
        n8458) );
  INV_X1 U10744 ( .A(n8458), .ZN(n8459) );
  INV_X1 U10745 ( .A(n11719), .ZN(n10189) );
  NAND2_X1 U10746 ( .A1(n7709), .A2(n10189), .ZN(n9242) );
  OAI21_X1 U10747 ( .B1(n9242), .B2(n13504), .A(n8460), .ZN(n8461) );
  INV_X1 U10748 ( .A(n8464), .ZN(n8494) );
  XNOR2_X1 U10749 ( .A(n13726), .B(n13430), .ZN(n8493) );
  NAND2_X1 U10750 ( .A1(n13742), .A2(n13336), .ZN(n9238) );
  OR2_X1 U10751 ( .A1(n13742), .A2(n13336), .ZN(n8466) );
  NAND2_X1 U10752 ( .A1(n9238), .A2(n8466), .ZN(n9290) );
  INV_X1 U10753 ( .A(n13605), .ZN(n8467) );
  NAND2_X1 U10754 ( .A1(n13747), .A2(n8467), .ZN(n9237) );
  OR2_X1 U10755 ( .A1(n13747), .A2(n8467), .ZN(n8468) );
  NAND2_X1 U10756 ( .A1(n9237), .A2(n8468), .ZN(n9236) );
  XNOR2_X1 U10757 ( .A(n13759), .B(n13606), .ZN(n9235) );
  XNOR2_X1 U10758 ( .A(n13777), .B(n13660), .ZN(n13674) );
  INV_X1 U10759 ( .A(n13435), .ZN(n13375) );
  XNOR2_X1 U10760 ( .A(n13782), .B(n13375), .ZN(n13692) );
  INV_X1 U10761 ( .A(n13436), .ZN(n9230) );
  XNOR2_X1 U10762 ( .A(n13787), .B(n9230), .ZN(n9278) );
  XNOR2_X1 U10763 ( .A(n12201), .B(n13437), .ZN(n12196) );
  NAND2_X1 U10764 ( .A1(n13811), .A2(n8469), .ZN(n9226) );
  OR2_X1 U10765 ( .A1(n13811), .A2(n8469), .ZN(n8470) );
  NAND2_X1 U10766 ( .A1(n9226), .A2(n8470), .ZN(n12117) );
  INV_X1 U10767 ( .A(n13442), .ZN(n11781) );
  XNOR2_X1 U10768 ( .A(n11917), .B(n11781), .ZN(n11906) );
  XNOR2_X1 U10769 ( .A(n12039), .B(n12119), .ZN(n12043) );
  XNOR2_X1 U10770 ( .A(n15286), .B(n13443), .ZN(n11807) );
  NAND2_X1 U10771 ( .A1(n15355), .A2(n11165), .ZN(n9216) );
  OR2_X1 U10772 ( .A1(n15355), .A2(n11165), .ZN(n8471) );
  NAND2_X1 U10773 ( .A1(n9216), .A2(n8471), .ZN(n11638) );
  INV_X1 U10774 ( .A(n13448), .ZN(n11130) );
  XNOR2_X1 U10775 ( .A(n11442), .B(n11130), .ZN(n11436) );
  INV_X1 U10776 ( .A(n13447), .ZN(n11164) );
  OR2_X1 U10777 ( .A1(n15348), .A2(n11164), .ZN(n9215) );
  NAND2_X1 U10778 ( .A1(n15348), .A2(n11164), .ZN(n8472) );
  NAND2_X1 U10779 ( .A1(n9215), .A2(n8472), .ZN(n11355) );
  OAI21_X1 U10780 ( .B1(n7176), .B2(n8474), .A(n10268), .ZN(n10695) );
  OR2_X1 U10781 ( .A1(n8475), .A2(n8476), .ZN(n9209) );
  NAND2_X1 U10782 ( .A1(n8475), .A2(n8476), .ZN(n8477) );
  NAND2_X1 U10783 ( .A1(n9209), .A2(n8477), .ZN(n10253) );
  INV_X1 U10784 ( .A(n10489), .ZN(n15316) );
  INV_X1 U10785 ( .A(n8478), .ZN(n9247) );
  NOR4_X1 U10786 ( .A1(n10695), .A2(n11719), .A3(n10253), .A4(n6663), .ZN(
        n8482) );
  INV_X1 U10787 ( .A(n8479), .ZN(n10778) );
  NAND2_X1 U10788 ( .A1(n10778), .A2(n8480), .ZN(n9210) );
  INV_X1 U10789 ( .A(n8480), .ZN(n15328) );
  NAND2_X1 U10790 ( .A1(n15328), .A2(n8479), .ZN(n8481) );
  XNOR2_X1 U10791 ( .A(n10780), .B(n13450), .ZN(n10855) );
  NAND4_X1 U10792 ( .A1(n8482), .A2(n10762), .A3(n10836), .A4(n10855), .ZN(
        n8483) );
  NOR4_X1 U10793 ( .A1(n11638), .A2(n11436), .A3(n11355), .A4(n8483), .ZN(
        n8484) );
  XNOR2_X1 U10794 ( .A(n11803), .B(n13444), .ZN(n11564) );
  XNOR2_X1 U10795 ( .A(n11484), .B(n13446), .ZN(n11421) );
  NAND4_X1 U10796 ( .A1(n11807), .A2(n8484), .A3(n11564), .A4(n11421), .ZN(
        n8485) );
  NOR4_X1 U10797 ( .A1(n12117), .A2(n11906), .A3(n12043), .A4(n8485), .ZN(
        n8486) );
  XNOR2_X1 U10798 ( .A(n13798), .B(n13438), .ZN(n12154) );
  XNOR2_X1 U10799 ( .A(n13805), .B(n13439), .ZN(n12167) );
  NAND4_X1 U10800 ( .A1(n12196), .A2(n8486), .A3(n12154), .A4(n12167), .ZN(
        n8487) );
  NOR4_X1 U10801 ( .A1(n13674), .A2(n13692), .A3(n9278), .A4(n8487), .ZN(n8488) );
  XNOR2_X1 U10802 ( .A(n13765), .B(n13432), .ZN(n13650) );
  XNOR2_X1 U10803 ( .A(n13772), .B(n13433), .ZN(n13655) );
  NAND4_X1 U10804 ( .A1(n9235), .A2(n8488), .A3(n13650), .A4(n13655), .ZN(
        n8489) );
  NOR4_X1 U10805 ( .A1(n9290), .A2(n9236), .A3(n13602), .A4(n8489), .ZN(n8491)
         );
  XNOR2_X1 U10806 ( .A(n13734), .B(n13575), .ZN(n13560) );
  NAND2_X1 U10807 ( .A1(n13729), .A2(n13551), .ZN(n9293) );
  OR2_X1 U10808 ( .A1(n13729), .A2(n13551), .ZN(n8490) );
  NAND2_X1 U10809 ( .A1(n9293), .A2(n8490), .ZN(n13534) );
  NAND4_X1 U10810 ( .A1(n9294), .A2(n8491), .A3(n13560), .A4(n13534), .ZN(
        n8492) );
  NAND2_X1 U10811 ( .A1(n8503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8500) );
  XNOR2_X1 U10812 ( .A(n8500), .B(n8499), .ZN(n10361) );
  INV_X1 U10813 ( .A(n10361), .ZN(n10352) );
  NAND2_X1 U10814 ( .A1(n10352), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12009) );
  NAND2_X1 U10815 ( .A1(n8510), .A2(n8506), .ZN(n8513) );
  NAND2_X1 U10816 ( .A1(n8513), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8507) );
  MUX2_X1 U10817 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8507), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8509) );
  NAND2_X1 U10818 ( .A1(n8509), .A2(n8508), .ZN(n13846) );
  INV_X1 U10819 ( .A(n8510), .ZN(n8511) );
  NAND2_X1 U10820 ( .A1(n8511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8512) );
  MUX2_X1 U10821 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8512), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8514) );
  NAND2_X1 U10822 ( .A1(n8514), .A2(n8513), .ZN(n13849) );
  NOR2_X1 U10823 ( .A1(n13846), .A2(n13849), .ZN(n8515) );
  NAND2_X1 U10824 ( .A1(n12187), .A2(n8515), .ZN(n10353) );
  NAND2_X1 U10825 ( .A1(n10353), .A2(n10361), .ZN(n9315) );
  INV_X1 U10826 ( .A(n8517), .ZN(n8518) );
  NOR4_X1 U10827 ( .A1(n15311), .A2(n10191), .A3(n12270), .A4(n13661), .ZN(
        n8520) );
  OAI21_X1 U10828 ( .B1(n12009), .B2(n11829), .A(P2_B_REG_SCAN_IN), .ZN(n8519)
         );
  NOR2_X1 U10829 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8525) );
  NOR2_X1 U10830 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n8531) );
  NOR2_X1 U10831 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8530) );
  NOR2_X1 U10832 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8529) );
  NOR2_X1 U10833 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n8534) );
  NAND2_X1 U10834 ( .A1(n8536), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8537) );
  MUX2_X1 U10835 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8537), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n8538) );
  NAND2_X1 U10836 ( .A1(n12292), .A2(n9154), .ZN(n8540) );
  INV_X2 U10837 ( .A(n8684), .ZN(n9163) );
  NAND2_X1 U10838 ( .A1(n9163), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8539) );
  XNOR2_X2 U10839 ( .A(n8546), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10840 ( .A1(n6678), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8558) );
  INV_X1 U10841 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8547) );
  OR2_X1 U10842 ( .A1(n9152), .A2(n8547), .ZN(n8557) );
  INV_X4 U10843 ( .A(n8851), .ZN(n8893) );
  INV_X1 U10844 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14660) );
  NAND2_X1 U10845 ( .A1(n8648), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8659) );
  NOR2_X1 U10846 ( .A1(n8659), .A2(n8658), .ZN(n8671) );
  NAND2_X1 U10847 ( .A1(n8671), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U10848 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n8550) );
  NAND2_X1 U10849 ( .A1(n8741), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8752) );
  INV_X1 U10850 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8751) );
  INV_X1 U10851 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13872) );
  NAND2_X1 U10852 ( .A1(n8872), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U10853 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8880), .ZN(n8890) );
  INV_X1 U10854 ( .A(n8890), .ZN(n8551) );
  NAND2_X1 U10855 ( .A1(n8551), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8892) );
  INV_X1 U10856 ( .A(n8892), .ZN(n8553) );
  AND2_X1 U10857 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n8552) );
  NAND2_X1 U10858 ( .A1(n8553), .A2(n8552), .ZN(n12253) );
  OR2_X1 U10859 ( .A1(n8893), .A2(n12253), .ZN(n8556) );
  INV_X1 U10860 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8554) );
  OR2_X1 U10861 ( .A1(n8873), .A2(n8554), .ZN(n8555) );
  AND4_X1 U10862 ( .A1(n8558), .A2(n8557), .A3(n8556), .A4(n8555), .ZN(n9003)
         );
  XNOR2_X1 U10863 ( .A(n9143), .B(n14070), .ZN(n9189) );
  NAND2_X1 U10864 ( .A1(n14387), .A2(n9154), .ZN(n8560) );
  NAND2_X1 U10865 ( .A1(n9163), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8559) );
  NAND2_X2 U10866 ( .A1(n8560), .A2(n8559), .ZN(n14279) );
  NAND2_X1 U10867 ( .A1(n6678), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8566) );
  INV_X1 U10868 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n14517) );
  OR2_X1 U10869 ( .A1(n9152), .A2(n14517), .ZN(n8565) );
  INV_X1 U10870 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8568) );
  INV_X1 U10871 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8561) );
  OAI21_X1 U10872 ( .B1(n8892), .B2(n8568), .A(n8561), .ZN(n8562) );
  NAND2_X1 U10873 ( .A1(n8562), .A2(n12253), .ZN(n14081) );
  OR2_X1 U10874 ( .A1(n8893), .A2(n14081), .ZN(n8564) );
  NAND2_X1 U10875 ( .A1(n8894), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8563) );
  NAND4_X1 U10876 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(n14095) );
  NAND2_X1 U10877 ( .A1(n9163), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U10878 ( .A1(n6678), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8572) );
  CLKBUF_X3 U10879 ( .A(n8593), .Z(n8889) );
  NAND2_X1 U10880 ( .A1(n8889), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8571) );
  XNOR2_X1 U10881 ( .A(n8892), .B(n8568), .ZN(n14101) );
  OR2_X1 U10882 ( .A1(n8893), .A2(n14101), .ZN(n8570) );
  NAND2_X1 U10883 ( .A1(n8894), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8569) );
  NAND4_X1 U10884 ( .A1(n8572), .A2(n8571), .A3(n8570), .A4(n8569), .ZN(n14069) );
  INV_X1 U10885 ( .A(n14069), .ZN(n12415) );
  NAND2_X1 U10886 ( .A1(n14285), .A2(n12415), .ZN(n8950) );
  OR2_X1 U10887 ( .A1(n14285), .A2(n12415), .ZN(n8573) );
  NAND2_X1 U10888 ( .A1(n8950), .A2(n8573), .ZN(n14090) );
  NAND2_X1 U10889 ( .A1(n8593), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U10890 ( .A1(n8851), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10891 ( .A1(n8796), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U10892 ( .A1(n8600), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8584) );
  INV_X1 U10893 ( .A(n10304), .ZN(n8577) );
  NAND2_X1 U10894 ( .A1(n9164), .A2(n8577), .ZN(n8583) );
  NAND2_X1 U10895 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8578) );
  MUX2_X1 U10896 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8578), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8581) );
  INV_X1 U10897 ( .A(n8579), .ZN(n8580) );
  NAND2_X1 U10898 ( .A1(n8581), .A2(n8580), .ZN(n10594) );
  INV_X1 U10899 ( .A(n10594), .ZN(n10499) );
  OR2_X2 U10900 ( .A1(n13966), .A2(n15124), .ZN(n9010) );
  NAND2_X1 U10901 ( .A1(n8593), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U10902 ( .A1(n8851), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8587) );
  INV_X1 U10903 ( .A(n8754), .ZN(n8796) );
  NAND2_X1 U10904 ( .A1(n8796), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8585) );
  INV_X1 U10905 ( .A(n6664), .ZN(n10716) );
  NAND2_X1 U10906 ( .A1(n10302), .A2(SI_0_), .ZN(n8589) );
  INV_X1 U10907 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U10908 ( .A1(n8589), .A2(n9575), .ZN(n8591) );
  NAND2_X1 U10909 ( .A1(n8591), .A2(n8590), .ZN(n14762) );
  MUX2_X1 U10910 ( .A(n10716), .B(n14762), .S(n6677), .Z(n14256) );
  NAND2_X1 U10911 ( .A1(n14262), .A2(n6858), .ZN(n14253) );
  NAND2_X1 U10912 ( .A1(n14264), .A2(n14253), .ZN(n14252) );
  INV_X1 U10913 ( .A(n15124), .ZN(n14254) );
  OR2_X1 U10914 ( .A1(n13966), .A2(n14254), .ZN(n8592) );
  NAND2_X1 U10915 ( .A1(n14252), .A2(n8592), .ZN(n11184) );
  NAND2_X1 U10916 ( .A1(n8593), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10917 ( .A1(n8851), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U10918 ( .A1(n8796), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8594) );
  NOR2_X1 U10919 ( .A1(n8579), .A2(n8787), .ZN(n8598) );
  MUX2_X1 U10920 ( .A(n8787), .B(n8598), .S(P1_IR_REG_2__SCAN_IN), .Z(n8599)
         );
  AOI22_X1 U10921 ( .A1(n8600), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n10477), 
        .B2(n10724), .ZN(n8603) );
  NAND2_X1 U10922 ( .A1(n8601), .A2(n9164), .ZN(n8602) );
  AND2_X2 U10923 ( .A1(n8603), .A2(n8602), .ZN(n15135) );
  NAND2_X1 U10924 ( .A1(n14267), .A2(n15135), .ZN(n9015) );
  AND2_X2 U10925 ( .A1(n9014), .A2(n9015), .ZN(n11191) );
  INV_X1 U10926 ( .A(n11191), .ZN(n11183) );
  NAND2_X1 U10927 ( .A1(n11184), .A2(n11183), .ZN(n11182) );
  INV_X1 U10928 ( .A(n15135), .ZN(n11188) );
  OR2_X1 U10929 ( .A1(n14267), .A2(n11188), .ZN(n8604) );
  NAND2_X1 U10930 ( .A1(n11182), .A2(n8604), .ZN(n11138) );
  NAND2_X1 U10931 ( .A1(n8605), .A2(n9164), .ZN(n8608) );
  OR2_X1 U10932 ( .A1(n6658), .A2(n8787), .ZN(n8606) );
  XNOR2_X1 U10933 ( .A(n8606), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U10934 ( .A1(n8600), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n10477), 
        .B2(n10511), .ZN(n8607) );
  NAND2_X1 U10935 ( .A1(n8889), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8611) );
  NAND2_X1 U10936 ( .A1(n8894), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U10937 ( .A1(n8796), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8609) );
  INV_X1 U10938 ( .A(n11142), .ZN(n11137) );
  NAND2_X1 U10939 ( .A1(n11138), .A2(n11137), .ZN(n11140) );
  INV_X1 U10940 ( .A(n13965), .ZN(n11193) );
  NAND2_X1 U10941 ( .A1(n6946), .A2(n11193), .ZN(n8613) );
  NAND2_X1 U10942 ( .A1(n8889), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8618) );
  INV_X1 U10943 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11178) );
  OR2_X1 U10944 ( .A1(n6679), .A2(n11178), .ZN(n8617) );
  XNOR2_X1 U10945 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11172) );
  OR2_X1 U10946 ( .A1(n8893), .A2(n11172), .ZN(n8616) );
  INV_X1 U10947 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8614) );
  OR2_X1 U10948 ( .A1(n8873), .A2(n8614), .ZN(n8615) );
  NAND2_X1 U10949 ( .A1(n10311), .A2(n9154), .ZN(n8623) );
  NAND2_X1 U10950 ( .A1(n6658), .A2(n8619), .ZN(n8627) );
  NAND2_X1 U10951 ( .A1(n8627), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8621) );
  XNOR2_X1 U10952 ( .A(n8621), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13991) );
  AOI22_X1 U10953 ( .A1(n9163), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n10477), 
        .B2(n13991), .ZN(n8622) );
  OAI21_X1 U10954 ( .B1(n11170), .B2(n11145), .A(n15149), .ZN(n8625) );
  NAND2_X1 U10955 ( .A1(n11170), .A2(n11145), .ZN(n8624) );
  NAND2_X1 U10956 ( .A1(n8625), .A2(n8624), .ZN(n15095) );
  NAND2_X1 U10957 ( .A1(n8626), .A2(n9164), .ZN(n8630) );
  NAND2_X1 U10958 ( .A1(n8638), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8628) );
  XNOR2_X1 U10959 ( .A(n8628), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U10960 ( .A1(n9163), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10477), 
        .B2(n10531), .ZN(n8629) );
  NAND2_X1 U10961 ( .A1(n8630), .A2(n8629), .ZN(n11519) );
  NAND2_X1 U10962 ( .A1(n8796), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U10963 ( .A1(n8889), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8634) );
  AOI21_X1 U10964 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8631) );
  NOR2_X1 U10965 ( .A1(n8631), .A2(n8648), .ZN(n15104) );
  NAND2_X1 U10966 ( .A1(n8851), .A2(n15104), .ZN(n8633) );
  NAND2_X1 U10967 ( .A1(n8894), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8632) );
  NAND4_X1 U10968 ( .A1(n8635), .A2(n8634), .A3(n8633), .A4(n8632), .ZN(n13963) );
  XNOR2_X1 U10969 ( .A(n11519), .B(n13963), .ZN(n15097) );
  INV_X1 U10970 ( .A(n15097), .ZN(n15094) );
  NAND2_X1 U10971 ( .A1(n15095), .A2(n15094), .ZN(n8637) );
  OR2_X1 U10972 ( .A1(n11519), .A2(n13963), .ZN(n8636) );
  NAND2_X1 U10973 ( .A1(n8637), .A2(n8636), .ZN(n11063) );
  NAND2_X1 U10974 ( .A1(n10340), .A2(n9154), .ZN(n8647) );
  INV_X1 U10975 ( .A(n8638), .ZN(n8640) );
  NAND2_X1 U10976 ( .A1(n8640), .A2(n8639), .ZN(n8642) );
  NAND2_X1 U10977 ( .A1(n8642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8641) );
  MUX2_X1 U10978 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8641), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n8645) );
  INV_X1 U10979 ( .A(n8642), .ZN(n8644) );
  NAND2_X1 U10980 ( .A1(n8644), .A2(n8643), .ZN(n8667) );
  AND2_X1 U10981 ( .A1(n8645), .A2(n8667), .ZN(n10533) );
  AOI22_X1 U10982 ( .A1(n9163), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10477), 
        .B2(n10533), .ZN(n8646) );
  NAND2_X1 U10983 ( .A1(n8647), .A2(n8646), .ZN(n11594) );
  NAND2_X1 U10984 ( .A1(n6678), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U10985 ( .A1(n8889), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8651) );
  OAI21_X1 U10986 ( .B1(n8648), .B2(P1_REG3_REG_6__SCAN_IN), .A(n8659), .ZN(
        n11597) );
  OR2_X1 U10987 ( .A1(n8893), .A2(n11597), .ZN(n8650) );
  NAND2_X1 U10988 ( .A1(n8894), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8649) );
  NAND4_X1 U10989 ( .A1(n8652), .A2(n8651), .A3(n8650), .A4(n8649), .ZN(n13962) );
  XNOR2_X1 U10990 ( .A(n11594), .B(n13962), .ZN(n11071) );
  INV_X1 U10991 ( .A(n11071), .ZN(n11062) );
  NAND2_X1 U10992 ( .A1(n11063), .A2(n11062), .ZN(n8654) );
  OR2_X1 U10993 ( .A1(n11594), .A2(n13962), .ZN(n8653) );
  NAND2_X1 U10994 ( .A1(n8654), .A2(n8653), .ZN(n15079) );
  NAND2_X1 U10995 ( .A1(n10345), .A2(n9154), .ZN(n8657) );
  NAND2_X1 U10996 ( .A1(n8667), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8655) );
  XNOR2_X1 U10997 ( .A(n8655), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U10998 ( .A1(n9163), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10477), 
        .B2(n10535), .ZN(n8656) );
  NAND2_X1 U10999 ( .A1(n8657), .A2(n8656), .ZN(n11773) );
  NAND2_X1 U11000 ( .A1(n6678), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U11001 ( .A1(n8889), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8663) );
  AND2_X1 U11002 ( .A1(n8659), .A2(n8658), .ZN(n8660) );
  OR2_X1 U11003 ( .A1(n8660), .A2(n8671), .ZN(n11777) );
  OR2_X1 U11004 ( .A1(n8893), .A2(n11777), .ZN(n8662) );
  NAND2_X1 U11005 ( .A1(n8894), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8661) );
  NAND4_X1 U11006 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), .ZN(n13961) );
  INV_X1 U11007 ( .A(n13961), .ZN(n11771) );
  XNOR2_X1 U11008 ( .A(n11773), .B(n11771), .ZN(n15081) );
  NAND2_X1 U11009 ( .A1(n15079), .A2(n15081), .ZN(n8666) );
  OR2_X1 U11010 ( .A1(n11773), .A2(n13961), .ZN(n8665) );
  NAND2_X1 U11011 ( .A1(n8666), .A2(n8665), .ZN(n11370) );
  NAND2_X1 U11012 ( .A1(n10350), .A2(n9154), .ZN(n8670) );
  NAND2_X1 U11013 ( .A1(n8678), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8668) );
  XNOR2_X1 U11014 ( .A(n8668), .B(P1_IR_REG_8__SCAN_IN), .ZN(n14012) );
  AOI22_X1 U11015 ( .A1(n9163), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n14012), 
        .B2(n10477), .ZN(n8669) );
  NAND2_X1 U11016 ( .A1(n6678), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U11017 ( .A1(n8889), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8675) );
  OR2_X1 U11018 ( .A1(n8671), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U11019 ( .A1(n8689), .A2(n8672), .ZN(n11876) );
  OR2_X1 U11020 ( .A1(n8893), .A2(n11876), .ZN(n8674) );
  NAND2_X1 U11021 ( .A1(n8894), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8673) );
  NAND4_X1 U11022 ( .A1(n8676), .A2(n8675), .A3(n8674), .A4(n8673), .ZN(n13960) );
  INV_X1 U11023 ( .A(n13960), .ZN(n8921) );
  OR2_X1 U11024 ( .A1(n15177), .A2(n13960), .ZN(n8677) );
  NAND2_X1 U11025 ( .A1(n10394), .A2(n9154), .ZN(n8687) );
  NAND2_X1 U11026 ( .A1(n8680), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8679) );
  MUX2_X1 U11027 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8679), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n8683) );
  INV_X1 U11028 ( .A(n8680), .ZN(n8682) );
  INV_X1 U11029 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11030 ( .A1(n8682), .A2(n8681), .ZN(n8707) );
  NAND2_X1 U11031 ( .A1(n8683), .A2(n8707), .ZN(n10638) );
  OAI22_X1 U11032 ( .A1(n10638), .A2(n8848), .B1(n8684), .B2(n10395), .ZN(
        n8685) );
  INV_X1 U11033 ( .A(n8685), .ZN(n8686) );
  NAND2_X1 U11034 ( .A1(n6678), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U11035 ( .A1(n8889), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U11036 ( .A1(n8689), .A2(n8688), .ZN(n8690) );
  NAND2_X1 U11037 ( .A1(n8698), .A2(n8690), .ZN(n12032) );
  OR2_X1 U11038 ( .A1(n8893), .A2(n12032), .ZN(n8692) );
  NAND2_X1 U11039 ( .A1(n8894), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8691) );
  NAND4_X1 U11040 ( .A1(n8694), .A2(n8693), .A3(n8692), .A4(n8691), .ZN(n14927) );
  XNOR2_X1 U11041 ( .A(n12029), .B(n14927), .ZN(n9178) );
  NAND2_X1 U11042 ( .A1(n10437), .A2(n9154), .ZN(n8697) );
  NAND2_X1 U11043 ( .A1(n8707), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8695) );
  XNOR2_X1 U11044 ( .A(n8695), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U11045 ( .A1(n10745), .A2(n10477), .B1(n9163), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U11046 ( .A1(n6678), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U11047 ( .A1(n8889), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U11048 ( .A1(n8698), .A2(n10645), .ZN(n8699) );
  NAND2_X1 U11049 ( .A1(n8725), .A2(n8699), .ZN(n14937) );
  OR2_X1 U11050 ( .A1(n8893), .A2(n14937), .ZN(n8701) );
  NAND2_X1 U11051 ( .A1(n8894), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8700) );
  NAND4_X1 U11052 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n14943) );
  INV_X1 U11053 ( .A(n14943), .ZN(n12209) );
  OR2_X1 U11054 ( .A1(n14925), .A2(n12209), .ZN(n8926) );
  NAND2_X1 U11055 ( .A1(n14925), .A2(n12209), .ZN(n8704) );
  NAND2_X1 U11056 ( .A1(n8926), .A2(n8704), .ZN(n11496) );
  NAND2_X1 U11057 ( .A1(n11492), .A2(n11496), .ZN(n8706) );
  OR2_X1 U11058 ( .A1(n14925), .A2(n14943), .ZN(n8705) );
  NAND2_X1 U11059 ( .A1(n8706), .A2(n8705), .ZN(n11539) );
  NAND2_X1 U11060 ( .A1(n10466), .A2(n9154), .ZN(n8712) );
  INV_X1 U11061 ( .A(n8707), .ZN(n8709) );
  INV_X1 U11062 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11063 ( .A1(n8709), .A2(n8708), .ZN(n8710) );
  NAND2_X1 U11064 ( .A1(n8710), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8721) );
  XNOR2_X1 U11065 ( .A(n8721), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U11066 ( .A1(n11022), .A2(n10477), .B1(n9163), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n8711) );
  NAND2_X1 U11067 ( .A1(n8889), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8717) );
  INV_X1 U11068 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8713) );
  XNOR2_X1 U11069 ( .A(n8725), .B(n8713), .ZN(n14949) );
  OR2_X1 U11070 ( .A1(n8893), .A2(n14949), .ZN(n8716) );
  NAND2_X1 U11071 ( .A1(n8894), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11072 ( .A1(n6678), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8714) );
  NAND4_X1 U11073 ( .A1(n8717), .A2(n8716), .A3(n8715), .A4(n8714), .ZN(n13959) );
  XNOR2_X1 U11074 ( .A(n12216), .B(n13959), .ZN(n11536) );
  INV_X1 U11075 ( .A(n11536), .ZN(n11540) );
  NAND2_X1 U11076 ( .A1(n11539), .A2(n11540), .ZN(n8719) );
  OR2_X1 U11077 ( .A1(n12216), .A2(n13959), .ZN(n8718) );
  NAND2_X1 U11078 ( .A1(n8719), .A2(n8718), .ZN(n11752) );
  NAND2_X1 U11079 ( .A1(n10558), .A2(n9154), .ZN(n8724) );
  INV_X1 U11080 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U11081 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  NAND2_X1 U11082 ( .A1(n8722), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8734) );
  XNOR2_X1 U11083 ( .A(n8734), .B(P1_IR_REG_12__SCAN_IN), .ZN(n15043) );
  AOI22_X1 U11084 ( .A1(n15043), .A2(n10477), .B1(n9163), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U11085 ( .A1(n6678), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11086 ( .A1(n8889), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8730) );
  INV_X1 U11087 ( .A(n8725), .ZN(n8726) );
  AOI21_X1 U11088 ( .B1(n8726), .B2(P1_REG3_REG_11__SCAN_IN), .A(
        P1_REG3_REG_12__SCAN_IN), .ZN(n8727) );
  OR2_X1 U11089 ( .A1(n8727), .A2(n8741), .ZN(n12231) );
  OR2_X1 U11090 ( .A1(n8893), .A2(n12231), .ZN(n8729) );
  NAND2_X1 U11091 ( .A1(n8894), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8728) );
  NAND4_X1 U11092 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n8728), .ZN(n14978) );
  XNOR2_X1 U11093 ( .A(n12227), .B(n14978), .ZN(n11751) );
  INV_X1 U11094 ( .A(n11751), .ZN(n11754) );
  OR2_X1 U11095 ( .A1(n12227), .A2(n14978), .ZN(n8732) );
  NAND2_X1 U11096 ( .A1(n10617), .A2(n9154), .ZN(n8740) );
  INV_X1 U11097 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11098 ( .A1(n8734), .A2(n8733), .ZN(n8735) );
  NAND2_X1 U11099 ( .A1(n8735), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8737) );
  INV_X1 U11100 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U11101 ( .A1(n8737), .A2(n8736), .ZN(n8747) );
  OR2_X1 U11102 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  AOI22_X1 U11103 ( .A1(n11024), .A2(n10477), .B1(n9163), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U11104 ( .A1(n6678), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U11105 ( .A1(n8889), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8745) );
  OR2_X1 U11106 ( .A1(n8741), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U11107 ( .A1(n8752), .A2(n8742), .ZN(n14802) );
  OR2_X1 U11108 ( .A1(n8893), .A2(n14802), .ZN(n8744) );
  NAND2_X1 U11109 ( .A1(n8894), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8743) );
  NAND4_X1 U11110 ( .A1(n8746), .A2(n8745), .A3(n8744), .A4(n8743), .ZN(n13958) );
  XNOR2_X1 U11111 ( .A(n14981), .B(n14911), .ZN(n14811) );
  INV_X1 U11112 ( .A(n11943), .ZN(n8759) );
  NAND2_X1 U11113 ( .A1(n10754), .A2(n9154), .ZN(n8750) );
  NAND2_X1 U11114 ( .A1(n8747), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8748) );
  XNOR2_X1 U11115 ( .A(n8748), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U11116 ( .A1(n11343), .A2(n10477), .B1(n9163), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U11117 ( .A1(n8894), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8758) );
  INV_X1 U11118 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11922) );
  OR2_X1 U11119 ( .A1(n9152), .A2(n11922), .ZN(n8757) );
  NAND2_X1 U11120 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  NAND2_X1 U11121 ( .A1(n8767), .A2(n8753), .ZN(n14924) );
  OR2_X1 U11122 ( .A1(n14924), .A2(n8893), .ZN(n8756) );
  INV_X1 U11123 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11344) );
  OR2_X1 U11124 ( .A1(n6679), .A2(n11344), .ZN(n8755) );
  OR2_X1 U11125 ( .A1(n14971), .A2(n12310), .ZN(n9069) );
  NAND2_X1 U11126 ( .A1(n14971), .A2(n12310), .ZN(n9064) );
  AND2_X2 U11127 ( .A1(n9069), .A2(n9064), .ZN(n11944) );
  NAND2_X1 U11128 ( .A1(n14971), .A2(n14955), .ZN(n8760) );
  NAND2_X1 U11129 ( .A1(n10990), .A2(n9154), .ZN(n8765) );
  NAND2_X1 U11130 ( .A1(n8761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8762) );
  MUX2_X1 U11131 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8762), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n8763) );
  OR2_X1 U11132 ( .A1(n8761), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n8775) );
  AOI22_X1 U11133 ( .A1(n9163), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10477), 
        .B2(n11928), .ZN(n8764) );
  AND2_X1 U11134 ( .A1(n8767), .A2(n8766), .ZN(n8768) );
  OR2_X1 U11135 ( .A1(n8768), .A2(n8780), .ZN(n14963) );
  NAND2_X1 U11136 ( .A1(n8894), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U11137 ( .A1(n6678), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8769) );
  AND2_X1 U11138 ( .A1(n8770), .A2(n8769), .ZN(n8772) );
  NAND2_X1 U11139 ( .A1(n8889), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8771) );
  OAI211_X1 U11140 ( .C1(n14963), .C2(n8893), .A(n8772), .B(n8771), .ZN(n13957) );
  INV_X1 U11141 ( .A(n13957), .ZN(n14908) );
  NAND2_X1 U11142 ( .A1(n14354), .A2(n14908), .ZN(n9078) );
  NAND2_X1 U11143 ( .A1(n9077), .A2(n9078), .ZN(n12092) );
  OR2_X1 U11144 ( .A1(n14354), .A2(n13957), .ZN(n8773) );
  NAND2_X1 U11145 ( .A1(n11135), .A2(n9154), .ZN(n8779) );
  NAND2_X1 U11146 ( .A1(n8775), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8774) );
  MUX2_X1 U11147 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8774), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8777) );
  NOR2_X1 U11148 ( .A1(n8775), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n8790) );
  INV_X1 U11149 ( .A(n8790), .ZN(n8776) );
  NAND2_X1 U11150 ( .A1(n8777), .A2(n8776), .ZN(n12060) );
  INV_X1 U11151 ( .A(n12060), .ZN(n12064) );
  AOI22_X1 U11152 ( .A1(n9163), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10477), 
        .B2(n12064), .ZN(n8778) );
  NOR2_X1 U11153 ( .A1(n8780), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8781) );
  OR2_X1 U11154 ( .A1(n8794), .A2(n8781), .ZN(n13899) );
  AOI22_X1 U11155 ( .A1(n8889), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6678), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n8783) );
  NAND2_X1 U11156 ( .A1(n8894), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8782) );
  OAI211_X1 U11157 ( .C1(n13899), .C2(n8893), .A(n8783), .B(n8782), .ZN(n14953) );
  INV_X1 U11158 ( .A(n14953), .ZN(n12328) );
  NAND2_X1 U11159 ( .A1(n12106), .A2(n12328), .ZN(n8934) );
  OR2_X1 U11160 ( .A1(n12106), .A2(n12328), .ZN(n8784) );
  AND2_X1 U11161 ( .A1(n14967), .A2(n12328), .ZN(n8785) );
  AOI21_X1 U11162 ( .B1(n12097), .B2(n12098), .A(n8785), .ZN(n12128) );
  NAND2_X1 U11163 ( .A1(n11226), .A2(n9154), .ZN(n8793) );
  NOR2_X1 U11164 ( .A1(n8790), .A2(n8787), .ZN(n8786) );
  MUX2_X1 U11165 ( .A(n8787), .B(n8786), .S(P1_IR_REG_17__SCAN_IN), .Z(n8788)
         );
  INV_X1 U11166 ( .A(n8788), .ZN(n8791) );
  INV_X1 U11167 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U11168 ( .A1(n8790), .A2(n8789), .ZN(n8799) );
  AND2_X1 U11169 ( .A1(n8791), .A2(n8799), .ZN(n14027) );
  AOI22_X1 U11170 ( .A1(n9163), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n14027), 
        .B2(n10477), .ZN(n8792) );
  OR2_X1 U11171 ( .A1(n8794), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11172 ( .A1(n8803), .A2(n8795), .ZN(n13910) );
  AOI22_X1 U11173 ( .A1(n8889), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n6678), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U11174 ( .A1(n8894), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U11175 ( .C1(n13910), .C2(n8893), .A(n8798), .B(n8797), .ZN(n14237) );
  INV_X1 U11176 ( .A(n14237), .ZN(n13943) );
  AND2_X1 U11177 ( .A1(n13912), .A2(n14237), .ZN(n9087) );
  INV_X1 U11178 ( .A(n9087), .ZN(n9182) );
  NAND2_X1 U11179 ( .A1(n11547), .A2(n9154), .ZN(n8802) );
  NAND2_X1 U11180 ( .A1(n8799), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8800) );
  XNOR2_X1 U11181 ( .A(n8800), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14041) );
  AOI22_X1 U11182 ( .A1(n9163), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10477), 
        .B2(n14041), .ZN(n8801) );
  NAND2_X1 U11183 ( .A1(n8803), .A2(n13940), .ZN(n8804) );
  AND2_X1 U11184 ( .A1(n8818), .A2(n8804), .ZN(n14245) );
  NAND2_X1 U11185 ( .A1(n14245), .A2(n8851), .ZN(n8809) );
  INV_X1 U11186 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14029) );
  NAND2_X1 U11187 ( .A1(n6678), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U11188 ( .A1(n8894), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8805) );
  OAI211_X1 U11189 ( .C1(n9152), .C2(n14029), .A(n8806), .B(n8805), .ZN(n8807)
         );
  INV_X1 U11190 ( .A(n8807), .ZN(n8808) );
  NAND2_X1 U11191 ( .A1(n8809), .A2(n8808), .ZN(n14222) );
  NAND2_X1 U11192 ( .A1(n8810), .A2(n8938), .ZN(n14218) );
  NAND2_X1 U11193 ( .A1(n8901), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8815) );
  AOI22_X1 U11194 ( .A1(n9163), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11942), 
        .B2(n10477), .ZN(n8816) );
  AND2_X1 U11195 ( .A1(n8818), .A2(n13872), .ZN(n8819) );
  NOR2_X1 U11196 ( .A1(n8819), .A2(n8827), .ZN(n14225) );
  INV_X1 U11197 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14635) );
  NAND2_X1 U11198 ( .A1(n6678), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U11199 ( .A1(n8889), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8820) );
  OAI211_X1 U11200 ( .C1(n14635), .C2(n8873), .A(n8821), .B(n8820), .ZN(n8822)
         );
  AOI21_X1 U11201 ( .B1(n14225), .B2(n8851), .A(n8822), .ZN(n14199) );
  NAND2_X1 U11202 ( .A1(n14229), .A2(n14199), .ZN(n9101) );
  NAND2_X1 U11203 ( .A1(n14218), .A2(n14217), .ZN(n8824) );
  INV_X1 U11204 ( .A(n14199), .ZN(n14238) );
  OR2_X1 U11205 ( .A1(n14229), .A2(n14238), .ZN(n8823) );
  NAND2_X1 U11206 ( .A1(n14759), .A2(n9154), .ZN(n8826) );
  NAND2_X1 U11207 ( .A1(n9163), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8825) );
  AND2_X2 U11208 ( .A1(n8826), .A2(n8825), .ZN(n14212) );
  NOR2_X1 U11209 ( .A1(n8827), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8828) );
  NOR2_X1 U11210 ( .A1(n8838), .A2(n8828), .ZN(n14205) );
  NAND2_X1 U11211 ( .A1(n14205), .A2(n8851), .ZN(n8833) );
  INV_X1 U11212 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14600) );
  NAND2_X1 U11213 ( .A1(n6678), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U11214 ( .A1(n8894), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8829) );
  OAI211_X1 U11215 ( .C1(n9152), .C2(n14600), .A(n8830), .B(n8829), .ZN(n8831)
         );
  INV_X1 U11216 ( .A(n8831), .ZN(n8832) );
  XNOR2_X1 U11217 ( .A(n14329), .B(n14221), .ZN(n14209) );
  INV_X1 U11218 ( .A(n14209), .ZN(n8834) );
  OR2_X1 U11219 ( .A1(n14212), .A2(n14221), .ZN(n8835) );
  NAND2_X1 U11220 ( .A1(n11832), .A2(n9154), .ZN(n8837) );
  NAND2_X1 U11221 ( .A1(n9163), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8836) );
  NOR2_X1 U11222 ( .A1(n8838), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8839) );
  OR2_X1 U11223 ( .A1(n8849), .A2(n8839), .ZN(n14188) );
  INV_X1 U11224 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U11225 ( .A1(n6678), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U11226 ( .A1(n8894), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8840) );
  OAI211_X1 U11227 ( .C1(n9152), .C2(n8842), .A(n8841), .B(n8840), .ZN(n8843)
         );
  INV_X1 U11228 ( .A(n8843), .ZN(n8844) );
  INV_X1 U11229 ( .A(n14175), .ZN(n14200) );
  XNOR2_X1 U11230 ( .A(n14324), .B(n14200), .ZN(n14184) );
  INV_X1 U11231 ( .A(n14184), .ZN(n14194) );
  OR2_X1 U11232 ( .A1(n14324), .A2(n14175), .ZN(n8845) );
  OR2_X1 U11233 ( .A1(n8846), .A2(n10286), .ZN(n8847) );
  XNOR2_X1 U11234 ( .A(n8847), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14399) );
  OR2_X1 U11235 ( .A1(n8849), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8850) );
  AND2_X1 U11236 ( .A1(n8850), .A2(n8862), .ZN(n14176) );
  NAND2_X1 U11237 ( .A1(n14176), .A2(n8851), .ZN(n8857) );
  INV_X1 U11238 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U11239 ( .A1(n6678), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U11240 ( .A1(n8894), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8852) );
  OAI211_X1 U11241 ( .C1(n9152), .C2(n8854), .A(n8853), .B(n8852), .ZN(n8855)
         );
  INV_X1 U11242 ( .A(n8855), .ZN(n8856) );
  NAND2_X1 U11243 ( .A1(n8857), .A2(n8856), .ZN(n14156) );
  XNOR2_X1 U11244 ( .A(n7369), .B(n13881), .ZN(n14170) );
  INV_X1 U11245 ( .A(n14170), .ZN(n14172) );
  NAND2_X1 U11246 ( .A1(n14171), .A2(n14172), .ZN(n8859) );
  OR2_X1 U11247 ( .A1(n12364), .A2(n14156), .ZN(n8858) );
  NAND2_X1 U11248 ( .A1(n12007), .A2(n9154), .ZN(n8861) );
  NAND2_X1 U11249 ( .A1(n9163), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U11250 ( .A1(n6678), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8868) );
  NAND2_X1 U11251 ( .A1(n8889), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8867) );
  INV_X1 U11252 ( .A(n8862), .ZN(n8864) );
  INV_X1 U11253 ( .A(n8872), .ZN(n8863) );
  OAI21_X1 U11254 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8864), .A(n8863), .ZN(
        n14160) );
  OR2_X1 U11255 ( .A1(n8893), .A2(n14160), .ZN(n8866) );
  NAND2_X1 U11256 ( .A1(n8894), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8865) );
  NAND4_X1 U11257 ( .A1(n8868), .A2(n8867), .A3(n8866), .A4(n8865), .ZN(n14174) );
  NAND2_X1 U11258 ( .A1(n12151), .A2(n9154), .ZN(n8870) );
  NAND2_X1 U11259 ( .A1(n9163), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U11260 ( .A1(n6678), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8877) );
  INV_X1 U11261 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14530) );
  OR2_X1 U11262 ( .A1(n9152), .A2(n14530), .ZN(n8876) );
  OAI21_X1 U11263 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8872), .A(n8871), .ZN(
        n14146) );
  OR2_X1 U11264 ( .A1(n8893), .A2(n14146), .ZN(n8875) );
  INV_X1 U11265 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14639) );
  OR2_X1 U11266 ( .A1(n8873), .A2(n14639), .ZN(n8874) );
  NAND4_X1 U11267 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .ZN(n14157) );
  INV_X1 U11268 ( .A(n14157), .ZN(n8945) );
  XNOR2_X1 U11269 ( .A(n14308), .B(n8945), .ZN(n14142) );
  NAND2_X1 U11270 ( .A1(n13847), .A2(n9154), .ZN(n8879) );
  NAND2_X1 U11271 ( .A1(n9163), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8878) );
  NAND2_X2 U11272 ( .A1(n8879), .A2(n8878), .ZN(n14131) );
  NAND2_X1 U11273 ( .A1(n6678), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U11274 ( .A1(n8889), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8883) );
  OAI21_X1 U11275 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8880), .A(n8890), .ZN(
        n14126) );
  OR2_X1 U11276 ( .A1(n8893), .A2(n14126), .ZN(n8882) );
  NAND2_X1 U11277 ( .A1(n8894), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8881) );
  NAND4_X1 U11278 ( .A1(n8884), .A2(n8883), .A3(n8882), .A4(n8881), .ZN(n13955) );
  NAND2_X1 U11279 ( .A1(n14131), .A2(n13955), .ZN(n8886) );
  OR2_X1 U11280 ( .A1(n14131), .A2(n13955), .ZN(n8885) );
  NAND2_X1 U11281 ( .A1(n8886), .A2(n8885), .ZN(n14123) );
  NAND2_X1 U11282 ( .A1(n13843), .A2(n9154), .ZN(n8888) );
  NAND2_X1 U11283 ( .A1(n9163), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U11284 ( .A1(n6678), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U11285 ( .A1(n8889), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8897) );
  INV_X1 U11286 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14599) );
  NAND2_X1 U11287 ( .A1(n8890), .A2(n14599), .ZN(n8891) );
  NAND2_X1 U11288 ( .A1(n8892), .A2(n8891), .ZN(n14113) );
  OR2_X1 U11289 ( .A1(n8893), .A2(n14113), .ZN(n8896) );
  NAND2_X1 U11290 ( .A1(n8894), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8895) );
  NAND4_X1 U11291 ( .A1(n8898), .A2(n8897), .A3(n8896), .A4(n8895), .ZN(n14094) );
  INV_X1 U11292 ( .A(n14094), .ZN(n13857) );
  XNOR2_X1 U11293 ( .A(n14112), .B(n13857), .ZN(n14107) );
  AND2_X1 U11294 ( .A1(n14112), .A2(n14094), .ZN(n8899) );
  INV_X1 U11295 ( .A(n14095), .ZN(n8960) );
  NAND2_X1 U11296 ( .A1(n14279), .A2(n8960), .ZN(n8951) );
  OR2_X1 U11297 ( .A1(n14279), .A2(n8960), .ZN(n8900) );
  NOR2_X1 U11298 ( .A1(n14076), .A2(n14077), .ZN(n14075) );
  NAND2_X1 U11299 ( .A1(n6752), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U11300 ( .A1(n14400), .A2(n14206), .ZN(n9001) );
  NAND2_X1 U11301 ( .A1(n8905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U11302 ( .A1(n6941), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8908) );
  OAI21_X1 U11303 ( .B1(n9001), .B2(n10206), .A(n10223), .ZN(n11120) );
  INV_X1 U11304 ( .A(n9170), .ZN(n8909) );
  NAND2_X1 U11305 ( .A1(n8909), .A2(n11942), .ZN(n14345) );
  NAND2_X1 U11306 ( .A1(n11189), .A2(n9014), .ZN(n11143) );
  NAND2_X1 U11307 ( .A1(n11143), .A2(n11142), .ZN(n11141) );
  NAND2_X1 U11308 ( .A1(n11193), .A2(n11150), .ZN(n8910) );
  NAND2_X1 U11309 ( .A1(n11141), .A2(n8910), .ZN(n11175) );
  NAND2_X1 U11310 ( .A1(n15149), .A2(n13964), .ZN(n8911) );
  NAND2_X1 U11311 ( .A1(n11175), .A2(n8911), .ZN(n8913) );
  OR2_X1 U11312 ( .A1(n15149), .A2(n13964), .ZN(n8912) );
  NAND2_X1 U11313 ( .A1(n8913), .A2(n8912), .ZN(n15096) );
  NAND2_X1 U11314 ( .A1(n15096), .A2(n15097), .ZN(n8915) );
  INV_X1 U11315 ( .A(n13963), .ZN(n11513) );
  NAND2_X1 U11316 ( .A1(n11519), .A2(n11513), .ZN(n8914) );
  NAND2_X1 U11317 ( .A1(n8915), .A2(n8914), .ZN(n11070) );
  NAND2_X1 U11318 ( .A1(n11070), .A2(n11071), .ZN(n8918) );
  INV_X1 U11319 ( .A(n13962), .ZN(n8916) );
  NAND2_X1 U11320 ( .A1(n11594), .A2(n8916), .ZN(n8917) );
  AND2_X1 U11321 ( .A1(n11773), .A2(n11771), .ZN(n8919) );
  OR2_X1 U11322 ( .A1(n11773), .A2(n11771), .ZN(n8920) );
  INV_X1 U11323 ( .A(n11371), .ZN(n8923) );
  NOR2_X1 U11324 ( .A1(n15177), .A2(n8921), .ZN(n8922) );
  NAND2_X1 U11325 ( .A1(n15066), .A2(n9178), .ZN(n8925) );
  INV_X1 U11326 ( .A(n14927), .ZN(n12027) );
  NAND2_X1 U11327 ( .A1(n12029), .A2(n12027), .ZN(n8924) );
  NAND2_X1 U11328 ( .A1(n11493), .A2(n8926), .ZN(n11537) );
  NAND2_X1 U11329 ( .A1(n11537), .A2(n11536), .ZN(n8928) );
  INV_X1 U11330 ( .A(n13959), .ZN(n12230) );
  OR2_X1 U11331 ( .A1(n12216), .A2(n12230), .ZN(n8927) );
  NAND2_X1 U11332 ( .A1(n8928), .A2(n8927), .ZN(n11753) );
  NAND2_X1 U11333 ( .A1(n11753), .A2(n11751), .ZN(n8930) );
  INV_X1 U11334 ( .A(n14978), .ZN(n12246) );
  OR2_X1 U11335 ( .A1(n12227), .A2(n12246), .ZN(n8929) );
  NAND2_X1 U11336 ( .A1(n14810), .A2(n7267), .ZN(n8932) );
  OR2_X1 U11337 ( .A1(n14981), .A2(n14911), .ZN(n8931) );
  NAND2_X1 U11338 ( .A1(n8932), .A2(n8931), .ZN(n11938) );
  AND2_X1 U11339 ( .A1(n13912), .A2(n13943), .ZN(n8936) );
  OR2_X1 U11340 ( .A1(n13912), .A2(n13943), .ZN(n8935) );
  NAND2_X1 U11341 ( .A1(n14236), .A2(n14235), .ZN(n8940) );
  INV_X1 U11342 ( .A(n14222), .ZN(n13907) );
  OR2_X1 U11343 ( .A1(n14342), .A2(n13907), .ZN(n8939) );
  INV_X1 U11344 ( .A(n14221), .ZN(n13956) );
  NAND2_X1 U11345 ( .A1(n14212), .A2(n13956), .ZN(n8941) );
  NAND2_X1 U11346 ( .A1(n14202), .A2(n8941), .ZN(n14185) );
  OR2_X1 U11347 ( .A1(n14324), .A2(n14200), .ZN(n8942) );
  NAND2_X1 U11348 ( .A1(n12364), .A2(n13881), .ZN(n8943) );
  XNOR2_X1 U11349 ( .A(n14313), .B(n14174), .ZN(n14154) );
  INV_X1 U11350 ( .A(n14174), .ZN(n14137) );
  NAND2_X1 U11351 ( .A1(n14313), .A2(n14137), .ZN(n8944) );
  OR2_X1 U11352 ( .A1(n14308), .A2(n8945), .ZN(n8946) );
  INV_X1 U11353 ( .A(n13955), .ZN(n14138) );
  NAND2_X1 U11354 ( .A1(n14131), .A2(n14138), .ZN(n8947) );
  NAND2_X1 U11355 ( .A1(n8948), .A2(n8947), .ZN(n14110) );
  NAND2_X1 U11356 ( .A1(n14112), .A2(n13857), .ZN(n8949) );
  NAND2_X1 U11357 ( .A1(n14400), .A2(n11942), .ZN(n8952) );
  NAND2_X1 U11358 ( .A1(n8961), .A2(n14757), .ZN(n9153) );
  NAND2_X1 U11359 ( .A1(n8953), .A2(n14206), .ZN(n8984) );
  AND2_X1 U11360 ( .A1(n11834), .A2(n8984), .ZN(n8954) );
  NAND2_X1 U11361 ( .A1(n14400), .A2(n8961), .ZN(n10236) );
  INV_X1 U11362 ( .A(n6661), .ZN(n10715) );
  NAND2_X1 U11363 ( .A1(n10478), .A2(n10715), .ZN(n14265) );
  NAND2_X1 U11364 ( .A1(n10478), .A2(n6661), .ZN(n14220) );
  INV_X1 U11365 ( .A(P1_B_REG_SCAN_IN), .ZN(n8955) );
  NOR2_X1 U11366 ( .A1(n15026), .A2(n8955), .ZN(n8956) );
  NOR2_X1 U11367 ( .A1(n14220), .A2(n8956), .ZN(n14057) );
  INV_X1 U11368 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U11369 ( .A1(n6678), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U11370 ( .A1(n8894), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8957) );
  OAI211_X1 U11371 ( .C1(n9152), .C2(n8959), .A(n8958), .B(n8957), .ZN(n13954)
         );
  NAND2_X1 U11372 ( .A1(n14057), .A2(n13954), .ZN(n12254) );
  OAI21_X1 U11373 ( .B1(n8960), .B2(n14265), .A(n12254), .ZN(n8962) );
  INV_X1 U11374 ( .A(n14131), .ZN(n14301) );
  INV_X1 U11375 ( .A(n11773), .ZN(n15171) );
  OR2_X1 U11376 ( .A1(n14342), .A2(n14244), .ZN(n14242) );
  NAND2_X1 U11377 ( .A1(n8976), .A2(P1_B_REG_SCAN_IN), .ZN(n8967) );
  MUX2_X1 U11378 ( .A(n8967), .B(P1_B_REG_SCAN_IN), .S(n8978), .Z(n8972) );
  INV_X1 U11379 ( .A(n8968), .ZN(n8969) );
  OAI21_X1 U11380 ( .B1(n6941), .B2(n8969), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8970) );
  MUX2_X1 U11381 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8970), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8971) );
  INV_X1 U11382 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10404) );
  INV_X1 U11383 ( .A(n8977), .ZN(n14394) );
  NAND2_X1 U11384 ( .A1(n15111), .A2(n11942), .ZN(n10239) );
  INV_X1 U11385 ( .A(n10239), .ZN(n11066) );
  NOR2_X1 U11386 ( .A1(n11064), .A2(n11066), .ZN(n8999) );
  INV_X1 U11387 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10401) );
  NAND2_X1 U11388 ( .A1(n10398), .A2(n10401), .ZN(n8975) );
  NOR2_X1 U11389 ( .A1(n8978), .A2(n8977), .ZN(n10400) );
  INV_X1 U11390 ( .A(n10400), .ZN(n8974) );
  NAND2_X1 U11391 ( .A1(n8975), .A2(n8974), .ZN(n8998) );
  NAND2_X1 U11392 ( .A1(n8963), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8981) );
  MUX2_X1 U11393 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8981), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8983) );
  NAND2_X1 U11394 ( .A1(n10478), .A2(n8984), .ZN(n10240) );
  NAND2_X1 U11395 ( .A1(n11067), .A2(n10240), .ZN(n10610) );
  INV_X1 U11396 ( .A(n10610), .ZN(n8997) );
  NOR4_X1 U11397 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8988) );
  NOR4_X1 U11398 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n8987) );
  NOR4_X1 U11399 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n8986) );
  NOR4_X1 U11400 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n8985) );
  NAND4_X1 U11401 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n8994)
         );
  NOR2_X1 U11402 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .ZN(
        n8992) );
  NOR4_X1 U11403 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n8991) );
  NOR4_X1 U11404 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n8990) );
  NOR4_X1 U11405 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n8989) );
  NAND4_X1 U11406 ( .A1(n8992), .A2(n8991), .A3(n8990), .A4(n8989), .ZN(n8993)
         );
  NOR2_X1 U11407 ( .A1(n8994), .A2(n8993), .ZN(n9202) );
  INV_X1 U11408 ( .A(n9202), .ZN(n8995) );
  NAND2_X1 U11409 ( .A1(n10398), .A2(n8995), .ZN(n8996) );
  NAND2_X1 U11410 ( .A1(n11079), .A2(n11942), .ZN(n9000) );
  NAND2_X1 U11411 ( .A1(n9001), .A2(n9000), .ZN(n9156) );
  MUX2_X1 U11412 ( .A(n14757), .B(n11834), .S(n9156), .Z(n9002) );
  INV_X1 U11413 ( .A(n9002), .ZN(n9070) );
  MUX2_X1 U11414 ( .A(n9003), .B(n12259), .S(n9142), .Z(n9145) );
  INV_X1 U11415 ( .A(n9145), .ZN(n9149) );
  NAND2_X1 U11416 ( .A1(n9175), .A2(n10206), .ZN(n9004) );
  NAND2_X1 U11417 ( .A1(n14262), .A2(n14256), .ZN(n9174) );
  NAND2_X1 U11418 ( .A1(n9004), .A2(n9174), .ZN(n9006) );
  INV_X1 U11419 ( .A(n9175), .ZN(n9005) );
  INV_X1 U11420 ( .A(n9070), .ZN(n9076) );
  MUX2_X1 U11421 ( .A(n9006), .B(n9005), .S(n9076), .Z(n9013) );
  INV_X1 U11422 ( .A(n9010), .ZN(n9007) );
  MUX2_X1 U11423 ( .A(n9008), .B(n9007), .S(n9076), .Z(n9012) );
  MUX2_X1 U11424 ( .A(n9010), .B(n9009), .S(n9076), .Z(n9011) );
  MUX2_X1 U11425 ( .A(n9015), .B(n9014), .S(n9076), .Z(n9016) );
  NAND2_X1 U11426 ( .A1(n9076), .A2(n13965), .ZN(n9019) );
  NAND2_X1 U11427 ( .A1(n9167), .A2(n11193), .ZN(n9018) );
  MUX2_X1 U11428 ( .A(n9019), .B(n9018), .S(n11150), .Z(n9020) );
  NAND2_X1 U11429 ( .A1(n9021), .A2(n9020), .ZN(n9024) );
  MUX2_X1 U11430 ( .A(n11145), .B(n15149), .S(n9076), .Z(n9023) );
  INV_X1 U11431 ( .A(n15149), .ZN(n11174) );
  MUX2_X1 U11432 ( .A(n11174), .B(n13964), .S(n9076), .Z(n9022) );
  OAI21_X1 U11433 ( .B1(n9024), .B2(n9023), .A(n9022), .ZN(n9026) );
  NAND2_X1 U11434 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  MUX2_X1 U11435 ( .A(n11519), .B(n13963), .S(n9076), .Z(n9028) );
  MUX2_X1 U11436 ( .A(n13963), .B(n11519), .S(n9076), .Z(n9027) );
  MUX2_X1 U11437 ( .A(n13962), .B(n11594), .S(n9142), .Z(n9032) );
  NAND2_X1 U11438 ( .A1(n9031), .A2(n9032), .ZN(n9030) );
  MUX2_X1 U11439 ( .A(n13962), .B(n11594), .S(n9167), .Z(n9029) );
  NAND2_X1 U11440 ( .A1(n9030), .A2(n9029), .ZN(n9036) );
  INV_X1 U11441 ( .A(n9031), .ZN(n9034) );
  INV_X1 U11442 ( .A(n9032), .ZN(n9033) );
  NAND2_X1 U11443 ( .A1(n9034), .A2(n9033), .ZN(n9035) );
  MUX2_X1 U11444 ( .A(n13961), .B(n11773), .S(n9167), .Z(n9038) );
  MUX2_X1 U11445 ( .A(n13961), .B(n11773), .S(n9142), .Z(n9037) );
  INV_X1 U11446 ( .A(n9038), .ZN(n9039) );
  MUX2_X1 U11447 ( .A(n13960), .B(n15177), .S(n9142), .Z(n9042) );
  NAND2_X1 U11448 ( .A1(n9043), .A2(n9042), .ZN(n9041) );
  MUX2_X1 U11449 ( .A(n13960), .B(n15177), .S(n9167), .Z(n9040) );
  NAND2_X1 U11450 ( .A1(n9041), .A2(n9040), .ZN(n9045) );
  OR2_X1 U11451 ( .A1(n9043), .A2(n9042), .ZN(n9044) );
  MUX2_X1 U11452 ( .A(n14927), .B(n12029), .S(n9167), .Z(n9047) );
  MUX2_X1 U11453 ( .A(n14927), .B(n12029), .S(n9142), .Z(n9046) );
  MUX2_X1 U11454 ( .A(n14943), .B(n14925), .S(n9142), .Z(n9051) );
  NAND2_X1 U11455 ( .A1(n9050), .A2(n9051), .ZN(n9049) );
  MUX2_X1 U11456 ( .A(n14943), .B(n14925), .S(n9167), .Z(n9048) );
  NAND2_X1 U11457 ( .A1(n9049), .A2(n9048), .ZN(n9055) );
  INV_X1 U11458 ( .A(n9050), .ZN(n9053) );
  INV_X1 U11459 ( .A(n9051), .ZN(n9052) );
  NAND2_X1 U11460 ( .A1(n9053), .A2(n9052), .ZN(n9054) );
  MUX2_X1 U11461 ( .A(n13959), .B(n12216), .S(n9167), .Z(n9057) );
  MUX2_X1 U11462 ( .A(n13959), .B(n12216), .S(n9142), .Z(n9056) );
  INV_X1 U11463 ( .A(n9057), .ZN(n9058) );
  MUX2_X1 U11464 ( .A(n14978), .B(n12227), .S(n9142), .Z(n9062) );
  MUX2_X1 U11465 ( .A(n13958), .B(n14981), .S(n9167), .Z(n9066) );
  NOR2_X1 U11466 ( .A1(n9142), .A2(n14911), .ZN(n9059) );
  AOI21_X1 U11467 ( .B1(n14981), .B2(n9142), .A(n9059), .ZN(n9065) );
  NAND2_X1 U11468 ( .A1(n9066), .A2(n9065), .ZN(n9060) );
  OAI211_X1 U11469 ( .C1(n9063), .C2(n9062), .A(n11944), .B(n9060), .ZN(n9075)
         );
  INV_X1 U11470 ( .A(n12227), .ZN(n14794) );
  MUX2_X1 U11471 ( .A(n12246), .B(n14794), .S(n9167), .Z(n9061) );
  AOI21_X1 U11472 ( .B1(n9063), .B2(n9062), .A(n9061), .ZN(n9074) );
  NAND2_X1 U11473 ( .A1(n9078), .A2(n9064), .ZN(n9068) );
  NOR2_X1 U11474 ( .A1(n9066), .A2(n9065), .ZN(n9067) );
  AOI22_X1 U11475 ( .A1(n9068), .A2(n9142), .B1(n11944), .B2(n9067), .ZN(n9073) );
  NAND2_X1 U11476 ( .A1(n9077), .A2(n9069), .ZN(n9071) );
  NAND2_X1 U11477 ( .A1(n9071), .A2(n9167), .ZN(n9072) );
  OAI211_X1 U11478 ( .C1(n9075), .C2(n9074), .A(n9073), .B(n9072), .ZN(n9082)
         );
  MUX2_X1 U11479 ( .A(n14237), .B(n13912), .S(n9076), .Z(n9092) );
  OR2_X1 U11480 ( .A1(n9092), .A2(n9089), .ZN(n9081) );
  MUX2_X1 U11481 ( .A(n12328), .B(n14967), .S(n9076), .Z(n9084) );
  MUX2_X1 U11482 ( .A(n14953), .B(n12106), .S(n9167), .Z(n9083) );
  NAND2_X1 U11483 ( .A1(n9084), .A2(n9083), .ZN(n9080) );
  MUX2_X1 U11484 ( .A(n9078), .B(n9077), .S(n9142), .Z(n9079) );
  NAND4_X1 U11485 ( .A1(n9082), .A2(n9081), .A3(n9080), .A4(n9079), .ZN(n9094)
         );
  INV_X1 U11486 ( .A(n9083), .ZN(n9086) );
  INV_X1 U11487 ( .A(n9084), .ZN(n9085) );
  NAND2_X1 U11488 ( .A1(n9086), .A2(n9085), .ZN(n9088) );
  NAND2_X1 U11489 ( .A1(n9088), .A2(n9087), .ZN(n9091) );
  INV_X1 U11490 ( .A(n9088), .ZN(n9090) );
  AOI22_X1 U11491 ( .A1(n9092), .A2(n9091), .B1(n9090), .B2(n9089), .ZN(n9093)
         );
  AND2_X1 U11492 ( .A1(n14342), .A2(n9167), .ZN(n9096) );
  NOR2_X1 U11493 ( .A1(n14342), .A2(n9167), .ZN(n9095) );
  MUX2_X1 U11494 ( .A(n9096), .B(n9095), .S(n14222), .Z(n9097) );
  INV_X1 U11495 ( .A(n9097), .ZN(n9099) );
  INV_X1 U11496 ( .A(n14217), .ZN(n9098) );
  NAND3_X1 U11497 ( .A1(n7656), .A2(n9099), .A3(n9098), .ZN(n9103) );
  MUX2_X1 U11498 ( .A(n9101), .B(n9100), .S(n9167), .Z(n9102) );
  MUX2_X1 U11499 ( .A(n14221), .B(n14212), .S(n9167), .Z(n9105) );
  MUX2_X1 U11500 ( .A(n13956), .B(n14329), .S(n9142), .Z(n9104) );
  MUX2_X1 U11501 ( .A(n14175), .B(n14324), .S(n9142), .Z(n9109) );
  MUX2_X1 U11502 ( .A(n14175), .B(n14324), .S(n9167), .Z(n9106) );
  NAND2_X1 U11503 ( .A1(n9107), .A2(n9106), .ZN(n9110) );
  MUX2_X1 U11504 ( .A(n14156), .B(n12364), .S(n9167), .Z(n9112) );
  MUX2_X1 U11505 ( .A(n14156), .B(n12364), .S(n9142), .Z(n9111) );
  INV_X1 U11506 ( .A(n9112), .ZN(n9113) );
  MUX2_X1 U11507 ( .A(n14174), .B(n14313), .S(n9142), .Z(n9117) );
  NAND2_X1 U11508 ( .A1(n9116), .A2(n9117), .ZN(n9115) );
  MUX2_X1 U11509 ( .A(n14174), .B(n14313), .S(n9167), .Z(n9114) );
  NAND2_X1 U11510 ( .A1(n9115), .A2(n9114), .ZN(n9121) );
  INV_X1 U11511 ( .A(n9116), .ZN(n9119) );
  INV_X1 U11512 ( .A(n9117), .ZN(n9118) );
  NAND2_X1 U11513 ( .A1(n9119), .A2(n9118), .ZN(n9120) );
  NAND2_X1 U11514 ( .A1(n9121), .A2(n9120), .ZN(n9124) );
  MUX2_X1 U11515 ( .A(n14157), .B(n14308), .S(n9167), .Z(n9125) );
  NAND2_X1 U11516 ( .A1(n9124), .A2(n9125), .ZN(n9123) );
  MUX2_X1 U11517 ( .A(n14157), .B(n14308), .S(n9142), .Z(n9122) );
  INV_X1 U11518 ( .A(n9124), .ZN(n9127) );
  INV_X1 U11519 ( .A(n9125), .ZN(n9126) );
  NAND2_X1 U11520 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  MUX2_X1 U11521 ( .A(n13955), .B(n14131), .S(n9142), .Z(n9130) );
  MUX2_X1 U11522 ( .A(n13955), .B(n14131), .S(n9167), .Z(n9129) );
  MUX2_X1 U11523 ( .A(n14094), .B(n14112), .S(n9167), .Z(n9134) );
  NAND2_X1 U11524 ( .A1(n9133), .A2(n9134), .ZN(n9132) );
  MUX2_X1 U11525 ( .A(n14094), .B(n14112), .S(n9142), .Z(n9131) );
  MUX2_X1 U11526 ( .A(n14069), .B(n14285), .S(n9142), .Z(n9137) );
  MUX2_X1 U11527 ( .A(n14069), .B(n14285), .S(n9167), .Z(n9136) );
  MUX2_X1 U11528 ( .A(n14095), .B(n14279), .S(n9167), .Z(n9140) );
  MUX2_X1 U11529 ( .A(n14095), .B(n14279), .S(n9142), .Z(n9138) );
  INV_X1 U11530 ( .A(n9140), .ZN(n9141) );
  MUX2_X1 U11531 ( .A(n9143), .B(n14070), .S(n9142), .Z(n9144) );
  OAI21_X1 U11532 ( .B1(n9149), .B2(n9148), .A(n9147), .ZN(n9161) );
  INV_X1 U11533 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14546) );
  NAND2_X1 U11534 ( .A1(n6678), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U11535 ( .A1(n8894), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9150) );
  OAI211_X1 U11536 ( .C1(n9152), .C2(n14546), .A(n9151), .B(n9150), .ZN(n14056) );
  OAI21_X1 U11537 ( .B1(n14056), .B2(n9153), .A(n13954), .ZN(n9155) );
  MUX2_X1 U11538 ( .A(n9155), .B(n14277), .S(n9142), .Z(n9160) );
  INV_X1 U11539 ( .A(n13954), .ZN(n9158) );
  AOI22_X1 U11540 ( .A1(n9142), .A2(n14056), .B1(n11834), .B2(n9156), .ZN(
        n9157) );
  OAI22_X1 U11541 ( .A1(n14277), .A2(n9142), .B1(n9158), .B2(n9157), .ZN(n9159) );
  NAND2_X1 U11542 ( .A1(n9161), .A2(n9160), .ZN(n9165) );
  XNOR2_X1 U11543 ( .A(n6685), .B(n14056), .ZN(n9193) );
  NOR3_X1 U11544 ( .A1(n6685), .A2(n14056), .A3(n9167), .ZN(n9169) );
  AND3_X1 U11545 ( .A1(n6685), .A2(n14056), .A3(n9167), .ZN(n9168) );
  NOR2_X1 U11546 ( .A1(n9169), .A2(n9168), .ZN(n9195) );
  INV_X1 U11547 ( .A(n10206), .ZN(n10205) );
  AND2_X1 U11548 ( .A1(n10205), .A2(n11942), .ZN(n11068) );
  AOI21_X1 U11549 ( .B1(n10236), .B2(n9170), .A(n11068), .ZN(n9171) );
  INV_X1 U11550 ( .A(n9171), .ZN(n9172) );
  NAND2_X1 U11551 ( .A1(n11834), .A2(n14757), .ZN(n11078) );
  INV_X1 U11552 ( .A(n14277), .ZN(n14054) );
  XNOR2_X1 U11553 ( .A(n14054), .B(n13954), .ZN(n9191) );
  INV_X1 U11554 ( .A(n11944), .ZN(n9181) );
  NAND2_X1 U11555 ( .A1(n9175), .A2(n9174), .ZN(n11121) );
  NOR4_X1 U11556 ( .A1(n11137), .A2(n11183), .A3(n14264), .A4(n11121), .ZN(
        n9176) );
  XNOR2_X1 U11557 ( .A(n11174), .B(n13964), .ZN(n11176) );
  NAND4_X1 U11558 ( .A1(n11071), .A2(n9176), .A3(n15097), .A4(n11176), .ZN(
        n9177) );
  NOR4_X1 U11559 ( .A1(n11496), .A2(n15081), .A3(n11371), .A4(n9177), .ZN(
        n9179) );
  NAND4_X1 U11560 ( .A1(n11751), .A2(n9179), .A3(n11536), .A4(n9178), .ZN(
        n9180) );
  NOR4_X1 U11561 ( .A1(n12092), .A2(n9181), .A3(n14811), .A4(n9180), .ZN(n9184) );
  NAND2_X1 U11562 ( .A1(n9183), .A2(n9182), .ZN(n12129) );
  NAND4_X1 U11563 ( .A1(n14235), .A2(n9185), .A3(n9184), .A4(n12129), .ZN(
        n9186) );
  NOR4_X1 U11564 ( .A1(n14184), .A2(n14209), .A3(n14217), .A4(n9186), .ZN(
        n9187) );
  NAND4_X1 U11565 ( .A1(n14123), .A2(n14170), .A3(n9187), .A4(n14154), .ZN(
        n9188) );
  NOR4_X1 U11566 ( .A1(n14090), .A2(n14142), .A3(n14107), .A4(n9188), .ZN(
        n9190) );
  NAND4_X1 U11567 ( .A1(n9191), .A2(n14077), .A3(n9190), .A4(n9189), .ZN(n9192) );
  NOR2_X1 U11568 ( .A1(n9193), .A2(n9192), .ZN(n9194) );
  INV_X1 U11569 ( .A(n9195), .ZN(n9197) );
  NAND2_X1 U11570 ( .A1(n9196), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12011) );
  AOI21_X1 U11571 ( .B1(n9197), .B2(n7642), .A(n12011), .ZN(n9198) );
  NOR3_X1 U11572 ( .A1(n10610), .A2(n14265), .A3(n15026), .ZN(n9200) );
  OAI21_X1 U11573 ( .B1(n12011), .B2(n14400), .A(P1_B_REG_SCAN_IN), .ZN(n9199)
         );
  OR2_X1 U11574 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  INV_X1 U11575 ( .A(n11064), .ZN(n9206) );
  NAND2_X1 U11576 ( .A1(n9202), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9203) );
  AOI21_X1 U11577 ( .B1(n10398), .B2(n9203), .A(n10400), .ZN(n10235) );
  NOR2_X1 U11578 ( .A1(n10610), .A2(n11066), .ZN(n9204) );
  AND2_X1 U11579 ( .A1(n10235), .A2(n9204), .ZN(n9205) );
  INV_X1 U11580 ( .A(n13551), .ZN(n9244) );
  INV_X1 U11581 ( .A(n13575), .ZN(n9239) );
  INV_X1 U11582 ( .A(n13606), .ZN(n13640) );
  INV_X1 U11583 ( .A(n13432), .ZN(n13662) );
  INV_X1 U11584 ( .A(n13782), .ZN(n13700) );
  NAND2_X1 U11585 ( .A1(n10270), .A2(n9208), .ZN(n10250) );
  NAND2_X1 U11586 ( .A1(n10249), .A2(n9209), .ZN(n10761) );
  NAND2_X1 U11587 ( .A1(n10780), .A2(n10838), .ZN(n9211) );
  INV_X1 U11588 ( .A(n13449), .ZN(n10885) );
  AND2_X1 U11589 ( .A1(n10848), .A2(n10885), .ZN(n9212) );
  OR2_X1 U11590 ( .A1(n10836), .A2(n10885), .ZN(n9213) );
  INV_X1 U11591 ( .A(n11436), .ZN(n11445) );
  AND2_X1 U11592 ( .A1(n11442), .A2(n11130), .ZN(n11353) );
  NOR2_X1 U11593 ( .A1(n11355), .A2(n11353), .ZN(n9214) );
  INV_X1 U11594 ( .A(n13446), .ZN(n11248) );
  NAND2_X1 U11595 ( .A1(n11639), .A2(n9216), .ZN(n11565) );
  INV_X1 U11596 ( .A(n13444), .ZN(n11785) );
  OR2_X1 U11597 ( .A1(n11803), .A2(n11785), .ZN(n9217) );
  NAND2_X1 U11598 ( .A1(n11565), .A2(n9217), .ZN(n9219) );
  NAND2_X1 U11599 ( .A1(n11803), .A2(n11785), .ZN(n9218) );
  NAND2_X1 U11600 ( .A1(n9219), .A2(n9218), .ZN(n11806) );
  NAND2_X1 U11601 ( .A1(n15286), .A2(n11907), .ZN(n9220) );
  OR2_X1 U11602 ( .A1(n11917), .A2(n11781), .ZN(n9221) );
  NAND2_X1 U11603 ( .A1(n11917), .A2(n11781), .ZN(n9222) );
  AND2_X1 U11604 ( .A1(n12039), .A2(n12119), .ZN(n9223) );
  INV_X1 U11605 ( .A(n12117), .ZN(n9224) );
  NAND2_X1 U11606 ( .A1(n12114), .A2(n9226), .ZN(n12168) );
  INV_X1 U11607 ( .A(n13439), .ZN(n13348) );
  NAND2_X1 U11608 ( .A1(n13805), .A2(n13348), .ZN(n9227) );
  OR2_X1 U11609 ( .A1(n13798), .A2(n9228), .ZN(n9229) );
  INV_X1 U11610 ( .A(n12196), .ZN(n12191) );
  INV_X1 U11611 ( .A(n12201), .ZN(n13792) );
  INV_X1 U11612 ( .A(n13787), .ZN(n13715) );
  NOR2_X1 U11613 ( .A1(n13715), .A2(n13436), .ZN(n9231) );
  OAI22_X1 U11614 ( .A1(n13704), .A2(n9231), .B1(n9230), .B2(n13787), .ZN(
        n13693) );
  AOI21_X1 U11615 ( .B1(n13700), .B2(n13435), .A(n13693), .ZN(n9232) );
  INV_X1 U11616 ( .A(n13777), .ZN(n9233) );
  INV_X1 U11617 ( .A(n13772), .ZN(n13669) );
  NOR2_X1 U11618 ( .A1(n13669), .A2(n13433), .ZN(n9234) );
  INV_X1 U11619 ( .A(n13433), .ZN(n13641) );
  NOR2_X1 U11620 ( .A1(n13616), .A2(n13584), .ZN(n13580) );
  INV_X1 U11621 ( .A(n13560), .ZN(n13549) );
  OAI21_X1 U11622 ( .B1(n9244), .B2(n13729), .A(n13533), .ZN(n9241) );
  INV_X1 U11623 ( .A(P2_B_REG_SCAN_IN), .ZN(n9301) );
  OAI21_X1 U11624 ( .B1(n12270), .B2(n9301), .A(n13604), .ZN(n13508) );
  OAI22_X1 U11625 ( .A1(n9244), .A2(n13661), .B1(n9243), .B2(n13508), .ZN(
        n9245) );
  INV_X1 U11626 ( .A(n10275), .ZN(n9246) );
  NAND2_X1 U11627 ( .A1(n10276), .A2(n9246), .ZN(n9249) );
  NAND2_X1 U11628 ( .A1(n9247), .A2(n15316), .ZN(n9248) );
  INV_X1 U11629 ( .A(n8475), .ZN(n10625) );
  NAND2_X1 U11630 ( .A1(n10625), .A2(n8476), .ZN(n9250) );
  NAND2_X1 U11631 ( .A1(n9251), .A2(n9250), .ZN(n10759) );
  INV_X1 U11632 ( .A(n10762), .ZN(n9252) );
  NAND2_X1 U11633 ( .A1(n10759), .A2(n9252), .ZN(n9254) );
  NAND2_X1 U11634 ( .A1(n10778), .A2(n15328), .ZN(n9253) );
  INV_X1 U11635 ( .A(n10855), .ZN(n9255) );
  OR2_X1 U11636 ( .A1(n10780), .A2(n13450), .ZN(n9256) );
  INV_X1 U11637 ( .A(n10836), .ZN(n9257) );
  OR2_X1 U11638 ( .A1(n10848), .A2(n13449), .ZN(n9258) );
  NAND2_X1 U11639 ( .A1(n9259), .A2(n9258), .ZN(n11437) );
  NAND2_X1 U11640 ( .A1(n11437), .A2(n11436), .ZN(n9261) );
  OR2_X1 U11641 ( .A1(n11442), .A2(n13448), .ZN(n9260) );
  OR2_X1 U11642 ( .A1(n15348), .A2(n13447), .ZN(n9262) );
  NAND2_X1 U11643 ( .A1(n11484), .A2(n13446), .ZN(n9264) );
  NAND2_X1 U11644 ( .A1(n15355), .A2(n13445), .ZN(n9265) );
  INV_X1 U11645 ( .A(n11564), .ZN(n11566) );
  NAND2_X1 U11646 ( .A1(n11567), .A2(n11566), .ZN(n11569) );
  NAND2_X1 U11647 ( .A1(n11803), .A2(n13444), .ZN(n9266) );
  NAND2_X1 U11648 ( .A1(n11569), .A2(n9266), .ZN(n11805) );
  OAI21_X1 U11649 ( .B1(n11805), .B2(n11807), .A(n15286), .ZN(n9268) );
  NAND2_X1 U11650 ( .A1(n11805), .A2(n13443), .ZN(n9267) );
  NAND2_X1 U11651 ( .A1(n9268), .A2(n9267), .ZN(n11904) );
  AND2_X1 U11652 ( .A1(n11917), .A2(n13442), .ZN(n9269) );
  OAI22_X1 U11653 ( .A1(n11904), .A2(n9269), .B1(n11917), .B2(n13442), .ZN(
        n12036) );
  NOR2_X1 U11654 ( .A1(n12039), .A2(n13441), .ZN(n9270) );
  NAND2_X1 U11655 ( .A1(n12039), .A2(n13441), .ZN(n9271) );
  AND2_X1 U11656 ( .A1(n13811), .A2(n13440), .ZN(n9272) );
  OR2_X1 U11657 ( .A1(n13811), .A2(n13440), .ZN(n9273) );
  INV_X1 U11658 ( .A(n12167), .ZN(n9275) );
  NOR2_X1 U11659 ( .A1(n13805), .A2(n13439), .ZN(n9274) );
  AOI21_X1 U11660 ( .B1(n12165), .B2(n9275), .A(n9274), .ZN(n12162) );
  INV_X1 U11661 ( .A(n12154), .ZN(n12161) );
  NAND2_X1 U11662 ( .A1(n13798), .A2(n13438), .ZN(n9276) );
  OR2_X1 U11663 ( .A1(n12201), .A2(n13437), .ZN(n9277) );
  OR2_X1 U11664 ( .A1(n13787), .A2(n13436), .ZN(n9279) );
  NAND2_X1 U11665 ( .A1(n13716), .A2(n9279), .ZN(n13691) );
  NOR2_X1 U11666 ( .A1(n13782), .A2(n13435), .ZN(n9280) );
  NAND2_X1 U11667 ( .A1(n13782), .A2(n13435), .ZN(n9281) );
  AND2_X1 U11668 ( .A1(n13777), .A2(n13434), .ZN(n9282) );
  OR2_X1 U11669 ( .A1(n13777), .A2(n13434), .ZN(n9283) );
  INV_X1 U11670 ( .A(n13655), .ZN(n13657) );
  OR2_X1 U11671 ( .A1(n13772), .A2(n13433), .ZN(n9284) );
  NAND2_X1 U11672 ( .A1(n13765), .A2(n13432), .ZN(n9286) );
  NAND2_X1 U11673 ( .A1(n13759), .A2(n13606), .ZN(n9287) );
  NAND2_X1 U11674 ( .A1(n13624), .A2(n9287), .ZN(n13598) );
  NAND2_X1 U11675 ( .A1(n13598), .A2(n13602), .ZN(n13600) );
  NAND2_X1 U11676 ( .A1(n13752), .A2(n13584), .ZN(n9288) );
  NAND2_X1 U11677 ( .A1(n13600), .A2(n9288), .ZN(n13593) );
  OR2_X1 U11678 ( .A1(n13747), .A2(n13605), .ZN(n9289) );
  NAND2_X1 U11679 ( .A1(n13591), .A2(n9289), .ZN(n13564) );
  NAND2_X1 U11680 ( .A1(n13564), .A2(n9290), .ZN(n9292) );
  OR2_X1 U11681 ( .A1(n13742), .A2(n13583), .ZN(n9291) );
  INV_X1 U11682 ( .A(n13534), .ZN(n13531) );
  NAND2_X1 U11683 ( .A1(n13532), .A2(n9293), .ZN(n9295) );
  XNOR2_X1 U11684 ( .A(n9296), .B(n9299), .ZN(n9297) );
  INV_X1 U11685 ( .A(n9298), .ZN(n13756) );
  INV_X1 U11686 ( .A(n13729), .ZN(n13545) );
  INV_X1 U11687 ( .A(n13742), .ZN(n13571) );
  INV_X1 U11688 ( .A(n12039), .ZN(n14896) );
  INV_X1 U11689 ( .A(n15355), .ZN(n11648) );
  NOR2_X1 U11690 ( .A1(n10489), .A2(n8474), .ZN(n10280) );
  NAND2_X1 U11691 ( .A1(n10280), .A2(n8476), .ZN(n10767) );
  OR2_X1 U11692 ( .A1(n10767), .A2(n8480), .ZN(n10860) );
  INV_X1 U11693 ( .A(n10848), .ZN(n11100) );
  INV_X1 U11694 ( .A(n11442), .ZN(n15343) );
  NAND2_X1 U11695 ( .A1(n14896), .A2(n12037), .ZN(n12120) );
  OR2_X1 U11696 ( .A1(n13787), .A2(n13707), .ZN(n13708) );
  OR2_X1 U11697 ( .A1(n13708), .A2(n13782), .ZN(n13696) );
  NAND2_X1 U11698 ( .A1(n13680), .A2(n13669), .ZN(n13665) );
  OR2_X2 U11699 ( .A1(n13665), .A2(n13765), .ZN(n13642) );
  NOR2_X1 U11700 ( .A1(n13734), .A2(n13565), .ZN(n13555) );
  NAND2_X1 U11701 ( .A1(n13545), .A2(n13555), .ZN(n13541) );
  AOI211_X1 U11702 ( .C1(n13521), .C2(n13541), .A(n10861), .B(n13515), .ZN(
        n13527) );
  XNOR2_X1 U11703 ( .A(n12187), .B(n9301), .ZN(n9302) );
  NAND2_X1 U11704 ( .A1(n9302), .A2(n13849), .ZN(n9303) );
  INV_X1 U11705 ( .A(n13846), .ZN(n9320) );
  NOR4_X1 U11706 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n9312) );
  INV_X1 U11707 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15304) );
  INV_X1 U11708 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15305) );
  INV_X1 U11709 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15303) );
  INV_X1 U11710 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15306) );
  NAND4_X1 U11711 ( .A1(n15304), .A2(n15305), .A3(n15303), .A4(n15306), .ZN(
        n9309) );
  NOR4_X1 U11712 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n9307) );
  NOR4_X1 U11713 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9306) );
  NOR4_X1 U11714 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9305) );
  NOR4_X1 U11715 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9304) );
  NAND4_X1 U11716 ( .A1(n9307), .A2(n9306), .A3(n9305), .A4(n9304), .ZN(n9308)
         );
  NOR4_X1 U11717 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        n9309), .A4(n9308), .ZN(n9311) );
  NOR4_X1 U11718 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9310) );
  NAND3_X1 U11719 ( .A1(n9312), .A2(n9311), .A3(n9310), .ZN(n9313) );
  AND2_X1 U11720 ( .A1(n15302), .A2(n9313), .ZN(n10195) );
  AND2_X1 U11721 ( .A1(n10360), .A2(n10191), .ZN(n9314) );
  NOR2_X1 U11722 ( .A1(n9315), .A2(n9314), .ZN(n10197) );
  INV_X1 U11723 ( .A(n10197), .ZN(n9316) );
  INV_X1 U11724 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U11725 ( .A1(n15302), .A2(n15312), .ZN(n9318) );
  NAND2_X1 U11726 ( .A1(n13846), .A2(n13849), .ZN(n9317) );
  NAND2_X1 U11727 ( .A1(n9318), .A2(n9317), .ZN(n15313) );
  NAND2_X1 U11728 ( .A1(n9298), .A2(n11835), .ZN(n10194) );
  NAND2_X1 U11729 ( .A1(n15313), .A2(n10194), .ZN(n9319) );
  INV_X1 U11730 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15309) );
  NAND2_X1 U11731 ( .A1(n15302), .A2(n15309), .ZN(n9322) );
  OR2_X1 U11732 ( .A1(n12187), .A2(n9320), .ZN(n9321) );
  INV_X1 U11733 ( .A(n15310), .ZN(n9323) );
  NAND2_X1 U11734 ( .A1(n13727), .A2(n15364), .ZN(n9326) );
  INV_X1 U11735 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9324) );
  XNOR2_X1 U11736 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n9424) );
  INV_X1 U11737 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n9362) );
  NOR2_X1 U11738 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9362), .ZN(n9361) );
  INV_X1 U11739 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9354) );
  INV_X1 U11740 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15048) );
  INV_X1 U11741 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U11742 ( .A1(n9327), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n9352) );
  INV_X1 U11743 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n9351) );
  INV_X1 U11744 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14572) );
  INV_X1 U11745 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14696) );
  XNOR2_X1 U11746 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), 
        .ZN(n9373) );
  INV_X1 U11747 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n9346) );
  XNOR2_X1 U11748 ( .A(n9330), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n9376) );
  NOR2_X1 U11749 ( .A1(n9377), .A2(n9376), .ZN(n9329) );
  NOR2_X1 U11750 ( .A1(n9331), .A2(n6862), .ZN(n9333) );
  NOR2_X1 U11751 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n9375), .ZN(n9332) );
  NOR2_X1 U11752 ( .A1(n9336), .A2(n9337), .ZN(n9339) );
  NOR2_X1 U11753 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9342), .ZN(n9344) );
  XOR2_X1 U11754 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n9342), .Z(n9397) );
  XNOR2_X1 U11755 ( .A(n9346), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n9402) );
  INV_X1 U11756 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n9348) );
  OAI22_X1 U11757 ( .A1(n9348), .A2(n14572), .B1(P1_ADDR_REG_10__SCAN_IN), 
        .B2(P3_ADDR_REG_10__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U11758 ( .A1(n9409), .A2(n9408), .ZN(n9349) );
  AND2_X1 U11759 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n9351), .ZN(n9350) );
  AND2_X1 U11760 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n9354), .ZN(n9353) );
  INV_X1 U11761 ( .A(n9419), .ZN(n9357) );
  INV_X1 U11762 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9355) );
  OR2_X1 U11763 ( .A1(n9355), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n9356) );
  INV_X1 U11764 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11765 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n9358), .ZN(n9359) );
  INV_X1 U11766 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15064) );
  AOI22_X1 U11767 ( .A1(n9368), .A2(n9359), .B1(P3_ADDR_REG_15__SCAN_IN), .B2(
        n15064), .ZN(n9366) );
  INV_X1 U11768 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n12891) );
  OR2_X1 U11769 ( .A1(n12891), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9360) );
  AOI22_X1 U11770 ( .A1(n9366), .A2(n9360), .B1(P1_ADDR_REG_16__SCAN_IN), .B2(
        n12891), .ZN(n9364) );
  INV_X1 U11771 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14566) );
  OAI22_X1 U11772 ( .A1(n9361), .A2(n9364), .B1(P3_ADDR_REG_17__SCAN_IN), .B2(
        n14566), .ZN(n9425) );
  XNOR2_X1 U11773 ( .A(n9424), .B(n9425), .ZN(n14766) );
  AOI22_X1 U11774 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n14566), .B2(n9362), .ZN(n9363) );
  XNOR2_X1 U11775 ( .A(n9364), .B(n9363), .ZN(n14821) );
  NAND2_X1 U11776 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n12891), .ZN(n9365) );
  OAI21_X1 U11777 ( .B1(n12891), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9365), .ZN(
        n9367) );
  XOR2_X1 U11778 ( .A(n9367), .B(n9366), .Z(n15022) );
  XNOR2_X1 U11779 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n9369) );
  XNOR2_X1 U11780 ( .A(n9369), .B(n9368), .ZN(n9420) );
  XNOR2_X1 U11781 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9371) );
  XNOR2_X1 U11782 ( .A(n9371), .B(n9370), .ZN(n15010) );
  XOR2_X1 U11783 ( .A(n9373), .B(n9372), .Z(n9406) );
  AND2_X1 U11784 ( .A1(n9386), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n9387) );
  XOR2_X1 U11785 ( .A(n9375), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15598) );
  XOR2_X1 U11786 ( .A(n9377), .B(n9376), .Z(n14772) );
  INV_X1 U11787 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9382) );
  NOR2_X1 U11788 ( .A1(n9381), .A2(n9382), .ZN(n9383) );
  OAI21_X1 U11789 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9380), .A(n9379), .ZN(
        n15592) );
  NAND2_X1 U11790 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15592), .ZN(n15603) );
  XNOR2_X1 U11791 ( .A(n9382), .B(n9381), .ZN(n15602) );
  NOR2_X1 U11792 ( .A1(n15603), .A2(n15602), .ZN(n15601) );
  NOR2_X1 U11793 ( .A1(n14772), .A2(n14771), .ZN(n9384) );
  NAND2_X1 U11794 ( .A1(n14772), .A2(n14771), .ZN(n14770) );
  NAND2_X1 U11795 ( .A1(n15598), .A2(n15597), .ZN(n9385) );
  NOR2_X1 U11796 ( .A1(n15598), .A2(n15597), .ZN(n15596) );
  XNOR2_X1 U11797 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n9386), .ZN(n15587) );
  NOR2_X1 U11798 ( .A1(n15588), .A2(n15587), .ZN(n15586) );
  NAND2_X1 U11799 ( .A1(n9389), .A2(n9390), .ZN(n9391) );
  INV_X1 U11800 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15590) );
  INV_X1 U11801 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9392) );
  NOR2_X1 U11802 ( .A1(n9393), .A2(n9392), .ZN(n9396) );
  XNOR2_X1 U11803 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n9395) );
  XNOR2_X1 U11804 ( .A(n9395), .B(n9394), .ZN(n14775) );
  INV_X1 U11805 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9399) );
  NOR2_X1 U11806 ( .A1(n9398), .A2(n9399), .ZN(n9400) );
  XNOR2_X1 U11807 ( .A(n9397), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15595) );
  NOR2_X1 U11808 ( .A1(n15595), .A2(n15594), .ZN(n15593) );
  XNOR2_X1 U11809 ( .A(n9402), .B(n9401), .ZN(n9404) );
  NAND2_X1 U11810 ( .A1(n9403), .A2(n9404), .ZN(n9405) );
  INV_X1 U11811 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14783) );
  INV_X1 U11812 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14787) );
  XNOR2_X1 U11813 ( .A(n9409), .B(n9408), .ZN(n14789) );
  XNOR2_X1 U11814 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9411) );
  XNOR2_X1 U11815 ( .A(n9411), .B(n9410), .ZN(n15001) );
  NAND2_X1 U11816 ( .A1(n15002), .A2(n15001), .ZN(n9412) );
  INV_X1 U11817 ( .A(n9413), .ZN(n9416) );
  XOR2_X1 U11818 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n9414) );
  XOR2_X1 U11819 ( .A(n9415), .B(n9414), .Z(n9417) );
  INV_X1 U11820 ( .A(n15005), .ZN(n15006) );
  INV_X1 U11821 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15008) );
  XOR2_X1 U11822 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n9418) );
  XNOR2_X1 U11823 ( .A(n9419), .B(n9418), .ZN(n15014) );
  INV_X1 U11824 ( .A(n15017), .ZN(n15018) );
  INV_X1 U11825 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15268) );
  NAND2_X1 U11826 ( .A1(n9421), .A2(n9420), .ZN(n15019) );
  NAND2_X1 U11827 ( .A1(n15268), .A2(n15019), .ZN(n15016) );
  NAND2_X1 U11828 ( .A1(n14821), .A2(n14822), .ZN(n14820) );
  INV_X1 U11829 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n9423) );
  INV_X1 U11830 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14627) );
  AND2_X1 U11831 ( .A1(n9425), .A2(n9424), .ZN(n9426) );
  AOI21_X1 U11832 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14627), .A(n9426), .ZN(
        n9428) );
  XNOR2_X1 U11833 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9427) );
  XNOR2_X1 U11834 ( .A(n9428), .B(n9427), .ZN(n9429) );
  NOR2_X1 U11835 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9616) );
  NAND2_X1 U11836 ( .A1(n9616), .A2(n14661), .ZN(n9629) );
  NAND2_X1 U11837 ( .A1(n9756), .A2(n11966), .ZN(n9769) );
  INV_X1 U11838 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n9430) );
  INV_X1 U11839 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n9434) );
  INV_X1 U11840 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12501) );
  INV_X1 U11841 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n9436) );
  INV_X1 U11842 ( .A(n9905), .ZN(n9439) );
  INV_X1 U11843 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9438) );
  INV_X1 U11844 ( .A(n9937), .ZN(n9441) );
  INV_X1 U11845 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U11846 ( .A1(n9441), .A2(n9440), .ZN(n9939) );
  NAND2_X1 U11847 ( .A1(n9939), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U11848 ( .A1(n9953), .A2(n9442), .ZN(n12979) );
  NOR2_X2 U11849 ( .A1(n9606), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9637) );
  NOR2_X1 U11850 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n9447) );
  NAND4_X1 U11851 ( .A1(n9447), .A2(n10002), .A3(n9446), .A4(n10003), .ZN(
        n9448) );
  NOR2_X1 U11852 ( .A1(n9448), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n9449) );
  AND2_X1 U11853 ( .A1(n9449), .A2(n9846), .ZN(n9452) );
  INV_X1 U11854 ( .A(n10009), .ZN(n9455) );
  INV_X1 U11855 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13234) );
  NAND2_X1 U11856 ( .A1(n9570), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U11857 ( .A1(n9692), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9462) );
  OAI211_X1 U11858 ( .C1(n13234), .C2(n9908), .A(n9463), .B(n9462), .ZN(n9464)
         );
  AOI21_X2 U11859 ( .B1(n12979), .B2(n9954), .A(n9464), .ZN(n12473) );
  AOI22_X1 U11860 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13851), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n14396), .ZN(n9531) );
  INV_X1 U11861 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10316) );
  INV_X1 U11862 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U11863 ( .A1(n9470), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U11864 ( .A1(n9611), .A2(n9610), .ZN(n9473) );
  NAND2_X1 U11865 ( .A1(n10318), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U11866 ( .A1(n9624), .A2(n9623), .ZN(n9476) );
  INV_X1 U11867 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U11868 ( .A1(n9474), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U11869 ( .A1(n10343), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9478) );
  NAND2_X1 U11870 ( .A1(n10348), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U11871 ( .A1(n9480), .A2(n9479), .ZN(n9668) );
  NAND2_X1 U11872 ( .A1(n9668), .A2(n9667), .ZN(n9483) );
  NAND2_X1 U11873 ( .A1(n9481), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U11874 ( .A1(n9483), .A2(n9482), .ZN(n9682) );
  XNOR2_X1 U11875 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9680) );
  NAND2_X1 U11876 ( .A1(n10395), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9484) );
  XNOR2_X1 U11877 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9700) );
  NAND2_X1 U11878 ( .A1(n10438), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U11879 ( .A1(n10469), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U11880 ( .A1(n10560), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U11881 ( .A1(n10559), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U11882 ( .A1(n9491), .A2(n9490), .ZN(n9738) );
  NAND2_X1 U11883 ( .A1(n10755), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9495) );
  INV_X1 U11884 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10756) );
  NAND2_X1 U11885 ( .A1(n10756), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9494) );
  NAND2_X1 U11886 ( .A1(n9765), .A2(n9764), .ZN(n9496) );
  NAND2_X1 U11887 ( .A1(n9496), .A2(n9495), .ZN(n9778) );
  NAND2_X1 U11888 ( .A1(n10991), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U11889 ( .A1(n10993), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11890 ( .A1(n9778), .A2(n9776), .ZN(n9499) );
  NAND2_X1 U11891 ( .A1(n14636), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U11892 ( .A1(n14648), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U11893 ( .A1(n9801), .A2(n9799), .ZN(n9502) );
  NAND2_X1 U11894 ( .A1(n9502), .A2(n9501), .ZN(n9814) );
  NAND2_X1 U11895 ( .A1(n11227), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U11896 ( .A1(n14610), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9504) );
  INV_X1 U11897 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U11898 ( .A1(n11548), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9506) );
  XNOR2_X1 U11899 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n9840) );
  NAND2_X1 U11900 ( .A1(n9842), .A2(n9840), .ZN(n9508) );
  NAND2_X1 U11901 ( .A1(n14521), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U11902 ( .A1(n9861), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9511) );
  INV_X1 U11903 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11721) );
  NAND2_X1 U11904 ( .A1(n9509), .A2(n11721), .ZN(n9510) );
  XNOR2_X1 U11905 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .ZN(n9874) );
  INV_X1 U11906 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11837) );
  NAND2_X1 U11907 ( .A1(n11837), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9512) );
  XNOR2_X1 U11908 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .ZN(n9887) );
  INV_X1 U11909 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9513) );
  XNOR2_X1 U11910 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9545) );
  NAND2_X1 U11911 ( .A1(n9546), .A2(n9545), .ZN(n9516) );
  INV_X1 U11912 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U11913 ( .A1(n9514), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U11914 ( .A1(n9517), .A2(n12190), .ZN(n9518) );
  NAND2_X1 U11915 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n14392), .ZN(n9522) );
  NAND2_X1 U11916 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n12271), .ZN(n9523) );
  INV_X1 U11917 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14390) );
  AOI22_X1 U11918 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(
        P2_DATAO_REG_28__SCAN_IN), .B1(n7129), .B2(n14552), .ZN(n9524) );
  INV_X1 U11919 ( .A(n9524), .ZN(n9525) );
  XNOR2_X1 U11920 ( .A(n9948), .B(n9525), .ZN(n12110) );
  NAND2_X1 U11921 ( .A1(n12110), .A2(n12602), .ZN(n9530) );
  OR2_X1 U11922 ( .A1(n6687), .A2(n12111), .ZN(n9529) );
  XNOR2_X1 U11923 ( .A(n9532), .B(n9531), .ZN(n11881) );
  NAND2_X1 U11924 ( .A1(n11881), .A2(n12602), .ZN(n9534) );
  OR2_X1 U11925 ( .A1(n9591), .A2(n14664), .ZN(n9533) );
  NAND2_X1 U11926 ( .A1(n9905), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U11927 ( .A1(n9920), .A2(n9535), .ZN(n13003) );
  NAND2_X1 U11928 ( .A1(n13003), .A2(n9954), .ZN(n9540) );
  INV_X1 U11929 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13241) );
  NAND2_X1 U11930 ( .A1(n9570), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U11931 ( .A1(n9692), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9536) );
  OAI211_X1 U11932 ( .C1(n9908), .C2(n13241), .A(n9537), .B(n9536), .ZN(n9538)
         );
  INV_X1 U11933 ( .A(n9538), .ZN(n9539) );
  NAND2_X1 U11934 ( .A1(n9894), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U11935 ( .A1(n9903), .A2(n9541), .ZN(n13036) );
  NAND2_X1 U11936 ( .A1(n13036), .A2(n9954), .ZN(n9544) );
  AOI22_X1 U11937 ( .A1(n6688), .A2(P3_REG0_REG_23__SCAN_IN), .B1(n9570), .B2(
        P3_REG1_REG_23__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U11938 ( .A1(n9692), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9542) );
  XNOR2_X1 U11939 ( .A(n9546), .B(n9545), .ZN(n11413) );
  NAND2_X1 U11940 ( .A1(n11413), .A2(n12602), .ZN(n9548) );
  INV_X1 U11941 ( .A(SI_23_), .ZN(n11415) );
  OR2_X1 U11942 ( .A1(n6687), .A2(n11415), .ZN(n9547) );
  NAND2_X1 U11943 ( .A1(n6688), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9553) );
  INV_X1 U11944 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11043) );
  OR2_X1 U11945 ( .A1(n9600), .A2(n11043), .ZN(n9551) );
  INV_X1 U11946 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9549) );
  OR2_X1 U11947 ( .A1(n6684), .A2(n9549), .ZN(n9550) );
  OR2_X1 U11948 ( .A1(n6687), .A2(SI_2_), .ZN(n9557) );
  XNOR2_X1 U11949 ( .A(n9555), .B(n9554), .ZN(n10322) );
  OAI211_X1 U11950 ( .C1(n10945), .C2(n10807), .A(n9557), .B(n9556), .ZN(
        n15497) );
  OR2_X1 U11951 ( .A1(n12826), .A2(n15497), .ZN(n12659) );
  NAND2_X1 U11952 ( .A1(n12826), .A2(n15497), .ZN(n12664) );
  INV_X1 U11953 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10898) );
  OR2_X1 U11954 ( .A1(n12609), .A2(n10898), .ZN(n9561) );
  INV_X1 U11955 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10826) );
  OR2_X1 U11956 ( .A1(n9867), .A2(n10826), .ZN(n9560) );
  INV_X1 U11957 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11014) );
  OR2_X1 U11958 ( .A1(n9600), .A2(n11014), .ZN(n9559) );
  NAND2_X1 U11959 ( .A1(n9569), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9558) );
  INV_X1 U11960 ( .A(n9577), .ZN(n9563) );
  XNOR2_X1 U11961 ( .A(n6676), .B(n9563), .ZN(n10295) );
  OR2_X1 U11962 ( .A1(n9742), .A2(n10295), .ZN(n9582) );
  NAND2_X1 U11963 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9565) );
  MUX2_X1 U11964 ( .A(n9565), .B(P3_IR_REG_31__SCAN_IN), .S(n9564), .Z(n9567)
         );
  OR2_X1 U11965 ( .A1(n10807), .A2(n10828), .ZN(n9581) );
  NAND2_X2 U11966 ( .A1(n12663), .A2(n12657), .ZN(n11008) );
  NAND2_X1 U11967 ( .A1(n6689), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9574) );
  INV_X1 U11968 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10827) );
  INV_X1 U11969 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10941) );
  INV_X1 U11970 ( .A(n6667), .ZN(n9570) );
  AND2_X1 U11971 ( .A1(n9575), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9576) );
  NOR2_X1 U11972 ( .A1(n9577), .A2(n9576), .ZN(n10288) );
  OR2_X1 U11973 ( .A1(n6687), .A2(n10287), .ZN(n9578) );
  AND2_X1 U11974 ( .A1(n9578), .A2(n7651), .ZN(n9579) );
  NAND2_X1 U11975 ( .A1(n10994), .A2(n10802), .ZN(n15506) );
  OR2_X1 U11976 ( .A1(n10788), .A2(n15503), .ZN(n15489) );
  NAND2_X1 U11977 ( .A1(n15505), .A2(n15489), .ZN(n9584) );
  NAND2_X1 U11978 ( .A1(n6688), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9588) );
  OR2_X1 U11979 ( .A1(n6667), .A2(n15574), .ZN(n9587) );
  OR2_X1 U11980 ( .A1(n9600), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9586) );
  INV_X1 U11981 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11388) );
  OR2_X1 U11982 ( .A1(n6684), .A2(n11388), .ZN(n9585) );
  OR3_X1 U11983 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n9589) );
  NAND2_X1 U11984 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n9589), .ZN(n9590) );
  XNOR2_X1 U11985 ( .A(n9590), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10987) );
  XNOR2_X1 U11986 ( .A(n9593), .B(n9592), .ZN(n10328) );
  OR2_X1 U11987 ( .A1(n9742), .A2(n10328), .ZN(n9594) );
  OAI211_X1 U11988 ( .C1(n10987), .C2(n10807), .A(n9595), .B(n9594), .ZN(
        n11389) );
  NAND2_X1 U11989 ( .A1(n12825), .A2(n11389), .ZN(n12668) );
  INV_X1 U11990 ( .A(n15497), .ZN(n11040) );
  OR2_X1 U11991 ( .A1(n12826), .A2(n11040), .ZN(n11383) );
  NAND2_X1 U11992 ( .A1(n15492), .A2(n9596), .ZN(n11382) );
  INV_X1 U11993 ( .A(n11389), .ZN(n11055) );
  NAND2_X1 U11994 ( .A1(n12825), .A2(n11055), .ZN(n9597) );
  NAND2_X1 U11995 ( .A1(n6688), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9605) );
  INV_X1 U11996 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9598) );
  OR2_X1 U11997 ( .A1(n6668), .A2(n9598), .ZN(n9604) );
  AND2_X1 U11998 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9599) );
  NOR2_X1 U11999 ( .A1(n9616), .A2(n9599), .ZN(n11857) );
  OR2_X1 U12000 ( .A1(n9600), .A2(n11857), .ZN(n9603) );
  INV_X1 U12001 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9601) );
  OR2_X1 U12002 ( .A1(n6683), .A2(n9601), .ZN(n9602) );
  NAND4_X1 U12003 ( .A1(n9605), .A2(n9604), .A3(n9603), .A4(n9602), .ZN(n12824) );
  NAND2_X1 U12004 ( .A1(n9607), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9608) );
  MUX2_X1 U12005 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9608), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9609) );
  AND2_X1 U12006 ( .A1(n9606), .A2(n9609), .ZN(n11288) );
  XNOR2_X1 U12007 ( .A(n9611), .B(n9610), .ZN(n10331) );
  OR2_X1 U12008 ( .A1(n9742), .A2(n10331), .ZN(n9613) );
  OR2_X1 U12009 ( .A1(n9591), .A2(SI_4_), .ZN(n9612) );
  OAI211_X1 U12010 ( .C1(n11288), .C2(n10807), .A(n9613), .B(n9612), .ZN(
        n15534) );
  XNOR2_X1 U12011 ( .A(n12824), .B(n15534), .ZN(n12630) );
  INV_X1 U12012 ( .A(n15534), .ZN(n11242) );
  NAND2_X1 U12013 ( .A1(n12824), .A2(n11242), .ZN(n9614) );
  NAND2_X1 U12014 ( .A1(n6689), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9621) );
  INV_X1 U12015 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15577) );
  OR2_X1 U12016 ( .A1(n6667), .A2(n15577), .ZN(n9620) );
  OR2_X1 U12017 ( .A1(n14661), .A2(n9616), .ZN(n9617) );
  AND2_X1 U12018 ( .A1(n9629), .A2(n9617), .ZN(n11559) );
  OR2_X1 U12019 ( .A1(n9600), .A2(n11559), .ZN(n9619) );
  INV_X1 U12020 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15374) );
  OR2_X1 U12021 ( .A1(n6684), .A2(n15374), .ZN(n9618) );
  NAND4_X1 U12022 ( .A1(n9621), .A2(n9620), .A3(n9619), .A4(n9618), .ZN(n11859) );
  NAND2_X1 U12023 ( .A1(n9606), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9622) );
  XNOR2_X1 U12024 ( .A(n9622), .B(P3_IR_REG_5__SCAN_IN), .ZN(n11293) );
  OR2_X1 U12025 ( .A1(n9591), .A2(SI_5_), .ZN(n9626) );
  XNOR2_X1 U12026 ( .A(n9624), .B(n9623), .ZN(n10325) );
  OR2_X1 U12027 ( .A1(n9742), .A2(n10325), .ZN(n9625) );
  OAI211_X1 U12028 ( .C1(n11293), .C2(n10807), .A(n9626), .B(n9625), .ZN(
        n11558) );
  NAND2_X1 U12029 ( .A1(n11859), .A2(n11558), .ZN(n12682) );
  INV_X1 U12030 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9628) );
  OR2_X1 U12031 ( .A1(n9908), .A2(n9628), .ZN(n9634) );
  INV_X1 U12032 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11295) );
  OR2_X1 U12033 ( .A1(n6668), .A2(n11295), .ZN(n9633) );
  NAND2_X1 U12034 ( .A1(n9629), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9630) );
  AND2_X1 U12035 ( .A1(n9644), .A2(n9630), .ZN(n11587) );
  OR2_X1 U12036 ( .A1(n9600), .A2(n11587), .ZN(n9632) );
  INV_X1 U12037 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11296) );
  OR2_X1 U12038 ( .A1(n6683), .A2(n11296), .ZN(n9631) );
  NAND4_X1 U12039 ( .A1(n9634), .A2(n9633), .A3(n9632), .A4(n9631), .ZN(n12823) );
  INV_X1 U12040 ( .A(SI_6_), .ZN(n10334) );
  OR2_X1 U12041 ( .A1(n9591), .A2(n10334), .ZN(n9641) );
  XNOR2_X1 U12042 ( .A(n10342), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n9635) );
  XNOR2_X1 U12043 ( .A(n9636), .B(n9635), .ZN(n10335) );
  OR2_X1 U12044 ( .A1(n9742), .A2(n10335), .ZN(n9640) );
  OR2_X1 U12045 ( .A1(n9637), .A2(n9720), .ZN(n9638) );
  XNOR2_X1 U12046 ( .A(n9638), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11297) );
  OR2_X1 U12047 ( .A1(n10807), .A2(n15397), .ZN(n9639) );
  NAND2_X1 U12048 ( .A1(n12823), .A2(n15546), .ZN(n12684) );
  NAND2_X1 U12049 ( .A1(n12686), .A2(n12684), .ZN(n12625) );
  INV_X1 U12050 ( .A(n11558), .ZN(n11460) );
  OR2_X1 U12051 ( .A1(n11859), .A2(n11460), .ZN(n11528) );
  AND2_X1 U12052 ( .A1(n12625), .A2(n11528), .ZN(n9642) );
  INV_X1 U12053 ( .A(n15546), .ZN(n11584) );
  NAND2_X1 U12054 ( .A1(n12823), .A2(n11584), .ZN(n9643) );
  NAND2_X1 U12055 ( .A1(n6689), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9649) );
  INV_X1 U12056 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11302) );
  OR2_X1 U12057 ( .A1(n6668), .A2(n11302), .ZN(n9648) );
  AND2_X1 U12058 ( .A1(n9644), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9645) );
  NOR2_X1 U12059 ( .A1(n9660), .A2(n9645), .ZN(n15480) );
  OR2_X1 U12060 ( .A1(n9600), .A2(n15480), .ZN(n9647) );
  INV_X1 U12061 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11303) );
  OR2_X1 U12062 ( .A1(n6683), .A2(n11303), .ZN(n9646) );
  NAND4_X1 U12063 ( .A1(n9649), .A2(n9648), .A3(n9647), .A4(n9646), .ZN(n12822) );
  OR2_X1 U12064 ( .A1(n9650), .A2(n9720), .ZN(n9652) );
  XNOR2_X1 U12065 ( .A(n9652), .B(n9651), .ZN(n15416) );
  INV_X1 U12066 ( .A(n15416), .ZN(n11304) );
  OR2_X1 U12067 ( .A1(n6687), .A2(SI_7_), .ZN(n9657) );
  INV_X1 U12068 ( .A(n9653), .ZN(n9654) );
  XNOR2_X1 U12069 ( .A(n6675), .B(n9654), .ZN(n10296) );
  OR2_X1 U12070 ( .A1(n9742), .A2(n10296), .ZN(n9656) );
  OAI211_X1 U12071 ( .C1(n11304), .C2(n10807), .A(n9657), .B(n9656), .ZN(
        n15478) );
  OR2_X1 U12072 ( .A1(n12822), .A2(n15478), .ZN(n12688) );
  NAND2_X1 U12073 ( .A1(n12822), .A2(n15478), .ZN(n12687) );
  NAND2_X1 U12074 ( .A1(n12688), .A2(n12687), .ZN(n15470) );
  INV_X1 U12075 ( .A(n15478), .ZN(n11613) );
  NAND2_X1 U12076 ( .A1(n12822), .A2(n11613), .ZN(n9658) );
  NAND2_X1 U12077 ( .A1(n6688), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9666) );
  INV_X1 U12078 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11309) );
  OR2_X1 U12079 ( .A1(n6667), .A2(n11309), .ZN(n9665) );
  NOR2_X1 U12080 ( .A1(n9660), .A2(n9659), .ZN(n9661) );
  OR2_X1 U12081 ( .A1(n9674), .A2(n9661), .ZN(n11826) );
  INV_X1 U12082 ( .A(n11826), .ZN(n9662) );
  OR2_X1 U12083 ( .A1(n9600), .A2(n9662), .ZN(n9664) );
  INV_X1 U12084 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11310) );
  OR2_X1 U12085 ( .A1(n6683), .A2(n11310), .ZN(n9663) );
  NAND4_X1 U12086 ( .A1(n9666), .A2(n9665), .A3(n9664), .A4(n9663), .ZN(n12821) );
  INV_X1 U12087 ( .A(SI_8_), .ZN(n10293) );
  OR2_X1 U12088 ( .A1(n6687), .A2(n10293), .ZN(n9673) );
  XNOR2_X1 U12089 ( .A(n9668), .B(n9667), .ZN(n10292) );
  OR2_X1 U12090 ( .A1(n9742), .A2(n10292), .ZN(n9672) );
  NAND2_X1 U12091 ( .A1(n9669), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9670) );
  XNOR2_X1 U12092 ( .A(n9670), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11311) );
  INV_X1 U12093 ( .A(n11311), .ZN(n15435) );
  OR2_X1 U12094 ( .A1(n10807), .A2(n15435), .ZN(n9671) );
  NAND2_X1 U12095 ( .A1(n12821), .A2(n11824), .ZN(n12693) );
  INV_X1 U12096 ( .A(n11824), .ZN(n11680) );
  NOR2_X1 U12097 ( .A1(n12821), .A2(n11680), .ZN(n11839) );
  NAND2_X1 U12098 ( .A1(n6688), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9679) );
  INV_X1 U12099 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11316) );
  OR2_X1 U12100 ( .A1(n6668), .A2(n11316), .ZN(n9678) );
  OR2_X1 U12101 ( .A1(n9674), .A2(n11700), .ZN(n9675) );
  AND2_X1 U12102 ( .A1(n9690), .A2(n9675), .ZN(n11699) );
  OR2_X1 U12103 ( .A1(n9600), .A2(n11699), .ZN(n9677) );
  INV_X1 U12104 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11851) );
  OR2_X1 U12105 ( .A1(n6684), .A2(n11851), .ZN(n9676) );
  NAND4_X1 U12106 ( .A1(n9679), .A2(n9678), .A3(n9677), .A4(n9676), .ZN(n12820) );
  INV_X1 U12107 ( .A(n9680), .ZN(n9681) );
  XNOR2_X1 U12108 ( .A(n9682), .B(n9681), .ZN(n10299) );
  OR2_X1 U12109 ( .A1(n9742), .A2(n10299), .ZN(n9686) );
  OR2_X1 U12110 ( .A1(n6687), .A2(SI_9_), .ZN(n9685) );
  OR2_X1 U12111 ( .A1(n9669), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9697) );
  NAND2_X1 U12112 ( .A1(n9697), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9683) );
  XNOR2_X1 U12113 ( .A(n9683), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11317) );
  OR2_X1 U12114 ( .A1(n10807), .A2(n11317), .ZN(n9684) );
  NAND2_X1 U12115 ( .A1(n12820), .A2(n12698), .ZN(n9689) );
  OR2_X1 U12116 ( .A1(n12820), .A2(n12698), .ZN(n9687) );
  NAND2_X1 U12117 ( .A1(n9689), .A2(n9687), .ZN(n12696) );
  NOR2_X1 U12118 ( .A1(n11839), .A2(n12696), .ZN(n9688) );
  NAND2_X1 U12119 ( .A1(n6689), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9696) );
  INV_X1 U12120 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11322) );
  OR2_X1 U12121 ( .A1(n6667), .A2(n11322), .ZN(n9695) );
  NAND2_X1 U12122 ( .A1(n9690), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9691) );
  AND2_X1 U12123 ( .A1(n9709), .A2(n9691), .ZN(n11985) );
  OR2_X1 U12124 ( .A1(n9600), .A2(n11985), .ZN(n9694) );
  INV_X1 U12125 ( .A(n6684), .ZN(n9692) );
  INV_X1 U12126 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11988) );
  OR2_X1 U12127 ( .A1(n6683), .A2(n11988), .ZN(n9693) );
  NAND4_X1 U12128 ( .A1(n9696), .A2(n9695), .A3(n9694), .A4(n9693), .ZN(n14852) );
  NAND2_X1 U12129 ( .A1(n9718), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9699) );
  XNOR2_X1 U12130 ( .A(n9699), .B(n9698), .ZN(n11470) );
  INV_X1 U12131 ( .A(n11470), .ZN(n11323) );
  OR2_X1 U12132 ( .A1(n6687), .A2(SI_10_), .ZN(n9704) );
  INV_X1 U12133 ( .A(n9700), .ZN(n9701) );
  XNOR2_X1 U12134 ( .A(n9702), .B(n9701), .ZN(n10306) );
  OR2_X1 U12135 ( .A1(n9742), .A2(n10306), .ZN(n9703) );
  OAI211_X1 U12136 ( .C1(n11323), .C2(n6680), .A(n9704), .B(n9703), .ZN(n11984) );
  OR2_X1 U12137 ( .A1(n14852), .A2(n11984), .ZN(n12704) );
  NAND2_X1 U12138 ( .A1(n14852), .A2(n11984), .ZN(n12710) );
  NAND2_X1 U12139 ( .A1(n12704), .A2(n12710), .ZN(n12701) );
  NAND2_X1 U12140 ( .A1(n11977), .A2(n12701), .ZN(n9706) );
  INV_X1 U12141 ( .A(n11984), .ZN(n11748) );
  NAND2_X1 U12142 ( .A1(n14852), .A2(n11748), .ZN(n9705) );
  NAND2_X1 U12143 ( .A1(n6688), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9715) );
  INV_X1 U12144 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n9707) );
  OR2_X1 U12145 ( .A1(n6667), .A2(n9707), .ZN(n9714) );
  INV_X1 U12146 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n9708) );
  OR2_X1 U12147 ( .A1(n6683), .A2(n9708), .ZN(n9713) );
  NAND2_X1 U12148 ( .A1(n9709), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9710) );
  NAND2_X1 U12149 ( .A1(n9732), .A2(n9710), .ZN(n14856) );
  INV_X1 U12150 ( .A(n14856), .ZN(n9711) );
  OR2_X1 U12151 ( .A1(n9600), .A2(n9711), .ZN(n9712) );
  NAND4_X1 U12152 ( .A1(n9715), .A2(n9714), .A3(n9713), .A4(n9712), .ZN(n12819) );
  XNOR2_X1 U12153 ( .A(n10469), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n9716) );
  XNOR2_X1 U12154 ( .A(n9717), .B(n9716), .ZN(n10319) );
  OR2_X1 U12155 ( .A1(n9742), .A2(n10319), .ZN(n9727) );
  OR2_X1 U12156 ( .A1(n6687), .A2(SI_11_), .ZN(n9726) );
  NOR2_X1 U12157 ( .A1(n9718), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n9722) );
  NOR2_X1 U12158 ( .A1(n9722), .A2(n9720), .ZN(n9719) );
  MUX2_X1 U12159 ( .A(n9720), .B(n9719), .S(P3_IR_REG_11__SCAN_IN), .Z(n9724)
         );
  NAND2_X1 U12160 ( .A1(n9722), .A2(n9721), .ZN(n9743) );
  INV_X1 U12161 ( .A(n9743), .ZN(n9723) );
  OR2_X1 U12162 ( .A1(n10807), .A2(n11667), .ZN(n9725) );
  AND2_X1 U12163 ( .A1(n12819), .A2(n11996), .ZN(n9729) );
  OR2_X1 U12164 ( .A1(n12819), .A2(n11996), .ZN(n9728) );
  OAI21_X1 U12165 ( .B1(n14850), .B2(n9729), .A(n9728), .ZN(n9730) );
  NAND2_X1 U12166 ( .A1(n9692), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9737) );
  INV_X1 U12167 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n9731) );
  OR2_X1 U12168 ( .A1(n6668), .A2(n9731), .ZN(n9736) );
  NOR2_X1 U12169 ( .A1(n9756), .A2(n7659), .ZN(n12080) );
  OR2_X1 U12170 ( .A1(n9600), .A2(n12080), .ZN(n9735) );
  INV_X1 U12171 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n9733) );
  OR2_X1 U12172 ( .A1(n9908), .A2(n9733), .ZN(n9734) );
  NAND4_X1 U12173 ( .A1(n9737), .A2(n9736), .A3(n9735), .A4(n9734), .ZN(n14854) );
  NAND2_X1 U12174 ( .A1(n9739), .A2(n9738), .ZN(n9740) );
  NAND2_X1 U12175 ( .A1(n9741), .A2(n9740), .ZN(n10338) );
  OR2_X1 U12176 ( .A1(n9742), .A2(n10338), .ZN(n9750) );
  OR2_X1 U12177 ( .A1(n9591), .A2(n10339), .ZN(n9749) );
  NAND2_X1 U12178 ( .A1(n9743), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9745) );
  MUX2_X1 U12179 ( .A(n9745), .B(P3_IR_REG_31__SCAN_IN), .S(n9744), .Z(n9747)
         );
  AND2_X1 U12180 ( .A1(n9747), .A2(n9843), .ZN(n11665) );
  OR2_X1 U12181 ( .A1(n10807), .A2(n11958), .ZN(n9748) );
  NAND2_X1 U12182 ( .A1(n14854), .A2(n12079), .ZN(n12709) );
  NAND2_X1 U12183 ( .A1(n12717), .A2(n12709), .ZN(n12073) );
  INV_X1 U12184 ( .A(n12079), .ZN(n12056) );
  NAND2_X1 U12185 ( .A1(n14854), .A2(n12056), .ZN(n9751) );
  XNOR2_X1 U12186 ( .A(n9752), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10432) );
  NAND2_X1 U12187 ( .A1(n10432), .A2(n12602), .ZN(n9755) );
  INV_X1 U12188 ( .A(n10807), .ZN(n9849) );
  NAND2_X1 U12189 ( .A1(n9843), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9753) );
  XNOR2_X1 U12190 ( .A(n9753), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12828) );
  AOI22_X1 U12191 ( .A1(n9850), .A2(SI_13_), .B1(n9849), .B2(n12828), .ZN(
        n9754) );
  NAND2_X1 U12192 ( .A1(n9755), .A2(n9754), .ZN(n14846) );
  NAND2_X1 U12193 ( .A1(n6688), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9763) );
  OR2_X1 U12194 ( .A1(n6668), .A2(n14875), .ZN(n9762) );
  INV_X1 U12195 ( .A(n9756), .ZN(n9757) );
  NAND2_X1 U12196 ( .A1(n9757), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U12197 ( .A1(n9769), .A2(n9758), .ZN(n14843) );
  INV_X1 U12198 ( .A(n14843), .ZN(n12147) );
  OR2_X1 U12199 ( .A1(n9600), .A2(n12147), .ZN(n9761) );
  INV_X1 U12200 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n9759) );
  OR2_X1 U12201 ( .A1(n6684), .A2(n9759), .ZN(n9760) );
  NAND4_X1 U12202 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n12818) );
  XNOR2_X1 U12203 ( .A(n9765), .B(n9764), .ZN(n14778) );
  NAND2_X1 U12204 ( .A1(n14778), .A2(n12602), .ZN(n9768) );
  OAI21_X1 U12205 ( .B1(n9843), .B2(P3_IR_REG_13__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9766) );
  INV_X1 U12206 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9779) );
  XNOR2_X1 U12207 ( .A(n9766), .B(n9779), .ZN(n14781) );
  AOI22_X1 U12208 ( .A1(n9850), .A2(n14777), .B1(n9849), .B2(n14781), .ZN(
        n9767) );
  NAND2_X1 U12209 ( .A1(n9768), .A2(n9767), .ZN(n13284) );
  NAND2_X1 U12210 ( .A1(n6689), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9775) );
  INV_X1 U12211 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13230) );
  OR2_X1 U12212 ( .A1(n6667), .A2(n13230), .ZN(n9774) );
  NAND2_X1 U12213 ( .A1(n9769), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9770) );
  AND2_X1 U12214 ( .A1(n9790), .A2(n9770), .ZN(n12181) );
  OR2_X1 U12215 ( .A1(n9600), .A2(n12181), .ZN(n9773) );
  INV_X1 U12216 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n9771) );
  OR2_X1 U12217 ( .A1(n6683), .A2(n9771), .ZN(n9772) );
  NAND4_X1 U12218 ( .A1(n9775), .A2(n9774), .A3(n9773), .A4(n9772), .ZN(n14841) );
  OR2_X1 U12219 ( .A1(n13284), .A2(n14841), .ZN(n12722) );
  NAND2_X1 U12220 ( .A1(n13284), .A2(n14841), .ZN(n12723) );
  NAND2_X1 U12221 ( .A1(n12722), .A2(n12723), .ZN(n13156) );
  INV_X1 U12222 ( .A(n14841), .ZN(n12429) );
  OR2_X1 U12223 ( .A1(n13284), .A2(n12429), .ZN(n13138) );
  INV_X1 U12224 ( .A(n9776), .ZN(n9777) );
  XNOR2_X1 U12225 ( .A(n9778), .B(n9777), .ZN(n10473) );
  NAND2_X1 U12226 ( .A1(n10473), .A2(n12602), .ZN(n9788) );
  NAND2_X1 U12227 ( .A1(n9780), .A2(n9779), .ZN(n9781) );
  NOR2_X1 U12228 ( .A1(n9843), .A2(n9781), .ZN(n9784) );
  NOR2_X1 U12229 ( .A1(n9784), .A2(n9720), .ZN(n9782) );
  MUX2_X1 U12230 ( .A(n9720), .B(n9782), .S(P3_IR_REG_15__SCAN_IN), .Z(n9786)
         );
  INV_X1 U12231 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9783) );
  NAND2_X1 U12232 ( .A1(n9784), .A2(n9783), .ZN(n9815) );
  INV_X1 U12233 ( .A(n9815), .ZN(n9785) );
  AOI22_X1 U12234 ( .A1(n9850), .A2(SI_15_), .B1(n9849), .B2(n12898), .ZN(
        n9787) );
  NAND2_X1 U12235 ( .A1(n9788), .A2(n9787), .ZN(n13278) );
  NAND2_X1 U12236 ( .A1(n6688), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9795) );
  INV_X1 U12237 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n9789) );
  OR2_X1 U12238 ( .A1(n6668), .A2(n9789), .ZN(n9794) );
  NAND2_X1 U12239 ( .A1(n9790), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9791) );
  AND2_X1 U12240 ( .A1(n9805), .A2(n9791), .ZN(n13145) );
  OR2_X1 U12241 ( .A1(n9600), .A2(n13145), .ZN(n9793) );
  INV_X1 U12242 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13146) );
  OR2_X1 U12243 ( .A1(n6684), .A2(n13146), .ZN(n9792) );
  INV_X1 U12244 ( .A(n13159), .ZN(n12817) );
  NAND2_X1 U12245 ( .A1(n13278), .A2(n12817), .ZN(n9796) );
  AND2_X1 U12246 ( .A1(n13138), .A2(n9796), .ZN(n9798) );
  INV_X1 U12247 ( .A(n9796), .ZN(n9797) );
  OR2_X1 U12248 ( .A1(n13278), .A2(n13159), .ZN(n12727) );
  NAND2_X1 U12249 ( .A1(n13278), .A2(n13159), .ZN(n12731) );
  NAND2_X1 U12250 ( .A1(n12727), .A2(n12731), .ZN(n9988) );
  INV_X1 U12251 ( .A(n9799), .ZN(n9800) );
  XNOR2_X1 U12252 ( .A(n9801), .B(n9800), .ZN(n10493) );
  NAND2_X1 U12253 ( .A1(n10493), .A2(n12602), .ZN(n9804) );
  NAND2_X1 U12254 ( .A1(n9815), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9802) );
  XNOR2_X1 U12255 ( .A(n9802), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12912) );
  AOI22_X1 U12256 ( .A1(n9850), .A2(SI_16_), .B1(n9849), .B2(n12912), .ZN(
        n9803) );
  NAND2_X1 U12257 ( .A1(n9804), .A2(n9803), .ZN(n12515) );
  NAND2_X1 U12258 ( .A1(n6688), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9810) );
  INV_X1 U12259 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13220) );
  OR2_X1 U12260 ( .A1(n6667), .A2(n13220), .ZN(n9809) );
  NAND2_X1 U12261 ( .A1(n9805), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9806) );
  AND2_X1 U12262 ( .A1(n9820), .A2(n9806), .ZN(n13131) );
  OR2_X1 U12263 ( .A1(n9600), .A2(n13131), .ZN(n9808) );
  INV_X1 U12264 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13132) );
  OR2_X1 U12265 ( .A1(n6683), .A2(n13132), .ZN(n9807) );
  OR2_X1 U12266 ( .A1(n12515), .A2(n13142), .ZN(n12733) );
  NAND2_X1 U12267 ( .A1(n12515), .A2(n13142), .ZN(n12732) );
  NAND2_X1 U12268 ( .A1(n12733), .A2(n12732), .ZN(n13128) );
  NAND2_X1 U12269 ( .A1(n13127), .A2(n13128), .ZN(n9812) );
  INV_X1 U12270 ( .A(n13142), .ZN(n12531) );
  NAND2_X1 U12271 ( .A1(n12515), .A2(n12531), .ZN(n9811) );
  XNOR2_X1 U12272 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n9813) );
  XNOR2_X1 U12273 ( .A(n9814), .B(n9813), .ZN(n10578) );
  NAND2_X1 U12274 ( .A1(n10578), .A2(n12602), .ZN(n9819) );
  OR2_X1 U12275 ( .A1(n9815), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U12276 ( .A1(n9830), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9817) );
  XNOR2_X1 U12277 ( .A(n9817), .B(n9816), .ZN(n14824) );
  AOI22_X1 U12278 ( .A1(n9850), .A2(n10579), .B1(n9849), .B2(n14824), .ZN(
        n9818) );
  NAND2_X1 U12279 ( .A1(n9570), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9825) );
  INV_X1 U12280 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14567) );
  OR2_X1 U12281 ( .A1(n9908), .A2(n14567), .ZN(n9824) );
  NAND2_X1 U12282 ( .A1(n9820), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9821) );
  AND2_X1 U12283 ( .A1(n9834), .A2(n9821), .ZN(n13119) );
  OR2_X1 U12284 ( .A1(n9600), .A2(n13119), .ZN(n9823) );
  INV_X1 U12285 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14834) );
  OR2_X1 U12286 ( .A1(n6684), .A2(n14834), .ZN(n9822) );
  NAND4_X1 U12287 ( .A1(n9825), .A2(n9824), .A3(n9823), .A4(n9822), .ZN(n13101) );
  NAND2_X1 U12288 ( .A1(n13271), .A2(n13101), .ZN(n12737) );
  NAND2_X1 U12289 ( .A1(n12736), .A2(n12737), .ZN(n13115) );
  OR2_X1 U12290 ( .A1(n13271), .A2(n13130), .ZN(n9826) );
  XNOR2_X1 U12291 ( .A(n11548), .B(P2_DATAO_REG_18__SCAN_IN), .ZN(n9828) );
  XNOR2_X1 U12292 ( .A(n9829), .B(n9828), .ZN(n10652) );
  NAND2_X1 U12293 ( .A1(n10652), .A2(n12602), .ZN(n9833) );
  OAI21_X1 U12294 ( .B1(n9830), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9831) );
  XNOR2_X1 U12295 ( .A(n9831), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12944) );
  AOI22_X1 U12296 ( .A1(n9850), .A2(SI_18_), .B1(n9849), .B2(n12944), .ZN(
        n9832) );
  NAND2_X1 U12297 ( .A1(n6689), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9838) );
  INV_X1 U12298 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12943) );
  OR2_X1 U12299 ( .A1(n6667), .A2(n12943), .ZN(n9837) );
  XNOR2_X1 U12300 ( .A(n9834), .B(n12564), .ZN(n13104) );
  OR2_X1 U12301 ( .A1(n9600), .A2(n13104), .ZN(n9836) );
  INV_X1 U12302 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13105) );
  OR2_X1 U12303 ( .A1(n6684), .A2(n13105), .ZN(n9835) );
  NAND2_X1 U12304 ( .A1(n13267), .A2(n13118), .ZN(n12743) );
  INV_X1 U12305 ( .A(n13118), .ZN(n13086) );
  OR2_X1 U12306 ( .A1(n13267), .A2(n13086), .ZN(n9839) );
  INV_X1 U12307 ( .A(n9840), .ZN(n9841) );
  XNOR2_X1 U12308 ( .A(n9842), .B(n9841), .ZN(n10712) );
  NAND2_X1 U12309 ( .A1(n10712), .A2(n12602), .ZN(n9852) );
  INV_X1 U12310 ( .A(n9847), .ZN(n9844) );
  NAND2_X1 U12311 ( .A1(n9844), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9845) );
  MUX2_X1 U12312 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9845), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n9848) );
  NAND2_X1 U12313 ( .A1(n9848), .A2(n9964), .ZN(n12942) );
  AOI22_X1 U12314 ( .A1(n9850), .A2(n10711), .B1(n9849), .B2(n12942), .ZN(
        n9851) );
  NAND2_X1 U12315 ( .A1(n6689), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9859) );
  INV_X1 U12316 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13206) );
  OR2_X1 U12317 ( .A1(n6668), .A2(n13206), .ZN(n9858) );
  INV_X1 U12318 ( .A(n9853), .ZN(n9854) );
  NAND2_X1 U12319 ( .A1(n9854), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9855) );
  AND2_X1 U12320 ( .A1(n9864), .A2(n9855), .ZN(n13089) );
  OR2_X1 U12321 ( .A1(n9600), .A2(n13089), .ZN(n9857) );
  INV_X1 U12322 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13090) );
  OR2_X1 U12323 ( .A1(n6684), .A2(n13090), .ZN(n9856) );
  NAND4_X1 U12324 ( .A1(n9859), .A2(n9858), .A3(n9857), .A4(n9856), .ZN(n13100) );
  NAND2_X1 U12325 ( .A1(n13264), .A2(n13100), .ZN(n12759) );
  INV_X1 U12326 ( .A(n13100), .ZN(n12549) );
  OR2_X1 U12327 ( .A1(n13264), .A2(n12549), .ZN(n9860) );
  XNOR2_X1 U12328 ( .A(n9861), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11058) );
  NAND2_X1 U12329 ( .A1(n11058), .A2(n12602), .ZN(n9863) );
  OR2_X1 U12330 ( .A1(n9591), .A2(n11059), .ZN(n9862) );
  NAND2_X1 U12331 ( .A1(n9864), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9865) );
  NAND2_X1 U12332 ( .A1(n9881), .A2(n9865), .ZN(n13072) );
  NAND2_X1 U12333 ( .A1(n9954), .A2(n13072), .ZN(n9871) );
  INV_X1 U12334 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n9866) );
  OR2_X1 U12335 ( .A1(n6668), .A2(n9866), .ZN(n9870) );
  INV_X1 U12336 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13074) );
  OR2_X1 U12337 ( .A1(n6683), .A2(n13074), .ZN(n9869) );
  INV_X1 U12338 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n14588) );
  OR2_X1 U12339 ( .A1(n9908), .A2(n14588), .ZN(n9868) );
  XNOR2_X1 U12340 ( .A(n13076), .B(n13058), .ZN(n13079) );
  NAND2_X1 U12341 ( .A1(n13076), .A2(n13085), .ZN(n9872) );
  XNOR2_X1 U12342 ( .A(n9875), .B(n9874), .ZN(n11205) );
  NAND2_X1 U12343 ( .A1(n11205), .A2(n12602), .ZN(n9877) );
  OR2_X1 U12344 ( .A1(n6687), .A2(n11206), .ZN(n9876) );
  INV_X1 U12345 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n9878) );
  OR2_X1 U12346 ( .A1(n9908), .A2(n9878), .ZN(n9880) );
  INV_X1 U12347 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n14663) );
  OR2_X1 U12348 ( .A1(n6668), .A2(n14663), .ZN(n9879) );
  AND2_X1 U12349 ( .A1(n9880), .A2(n9879), .ZN(n9885) );
  NAND2_X1 U12350 ( .A1(n9881), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U12351 ( .A1(n9892), .A2(n9882), .ZN(n13061) );
  NAND2_X1 U12352 ( .A1(n13061), .A2(n9954), .ZN(n9884) );
  NAND2_X1 U12353 ( .A1(n9692), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U12354 ( .A1(n13258), .A2(n13042), .ZN(n12750) );
  OR2_X1 U12355 ( .A1(n13258), .A2(n13070), .ZN(n9886) );
  XNOR2_X1 U12356 ( .A(n9888), .B(n9887), .ZN(n11260) );
  NAND2_X1 U12357 ( .A1(n11260), .A2(n12602), .ZN(n9891) );
  INV_X1 U12358 ( .A(SI_22_), .ZN(n9889) );
  OR2_X1 U12359 ( .A1(n6687), .A2(n9889), .ZN(n9890) );
  INV_X1 U12360 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U12361 ( .A1(n9892), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9893) );
  NAND2_X1 U12362 ( .A1(n9894), .A2(n9893), .ZN(n13048) );
  NAND2_X1 U12363 ( .A1(n13048), .A2(n9954), .ZN(n9896) );
  AOI22_X1 U12364 ( .A1(n6689), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n9570), .B2(
        P3_REG1_REG_22__SCAN_IN), .ZN(n9895) );
  OAI211_X1 U12365 ( .C1(n6683), .C2(n9897), .A(n9896), .B(n9895), .ZN(n13056)
         );
  NAND2_X1 U12366 ( .A1(n12453), .A2(n13056), .ZN(n9898) );
  NAND2_X1 U12367 ( .A1(n12767), .A2(n13043), .ZN(n9899) );
  NAND2_X1 U12368 ( .A1(n13009), .A2(n9899), .ZN(n13031) );
  XNOR2_X1 U12369 ( .A(n9900), .B(n7157), .ZN(n12265) );
  NAND2_X1 U12370 ( .A1(n12265), .A2(n12602), .ZN(n9902) );
  INV_X1 U12371 ( .A(SI_24_), .ZN(n12266) );
  OR2_X1 U12372 ( .A1(n6687), .A2(n12266), .ZN(n9901) );
  NAND2_X1 U12373 ( .A1(n9903), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U12374 ( .A1(n9905), .A2(n9904), .ZN(n13021) );
  NAND2_X1 U12375 ( .A1(n13021), .A2(n9954), .ZN(n9911) );
  INV_X1 U12376 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13245) );
  NAND2_X1 U12377 ( .A1(n9692), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9907) );
  NAND2_X1 U12378 ( .A1(n9570), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9906) );
  OAI211_X1 U12379 ( .C1(n9908), .C2(n13245), .A(n9907), .B(n9906), .ZN(n9909)
         );
  INV_X1 U12380 ( .A(n9909), .ZN(n9910) );
  NAND2_X1 U12381 ( .A1(n13017), .A2(n13016), .ZN(n13015) );
  OR2_X1 U12382 ( .A1(n13013), .A2(n9914), .ZN(n12776) );
  NAND2_X1 U12383 ( .A1(n9914), .A2(n13013), .ZN(n12777) );
  NAND2_X1 U12384 ( .A1(n12776), .A2(n12777), .ZN(n12998) );
  NAND2_X1 U12385 ( .A1(n12999), .A2(n12998), .ZN(n12997) );
  AOI22_X1 U12386 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n13845), .B2(n14392), .ZN(n9915) );
  INV_X1 U12387 ( .A(n9915), .ZN(n9916) );
  XNOR2_X1 U12388 ( .A(n9917), .B(n9916), .ZN(n11973) );
  NAND2_X1 U12389 ( .A1(n11973), .A2(n12602), .ZN(n9919) );
  INV_X1 U12390 ( .A(SI_26_), .ZN(n11975) );
  NAND2_X1 U12391 ( .A1(n9920), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U12392 ( .A1(n9937), .A2(n9921), .ZN(n12989) );
  NAND2_X1 U12393 ( .A1(n12989), .A2(n9954), .ZN(n9926) );
  INV_X1 U12394 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13238) );
  NAND2_X1 U12395 ( .A1(n9692), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U12396 ( .A1(n9570), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9922) );
  OAI211_X1 U12397 ( .C1(n9908), .C2(n13238), .A(n9923), .B(n9922), .ZN(n9924)
         );
  INV_X1 U12398 ( .A(n9924), .ZN(n9925) );
  NAND2_X1 U12399 ( .A1(n12984), .A2(n9929), .ZN(n9931) );
  NAND2_X1 U12400 ( .A1(n12467), .A2(n12996), .ZN(n9930) );
  AOI22_X1 U12401 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n12271), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n14390), .ZN(n9932) );
  INV_X1 U12402 ( .A(n9932), .ZN(n9933) );
  XNOR2_X1 U12403 ( .A(n9934), .B(n9933), .ZN(n12303) );
  NAND2_X1 U12404 ( .A1(n12303), .A2(n12602), .ZN(n9936) );
  INV_X1 U12405 ( .A(SI_27_), .ZN(n12304) );
  NAND2_X1 U12406 ( .A1(n9937), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U12407 ( .A1(n9939), .A2(n9938), .ZN(n12475) );
  NAND2_X1 U12408 ( .A1(n12475), .A2(n9954), .ZN(n9944) );
  INV_X1 U12409 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n14580) );
  NAND2_X1 U12410 ( .A1(n6689), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9941) );
  INV_X1 U12411 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12285) );
  OR2_X1 U12412 ( .A1(n6683), .A2(n12285), .ZN(n9940) );
  OAI211_X1 U12413 ( .C1(n6668), .C2(n14580), .A(n9941), .B(n9940), .ZN(n9942)
         );
  INV_X1 U12414 ( .A(n9942), .ZN(n9943) );
  NAND2_X1 U12415 ( .A1(n12470), .A2(n12986), .ZN(n9993) );
  NAND2_X1 U12416 ( .A1(n9947), .A2(n12473), .ZN(n12790) );
  NOR2_X1 U12417 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n7129), .ZN(n9949) );
  OAI22_X1 U12418 ( .A1(n14597), .A2(n12294), .B1(P1_DATAO_REG_29__SCAN_IN), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12421) );
  INV_X1 U12419 ( .A(n12421), .ZN(n9950) );
  XNOR2_X1 U12420 ( .A(n12420), .B(n9950), .ZN(n12295) );
  NAND2_X1 U12421 ( .A1(n12295), .A2(n12602), .ZN(n9952) );
  OR2_X1 U12422 ( .A1(n9591), .A2(n12297), .ZN(n9951) );
  NAND2_X1 U12423 ( .A1(n12960), .A2(n9954), .ZN(n12612) );
  INV_X1 U12424 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12966) );
  NAND2_X1 U12425 ( .A1(n6688), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U12426 ( .A1(n9570), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9955) );
  OAI211_X1 U12427 ( .C1(n6684), .C2(n12966), .A(n9956), .B(n9955), .ZN(n9957)
         );
  INV_X1 U12428 ( .A(n9957), .ZN(n9958) );
  NAND2_X1 U12429 ( .A1(n12968), .A2(n12977), .ZN(n12617) );
  NAND2_X1 U12430 ( .A1(n12792), .A2(n12617), .ZN(n12648) );
  XNOR2_X1 U12431 ( .A(n9959), .B(n12648), .ZN(n9977) );
  NAND2_X1 U12432 ( .A1(n9960), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9961) );
  NAND2_X1 U12433 ( .A1(n12810), .A2(n12649), .ZN(n10047) );
  NAND2_X1 U12434 ( .A1(n9966), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9963) );
  NAND2_X1 U12435 ( .A1(n9964), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9965) );
  MUX2_X1 U12436 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9965), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9967) );
  INV_X1 U12437 ( .A(n11061), .ZN(n10033) );
  NAND2_X1 U12438 ( .A1(n11381), .A2(n10033), .ZN(n12622) );
  INV_X1 U12439 ( .A(n9968), .ZN(n12807) );
  NAND2_X1 U12440 ( .A1(n12807), .A2(n10825), .ZN(n10817) );
  NAND2_X1 U12441 ( .A1(n6669), .A2(n10817), .ZN(n10995) );
  AND2_X2 U12442 ( .A1(n12810), .A2(n11381), .ZN(n12780) );
  INV_X1 U12443 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14870) );
  NAND2_X1 U12444 ( .A1(n6689), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U12445 ( .A1(n9692), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9969) );
  OAI211_X1 U12446 ( .C1(n6668), .C2(n14870), .A(n9970), .B(n9969), .ZN(n9971)
         );
  INV_X1 U12447 ( .A(n9971), .ZN(n9972) );
  AND2_X1 U12448 ( .A1(n12807), .A2(P3_B_REG_SCAN_IN), .ZN(n9973) );
  OR2_X1 U12449 ( .A1(n15507), .A2(n9973), .ZN(n12957) );
  INV_X1 U12450 ( .A(n10994), .ZN(n9978) );
  INV_X1 U12451 ( .A(n9979), .ZN(n12627) );
  NAND2_X1 U12452 ( .A1(n15487), .A2(n12627), .ZN(n15486) );
  NAND2_X1 U12453 ( .A1(n15486), .A2(n12659), .ZN(n11379) );
  INV_X1 U12454 ( .A(n12626), .ZN(n11380) );
  NAND2_X1 U12455 ( .A1(n11379), .A2(n11380), .ZN(n9980) );
  NAND2_X1 U12456 ( .A1(n9980), .A2(n12669), .ZN(n11854) );
  INV_X1 U12457 ( .A(n12630), .ZN(n12671) );
  OR2_X1 U12458 ( .A1(n12824), .A2(n15534), .ZN(n9981) );
  INV_X1 U12459 ( .A(n12625), .ZN(n9982) );
  NAND2_X1 U12460 ( .A1(n11527), .A2(n9982), .ZN(n9983) );
  NAND2_X1 U12461 ( .A1(n9983), .A2(n12686), .ZN(n15469) );
  NAND2_X1 U12462 ( .A1(n12820), .A2(n11703), .ZN(n9984) );
  OR2_X1 U12463 ( .A1(n12820), .A2(n11703), .ZN(n9985) );
  XNOR2_X1 U12464 ( .A(n12819), .B(n14859), .ZN(n12711) );
  OR2_X1 U12465 ( .A1(n12819), .A2(n14859), .ZN(n12703) );
  AND2_X1 U12466 ( .A1(n13158), .A2(n14846), .ZN(n12636) );
  OR2_X1 U12467 ( .A1(n13158), .A2(n14846), .ZN(n12719) );
  NAND2_X1 U12468 ( .A1(n13160), .A2(n12722), .ZN(n13150) );
  INV_X1 U12469 ( .A(n13128), .ZN(n13125) );
  INV_X1 U12470 ( .A(n13115), .ZN(n13114) );
  NAND2_X1 U12471 ( .A1(n13113), .A2(n13114), .ZN(n9989) );
  OR2_X1 U12472 ( .A1(n13076), .A2(n13058), .ZN(n9990) );
  NAND2_X1 U12473 ( .A1(n13066), .A2(n12750), .ZN(n9991) );
  NAND2_X1 U12474 ( .A1(n9991), .A2(n12749), .ZN(n13047) );
  NAND2_X1 U12475 ( .A1(n12453), .A2(n12554), .ZN(n12757) );
  NAND2_X1 U12476 ( .A1(n13047), .A2(n12757), .ZN(n9992) );
  INV_X1 U12477 ( .A(n13031), .ZN(n13026) );
  INV_X2 U12478 ( .A(n13016), .ZN(n13008) );
  INV_X1 U12479 ( .A(n9993), .ZN(n12788) );
  INV_X1 U12480 ( .A(n12787), .ZN(n9994) );
  OAI21_X1 U12481 ( .B1(n10032), .B2(n10033), .A(n12649), .ZN(n9995) );
  NAND2_X1 U12482 ( .A1(n9995), .A2(n12651), .ZN(n9997) );
  OAI21_X1 U12483 ( .B1(n10033), .B2(n11381), .A(n10032), .ZN(n9996) );
  NAND2_X1 U12484 ( .A1(n9997), .A2(n9996), .ZN(n10916) );
  NAND2_X1 U12485 ( .A1(n11061), .A2(n12942), .ZN(n11002) );
  INV_X1 U12486 ( .A(n11002), .ZN(n12803) );
  AND2_X1 U12487 ( .A1(n15545), .A2(n12803), .ZN(n9998) );
  NAND2_X1 U12488 ( .A1(n10916), .A2(n9998), .ZN(n10000) );
  NOR2_X1 U12489 ( .A1(n11061), .A2(n12649), .ZN(n9999) );
  NAND2_X1 U12490 ( .A1(n12810), .A2(n9999), .ZN(n10036) );
  AND2_X1 U12491 ( .A1(n11061), .A2(n12649), .ZN(n12804) );
  XNOR2_X1 U12492 ( .A(n12268), .B(P3_B_REG_SCAN_IN), .ZN(n10008) );
  NAND2_X1 U12493 ( .A1(n10008), .A2(n11883), .ZN(n10013) );
  NAND2_X1 U12494 ( .A1(n10009), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10010) );
  MUX2_X1 U12495 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10010), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n10012) );
  OR2_X1 U12496 ( .A1(n10472), .A2(P3_D_REG_1__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U12497 ( .A1(n11883), .A2(n11976), .ZN(n10015) );
  NAND2_X1 U12498 ( .A1(n12268), .A2(n11976), .ZN(n10017) );
  NOR4_X1 U12499 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n10027) );
  INV_X1 U12500 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10482) );
  INV_X1 U12501 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n14694) );
  INV_X1 U12502 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n14585) );
  INV_X1 U12503 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n14608) );
  NAND4_X1 U12504 ( .A1(n10482), .A2(n14694), .A3(n14585), .A4(n14608), .ZN(
        n10024) );
  NOR4_X1 U12505 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n10022) );
  NOR4_X1 U12506 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n10021) );
  NOR4_X1 U12507 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n10020) );
  NOR4_X1 U12508 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n10019) );
  NAND4_X1 U12509 ( .A1(n10022), .A2(n10021), .A3(n10020), .A4(n10019), .ZN(
        n10023) );
  NOR4_X1 U12510 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        n10024), .A4(n10023), .ZN(n10026) );
  NOR4_X1 U12511 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n10025) );
  AND3_X1 U12512 ( .A1(n10027), .A2(n10026), .A3(n10025), .ZN(n10028) );
  NAND2_X1 U12513 ( .A1(n6822), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10030) );
  AND2_X1 U12514 ( .A1(n10049), .A2(n10932), .ZN(n10031) );
  OAI22_X1 U12515 ( .A1(n15545), .A2(n10033), .B1(n12649), .B2(n10032), .ZN(
        n10034) );
  NAND2_X1 U12516 ( .A1(n10034), .A2(n11002), .ZN(n10035) );
  NAND2_X1 U12517 ( .A1(n10035), .A2(n12794), .ZN(n10038) );
  AND2_X1 U12518 ( .A1(n12794), .A2(n10036), .ZN(n10793) );
  AND2_X1 U12519 ( .A1(n12780), .A2(n11002), .ZN(n10920) );
  OAI21_X1 U12520 ( .B1(n11001), .B2(n10038), .A(n10037), .ZN(n10039) );
  OR2_X1 U12521 ( .A1(n10053), .A2(n15583), .ZN(n10044) );
  INV_X1 U12522 ( .A(n12968), .ZN(n10054) );
  INV_X1 U12523 ( .A(n15545), .ZN(n11848) );
  NAND2_X1 U12524 ( .A1(n15585), .A2(n11848), .ZN(n13232) );
  INV_X1 U12525 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U12526 ( .A1(n10044), .A2(n10043), .ZN(P3_U3488) );
  INV_X1 U12527 ( .A(n10049), .ZN(n10045) );
  NAND2_X1 U12528 ( .A1(n10917), .A2(n10932), .ZN(n10935) );
  AND2_X1 U12529 ( .A1(n12780), .A2(n12803), .ZN(n10048) );
  AND2_X1 U12530 ( .A1(n10932), .A2(n10048), .ZN(n12808) );
  AND2_X1 U12531 ( .A1(n10932), .A2(n10916), .ZN(n10050) );
  AOI22_X1 U12532 ( .A1(n10917), .A2(n12808), .B1(n10998), .B2(n10050), .ZN(
        n10051) );
  OR2_X1 U12533 ( .A1(n10053), .A2(n15568), .ZN(n10059) );
  INV_X1 U12534 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U12535 ( .A1(n15570), .A2(n10056), .ZN(n10057) );
  NAND2_X1 U12536 ( .A1(n10059), .A2(n10058), .ZN(P3_U3456) );
  NAND2_X4 U12537 ( .A1(n10061), .A2(n10060), .ZN(n13316) );
  NAND2_X1 U12538 ( .A1(n10062), .A2(n10861), .ZN(n10065) );
  NAND2_X1 U12539 ( .A1(n10275), .A2(n10861), .ZN(n10656) );
  NAND2_X1 U12540 ( .A1(n10161), .A2(n10655), .ZN(n10063) );
  NAND2_X1 U12541 ( .A1(n10064), .A2(n10065), .ZN(n10066) );
  XNOR2_X1 U12542 ( .A(n10067), .B(n13316), .ZN(n10068) );
  NAND2_X1 U12543 ( .A1(n8475), .A2(n10861), .ZN(n10069) );
  XNOR2_X1 U12544 ( .A(n10068), .B(n10069), .ZN(n10680) );
  INV_X1 U12545 ( .A(n10068), .ZN(n10070) );
  NAND2_X1 U12546 ( .A1(n10070), .A2(n10069), .ZN(n10071) );
  XNOR2_X1 U12547 ( .A(n8480), .B(n13316), .ZN(n10776) );
  AND2_X1 U12548 ( .A1(n8479), .A2(n10861), .ZN(n10072) );
  NAND2_X1 U12549 ( .A1(n10776), .A2(n10072), .ZN(n10076) );
  INV_X1 U12550 ( .A(n10776), .ZN(n10074) );
  INV_X1 U12551 ( .A(n10072), .ZN(n10073) );
  NAND2_X1 U12552 ( .A1(n10074), .A2(n10073), .ZN(n10075) );
  AND2_X1 U12553 ( .A1(n10076), .A2(n10075), .ZN(n10628) );
  XNOR2_X1 U12554 ( .A(n10780), .B(n13316), .ZN(n10077) );
  NAND2_X1 U12555 ( .A1(n13450), .A2(n10861), .ZN(n10078) );
  XNOR2_X1 U12556 ( .A(n10077), .B(n10078), .ZN(n10775) );
  NAND3_X1 U12557 ( .A1(n10774), .A2(n10775), .A3(n10076), .ZN(n10773) );
  INV_X1 U12558 ( .A(n10077), .ZN(n10702) );
  NAND2_X1 U12559 ( .A1(n10702), .A2(n10078), .ZN(n10079) );
  NAND2_X1 U12560 ( .A1(n10773), .A2(n10079), .ZN(n10080) );
  XNOR2_X1 U12561 ( .A(n10848), .B(n13316), .ZN(n10081) );
  NAND2_X1 U12562 ( .A1(n13449), .A2(n10861), .ZN(n10082) );
  XNOR2_X1 U12563 ( .A(n10081), .B(n10082), .ZN(n10701) );
  INV_X1 U12564 ( .A(n10081), .ZN(n10083) );
  NAND2_X1 U12565 ( .A1(n10083), .A2(n10082), .ZN(n10084) );
  XNOR2_X1 U12566 ( .A(n11442), .B(n13316), .ZN(n10085) );
  AND2_X1 U12567 ( .A1(n13448), .A2(n10861), .ZN(n10086) );
  NAND2_X1 U12568 ( .A1(n10085), .A2(n10086), .ZN(n10090) );
  INV_X1 U12569 ( .A(n10085), .ZN(n11127) );
  INV_X1 U12570 ( .A(n10086), .ZN(n10087) );
  NAND2_X1 U12571 ( .A1(n11127), .A2(n10087), .ZN(n10088) );
  NAND2_X1 U12572 ( .A1(n10090), .A2(n10088), .ZN(n10888) );
  INV_X1 U12573 ( .A(n10888), .ZN(n10089) );
  XNOR2_X1 U12574 ( .A(n15348), .B(n13316), .ZN(n11157) );
  AND2_X1 U12575 ( .A1(n13447), .A2(n10861), .ZN(n10091) );
  NAND2_X1 U12576 ( .A1(n11157), .A2(n10091), .ZN(n10095) );
  INV_X1 U12577 ( .A(n11157), .ZN(n10093) );
  INV_X1 U12578 ( .A(n10091), .ZN(n10092) );
  NAND2_X1 U12579 ( .A1(n10093), .A2(n10092), .ZN(n10094) );
  AND2_X1 U12580 ( .A1(n10095), .A2(n10094), .ZN(n11124) );
  XNOR2_X1 U12581 ( .A(n11484), .B(n13316), .ZN(n11246) );
  NAND2_X1 U12582 ( .A1(n13446), .A2(n10861), .ZN(n10096) );
  XNOR2_X1 U12583 ( .A(n11246), .B(n10096), .ZN(n11160) );
  NAND3_X1 U12584 ( .A1(n11159), .A2(n11160), .A3(n10095), .ZN(n11251) );
  INV_X1 U12585 ( .A(n11246), .ZN(n10097) );
  NAND2_X1 U12586 ( .A1(n10097), .A2(n10096), .ZN(n10098) );
  NAND2_X1 U12587 ( .A1(n11251), .A2(n10098), .ZN(n10099) );
  XNOR2_X1 U12588 ( .A(n15355), .B(n13316), .ZN(n10100) );
  NAND2_X1 U12589 ( .A1(n13445), .A2(n10861), .ZN(n10101) );
  XNOR2_X1 U12590 ( .A(n10100), .B(n10101), .ZN(n11245) );
  INV_X1 U12591 ( .A(n10100), .ZN(n10102) );
  NAND2_X1 U12592 ( .A1(n10102), .A2(n10101), .ZN(n10103) );
  XNOR2_X1 U12593 ( .A(n11803), .B(n13316), .ZN(n10104) );
  AND2_X1 U12594 ( .A1(n13444), .A2(n10861), .ZN(n10105) );
  NAND2_X1 U12595 ( .A1(n10104), .A2(n10105), .ZN(n10109) );
  INV_X1 U12596 ( .A(n10104), .ZN(n11786) );
  INV_X1 U12597 ( .A(n10105), .ZN(n10106) );
  NAND2_X1 U12598 ( .A1(n11786), .A2(n10106), .ZN(n10107) );
  NAND2_X1 U12599 ( .A1(n10109), .A2(n10107), .ZN(n11800) );
  XNOR2_X1 U12600 ( .A(n15286), .B(n13316), .ZN(n10111) );
  NAND2_X1 U12601 ( .A1(n13443), .A2(n10861), .ZN(n10112) );
  XNOR2_X1 U12602 ( .A(n10111), .B(n10112), .ZN(n11788) );
  AND2_X1 U12603 ( .A1(n11788), .A2(n10109), .ZN(n10110) );
  INV_X1 U12604 ( .A(n10111), .ZN(n10113) );
  NAND2_X1 U12605 ( .A1(n10113), .A2(n10112), .ZN(n10114) );
  XNOR2_X1 U12606 ( .A(n11917), .B(n10161), .ZN(n10116) );
  NAND2_X1 U12607 ( .A1(n13442), .A2(n10861), .ZN(n10117) );
  AND2_X1 U12608 ( .A1(n10116), .A2(n10117), .ZN(n11722) );
  INV_X1 U12609 ( .A(n11722), .ZN(n10115) );
  INV_X1 U12610 ( .A(n10116), .ZN(n10119) );
  INV_X1 U12611 ( .A(n10117), .ZN(n10118) );
  NAND2_X1 U12612 ( .A1(n10119), .A2(n10118), .ZN(n11723) );
  XNOR2_X1 U12613 ( .A(n12039), .B(n13316), .ZN(n10122) );
  NAND2_X1 U12614 ( .A1(n13441), .A2(n10861), .ZN(n10120) );
  XNOR2_X1 U12615 ( .A(n10122), .B(n10120), .ZN(n11884) );
  INV_X1 U12616 ( .A(n10120), .ZN(n10121) );
  AND2_X1 U12617 ( .A1(n10122), .A2(n10121), .ZN(n10123) );
  XNOR2_X1 U12618 ( .A(n13811), .B(n10161), .ZN(n10124) );
  NAND2_X1 U12619 ( .A1(n13440), .A2(n10861), .ZN(n10125) );
  NAND2_X1 U12620 ( .A1(n10124), .A2(n10125), .ZN(n10129) );
  INV_X1 U12621 ( .A(n10124), .ZN(n10127) );
  INV_X1 U12622 ( .A(n10125), .ZN(n10126) );
  NAND2_X1 U12623 ( .A1(n10127), .A2(n10126), .ZN(n10128) );
  AND2_X1 U12624 ( .A1(n10129), .A2(n10128), .ZN(n12016) );
  NAND2_X1 U12625 ( .A1(n12015), .A2(n12016), .ZN(n12014) );
  NAND2_X1 U12626 ( .A1(n12014), .A2(n10129), .ZN(n10132) );
  XNOR2_X1 U12627 ( .A(n13805), .B(n13316), .ZN(n10130) );
  AND2_X1 U12628 ( .A1(n13439), .A2(n10861), .ZN(n13416) );
  INV_X1 U12629 ( .A(n10130), .ZN(n10131) );
  OR2_X1 U12630 ( .A1(n10132), .A2(n10131), .ZN(n10133) );
  XNOR2_X1 U12631 ( .A(n13798), .B(n10161), .ZN(n10134) );
  NAND2_X1 U12632 ( .A1(n13438), .A2(n10861), .ZN(n10135) );
  NAND2_X1 U12633 ( .A1(n10134), .A2(n10135), .ZN(n10139) );
  INV_X1 U12634 ( .A(n10134), .ZN(n10137) );
  INV_X1 U12635 ( .A(n10135), .ZN(n10136) );
  NAND2_X1 U12636 ( .A1(n10137), .A2(n10136), .ZN(n10138) );
  NAND2_X1 U12637 ( .A1(n10139), .A2(n10138), .ZN(n13345) );
  XNOR2_X1 U12638 ( .A(n12201), .B(n10161), .ZN(n10140) );
  NAND2_X1 U12639 ( .A1(n13437), .A2(n10861), .ZN(n10141) );
  NAND2_X1 U12640 ( .A1(n10140), .A2(n10141), .ZN(n10145) );
  INV_X1 U12641 ( .A(n10140), .ZN(n10143) );
  INV_X1 U12642 ( .A(n10141), .ZN(n10142) );
  NAND2_X1 U12643 ( .A1(n10143), .A2(n10142), .ZN(n10144) );
  AND2_X1 U12644 ( .A1(n10145), .A2(n10144), .ZN(n13355) );
  XNOR2_X1 U12645 ( .A(n13787), .B(n10161), .ZN(n10147) );
  NAND2_X1 U12646 ( .A1(n13436), .A2(n10861), .ZN(n10148) );
  XNOR2_X1 U12647 ( .A(n10147), .B(n10148), .ZN(n13395) );
  INV_X1 U12648 ( .A(n10147), .ZN(n10150) );
  INV_X1 U12649 ( .A(n10148), .ZN(n10149) );
  NAND2_X1 U12650 ( .A1(n10150), .A2(n10149), .ZN(n10151) );
  XNOR2_X1 U12651 ( .A(n13782), .B(n13316), .ZN(n13302) );
  AND2_X1 U12652 ( .A1(n13435), .A2(n10861), .ZN(n13303) );
  NAND2_X1 U12653 ( .A1(n13372), .A2(n13303), .ZN(n10153) );
  XNOR2_X1 U12654 ( .A(n13777), .B(n10161), .ZN(n10155) );
  NAND2_X1 U12655 ( .A1(n13434), .A2(n10861), .ZN(n10154) );
  XNOR2_X1 U12656 ( .A(n10155), .B(n10154), .ZN(n13377) );
  NAND2_X1 U12657 ( .A1(n10155), .A2(n10154), .ZN(n10156) );
  XNOR2_X1 U12658 ( .A(n13772), .B(n13316), .ZN(n10159) );
  NAND2_X1 U12659 ( .A1(n13433), .A2(n10861), .ZN(n10157) );
  XNOR2_X1 U12660 ( .A(n10159), .B(n10157), .ZN(n13326) );
  INV_X1 U12661 ( .A(n10157), .ZN(n10158) );
  NAND2_X1 U12662 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  XNOR2_X1 U12663 ( .A(n13765), .B(n10161), .ZN(n10162) );
  NAND2_X1 U12664 ( .A1(n13432), .A2(n10861), .ZN(n13385) );
  INV_X1 U12665 ( .A(n10162), .ZN(n10163) );
  NOR2_X1 U12666 ( .A1(n10164), .A2(n10163), .ZN(n10165) );
  AOI21_X1 U12667 ( .B1(n13386), .B2(n13385), .A(n10165), .ZN(n10167) );
  XNOR2_X1 U12668 ( .A(n13759), .B(n13316), .ZN(n10166) );
  AND2_X1 U12669 ( .A1(n10167), .A2(n10166), .ZN(n10168) );
  XNOR2_X1 U12670 ( .A(n13752), .B(n13316), .ZN(n13332) );
  AND2_X1 U12671 ( .A1(n13584), .A2(n10861), .ZN(n10169) );
  NAND2_X1 U12672 ( .A1(n13332), .A2(n10169), .ZN(n10170) );
  OAI21_X1 U12673 ( .B1(n13332), .B2(n10169), .A(n10170), .ZN(n13365) );
  INV_X1 U12674 ( .A(n10170), .ZN(n10175) );
  XNOR2_X1 U12675 ( .A(n13747), .B(n13316), .ZN(n10171) );
  AND2_X1 U12676 ( .A1(n13605), .A2(n10861), .ZN(n10172) );
  NAND2_X1 U12677 ( .A1(n10171), .A2(n10172), .ZN(n10176) );
  INV_X1 U12678 ( .A(n10171), .ZN(n13409) );
  INV_X1 U12679 ( .A(n10172), .ZN(n10173) );
  NAND2_X1 U12680 ( .A1(n13409), .A2(n10173), .ZN(n10174) );
  AND2_X1 U12681 ( .A1(n10176), .A2(n10174), .ZN(n13331) );
  XNOR2_X1 U12682 ( .A(n13742), .B(n13316), .ZN(n10179) );
  NAND2_X1 U12683 ( .A1(n13583), .A2(n10861), .ZN(n10177) );
  XNOR2_X1 U12684 ( .A(n10179), .B(n10177), .ZN(n13410) );
  INV_X1 U12685 ( .A(n10177), .ZN(n10178) );
  XNOR2_X1 U12686 ( .A(n13734), .B(n13316), .ZN(n10182) );
  AND2_X1 U12687 ( .A1(n13575), .A2(n10861), .ZN(n10181) );
  NAND2_X1 U12688 ( .A1(n10182), .A2(n10181), .ZN(n13312) );
  OAI21_X1 U12689 ( .B1(n10182), .B2(n10181), .A(n13312), .ZN(n10183) );
  OR2_X1 U12690 ( .A1(n15310), .A2(n15313), .ZN(n10196) );
  INV_X1 U12691 ( .A(n10360), .ZN(n10185) );
  NAND2_X1 U12692 ( .A1(n15342), .A2(n10185), .ZN(n10186) );
  INV_X1 U12693 ( .A(n13734), .ZN(n13558) );
  NAND2_X1 U12694 ( .A1(n10696), .A2(n10189), .ZN(n10263) );
  OR2_X1 U12695 ( .A1(n10192), .A2(n10263), .ZN(n10190) );
  INV_X1 U12696 ( .A(n13604), .ZN(n13663) );
  NOR2_X2 U12697 ( .A1(n13397), .A2(n13663), .ZN(n13422) );
  AOI22_X1 U12698 ( .A1(n13422), .A2(n13551), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10200) );
  INV_X1 U12699 ( .A(n10193), .ZN(n13556) );
  OAI21_X1 U12700 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10198) );
  NAND2_X1 U12701 ( .A1(n10198), .A2(n10197), .ZN(n10487) );
  INV_X1 U12702 ( .A(n13406), .ZN(n13424) );
  AOI22_X1 U12703 ( .A1(n13556), .A2(n13424), .B1(n13421), .B2(n13583), .ZN(
        n10199) );
  OAI211_X1 U12704 ( .C1(n13558), .C2(n13369), .A(n10200), .B(n10199), .ZN(
        n10201) );
  OAI21_X1 U12705 ( .B1(n13314), .B2(n10203), .A(n10202), .ZN(P2_U3186) );
  INV_X1 U12706 ( .A(n10207), .ZN(n10212) );
  NAND2_X1 U12707 ( .A1(n11511), .A2(n14262), .ZN(n10214) );
  NAND2_X1 U12708 ( .A1(n10212), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10213) );
  OAI211_X1 U12709 ( .C1(n12353), .C2(n14256), .A(n10214), .B(n10213), .ZN(
        n10613) );
  INV_X1 U12710 ( .A(n10613), .ZN(n10215) );
  NAND2_X1 U12711 ( .A1(n10612), .A2(n10216), .ZN(n10688) );
  NOR2_X1 U12712 ( .A1(n10219), .A2(n10218), .ZN(n10221) );
  NOR2_X1 U12713 ( .A1(n10221), .A2(n10220), .ZN(n10689) );
  NAND2_X1 U12714 ( .A1(n10688), .A2(n10689), .ZN(n10687) );
  INV_X1 U12715 ( .A(n10221), .ZN(n10222) );
  NAND2_X1 U12716 ( .A1(n10687), .A2(n10222), .ZN(n10732) );
  INV_X1 U12717 ( .A(n14267), .ZN(n11106) );
  OAI22_X1 U12718 ( .A1(n10229), .A2(n11106), .B1(n15135), .B2(n12363), .ZN(
        n10225) );
  OAI22_X1 U12719 ( .A1(n15135), .A2(n12353), .B1(n12363), .B2(n11106), .ZN(
        n10224) );
  XNOR2_X1 U12720 ( .A(n10224), .B(n10223), .ZN(n10226) );
  XOR2_X1 U12721 ( .A(n10225), .B(n10226), .Z(n10733) );
  AOI22_X1 U12722 ( .A1(n10208), .A2(n11150), .B1(n12404), .B2(n13965), .ZN(
        n10228) );
  XNOR2_X1 U12723 ( .A(n10228), .B(n10223), .ZN(n10230) );
  INV_X2 U12724 ( .A(n10229), .ZN(n12408) );
  AOI22_X1 U12725 ( .A1(n12408), .A2(n13965), .B1(n12404), .B2(n11150), .ZN(
        n10231) );
  XNOR2_X1 U12726 ( .A(n10230), .B(n10231), .ZN(n11112) );
  INV_X1 U12727 ( .A(n10230), .ZN(n10233) );
  INV_X1 U12728 ( .A(n10231), .ZN(n10232) );
  OAI22_X1 U12729 ( .A1(n10229), .A2(n11145), .B1(n15149), .B2(n12363), .ZN(
        n11507) );
  XNOR2_X1 U12730 ( .A(n11506), .B(n11507), .ZN(n11510) );
  OAI22_X1 U12731 ( .A1(n15149), .A2(n12353), .B1(n12363), .B2(n11145), .ZN(
        n10234) );
  XNOR2_X1 U12732 ( .A(n10234), .B(n10223), .ZN(n11509) );
  XNOR2_X1 U12733 ( .A(n11510), .B(n11509), .ZN(n10238) );
  NAND2_X1 U12734 ( .A1(n11064), .A2(n10235), .ZN(n10243) );
  NAND3_X1 U12735 ( .A1(n11067), .A2(n10236), .A3(n15185), .ZN(n10237) );
  NOR2_X1 U12736 ( .A1(n10238), .A2(n14916), .ZN(n10248) );
  NAND2_X1 U12737 ( .A1(n10243), .A2(n10239), .ZN(n10609) );
  NAND3_X1 U12738 ( .A1(n10609), .A2(n10240), .A3(n10207), .ZN(n10241) );
  NAND2_X1 U12739 ( .A1(n10241), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10242) );
  NOR2_X1 U12740 ( .A1(n14964), .A2(n11172), .ZN(n10247) );
  AND2_X1 U12741 ( .A1(n10609), .A2(n11067), .ZN(n14926) );
  AND2_X1 U12742 ( .A1(n14921), .A2(n11174), .ZN(n10246) );
  INV_X1 U12743 ( .A(n14910), .ZN(n14956) );
  NAND2_X1 U12744 ( .A1(n14956), .A2(n13965), .ZN(n10244) );
  NAND2_X1 U12745 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13982) );
  OAI211_X1 U12746 ( .C1(n11513), .C2(n14909), .A(n10244), .B(n13982), .ZN(
        n10245) );
  OR4_X1 U12747 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        P1_U3230) );
  OAI21_X1 U12748 ( .B1(n10251), .B2(n10250), .A(n10249), .ZN(n10252) );
  NAND2_X1 U12749 ( .A1(n10252), .A2(n13705), .ZN(n10256) );
  INV_X1 U12750 ( .A(n10061), .ZN(n13611) );
  NAND2_X1 U12751 ( .A1(n15324), .A2(n13611), .ZN(n10255) );
  AOI22_X1 U12752 ( .A1(n13607), .A2(n10062), .B1(n8479), .B2(n13604), .ZN(
        n10254) );
  NAND3_X1 U12753 ( .A1(n10256), .A2(n10255), .A3(n10254), .ZN(n15322) );
  INV_X1 U12754 ( .A(n10257), .ZN(n10259) );
  INV_X1 U12755 ( .A(n15313), .ZN(n10258) );
  NAND3_X1 U12756 ( .A1(n10259), .A2(n10258), .A3(n15310), .ZN(n10260) );
  MUX2_X1 U12757 ( .A(n15322), .B(P2_REG2_REG_2__SCAN_IN), .S(n15301), .Z(
        n10267) );
  NAND2_X1 U12758 ( .A1(n7709), .A2(n10911), .ZN(n10851) );
  INV_X1 U12759 ( .A(n15324), .ZN(n10261) );
  NOR2_X1 U12760 ( .A1(n13618), .A2(n10261), .ZN(n10266) );
  OAI211_X1 U12761 ( .C1(n10280), .C2(n8476), .A(n10146), .B(n10767), .ZN(
        n15321) );
  NOR2_X1 U12762 ( .A1(n13519), .A2(n15321), .ZN(n10265) );
  OR2_X2 U12763 ( .A1(n15301), .A2(n10263), .ZN(n15292) );
  OAI22_X1 U12764 ( .A1(n15292), .A2(n8476), .B1(n13683), .B2(n10676), .ZN(
        n10264) );
  OR4_X1 U12765 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        P2_U3263) );
  NAND2_X1 U12766 ( .A1(n6663), .A2(n10268), .ZN(n10269) );
  NAND2_X1 U12767 ( .A1(n10270), .A2(n10269), .ZN(n10274) );
  NAND2_X1 U12768 ( .A1(n8473), .A2(n13607), .ZN(n10272) );
  NAND2_X1 U12769 ( .A1(n8475), .A2(n13604), .ZN(n10271) );
  NAND2_X1 U12770 ( .A1(n10272), .A2(n10271), .ZN(n10273) );
  AOI21_X1 U12771 ( .B1(n10274), .B2(n13705), .A(n10273), .ZN(n10278) );
  XNOR2_X1 U12772 ( .A(n6663), .B(n10275), .ZN(n10282) );
  INV_X1 U12773 ( .A(n10282), .ZN(n15319) );
  NAND2_X1 U12774 ( .A1(n15319), .A2(n13611), .ZN(n10277) );
  NAND2_X1 U12775 ( .A1(n10278), .A2(n10277), .ZN(n15317) );
  MUX2_X1 U12776 ( .A(n15317), .B(P2_REG2_REG_1__SCAN_IN), .S(n15290), .Z(
        n10285) );
  OAI22_X1 U12777 ( .A1(n15292), .A2(n15316), .B1(n10279), .B2(n13683), .ZN(
        n10284) );
  INV_X1 U12778 ( .A(n10280), .ZN(n10281) );
  OAI211_X1 U12779 ( .C1(n15316), .C2(n10655), .A(n10281), .B(n10146), .ZN(
        n15315) );
  OAI22_X1 U12780 ( .A1(n10282), .A2(n13618), .B1(n13519), .B2(n15315), .ZN(
        n10283) );
  OR3_X1 U12781 ( .A1(n10285), .A2(n10284), .A3(n10283), .ZN(P2_U3264) );
  AND2_X1 U12782 ( .A1(n7731), .A2(P3_U3151), .ZN(n13291) );
  INV_X2 U12783 ( .A(n13291), .ZN(n12306) );
  NAND2_X2 U12784 ( .A1(n10286), .A2(P3_U3151), .ZN(n12423) );
  OAI222_X1 U12785 ( .A1(P3_U3151), .A2(n10809), .B1(n12306), .B2(n10288), 
        .C1(n10287), .C2(n12423), .ZN(P3_U3295) );
  NOR2_X1 U12786 ( .A1(n10302), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14756) );
  INV_X1 U12787 ( .A(n14756), .ZN(n14395) );
  INV_X1 U12788 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10289) );
  NAND2_X1 U12789 ( .A1(n10302), .A2(P1_U3086), .ZN(n14398) );
  OAI222_X1 U12790 ( .A1(n10594), .A2(P1_U3086), .B1(n14395), .B2(n10289), 
        .C1(n14398), .C2(n10304), .ZN(P1_U3354) );
  INV_X1 U12791 ( .A(n10724), .ZN(n10291) );
  INV_X1 U12792 ( .A(n8601), .ZN(n10315) );
  INV_X1 U12793 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10290) );
  OAI222_X1 U12794 ( .A1(n10291), .A2(P1_U3086), .B1(n14398), .B2(n10315), 
        .C1(n10290), .C2(n14395), .ZN(P1_U3353) );
  OAI222_X1 U12795 ( .A1(P3_U3151), .A2(n15435), .B1(n12423), .B2(n10293), 
        .C1(n12306), .C2(n10292), .ZN(P3_U3287) );
  OAI222_X1 U12796 ( .A1(n12306), .A2(n10295), .B1(n12423), .B2(n10294), .C1(
        P3_U3151), .C2(n10828), .ZN(P3_U3294) );
  INV_X1 U12797 ( .A(n10296), .ZN(n10298) );
  INV_X1 U12798 ( .A(SI_7_), .ZN(n10297) );
  OAI222_X1 U12799 ( .A1(n12306), .A2(n10298), .B1(n12423), .B2(n10297), .C1(
        P3_U3151), .C2(n15416), .ZN(P3_U3288) );
  INV_X1 U12800 ( .A(SI_9_), .ZN(n10301) );
  INV_X1 U12801 ( .A(n10299), .ZN(n10300) );
  OAI222_X1 U12802 ( .A1(P3_U3151), .A2(n15455), .B1(n12423), .B2(n10301), 
        .C1(n12306), .C2(n10300), .ZN(P3_U3286) );
  NOR2_X1 U12803 ( .A1(n10302), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13840) );
  INV_X2 U12804 ( .A(n13840), .ZN(n13850) );
  NAND2_X1 U12805 ( .A1(n10302), .A2(P2_U3088), .ZN(n13852) );
  NOR2_X1 U12806 ( .A1(n10374), .A2(P2_U3088), .ZN(n15219) );
  AOI21_X1 U12807 ( .B1(n12008), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n15219), 
        .ZN(n10303) );
  OAI21_X1 U12808 ( .B1(n10304), .B2(n13850), .A(n10303), .ZN(P2_U3326) );
  INV_X1 U12809 ( .A(n8605), .ZN(n10310) );
  AOI22_X1 U12810 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n12008), .B1(n15251), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n10305) );
  OAI21_X1 U12811 ( .B1(n10310), .B2(n13850), .A(n10305), .ZN(P2_U3324) );
  INV_X1 U12812 ( .A(n10306), .ZN(n10307) );
  OAI222_X1 U12813 ( .A1(P3_U3151), .A2(n11470), .B1(n12423), .B2(n10308), 
        .C1(n12306), .C2(n10307), .ZN(P3_U3285) );
  INV_X1 U12814 ( .A(n10511), .ZN(n13968) );
  INV_X1 U12815 ( .A(n14398), .ZN(n14758) );
  INV_X1 U12816 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10309) );
  OAI222_X1 U12817 ( .A1(n13968), .A2(P1_U3086), .B1(n14383), .B2(n10310), 
        .C1(n10309), .C2(n14395), .ZN(P1_U3352) );
  INV_X1 U12818 ( .A(n13991), .ZN(n10313) );
  INV_X1 U12819 ( .A(n10311), .ZN(n10317) );
  INV_X1 U12820 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10312) );
  OAI222_X1 U12821 ( .A1(n10313), .A2(P1_U3086), .B1(n14383), .B2(n10317), 
        .C1(n10312), .C2(n14395), .ZN(P1_U3351) );
  INV_X1 U12822 ( .A(n8626), .ZN(n10337) );
  AOI22_X1 U12823 ( .A1(n10429), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n12008), .ZN(n10314) );
  OAI21_X1 U12824 ( .B1(n10337), .B2(n13850), .A(n10314), .ZN(P2_U3322) );
  OAI222_X1 U12825 ( .A1(n13844), .A2(n10316), .B1(n13850), .B2(n10315), .C1(
        P2_U3088), .C2(n15235), .ZN(P2_U3325) );
  OAI222_X1 U12826 ( .A1(n13844), .A2(n10318), .B1(n13850), .B2(n10317), .C1(
        P2_U3088), .C2(n10408), .ZN(P2_U3323) );
  INV_X1 U12827 ( .A(n10319), .ZN(n10320) );
  OAI222_X1 U12828 ( .A1(P3_U3151), .A2(n11658), .B1(n12423), .B2(n10321), 
        .C1(n12306), .C2(n10320), .ZN(P3_U3284) );
  INV_X1 U12829 ( .A(n10945), .ZN(n10961) );
  INV_X1 U12830 ( .A(n10322), .ZN(n10324) );
  INV_X1 U12831 ( .A(SI_2_), .ZN(n10323) );
  OAI222_X1 U12832 ( .A1(P3_U3151), .A2(n10961), .B1(n12306), .B2(n10324), 
        .C1(n10323), .C2(n12423), .ZN(P3_U3293) );
  INV_X1 U12833 ( .A(n10325), .ZN(n10327) );
  INV_X1 U12834 ( .A(SI_5_), .ZN(n10326) );
  OAI222_X1 U12835 ( .A1(P3_U3151), .A2(n7028), .B1(n12306), .B2(n10327), .C1(
        n10326), .C2(n12423), .ZN(P3_U3290) );
  INV_X1 U12836 ( .A(n10987), .ZN(n10964) );
  INV_X1 U12837 ( .A(n10328), .ZN(n10330) );
  INV_X1 U12838 ( .A(SI_3_), .ZN(n10329) );
  OAI222_X1 U12839 ( .A1(P3_U3151), .A2(n10964), .B1(n12306), .B2(n10330), 
        .C1(n10329), .C2(n12423), .ZN(P3_U3292) );
  INV_X1 U12840 ( .A(n11288), .ZN(n11264) );
  INV_X1 U12841 ( .A(n10331), .ZN(n10333) );
  INV_X1 U12842 ( .A(SI_4_), .ZN(n10332) );
  OAI222_X1 U12843 ( .A1(n11264), .A2(P3_U3151), .B1(n12306), .B2(n10333), 
        .C1(n10332), .C2(n12423), .ZN(P3_U3291) );
  OAI222_X1 U12844 ( .A1(P3_U3151), .A2(n15397), .B1(n12306), .B2(n10335), 
        .C1(n10334), .C2(n12423), .ZN(P3_U3289) );
  INV_X1 U12845 ( .A(n10531), .ZN(n10522) );
  INV_X1 U12846 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10336) );
  OAI222_X1 U12847 ( .A1(n10522), .A2(P1_U3086), .B1(n14383), .B2(n10337), 
        .C1(n10336), .C2(n14395), .ZN(P1_U3350) );
  OAI222_X1 U12848 ( .A1(P3_U3151), .A2(n11958), .B1(n12423), .B2(n10339), 
        .C1(n12306), .C2(n10338), .ZN(P3_U3283) );
  INV_X1 U12849 ( .A(n10340), .ZN(n10344) );
  INV_X1 U12850 ( .A(n10454), .ZN(n10341) );
  OAI222_X1 U12851 ( .A1(n13844), .A2(n10342), .B1(n13850), .B2(n10344), .C1(
        P2_U3088), .C2(n10341), .ZN(P2_U3321) );
  INV_X1 U12852 ( .A(n10533), .ZN(n10549) );
  OAI222_X1 U12853 ( .A1(n10549), .A2(P1_U3086), .B1(n14383), .B2(n10344), 
        .C1(n10343), .C2(n14395), .ZN(P1_U3349) );
  INV_X1 U12854 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10347) );
  INV_X1 U12855 ( .A(n10345), .ZN(n10349) );
  INV_X1 U12856 ( .A(n10565), .ZN(n10346) );
  OAI222_X1 U12857 ( .A1(n13844), .A2(n10347), .B1(n13850), .B2(n10349), .C1(
        P2_U3088), .C2(n10346), .ZN(P2_U3320) );
  INV_X1 U12858 ( .A(n10535), .ZN(n10606) );
  OAI222_X1 U12859 ( .A1(n10606), .A2(P1_U3086), .B1(n14383), .B2(n10349), 
        .C1(n10348), .C2(n14395), .ZN(P1_U3348) );
  INV_X1 U12860 ( .A(n10350), .ZN(n10354) );
  AOI22_X1 U12861 ( .A1(n14012), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n14756), .ZN(n10351) );
  OAI21_X1 U12862 ( .B1(n10354), .B2(n14383), .A(n10351), .ZN(P1_U3347) );
  INV_X1 U12863 ( .A(n13451), .ZN(P2_U3947) );
  INV_X1 U12864 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10355) );
  OAI222_X1 U12865 ( .A1(n13852), .A2(n10355), .B1(n13850), .B2(n10354), .C1(
        P2_U3088), .C2(n7103), .ZN(P2_U3319) );
  MUX2_X1 U12866 ( .A(n10357), .B(P2_REG1_REG_2__SCAN_IN), .S(n15235), .Z(
        n15233) );
  MUX2_X1 U12867 ( .A(n10356), .B(P2_REG1_REG_1__SCAN_IN), .S(n10374), .Z(
        n15218) );
  AND2_X1 U12868 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15217) );
  NAND2_X1 U12869 ( .A1(n15218), .A2(n15217), .ZN(n15216) );
  OAI21_X1 U12870 ( .B1(n10374), .B2(n10356), .A(n15216), .ZN(n15232) );
  NAND2_X1 U12871 ( .A1(n15233), .A2(n15232), .ZN(n15230) );
  OAI21_X1 U12872 ( .B1(n10357), .B2(n15235), .A(n15230), .ZN(n15246) );
  MUX2_X1 U12873 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7780), .S(n15251), .Z(
        n15245) );
  MUX2_X1 U12874 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7811), .S(n10408), .Z(
        n10406) );
  MUX2_X1 U12875 ( .A(n10358), .B(P2_REG1_REG_5__SCAN_IN), .S(n10429), .Z(
        n10420) );
  NOR2_X1 U12876 ( .A1(n6731), .A2(n10420), .ZN(n10419) );
  AOI21_X1 U12877 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n10429), .A(n10419), .ZN(
        n10368) );
  INV_X1 U12878 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10359) );
  MUX2_X1 U12879 ( .A(n10359), .B(P2_REG1_REG_6__SCAN_IN), .S(n10454), .Z(
        n10367) );
  NAND2_X1 U12880 ( .A1(n10361), .A2(n10360), .ZN(n10363) );
  NAND2_X1 U12881 ( .A1(n10363), .A2(n10362), .ZN(n10364) );
  AND2_X1 U12882 ( .A1(n10365), .A2(n10364), .ZN(n15221) );
  OR2_X1 U12883 ( .A1(n8517), .A2(P2_U3088), .ZN(n13841) );
  INV_X1 U12884 ( .A(n13841), .ZN(n10366) );
  NAND2_X1 U12885 ( .A1(n10389), .A2(n10366), .ZN(n10369) );
  INV_X1 U12886 ( .A(n12270), .ZN(n10370) );
  NOR2_X1 U12887 ( .A1(n10368), .A2(n10367), .ZN(n10450) );
  AOI211_X1 U12888 ( .C1(n10368), .C2(n10367), .A(n15271), .B(n10450), .ZN(
        n10393) );
  AND2_X1 U12889 ( .A1(n15221), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15275) );
  INV_X1 U12890 ( .A(n10369), .ZN(n10371) );
  MUX2_X1 U12891 ( .A(n10372), .B(P2_REG2_REG_2__SCAN_IN), .S(n15235), .Z(
        n15240) );
  MUX2_X1 U12892 ( .A(n10373), .B(P2_REG2_REG_1__SCAN_IN), .S(n10374), .Z(
        n15225) );
  AND2_X1 U12893 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n15226) );
  NAND2_X1 U12894 ( .A1(n15225), .A2(n15226), .ZN(n15224) );
  OAI21_X1 U12895 ( .B1(n10373), .B2(n10374), .A(n15224), .ZN(n15241) );
  NAND2_X1 U12896 ( .A1(n15240), .A2(n15241), .ZN(n15239) );
  OR2_X1 U12897 ( .A1(n15235), .A2(n10372), .ZN(n10375) );
  NAND2_X1 U12898 ( .A1(n15239), .A2(n10375), .ZN(n15254) );
  MUX2_X1 U12899 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10376), .S(n15251), .Z(
        n15253) );
  NAND2_X1 U12900 ( .A1(n15254), .A2(n15253), .ZN(n15252) );
  NAND2_X1 U12901 ( .A1(n15251), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10409) );
  NAND2_X1 U12902 ( .A1(n15252), .A2(n10409), .ZN(n10378) );
  MUX2_X1 U12903 ( .A(n10858), .B(P2_REG2_REG_4__SCAN_IN), .S(n10408), .Z(
        n10377) );
  NAND2_X1 U12904 ( .A1(n10378), .A2(n10377), .ZN(n10422) );
  NAND2_X1 U12905 ( .A1(n10415), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10421) );
  NAND2_X1 U12906 ( .A1(n10422), .A2(n10421), .ZN(n10381) );
  MUX2_X1 U12907 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10379), .S(n10429), .Z(
        n10380) );
  NAND2_X1 U12908 ( .A1(n10381), .A2(n10380), .ZN(n10425) );
  NAND2_X1 U12909 ( .A1(n10429), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10386) );
  NAND2_X1 U12910 ( .A1(n10425), .A2(n10386), .ZN(n10384) );
  MUX2_X1 U12911 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10382), .S(n10454), .Z(
        n10383) );
  NAND2_X1 U12912 ( .A1(n10384), .A2(n10383), .ZN(n10460) );
  MUX2_X1 U12913 ( .A(n10382), .B(P2_REG2_REG_6__SCAN_IN), .S(n10454), .Z(
        n10385) );
  NAND3_X1 U12914 ( .A1(n10425), .A2(n10386), .A3(n10385), .ZN(n10387) );
  NAND3_X1 U12915 ( .A1(n15277), .A2(n10460), .A3(n10387), .ZN(n10391) );
  AND2_X1 U12916 ( .A1(n8517), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10388) );
  NAND2_X1 U12917 ( .A1(n10389), .A2(n10388), .ZN(n15236) );
  AND2_X1 U12918 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10887) );
  AOI21_X1 U12919 ( .B1(n15281), .B2(n10454), .A(n10887), .ZN(n10390) );
  OAI211_X1 U12920 ( .C1(n15269), .C2(n9392), .A(n10391), .B(n10390), .ZN(
        n10392) );
  OR2_X1 U12921 ( .A1(n10393), .A2(n10392), .ZN(P2_U3220) );
  INV_X1 U12922 ( .A(n10394), .ZN(n10396) );
  OAI222_X1 U12923 ( .A1(n10638), .A2(P1_U3086), .B1(n14398), .B2(n10396), 
        .C1(n10395), .C2(n14395), .ZN(P1_U3346) );
  INV_X1 U12924 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10397) );
  INV_X1 U12925 ( .A(n10869), .ZN(n10872) );
  OAI222_X1 U12926 ( .A1(n13852), .A2(n10397), .B1(n13850), .B2(n10396), .C1(
        P2_U3088), .C2(n10872), .ZN(P2_U3318) );
  INV_X1 U12927 ( .A(n10398), .ZN(n10399) );
  NAND2_X1 U12928 ( .A1(n10399), .A2(n11067), .ZN(n15123) );
  AOI22_X1 U12929 ( .A1(n15123), .A2(n10401), .B1(n10403), .B2(n10400), .ZN(
        P1_U3445) );
  AOI22_X1 U12930 ( .A1(n15123), .A2(n10404), .B1(n10403), .B2(n10402), .ZN(
        P1_U3446) );
  INV_X1 U12931 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10418) );
  AOI211_X1 U12932 ( .C1(n10407), .C2(n10406), .A(n10405), .B(n15271), .ZN(
        n10413) );
  MUX2_X1 U12933 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10858), .S(n10408), .Z(
        n10410) );
  NAND3_X1 U12934 ( .A1(n10410), .A2(n15252), .A3(n10409), .ZN(n10411) );
  AND3_X1 U12935 ( .A1(n15277), .A2(n10422), .A3(n10411), .ZN(n10412) );
  NOR2_X1 U12936 ( .A1(n10413), .A2(n10412), .ZN(n10417) );
  NAND2_X1 U12937 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10782) );
  INV_X1 U12938 ( .A(n10782), .ZN(n10414) );
  AOI21_X1 U12939 ( .B1(n15281), .B2(n10415), .A(n10414), .ZN(n10416) );
  OAI211_X1 U12940 ( .C1(n15269), .C2(n10418), .A(n10417), .B(n10416), .ZN(
        P2_U3218) );
  AOI211_X1 U12941 ( .C1(n6731), .C2(n10420), .A(n15271), .B(n10419), .ZN(
        n10427) );
  MUX2_X1 U12942 ( .A(n10379), .B(P2_REG2_REG_5__SCAN_IN), .S(n10429), .Z(
        n10423) );
  NAND3_X1 U12943 ( .A1(n10423), .A2(n10422), .A3(n10421), .ZN(n10424) );
  AND3_X1 U12944 ( .A1(n15277), .A2(n10425), .A3(n10424), .ZN(n10426) );
  NOR2_X1 U12945 ( .A1(n10427), .A2(n10426), .ZN(n10431) );
  NAND2_X1 U12946 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10698) );
  INV_X1 U12947 ( .A(n10698), .ZN(n10428) );
  AOI21_X1 U12948 ( .B1(n15281), .B2(n10429), .A(n10428), .ZN(n10430) );
  OAI211_X1 U12949 ( .C1(n15269), .C2(n15590), .A(n10431), .B(n10430), .ZN(
        P2_U3219) );
  INV_X1 U12950 ( .A(n12828), .ZN(n12836) );
  INV_X1 U12951 ( .A(n10432), .ZN(n10433) );
  OAI222_X1 U12952 ( .A1(P3_U3151), .A2(n12836), .B1(n12423), .B2(n10434), 
        .C1(n12306), .C2(n10433), .ZN(P3_U3282) );
  NAND2_X1 U12953 ( .A1(n10436), .A2(P3_D_REG_1__SCAN_IN), .ZN(n10435) );
  OAI21_X1 U12954 ( .B1(n10792), .B2(n10436), .A(n10435), .ZN(P3_U3377) );
  INV_X1 U12955 ( .A(n10745), .ZN(n10649) );
  INV_X1 U12956 ( .A(n10437), .ZN(n10440) );
  OAI222_X1 U12957 ( .A1(n10649), .A2(P1_U3086), .B1(n14383), .B2(n10440), 
        .C1(n10438), .C2(n14395), .ZN(P1_U3345) );
  INV_X1 U12958 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10441) );
  INV_X1 U12959 ( .A(n11219), .ZN(n10439) );
  OAI222_X1 U12960 ( .A1(n13844), .A2(n10441), .B1(n13850), .B2(n10440), .C1(
        P2_U3088), .C2(n10439), .ZN(P2_U3317) );
  INV_X1 U12961 ( .A(n15271), .ZN(n15231) );
  AOI22_X1 U12962 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15231), .B1(n15277), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10446) );
  NAND2_X1 U12963 ( .A1(n15277), .A2(n10442), .ZN(n10443) );
  OAI211_X1 U12964 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15271), .A(n10443), .B(
        n15236), .ZN(n10444) );
  INV_X1 U12965 ( .A(n10444), .ZN(n10445) );
  MUX2_X1 U12966 ( .A(n10446), .B(n10445), .S(P2_IR_REG_0__SCAN_IN), .Z(n10449) );
  NOR2_X1 U12967 ( .A1(n10660), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10447) );
  AOI21_X1 U12968 ( .B1(n15275), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n10447), .ZN(
        n10448) );
  NAND2_X1 U12969 ( .A1(n10449), .A2(n10448), .ZN(P2_U3214) );
  AOI21_X1 U12970 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n10454), .A(n10450), .ZN(
        n10453) );
  INV_X1 U12971 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10451) );
  MUX2_X1 U12972 ( .A(n10451), .B(P2_REG1_REG_7__SCAN_IN), .S(n10565), .Z(
        n10452) );
  NOR2_X1 U12973 ( .A1(n10453), .A2(n10452), .ZN(n10562) );
  AOI211_X1 U12974 ( .C1(n10453), .C2(n10452), .A(n15271), .B(n10562), .ZN(
        n10465) );
  NAND2_X1 U12975 ( .A1(n10454), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10459) );
  NAND2_X1 U12976 ( .A1(n10460), .A2(n10459), .ZN(n10457) );
  MUX2_X1 U12977 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10455), .S(n10565), .Z(
        n10456) );
  NAND2_X1 U12978 ( .A1(n10457), .A2(n10456), .ZN(n10571) );
  MUX2_X1 U12979 ( .A(n10455), .B(P2_REG2_REG_7__SCAN_IN), .S(n10565), .Z(
        n10458) );
  NAND3_X1 U12980 ( .A1(n10460), .A2(n10459), .A3(n10458), .ZN(n10461) );
  NAND3_X1 U12981 ( .A1(n15277), .A2(n10571), .A3(n10461), .ZN(n10463) );
  AND2_X1 U12982 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11132) );
  AOI21_X1 U12983 ( .B1(n15281), .B2(n10565), .A(n11132), .ZN(n10462) );
  OAI211_X1 U12984 ( .C1(n15269), .C2(n9399), .A(n10463), .B(n10462), .ZN(
        n10464) );
  OR2_X1 U12985 ( .A1(n10465), .A2(n10464), .ZN(P2_U3221) );
  INV_X1 U12986 ( .A(n11022), .ZN(n11016) );
  INV_X1 U12987 ( .A(n10466), .ZN(n10468) );
  OAI222_X1 U12988 ( .A1(n11016), .A2(P1_U3086), .B1(n14398), .B2(n10468), 
        .C1(n10467), .C2(n14395), .ZN(P1_U3344) );
  INV_X1 U12989 ( .A(n11396), .ZN(n11400) );
  OAI222_X1 U12990 ( .A1(n13852), .A2(n10469), .B1(n13850), .B2(n10468), .C1(
        P2_U3088), .C2(n11400), .ZN(P2_U3316) );
  NAND2_X1 U12991 ( .A1(n7253), .A2(n10471), .ZN(n10470) );
  OAI21_X1 U12992 ( .B1(n10471), .B2(n7213), .A(n10470), .ZN(P3_U3376) );
  AND2_X1 U12993 ( .A1(n10481), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12994 ( .A1(n10481), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12995 ( .A1(n10481), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12996 ( .A1(n10481), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12997 ( .A1(n10481), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12998 ( .A1(n10481), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12999 ( .A1(n10481), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13000 ( .A1(n10481), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13001 ( .A1(n10481), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U13002 ( .A1(n10481), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13003 ( .A1(n10481), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13004 ( .A1(n10481), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13005 ( .A1(n10481), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U13006 ( .A1(n10481), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U13007 ( .A1(n10481), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13008 ( .A1(n10481), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13009 ( .A1(n10481), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13010 ( .A1(n10481), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U13011 ( .A1(n10481), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U13012 ( .A1(n10481), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U13013 ( .A1(n10481), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U13014 ( .A1(n10481), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13015 ( .A1(n10481), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13016 ( .A1(n10481), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13017 ( .A1(n10481), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  INV_X1 U13018 ( .A(n12898), .ZN(n12884) );
  INV_X1 U13019 ( .A(n10473), .ZN(n10475) );
  OAI222_X1 U13020 ( .A1(n12884), .A2(P3_U3151), .B1(n12306), .B2(n10475), 
        .C1(n10474), .C2(n12423), .ZN(P3_U3280) );
  INV_X1 U13021 ( .A(n11067), .ZN(n10476) );
  NAND2_X1 U13022 ( .A1(n10476), .A2(n12011), .ZN(n10497) );
  AOI21_X1 U13023 ( .B1(n10479), .B2(n10478), .A(n10477), .ZN(n10496) );
  INV_X1 U13024 ( .A(n10496), .ZN(n10480) );
  AND2_X1 U13025 ( .A1(n10497), .A2(n10480), .ZN(n15031) );
  CLKBUF_X2 U13026 ( .A(P1_U4016), .Z(n13967) );
  NOR2_X1 U13027 ( .A1(n15031), .A2(n13967), .ZN(P1_U3085) );
  INV_X1 U13028 ( .A(n10481), .ZN(n10483) );
  NOR2_X1 U13029 ( .A1(n10483), .A2(n14608), .ZN(P3_U3257) );
  NOR2_X1 U13030 ( .A1(n10483), .A2(n14585), .ZN(P3_U3251) );
  NOR2_X1 U13031 ( .A1(n10483), .A2(n10482), .ZN(P3_U3246) );
  INV_X1 U13032 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n14658) );
  NOR2_X1 U13033 ( .A1(n10483), .A2(n14658), .ZN(P3_U3248) );
  NOR2_X1 U13034 ( .A1(n10483), .A2(n14694), .ZN(P3_U3262) );
  INV_X1 U13035 ( .A(n10681), .ZN(n10484) );
  AOI21_X1 U13036 ( .B1(n10486), .B2(n10485), .A(n10484), .ZN(n10492) );
  NOR2_X1 U13037 ( .A1(n10487), .A2(P2_U3088), .ZN(n10677) );
  INV_X1 U13038 ( .A(n10677), .ZN(n10488) );
  AOI22_X1 U13039 ( .A1(n10488), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n13421), 
        .B2(n8473), .ZN(n10491) );
  AOI22_X1 U13040 ( .A1(n13422), .A2(n8475), .B1(n10489), .B2(n13425), .ZN(
        n10490) );
  OAI211_X1 U13041 ( .C1(n10492), .C2(n13417), .A(n10491), .B(n10490), .ZN(
        P2_U3194) );
  INV_X1 U13042 ( .A(n12912), .ZN(n12889) );
  INV_X1 U13043 ( .A(n10493), .ZN(n10495) );
  OAI222_X1 U13044 ( .A1(n12889), .A2(P3_U3151), .B1(n12306), .B2(n10495), 
        .C1(n10494), .C2(n12423), .ZN(P3_U3279) );
  NAND2_X1 U13045 ( .A1(n10497), .A2(n10496), .ZN(n15029) );
  INV_X1 U13046 ( .A(n15026), .ZN(n10508) );
  INV_X1 U13047 ( .A(n12065), .ZN(n15059) );
  INV_X1 U13048 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15204) );
  MUX2_X1 U13049 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n15204), .S(n10724), .Z(
        n10723) );
  INV_X1 U13050 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15202) );
  MUX2_X1 U13051 ( .A(n15202), .B(P1_REG1_REG_1__SCAN_IN), .S(n10594), .Z(
        n10580) );
  NAND2_X1 U13052 ( .A1(n6664), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10584) );
  INV_X1 U13053 ( .A(n10584), .ZN(n10498) );
  NAND2_X1 U13054 ( .A1(n10580), .A2(n10498), .ZN(n10581) );
  NAND2_X1 U13055 ( .A1(n10499), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10500) );
  NAND2_X1 U13056 ( .A1(n10581), .A2(n10500), .ZN(n10722) );
  NAND2_X1 U13057 ( .A1(n10723), .A2(n10722), .ZN(n10721) );
  NAND2_X1 U13058 ( .A1(n10724), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10501) );
  NAND2_X1 U13059 ( .A1(n10721), .A2(n10501), .ZN(n13972) );
  INV_X1 U13060 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10502) );
  XNOR2_X1 U13061 ( .A(n10511), .B(n10502), .ZN(n13973) );
  NAND2_X1 U13062 ( .A1(n13972), .A2(n13973), .ZN(n13971) );
  NAND2_X1 U13063 ( .A1(n10511), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10503) );
  NAND2_X1 U13064 ( .A1(n13971), .A2(n10503), .ZN(n13994) );
  INV_X1 U13065 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10504) );
  XNOR2_X1 U13066 ( .A(n13991), .B(n10504), .ZN(n13995) );
  AND2_X1 U13067 ( .A1(n13994), .A2(n13995), .ZN(n13992) );
  INV_X1 U13068 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10505) );
  MUX2_X1 U13069 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10505), .S(n10531), .Z(
        n10506) );
  NAND2_X1 U13070 ( .A1(n10507), .A2(n10506), .ZN(n10530) );
  OAI21_X1 U13071 ( .B1(n10507), .B2(n10506), .A(n10530), .ZN(n10517) );
  NAND2_X1 U13072 ( .A1(n10715), .A2(n10508), .ZN(n10509) );
  INV_X1 U13073 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11198) );
  MUX2_X1 U13074 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n11198), .S(n10724), .Z(
        n10720) );
  INV_X1 U13075 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10586) );
  MUX2_X1 U13076 ( .A(n10586), .B(P1_REG2_REG_1__SCAN_IN), .S(n10594), .Z(
        n10510) );
  AND2_X1 U13077 ( .A1(n6664), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13078 ( .A1(n10510), .A2(n10585), .ZN(n10587) );
  OAI21_X1 U13079 ( .B1(n10586), .B2(n10594), .A(n10587), .ZN(n10719) );
  NAND2_X1 U13080 ( .A1(n10720), .A2(n10719), .ZN(n13976) );
  NAND2_X1 U13081 ( .A1(n10724), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13975) );
  INV_X1 U13082 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10512) );
  MUX2_X1 U13083 ( .A(n10512), .B(P1_REG2_REG_3__SCAN_IN), .S(n10511), .Z(
        n13974) );
  AOI21_X1 U13084 ( .B1(n13976), .B2(n13975), .A(n13974), .ZN(n13986) );
  NOR2_X1 U13085 ( .A1(n13968), .A2(n10512), .ZN(n13985) );
  MUX2_X1 U13086 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11178), .S(n13991), .Z(
        n13984) );
  OAI21_X1 U13087 ( .B1(n13986), .B2(n13985), .A(n13984), .ZN(n13983) );
  NAND2_X1 U13088 ( .A1(n13991), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10514) );
  INV_X1 U13089 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10521) );
  MUX2_X1 U13090 ( .A(n10521), .B(P1_REG2_REG_5__SCAN_IN), .S(n10531), .Z(
        n10513) );
  AOI21_X1 U13091 ( .B1(n13983), .B2(n10514), .A(n10513), .ZN(n10552) );
  AND3_X1 U13092 ( .A1(n13983), .A2(n10514), .A3(n10513), .ZN(n10515) );
  NOR3_X1 U13093 ( .A1(n15056), .A2(n10552), .A3(n10515), .ZN(n10516) );
  AOI21_X1 U13094 ( .B1(n15059), .B2(n10517), .A(n10516), .ZN(n10520) );
  AND2_X1 U13095 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10518) );
  AOI21_X1 U13096 ( .B1(n15031), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10518), .ZN(
        n10519) );
  OAI211_X1 U13097 ( .C1(n10522), .C2(n15054), .A(n10520), .B(n10519), .ZN(
        P1_U3248) );
  NOR2_X1 U13098 ( .A1(n10522), .A2(n10521), .ZN(n10551) );
  INV_X1 U13099 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11075) );
  MUX2_X1 U13100 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11075), .S(n10533), .Z(
        n10550) );
  OAI21_X1 U13101 ( .B1(n10552), .B2(n10551), .A(n10550), .ZN(n10601) );
  NAND2_X1 U13102 ( .A1(n10533), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10600) );
  INV_X1 U13103 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10523) );
  MUX2_X1 U13104 ( .A(n10523), .B(P1_REG2_REG_7__SCAN_IN), .S(n10535), .Z(
        n10599) );
  AOI21_X1 U13105 ( .B1(n10601), .B2(n10600), .A(n10599), .ZN(n10598) );
  NOR2_X1 U13106 ( .A1(n10606), .A2(n10523), .ZN(n14006) );
  INV_X1 U13107 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10524) );
  MUX2_X1 U13108 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10524), .S(n14012), .Z(
        n10525) );
  OAI21_X1 U13109 ( .B1(n10598), .B2(n14006), .A(n10525), .ZN(n14011) );
  NAND2_X1 U13110 ( .A1(n14012), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10527) );
  INV_X1 U13111 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10637) );
  MUX2_X1 U13112 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10637), .S(n10638), .Z(
        n10526) );
  AOI21_X1 U13113 ( .B1(n14011), .B2(n10527), .A(n10526), .ZN(n10644) );
  NAND3_X1 U13114 ( .A1(n14011), .A2(n10527), .A3(n10526), .ZN(n10528) );
  NAND2_X1 U13115 ( .A1(n15044), .A2(n10528), .ZN(n10544) );
  INV_X1 U13116 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10529) );
  MUX2_X1 U13117 ( .A(n10529), .B(P1_REG1_REG_9__SCAN_IN), .S(n10638), .Z(
        n10538) );
  OAI21_X1 U13118 ( .B1(n10531), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10530), .ZN(
        n10546) );
  INV_X1 U13119 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10532) );
  MUX2_X1 U13120 ( .A(n10532), .B(P1_REG1_REG_6__SCAN_IN), .S(n10533), .Z(
        n10547) );
  NOR2_X1 U13121 ( .A1(n10546), .A2(n10547), .ZN(n10545) );
  INV_X1 U13122 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10534) );
  MUX2_X1 U13123 ( .A(n10534), .B(P1_REG1_REG_7__SCAN_IN), .S(n10535), .Z(
        n10596) );
  NOR2_X1 U13124 ( .A1(n10597), .A2(n10596), .ZN(n10595) );
  INV_X1 U13125 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10536) );
  MUX2_X1 U13126 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10536), .S(n14012), .Z(
        n14001) );
  NAND2_X1 U13127 ( .A1(n14002), .A2(n14001), .ZN(n14000) );
  OAI21_X1 U13128 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n14012), .A(n14000), .ZN(
        n10537) );
  NAND2_X1 U13129 ( .A1(n10537), .A2(n10538), .ZN(n10633) );
  OAI21_X1 U13130 ( .B1(n10538), .B2(n10537), .A(n10633), .ZN(n10539) );
  NAND2_X1 U13131 ( .A1(n10539), .A2(n15059), .ZN(n10543) );
  NOR2_X1 U13132 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8688), .ZN(n10541) );
  NOR2_X1 U13133 ( .A1(n15054), .A2(n10638), .ZN(n10540) );
  AOI211_X1 U13134 ( .C1(n15031), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10541), .B(
        n10540), .ZN(n10542) );
  OAI211_X1 U13135 ( .C1(n10644), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        P1_U3252) );
  AOI211_X1 U13136 ( .C1(n10547), .C2(n10546), .A(n10545), .B(n12065), .ZN(
        n10557) );
  NAND2_X1 U13137 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11598) );
  NAND2_X1 U13138 ( .A1(n15031), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10548) );
  OAI211_X1 U13139 ( .C1(n15054), .C2(n10549), .A(n11598), .B(n10548), .ZN(
        n10556) );
  INV_X1 U13140 ( .A(n10601), .ZN(n10554) );
  NOR3_X1 U13141 ( .A1(n10552), .A2(n10551), .A3(n10550), .ZN(n10553) );
  NOR3_X1 U13142 ( .A1(n15056), .A2(n10554), .A3(n10553), .ZN(n10555) );
  OR3_X1 U13143 ( .A1(n10557), .A2(n10556), .A3(n10555), .ZN(P1_U3249) );
  INV_X1 U13144 ( .A(n10558), .ZN(n10561) );
  INV_X1 U13145 ( .A(n11618), .ZN(n11621) );
  OAI222_X1 U13146 ( .A1(n13852), .A2(n10559), .B1(n13850), .B2(n10561), .C1(
        n11621), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U13147 ( .A(n15043), .ZN(n11017) );
  OAI222_X1 U13148 ( .A1(P1_U3086), .A2(n11017), .B1(n14383), .B2(n10561), 
        .C1(n10560), .C2(n14395), .ZN(P1_U3343) );
  MUX2_X1 U13149 ( .A(n7102), .B(P2_REG1_REG_8__SCAN_IN), .S(n10667), .Z(
        n10563) );
  AOI211_X1 U13150 ( .C1(n10564), .C2(n10563), .A(n15271), .B(n10666), .ZN(
        n10577) );
  NAND2_X1 U13151 ( .A1(n10565), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10570) );
  NAND2_X1 U13152 ( .A1(n10571), .A2(n10570), .ZN(n10568) );
  MUX2_X1 U13153 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10566), .S(n10667), .Z(
        n10567) );
  NAND2_X1 U13154 ( .A1(n10568), .A2(n10567), .ZN(n10662) );
  MUX2_X1 U13155 ( .A(n10566), .B(P2_REG2_REG_8__SCAN_IN), .S(n10667), .Z(
        n10569) );
  NAND3_X1 U13156 ( .A1(n10571), .A2(n10570), .A3(n10569), .ZN(n10572) );
  NAND3_X1 U13157 ( .A1(n15277), .A2(n10662), .A3(n10572), .ZN(n10575) );
  NAND2_X1 U13158 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11163) );
  INV_X1 U13159 ( .A(n11163), .ZN(n10573) );
  AOI21_X1 U13160 ( .B1(n15281), .B2(n10667), .A(n10573), .ZN(n10574) );
  OAI211_X1 U13161 ( .C1(n15269), .C2(n14783), .A(n10575), .B(n10574), .ZN(
        n10576) );
  OR2_X1 U13162 ( .A1(n10577), .A2(n10576), .ZN(P2_U3222) );
  OAI222_X1 U13163 ( .A1(P3_U3151), .A2(n14824), .B1(n12423), .B2(n10579), 
        .C1(n12306), .C2(n10578), .ZN(P3_U3278) );
  INV_X1 U13164 ( .A(n10580), .ZN(n10583) );
  INV_X1 U13165 ( .A(n10581), .ZN(n10582) );
  AOI211_X1 U13166 ( .C1(n10584), .C2(n10583), .A(n10582), .B(n12065), .ZN(
        n10591) );
  INV_X1 U13167 ( .A(n10585), .ZN(n10714) );
  MUX2_X1 U13168 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10586), .S(n10594), .Z(
        n10589) );
  INV_X1 U13169 ( .A(n10587), .ZN(n10588) );
  AOI211_X1 U13170 ( .C1(n10714), .C2(n10589), .A(n10588), .B(n15056), .ZN(
        n10590) );
  NOR2_X1 U13171 ( .A1(n10591), .A2(n10590), .ZN(n10593) );
  AOI22_X1 U13172 ( .A1(n15031), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10592) );
  OAI211_X1 U13173 ( .C1(n10594), .C2(n15054), .A(n10593), .B(n10592), .ZN(
        P1_U3244) );
  AOI211_X1 U13174 ( .C1(n10597), .C2(n10596), .A(n12065), .B(n10595), .ZN(
        n10608) );
  INV_X1 U13175 ( .A(n10598), .ZN(n14009) );
  NAND3_X1 U13176 ( .A1(n10601), .A2(n10600), .A3(n10599), .ZN(n10602) );
  NAND3_X1 U13177 ( .A1(n15044), .A2(n14009), .A3(n10602), .ZN(n10605) );
  NOR2_X1 U13178 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8658), .ZN(n10603) );
  AOI21_X1 U13179 ( .B1(n15031), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10603), .ZN(
        n10604) );
  OAI211_X1 U13180 ( .C1(n15054), .C2(n10606), .A(n10605), .B(n10604), .ZN(
        n10607) );
  OR2_X1 U13181 ( .A1(n10608), .A2(n10607), .ZN(P1_U3250) );
  INV_X1 U13182 ( .A(n10609), .ZN(n10611) );
  NOR2_X1 U13183 ( .A1(n10611), .A2(n10610), .ZN(n10735) );
  INV_X1 U13184 ( .A(n10735), .ZN(n10691) );
  OAI21_X1 U13185 ( .B1(n10614), .B2(n10613), .A(n10612), .ZN(n10713) );
  AOI22_X1 U13186 ( .A1(n10691), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n10713), 
        .B2(n14960), .ZN(n10616) );
  NAND2_X1 U13187 ( .A1(n14921), .A2(n6858), .ZN(n10615) );
  OAI211_X1 U13188 ( .C1(n14261), .C2(n14909), .A(n10616), .B(n10615), .ZN(
        P1_U3232) );
  INV_X1 U13189 ( .A(n10617), .ZN(n10619) );
  OAI222_X1 U13190 ( .A1(P1_U3086), .A2(n11342), .B1(n14398), .B2(n10619), 
        .C1(n10618), .C2(n14395), .ZN(P1_U3342) );
  OAI222_X1 U13191 ( .A1(n13844), .A2(n10620), .B1(n13850), .B2(n10619), .C1(
        n11629), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U13192 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10624) );
  OAI21_X1 U13193 ( .B1(n15198), .B2(n15098), .A(n11121), .ZN(n10622) );
  NAND2_X1 U13194 ( .A1(n14812), .A2(n13966), .ZN(n11117) );
  NAND3_X1 U13195 ( .A1(n6858), .A2(n11079), .A3(n11834), .ZN(n10621) );
  NAND3_X1 U13196 ( .A1(n10622), .A2(n11117), .A3(n10621), .ZN(n14360) );
  NAND2_X1 U13197 ( .A1(n15201), .A2(n14360), .ZN(n10623) );
  OAI21_X1 U13198 ( .B1(n15201), .B2(n10624), .A(n10623), .ZN(P1_U3459) );
  INV_X1 U13199 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15244) );
  OAI22_X1 U13200 ( .A1(n13369), .A2(n15328), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15244), .ZN(n10627) );
  OAI22_X1 U13201 ( .A1(n10625), .A2(n13389), .B1(n13390), .B2(n10838), .ZN(
        n10626) );
  AOI211_X1 U13202 ( .C1(n13424), .C2(n15244), .A(n10627), .B(n10626), .ZN(
        n10631) );
  OAI211_X1 U13203 ( .C1(n10629), .C2(n10628), .A(n10774), .B(n10187), .ZN(
        n10630) );
  NAND2_X1 U13204 ( .A1(n10631), .A2(n10630), .ZN(P2_U3190) );
  INV_X1 U13205 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10632) );
  MUX2_X1 U13206 ( .A(n10632), .B(P1_REG1_REG_10__SCAN_IN), .S(n10745), .Z(
        n10636) );
  INV_X1 U13207 ( .A(n10638), .ZN(n10634) );
  OAI21_X1 U13208 ( .B1(n10634), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10633), .ZN(
        n10635) );
  NOR2_X1 U13209 ( .A1(n10635), .A2(n10636), .ZN(n10744) );
  AOI211_X1 U13210 ( .C1(n10636), .C2(n10635), .A(n12065), .B(n10744), .ZN(
        n10651) );
  INV_X1 U13211 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11498) );
  MUX2_X1 U13212 ( .A(n11498), .B(P1_REG2_REG_10__SCAN_IN), .S(n10745), .Z(
        n10640) );
  NOR2_X1 U13213 ( .A1(n10638), .A2(n10637), .ZN(n10642) );
  INV_X1 U13214 ( .A(n10642), .ZN(n10639) );
  NAND2_X1 U13215 ( .A1(n10640), .A2(n10639), .ZN(n10643) );
  MUX2_X1 U13216 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11498), .S(n10745), .Z(
        n10641) );
  OAI21_X1 U13217 ( .B1(n10644), .B2(n10642), .A(n10641), .ZN(n10742) );
  OAI211_X1 U13218 ( .C1(n10644), .C2(n10643), .A(n10742), .B(n15044), .ZN(
        n10648) );
  NOR2_X1 U13219 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10645), .ZN(n10646) );
  AOI21_X1 U13220 ( .B1(n15031), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10646), 
        .ZN(n10647) );
  OAI211_X1 U13221 ( .C1(n15054), .C2(n10649), .A(n10648), .B(n10647), .ZN(
        n10650) );
  OR2_X1 U13222 ( .A1(n10651), .A2(n10650), .ZN(P1_U3253) );
  INV_X1 U13223 ( .A(n12944), .ZN(n12920) );
  INV_X1 U13224 ( .A(n10652), .ZN(n10653) );
  OAI222_X1 U13225 ( .A1(P3_U3151), .A2(n12920), .B1(n12423), .B2(n10654), 
        .C1(n12306), .C2(n10653), .ZN(P3_U3277) );
  NAND2_X1 U13226 ( .A1(n10187), .A2(n10861), .ZN(n13408) );
  OAI22_X1 U13227 ( .A1(n13408), .A2(n7176), .B1(n13417), .B2(n10655), .ZN(
        n10657) );
  NAND2_X1 U13228 ( .A1(n10657), .A2(n10656), .ZN(n10659) );
  AOI22_X1 U13229 ( .A1(n13422), .A2(n10062), .B1(n8474), .B2(n13425), .ZN(
        n10658) );
  OAI211_X1 U13230 ( .C1(n10677), .C2(n10660), .A(n10659), .B(n10658), .ZN(
        P2_U3204) );
  NAND2_X1 U13231 ( .A1(n10667), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10661) );
  NAND2_X1 U13232 ( .A1(n10662), .A2(n10661), .ZN(n10665) );
  MUX2_X1 U13233 ( .A(n11642), .B(P2_REG2_REG_9__SCAN_IN), .S(n10869), .Z(
        n10664) );
  OR2_X1 U13234 ( .A1(n10665), .A2(n10664), .ZN(n10874) );
  INV_X1 U13235 ( .A(n10874), .ZN(n10663) );
  AOI21_X1 U13236 ( .B1(n10665), .B2(n10664), .A(n10663), .ZN(n10675) );
  INV_X1 U13237 ( .A(n15277), .ZN(n13489) );
  MUX2_X1 U13238 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10668), .S(n10869), .Z(
        n10669) );
  OAI21_X1 U13239 ( .B1(n10670), .B2(n10669), .A(n10868), .ZN(n10671) );
  NAND2_X1 U13240 ( .A1(n10671), .A2(n15231), .ZN(n10674) );
  AND2_X1 U13241 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11252) );
  NOR2_X1 U13242 ( .A1(n15236), .A2(n10872), .ZN(n10672) );
  AOI211_X1 U13243 ( .C1(n15275), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n11252), .B(
        n10672), .ZN(n10673) );
  OAI211_X1 U13244 ( .C1(n10675), .C2(n13489), .A(n10674), .B(n10673), .ZN(
        P2_U3223) );
  OAI22_X1 U13245 ( .A1(n13390), .A2(n10778), .B1(n8476), .B2(n13369), .ZN(
        n10679) );
  OAI22_X1 U13246 ( .A1(n13389), .A2(n9247), .B1(n10677), .B2(n10676), .ZN(
        n10678) );
  NOR2_X1 U13247 ( .A1(n10679), .A2(n10678), .ZN(n10685) );
  OAI22_X1 U13248 ( .A1(n13408), .A2(n9247), .B1(n10064), .B2(n13417), .ZN(
        n10683) );
  INV_X1 U13249 ( .A(n10680), .ZN(n10682) );
  NAND3_X1 U13250 ( .A1(n10683), .A2(n10682), .A3(n10681), .ZN(n10684) );
  OAI211_X1 U13251 ( .C1(n13417), .C2(n10686), .A(n10685), .B(n10684), .ZN(
        P2_U3209) );
  OAI21_X1 U13252 ( .B1(n10689), .B2(n10688), .A(n10687), .ZN(n10690) );
  AOI22_X1 U13253 ( .A1(n10690), .A2(n14960), .B1(n14921), .B2(n14254), .ZN(
        n10693) );
  AOI22_X1 U13254 ( .A1(n10691), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n14956), 
        .B2(n14262), .ZN(n10692) );
  OAI211_X1 U13255 ( .C1(n11106), .C2(n14909), .A(n10693), .B(n10692), .ZN(
        P1_U3222) );
  INV_X1 U13256 ( .A(n10695), .ZN(n10915) );
  NAND2_X1 U13257 ( .A1(n13676), .A2(n10061), .ZN(n10694) );
  AOI22_X1 U13258 ( .A1(n10695), .A2(n10694), .B1(n13604), .B2(n10062), .ZN(
        n10909) );
  NAND2_X1 U13259 ( .A1(n8474), .A2(n10696), .ZN(n10910) );
  OAI211_X1 U13260 ( .C1(n10915), .C2(n13756), .A(n10909), .B(n10910), .ZN(
        n13816) );
  NAND2_X1 U13261 ( .A1(n13816), .A2(n15364), .ZN(n10697) );
  OAI21_X1 U13262 ( .B1(n15364), .B2(n7681), .A(n10697), .ZN(P2_U3430) );
  OAI21_X1 U13263 ( .B1(n13389), .B2(n10838), .A(n10698), .ZN(n10700) );
  OAI22_X1 U13264 ( .A1(n13390), .A2(n11130), .B1(n11100), .B2(n13369), .ZN(
        n10699) );
  AOI211_X1 U13265 ( .C1(n10844), .C2(n13424), .A(n10700), .B(n10699), .ZN(
        n10705) );
  OAI22_X1 U13266 ( .A1(n13408), .A2(n10838), .B1(n10702), .B2(n13417), .ZN(
        n10703) );
  NAND3_X1 U13267 ( .A1(n10773), .A2(n6981), .A3(n10703), .ZN(n10704) );
  OAI211_X1 U13268 ( .C1(n13417), .C2(n10706), .A(n10705), .B(n10704), .ZN(
        P2_U3199) );
  INV_X1 U13269 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n14646) );
  NAND2_X1 U13270 ( .A1(n11859), .A2(P3_U3897), .ZN(n10707) );
  OAI21_X1 U13271 ( .B1(P3_U3897), .B2(n14646), .A(n10707), .ZN(P3_U3496) );
  INV_X1 U13272 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n14569) );
  NAND2_X1 U13273 ( .A1(n12531), .A2(P3_U3897), .ZN(n10708) );
  OAI21_X1 U13274 ( .B1(P3_U3897), .B2(n14569), .A(n10708), .ZN(P3_U3507) );
  INV_X1 U13275 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n10710) );
  NAND2_X1 U13276 ( .A1(n10994), .A2(P3_U3897), .ZN(n10709) );
  OAI21_X1 U13277 ( .B1(P3_U3897), .B2(n10710), .A(n10709), .ZN(P3_U3491) );
  OAI222_X1 U13278 ( .A1(P3_U3151), .A2(n12942), .B1(n12306), .B2(n10712), 
        .C1(n10711), .C2(n12423), .ZN(P3_U3276) );
  MUX2_X1 U13279 ( .A(n10714), .B(n10713), .S(n15026), .Z(n10718) );
  OAI21_X1 U13280 ( .B1(n15026), .B2(P1_REG2_REG_0__SCAN_IN), .A(n10715), .ZN(
        n15024) );
  NAND2_X1 U13281 ( .A1(n15024), .A2(n10716), .ZN(n10717) );
  OAI211_X1 U13282 ( .C1(n10718), .C2(n6661), .A(n13967), .B(n10717), .ZN(
        n13999) );
  INV_X1 U13283 ( .A(n13999), .ZN(n10730) );
  OAI211_X1 U13284 ( .C1(n10720), .C2(n10719), .A(n15044), .B(n13976), .ZN(
        n10728) );
  OAI211_X1 U13285 ( .C1(n10723), .C2(n10722), .A(n15059), .B(n10721), .ZN(
        n10727) );
  AOI22_X1 U13286 ( .A1(n15031), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10726) );
  INV_X1 U13287 ( .A(n15054), .ZN(n15042) );
  NAND2_X1 U13288 ( .A1(n15042), .A2(n10724), .ZN(n10725) );
  NAND4_X1 U13289 ( .A1(n10728), .A2(n10727), .A3(n10726), .A4(n10725), .ZN(
        n10729) );
  OR2_X1 U13290 ( .A1(n10730), .A2(n10729), .ZN(P1_U3245) );
  OAI21_X1 U13291 ( .B1(n10733), .B2(n10732), .A(n10731), .ZN(n10734) );
  NAND2_X1 U13292 ( .A1(n10734), .A2(n14960), .ZN(n10738) );
  INV_X1 U13293 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11186) );
  OAI22_X1 U13294 ( .A1(n10735), .A2(n11186), .B1(n14261), .B2(n14910), .ZN(
        n10736) );
  AOI21_X1 U13295 ( .B1(n14954), .B2(n13965), .A(n10736), .ZN(n10737) );
  OAI211_X1 U13296 ( .C1(n15135), .C2(n14958), .A(n10738), .B(n10737), .ZN(
        P1_U3237) );
  NAND2_X1 U13297 ( .A1(n10745), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10741) );
  INV_X1 U13298 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10739) );
  MUX2_X1 U13299 ( .A(n10739), .B(P1_REG2_REG_11__SCAN_IN), .S(n11022), .Z(
        n10740) );
  AOI21_X1 U13300 ( .B1(n10742), .B2(n10741), .A(n10740), .ZN(n11021) );
  NAND3_X1 U13301 ( .A1(n10742), .A2(n10741), .A3(n10740), .ZN(n10743) );
  NAND2_X1 U13302 ( .A1(n10743), .A2(n15044), .ZN(n10753) );
  INV_X1 U13303 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11015) );
  MUX2_X1 U13304 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11015), .S(n11022), .Z(
        n10746) );
  NAND2_X1 U13305 ( .A1(n10747), .A2(n10746), .ZN(n15038) );
  OAI21_X1 U13306 ( .B1(n10747), .B2(n10746), .A(n15038), .ZN(n10748) );
  NAND2_X1 U13307 ( .A1(n10748), .A2(n15059), .ZN(n10752) );
  NAND2_X1 U13308 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14947)
         );
  INV_X1 U13309 ( .A(n14947), .ZN(n10750) );
  NOR2_X1 U13310 ( .A1(n15054), .A2(n11016), .ZN(n10749) );
  AOI211_X1 U13311 ( .C1(n15031), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10750), 
        .B(n10749), .ZN(n10751) );
  OAI211_X1 U13312 ( .C1(n11021), .C2(n10753), .A(n10752), .B(n10751), .ZN(
        P1_U3254) );
  INV_X1 U13313 ( .A(n11343), .ZN(n11927) );
  INV_X1 U13314 ( .A(n10754), .ZN(n10757) );
  OAI222_X1 U13315 ( .A1(P1_U3086), .A2(n11927), .B1(n14383), .B2(n10757), 
        .C1(n10755), .C2(n14395), .ZN(P1_U3341) );
  INV_X1 U13316 ( .A(n13467), .ZN(n10758) );
  OAI222_X1 U13317 ( .A1(P2_U3088), .A2(n10758), .B1(n13850), .B2(n10757), 
        .C1(n10756), .C2(n13844), .ZN(P2_U3313) );
  XNOR2_X1 U13318 ( .A(n10759), .B(n10762), .ZN(n15326) );
  AOI22_X1 U13319 ( .A1(n13607), .A2(n8475), .B1(n13450), .B2(n13604), .ZN(
        n10765) );
  OAI21_X1 U13320 ( .B1(n10762), .B2(n10761), .A(n10760), .ZN(n10763) );
  NAND2_X1 U13321 ( .A1(n10763), .A2(n13705), .ZN(n10764) );
  OAI211_X1 U13322 ( .C1(n15326), .C2(n10061), .A(n10765), .B(n10764), .ZN(
        n15329) );
  MUX2_X1 U13323 ( .A(n15329), .B(P2_REG2_REG_3__SCAN_IN), .S(n15301), .Z(
        n10766) );
  INV_X1 U13324 ( .A(n10766), .ZN(n10772) );
  OAI22_X1 U13325 ( .A1(n15292), .A2(n15328), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13683), .ZN(n10770) );
  AOI21_X1 U13326 ( .B1(n10767), .B2(n8480), .A(n10861), .ZN(n10768) );
  NAND2_X1 U13327 ( .A1(n10768), .A2(n10860), .ZN(n15327) );
  NOR2_X1 U13328 ( .A1(n13519), .A2(n15327), .ZN(n10769) );
  NOR2_X1 U13329 ( .A1(n10770), .A2(n10769), .ZN(n10771) );
  OAI211_X1 U13330 ( .C1(n15326), .C2(n13618), .A(n10772), .B(n10771), .ZN(
        P2_U3262) );
  OAI21_X1 U13331 ( .B1(n10774), .B2(n10775), .A(n10773), .ZN(n10786) );
  INV_X1 U13332 ( .A(n13408), .ZN(n13415) );
  INV_X1 U13333 ( .A(n10775), .ZN(n10777) );
  NAND3_X1 U13334 ( .A1(n13415), .A2(n10777), .A3(n10776), .ZN(n10779) );
  AOI21_X1 U13335 ( .B1(n10779), .B2(n13389), .A(n10778), .ZN(n10785) );
  INV_X1 U13336 ( .A(n10780), .ZN(n15336) );
  INV_X1 U13337 ( .A(n10859), .ZN(n10781) );
  AOI22_X1 U13338 ( .A1(n13424), .A2(n10781), .B1(n13422), .B2(n13449), .ZN(
        n10783) );
  OAI211_X1 U13339 ( .C1(n15336), .C2(n13369), .A(n10783), .B(n10782), .ZN(
        n10784) );
  AOI211_X1 U13340 ( .C1(n10187), .C2(n10786), .A(n10785), .B(n10784), .ZN(
        n10787) );
  INV_X1 U13341 ( .A(n10787), .ZN(P2_U3202) );
  NAND2_X1 U13342 ( .A1(n10994), .A2(n10790), .ZN(n12653) );
  AND2_X1 U13343 ( .A1(n10789), .A2(n12653), .ZN(n12632) );
  NOR3_X1 U13344 ( .A1(n12632), .A2(n11848), .A3(n12780), .ZN(n10791) );
  AOI21_X1 U13345 ( .B1(n14853), .B2(n10788), .A(n10791), .ZN(n12300) );
  NAND2_X1 U13346 ( .A1(n10792), .A2(n10793), .ZN(n10797) );
  INV_X1 U13347 ( .A(n10793), .ZN(n10794) );
  NAND2_X1 U13348 ( .A1(n11001), .A2(n10794), .ZN(n10796) );
  INV_X1 U13349 ( .A(n10920), .ZN(n10795) );
  NAND2_X1 U13350 ( .A1(n10799), .A2(n10798), .ZN(n10801) );
  INV_X1 U13351 ( .A(n12804), .ZN(n15515) );
  NOR2_X1 U13352 ( .A1(n15545), .A2(n15515), .ZN(n10800) );
  MUX2_X1 U13353 ( .A(n10827), .B(n12300), .S(n15501), .Z(n10804) );
  OR2_X1 U13354 ( .A1(n10801), .A2(n12804), .ZN(n15482) );
  AOI22_X1 U13355 ( .A1(n13148), .A2(n10802), .B1(n15517), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10803) );
  NAND2_X1 U13356 ( .A1(n10804), .A2(n10803), .ZN(P3_U3233) );
  INV_X1 U13357 ( .A(n10932), .ZN(n10805) );
  OR2_X1 U13358 ( .A1(n10918), .A2(P3_U3151), .ZN(n12812) );
  NAND2_X1 U13359 ( .A1(n10805), .A2(n12812), .ZN(n10815) );
  NAND2_X1 U13360 ( .A1(n12780), .A2(n10918), .ZN(n10806) );
  AND2_X1 U13361 ( .A1(n10807), .A2(n10806), .ZN(n10813) );
  INV_X1 U13362 ( .A(n10819), .ZN(n10808) );
  MUX2_X1 U13363 ( .A(n12816), .B(n10808), .S(n9968), .Z(n15454) );
  NAND2_X1 U13364 ( .A1(n10819), .A2(n12936), .ZN(n12949) );
  MUX2_X1 U13365 ( .A(n15572), .B(P3_REG1_REG_2__SCAN_IN), .S(n10945), .Z(
        n10812) );
  NAND2_X1 U13366 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10809), .ZN(n11091) );
  INV_X1 U13367 ( .A(n11091), .ZN(n10810) );
  OAI21_X1 U13368 ( .B1(n10828), .B2(n10810), .A(n7655), .ZN(n10897) );
  OR2_X1 U13369 ( .A1(n10897), .A2(n10898), .ZN(n10895) );
  NAND2_X1 U13370 ( .A1(n10895), .A2(n7655), .ZN(n10811) );
  NAND2_X1 U13371 ( .A1(n10811), .A2(n10812), .ZN(n10954) );
  OAI21_X1 U13372 ( .B1(n10812), .B2(n10811), .A(n10954), .ZN(n10824) );
  INV_X1 U13373 ( .A(n10813), .ZN(n10814) );
  INV_X1 U13374 ( .A(n15460), .ZN(n12892) );
  INV_X1 U13375 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10816) );
  OAI22_X1 U13376 ( .A1(n12892), .A2(n10816), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11043), .ZN(n10823) );
  INV_X1 U13377 ( .A(n10817), .ZN(n10818) );
  NOR2_X1 U13378 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10827), .ZN(n11093) );
  AND2_X1 U13379 ( .A1(n14832), .A2(n10821), .ZN(n10822) );
  AOI211_X1 U13380 ( .C1(n15463), .C2(n10824), .A(n10823), .B(n10822), .ZN(
        n10834) );
  INV_X2 U13381 ( .A(n10825), .ZN(n12913) );
  MUX2_X1 U13382 ( .A(n10826), .B(n10898), .S(n12913), .Z(n10829) );
  XNOR2_X1 U13383 ( .A(n10829), .B(n10828), .ZN(n10894) );
  INV_X1 U13384 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n12301) );
  MUX2_X1 U13385 ( .A(n10827), .B(n12301), .S(n12913), .Z(n11087) );
  AND2_X1 U13386 ( .A1(n11087), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U13387 ( .A1(n10894), .A2(n10893), .ZN(n10831) );
  INV_X1 U13388 ( .A(n10828), .ZN(n10906) );
  NAND2_X1 U13389 ( .A1(n10829), .A2(n10906), .ZN(n10830) );
  NAND2_X1 U13390 ( .A1(n10831), .A2(n10830), .ZN(n10943) );
  MUX2_X1 U13391 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12913), .Z(n10944) );
  XNOR2_X1 U13392 ( .A(n10944), .B(n10945), .ZN(n10942) );
  XNOR2_X1 U13393 ( .A(n10943), .B(n10942), .ZN(n10832) );
  NAND2_X1 U13394 ( .A1(n10832), .A2(n12954), .ZN(n10833) );
  OAI211_X1 U13395 ( .C1(n15454), .C2(n10961), .A(n10834), .B(n10833), .ZN(
        P3_U3184) );
  XNOR2_X1 U13396 ( .A(n10835), .B(n10836), .ZN(n11098) );
  XNOR2_X1 U13397 ( .A(n10837), .B(n10836), .ZN(n10840) );
  OAI22_X1 U13398 ( .A1(n10838), .A2(n13661), .B1(n11130), .B2(n13663), .ZN(
        n10839) );
  AOI21_X1 U13399 ( .B1(n10840), .B2(n13705), .A(n10839), .ZN(n10841) );
  OAI21_X1 U13400 ( .B1(n10061), .B2(n11098), .A(n10841), .ZN(n11101) );
  NAND2_X1 U13401 ( .A1(n11101), .A2(n13689), .ZN(n10850) );
  INV_X1 U13402 ( .A(n15292), .ZN(n13685) );
  INV_X1 U13403 ( .A(n11439), .ZN(n10842) );
  OAI211_X1 U13404 ( .C1(n11100), .C2(n10843), .A(n10842), .B(n10146), .ZN(
        n11099) );
  NOR2_X1 U13405 ( .A1(n13519), .A2(n11099), .ZN(n10847) );
  INV_X1 U13406 ( .A(n10844), .ZN(n10845) );
  OAI22_X1 U13407 ( .A1(n13689), .A2(n10379), .B1(n10845), .B2(n13683), .ZN(
        n10846) );
  AOI211_X1 U13408 ( .C1(n13685), .C2(n10848), .A(n10847), .B(n10846), .ZN(
        n10849) );
  OAI211_X1 U13409 ( .C1(n11098), .C2(n13618), .A(n10850), .B(n10849), .ZN(
        P2_U3260) );
  AND2_X1 U13410 ( .A1(n10061), .A2(n10851), .ZN(n10852) );
  XNOR2_X1 U13411 ( .A(n10853), .B(n10855), .ZN(n15333) );
  OAI21_X1 U13412 ( .B1(n10856), .B2(n10855), .A(n10854), .ZN(n10857) );
  AOI222_X1 U13413 ( .A1(n13705), .A2(n10857), .B1(n13449), .B2(n13604), .C1(
        n8479), .C2(n13607), .ZN(n15335) );
  INV_X1 U13414 ( .A(n15301), .ZN(n13689) );
  MUX2_X1 U13415 ( .A(n10858), .B(n15335), .S(n13689), .Z(n10866) );
  OAI22_X1 U13416 ( .A1(n15292), .A2(n15336), .B1(n13683), .B2(n10859), .ZN(
        n10864) );
  XNOR2_X1 U13417 ( .A(n15336), .B(n10860), .ZN(n10862) );
  NAND2_X1 U13418 ( .A1(n10862), .A2(n10146), .ZN(n15334) );
  NOR2_X1 U13419 ( .A1(n13519), .A2(n15334), .ZN(n10863) );
  NOR2_X1 U13420 ( .A1(n10864), .A2(n10863), .ZN(n10865) );
  OAI211_X1 U13421 ( .C1(n15293), .C2(n15333), .A(n10866), .B(n10865), .ZN(
        P2_U3261) );
  INV_X1 U13422 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10867) );
  MUX2_X1 U13423 ( .A(n10867), .B(P2_REG1_REG_10__SCAN_IN), .S(n11219), .Z(
        n10871) );
  OAI21_X1 U13424 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n10869), .A(n10868), .ZN(
        n10870) );
  AOI211_X1 U13425 ( .C1(n10871), .C2(n10870), .A(n15271), .B(n11218), .ZN(
        n10884) );
  NAND2_X1 U13426 ( .A1(n10872), .A2(n11642), .ZN(n10873) );
  NAND2_X1 U13427 ( .A1(n10874), .A2(n10873), .ZN(n10877) );
  INV_X1 U13428 ( .A(n10877), .ZN(n10879) );
  MUX2_X1 U13429 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10875), .S(n11219), .Z(
        n10878) );
  MUX2_X1 U13430 ( .A(n10875), .B(P2_REG2_REG_10__SCAN_IN), .S(n11219), .Z(
        n10876) );
  OR2_X1 U13431 ( .A1(n10877), .A2(n10876), .ZN(n11209) );
  OAI211_X1 U13432 ( .C1(n10879), .C2(n10878), .A(n15277), .B(n11209), .ZN(
        n10882) );
  AND2_X1 U13433 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10880) );
  AOI21_X1 U13434 ( .B1(n15281), .B2(n11219), .A(n10880), .ZN(n10881) );
  OAI211_X1 U13435 ( .C1(n15269), .C2(n7389), .A(n10882), .B(n10881), .ZN(
        n10883) );
  OR2_X1 U13436 ( .A1(n10884), .A2(n10883), .ZN(P2_U3224) );
  OAI22_X1 U13437 ( .A1(n13389), .A2(n10885), .B1(n11440), .B2(n13406), .ZN(
        n10886) );
  AOI211_X1 U13438 ( .C1(n13422), .C2(n13447), .A(n10887), .B(n10886), .ZN(
        n10892) );
  AOI21_X1 U13439 ( .B1(n10889), .B2(n10888), .A(n13417), .ZN(n10890) );
  NAND2_X1 U13440 ( .A1(n10890), .A2(n11126), .ZN(n10891) );
  OAI211_X1 U13441 ( .C1(n15343), .C2(n13369), .A(n10892), .B(n10891), .ZN(
        P2_U3211) );
  INV_X1 U13442 ( .A(n10893), .ZN(n11096) );
  XNOR2_X1 U13443 ( .A(n10894), .B(n11096), .ZN(n10908) );
  INV_X1 U13444 ( .A(n10895), .ZN(n10896) );
  AOI21_X1 U13445 ( .B1(n10898), .B2(n10897), .A(n10896), .ZN(n10900) );
  AOI22_X1 U13446 ( .A1(n15460), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10899) );
  OAI21_X1 U13447 ( .B1(n10900), .B2(n12949), .A(n10899), .ZN(n10905) );
  NAND2_X1 U13448 ( .A1(n10901), .A2(n10826), .ZN(n10902) );
  AOI21_X1 U13449 ( .B1(n10903), .B2(n10902), .A(n15467), .ZN(n10904) );
  AOI211_X1 U13450 ( .C1(n14825), .C2(n10906), .A(n10905), .B(n10904), .ZN(
        n10907) );
  OAI21_X1 U13451 ( .B1(n15456), .B2(n10908), .A(n10907), .ZN(P3_U3183) );
  OAI21_X1 U13452 ( .B1(n10911), .B2(n10910), .A(n10909), .ZN(n10912) );
  INV_X1 U13453 ( .A(n13683), .ZN(n15288) );
  AOI22_X1 U13454 ( .A1(n13689), .A2(n10912), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n15288), .ZN(n10914) );
  NAND2_X1 U13455 ( .A1(n15290), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10913) );
  OAI211_X1 U13456 ( .C1(n10915), .C2(n13618), .A(n10914), .B(n10913), .ZN(
        P2_U3265) );
  INV_X1 U13457 ( .A(n10916), .ZN(n10929) );
  OR2_X1 U13458 ( .A1(n10917), .A2(n10929), .ZN(n10924) );
  INV_X1 U13459 ( .A(n10918), .ZN(n10919) );
  NOR2_X1 U13460 ( .A1(n10920), .A2(n10919), .ZN(n10923) );
  OR2_X1 U13461 ( .A1(n10998), .A2(n10930), .ZN(n10921) );
  NAND4_X1 U13462 ( .A1(n10924), .A2(n10923), .A3(n10922), .A4(n10921), .ZN(
        n10925) );
  NAND2_X1 U13463 ( .A1(n10925), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10928) );
  INV_X1 U13464 ( .A(n12808), .ZN(n10926) );
  OR2_X1 U13465 ( .A1(n10998), .A2(n10926), .ZN(n10927) );
  NOR2_X1 U13466 ( .A1(n12578), .A2(P3_U3151), .ZN(n11044) );
  OR3_X1 U13467 ( .A1(n10935), .A2(n10929), .A3(n11848), .ZN(n10934) );
  INV_X1 U13468 ( .A(n10930), .ZN(n10931) );
  NAND3_X1 U13469 ( .A1(n10998), .A2(n10932), .A3(n10931), .ZN(n10933) );
  INV_X1 U13470 ( .A(n12632), .ZN(n10939) );
  OR2_X1 U13471 ( .A1(n10935), .A2(n15545), .ZN(n10936) );
  AND2_X1 U13472 ( .A1(n12808), .A2(n10995), .ZN(n10937) );
  OAI22_X1 U13473 ( .A1(n12581), .A2(n10790), .B1(n6848), .B2(n12584), .ZN(
        n10938) );
  AOI21_X1 U13474 ( .B1(n12572), .B2(n10939), .A(n10938), .ZN(n10940) );
  OAI21_X1 U13475 ( .B1(n11044), .B2(n10941), .A(n10940), .ZN(P3_U3172) );
  MUX2_X1 U13476 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12913), .Z(n11287) );
  XNOR2_X1 U13477 ( .A(n11287), .B(n11288), .ZN(n11285) );
  NAND2_X1 U13478 ( .A1(n10943), .A2(n10942), .ZN(n10948) );
  INV_X1 U13479 ( .A(n10944), .ZN(n10946) );
  NAND2_X1 U13480 ( .A1(n10946), .A2(n10945), .ZN(n10947) );
  NAND2_X1 U13481 ( .A1(n10948), .A2(n10947), .ZN(n10977) );
  MUX2_X1 U13482 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12913), .Z(n10949) );
  XNOR2_X1 U13483 ( .A(n10949), .B(n10987), .ZN(n10978) );
  NAND2_X1 U13484 ( .A1(n10977), .A2(n10978), .ZN(n10952) );
  INV_X1 U13485 ( .A(n10949), .ZN(n10950) );
  NAND2_X1 U13486 ( .A1(n10950), .A2(n10987), .ZN(n10951) );
  NAND2_X1 U13487 ( .A1(n10952), .A2(n10951), .ZN(n11286) );
  XOR2_X1 U13488 ( .A(n11285), .B(n11286), .Z(n10976) );
  NAND2_X1 U13489 ( .A1(n10961), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10953) );
  NAND2_X1 U13490 ( .A1(n10954), .A2(n10953), .ZN(n10955) );
  XNOR2_X1 U13491 ( .A(n10955), .B(n10987), .ZN(n10981) );
  MUX2_X1 U13492 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n9598), .S(n11288), .Z(
        n10957) );
  NAND2_X1 U13493 ( .A1(n10956), .A2(n10957), .ZN(n10960) );
  INV_X1 U13494 ( .A(n10957), .ZN(n10958) );
  NAND2_X1 U13495 ( .A1(n10959), .A2(n10958), .ZN(n11273) );
  AND2_X1 U13496 ( .A1(n10960), .A2(n11273), .ZN(n10973) );
  MUX2_X1 U13497 ( .A(n9601), .B(P3_REG2_REG_4__SCAN_IN), .S(n11288), .Z(
        n10968) );
  NAND2_X1 U13498 ( .A1(n10961), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U13499 ( .A1(n10963), .A2(n10962), .ZN(n10965) );
  NAND2_X1 U13500 ( .A1(n10965), .A2(n10964), .ZN(n10966) );
  OAI21_X1 U13501 ( .B1(n10968), .B2(n10967), .A(n11263), .ZN(n10969) );
  NAND2_X1 U13502 ( .A1(n14832), .A2(n10969), .ZN(n10972) );
  INV_X1 U13503 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10970) );
  NOR2_X1 U13504 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10970), .ZN(n11239) );
  AOI21_X1 U13505 ( .B1(n15460), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11239), .ZN(
        n10971) );
  OAI211_X1 U13506 ( .C1(n10973), .C2(n12949), .A(n10972), .B(n10971), .ZN(
        n10974) );
  AOI21_X1 U13507 ( .B1(n14825), .B2(n11288), .A(n10974), .ZN(n10975) );
  OAI21_X1 U13508 ( .B1(n10976), .B2(n15456), .A(n10975), .ZN(P3_U3186) );
  XOR2_X1 U13509 ( .A(n10978), .B(n10977), .Z(n10989) );
  XOR2_X1 U13510 ( .A(n11388), .B(n10979), .Z(n10985) );
  INV_X1 U13511 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11390) );
  NOR2_X1 U13512 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11390), .ZN(n11052) );
  AOI21_X1 U13513 ( .B1(n15460), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11052), .ZN(
        n10984) );
  OAI21_X1 U13514 ( .B1(n10981), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10980), .ZN(
        n10982) );
  NAND2_X1 U13515 ( .A1(n15463), .A2(n10982), .ZN(n10983) );
  OAI211_X1 U13516 ( .C1(n15467), .C2(n10985), .A(n10984), .B(n10983), .ZN(
        n10986) );
  AOI21_X1 U13517 ( .B1(n10987), .B2(n14825), .A(n10986), .ZN(n10988) );
  OAI21_X1 U13518 ( .B1(n10989), .B2(n15456), .A(n10988), .ZN(P3_U3185) );
  INV_X1 U13519 ( .A(n11928), .ZN(n15055) );
  INV_X1 U13520 ( .A(n10990), .ZN(n10992) );
  OAI222_X1 U13521 ( .A1(P1_U3086), .A2(n15055), .B1(n14383), .B2(n10992), 
        .C1(n10991), .C2(n14395), .ZN(P1_U3340) );
  OAI222_X1 U13522 ( .A1(n13844), .A2(n10993), .B1(n13850), .B2(n10992), .C1(
        n13468), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U13523 ( .A(n10995), .ZN(n10996) );
  AND2_X1 U13524 ( .A1(n12808), .A2(n10996), .ZN(n10997) );
  INV_X1 U13525 ( .A(n12826), .ZN(n15508) );
  OAI22_X1 U13526 ( .A1(n9978), .A2(n12576), .B1(n12584), .B2(n15508), .ZN(
        n10999) );
  AOI21_X1 U13527 ( .B1(n12590), .B2(n15503), .A(n10999), .ZN(n11013) );
  NAND2_X1 U13528 ( .A1(n10788), .A2(n15503), .ZN(n11000) );
  AND2_X1 U13529 ( .A1(n15489), .A2(n11000), .ZN(n11005) );
  NAND2_X1 U13530 ( .A1(n11381), .A2(n11061), .ZN(n11003) );
  AND2_X1 U13531 ( .A1(n11003), .A2(n11002), .ZN(n11004) );
  INV_X2 U13532 ( .A(n12452), .ZN(n12469) );
  NAND3_X1 U13533 ( .A1(n11008), .A2(n10789), .A3(n12469), .ZN(n11009) );
  OAI211_X1 U13534 ( .C1(n11010), .C2(n15506), .A(n11035), .B(n11009), .ZN(
        n11011) );
  NAND2_X1 U13535 ( .A1(n11011), .A2(n12572), .ZN(n11012) );
  OAI211_X1 U13536 ( .C1(n11044), .C2(n11014), .A(n11013), .B(n11012), .ZN(
        P3_U3162) );
  INV_X1 U13537 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U13538 ( .A1(n11016), .A2(n11015), .ZN(n15037) );
  MUX2_X1 U13539 ( .A(n11018), .B(P1_REG1_REG_12__SCAN_IN), .S(n15043), .Z(
        n15036) );
  AOI21_X1 U13540 ( .B1(n15038), .B2(n15037), .A(n15036), .ZN(n15035) );
  AOI21_X1 U13541 ( .B1(n11018), .B2(n11017), .A(n15035), .ZN(n11020) );
  INV_X1 U13542 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14987) );
  MUX2_X1 U13543 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n14987), .S(n11024), .Z(
        n11019) );
  NAND2_X1 U13544 ( .A1(n11020), .A2(n11019), .ZN(n11337) );
  OAI211_X1 U13545 ( .C1(n11020), .C2(n11019), .A(n11337), .B(n15059), .ZN(
        n11032) );
  AOI21_X1 U13546 ( .B1(n11022), .B2(P1_REG2_REG_11__SCAN_IN), .A(n11021), 
        .ZN(n15033) );
  INV_X1 U13547 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11023) );
  MUX2_X1 U13548 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11023), .S(n15043), .Z(
        n15034) );
  NAND2_X1 U13549 ( .A1(n15033), .A2(n15034), .ZN(n15032) );
  OAI21_X1 U13550 ( .B1(n15043), .B2(P1_REG2_REG_12__SCAN_IN), .A(n15032), 
        .ZN(n11026) );
  INV_X1 U13551 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n14803) );
  MUX2_X1 U13552 ( .A(n14803), .B(P1_REG2_REG_13__SCAN_IN), .S(n11024), .Z(
        n11025) );
  NOR2_X1 U13553 ( .A1(n11026), .A2(n11025), .ZN(n11347) );
  AOI211_X1 U13554 ( .C1(n11026), .C2(n11025), .A(n15056), .B(n11347), .ZN(
        n11030) );
  INV_X1 U13555 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n12245) );
  NOR2_X1 U13556 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12245), .ZN(n11027) );
  AOI21_X1 U13557 ( .B1(n15031), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11027), 
        .ZN(n11028) );
  OAI21_X1 U13558 ( .B1(n15054), .B2(n11342), .A(n11028), .ZN(n11029) );
  NOR2_X1 U13559 ( .A1(n11030), .A2(n11029), .ZN(n11031) );
  NAND2_X1 U13560 ( .A1(n11032), .A2(n11031), .ZN(P1_U3256) );
  XNOR2_X1 U13561 ( .A(n11045), .B(n12826), .ZN(n11037) );
  XNOR2_X1 U13562 ( .A(n11046), .B(n15503), .ZN(n11033) );
  NAND2_X1 U13563 ( .A1(n11033), .A2(n6848), .ZN(n11034) );
  NAND2_X1 U13564 ( .A1(n11035), .A2(n11034), .ZN(n11036) );
  NAND2_X1 U13565 ( .A1(n11036), .A2(n11037), .ZN(n11049) );
  OAI21_X1 U13566 ( .B1(n11037), .B2(n11036), .A(n11049), .ZN(n11038) );
  NAND2_X1 U13567 ( .A1(n11038), .A2(n12572), .ZN(n11042) );
  INV_X1 U13568 ( .A(n12825), .ZN(n15488) );
  OAI22_X1 U13569 ( .A1(n6848), .A2(n12576), .B1(n12584), .B2(n15488), .ZN(
        n11039) );
  AOI21_X1 U13570 ( .B1(n12590), .B2(n11040), .A(n11039), .ZN(n11041) );
  OAI211_X1 U13571 ( .C1(n11044), .C2(n11043), .A(n11042), .B(n11041), .ZN(
        P3_U3177) );
  NAND2_X1 U13572 ( .A1(n11045), .A2(n15508), .ZN(n11047) );
  AND2_X1 U13573 ( .A1(n11049), .A2(n11047), .ZN(n11051) );
  XNOR2_X1 U13574 ( .A(n11046), .B(n11055), .ZN(n11229) );
  XNOR2_X1 U13575 ( .A(n11229), .B(n12825), .ZN(n11050) );
  AND2_X1 U13576 ( .A1(n11050), .A2(n11047), .ZN(n11048) );
  NAND2_X1 U13577 ( .A1(n11049), .A2(n11048), .ZN(n11232) );
  OAI211_X1 U13578 ( .C1(n11051), .C2(n11050), .A(n12572), .B(n11232), .ZN(
        n11057) );
  INV_X1 U13579 ( .A(n12584), .ZN(n12574) );
  AOI21_X1 U13580 ( .B1(n12574), .B2(n12824), .A(n11052), .ZN(n11053) );
  OAI21_X1 U13581 ( .B1(n15508), .B2(n12576), .A(n11053), .ZN(n11054) );
  AOI21_X1 U13582 ( .B1(n12590), .B2(n11055), .A(n11054), .ZN(n11056) );
  OAI211_X1 U13583 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12588), .A(n11057), .B(
        n11056), .ZN(P3_U3158) );
  INV_X1 U13584 ( .A(n11058), .ZN(n11060) );
  OAI222_X1 U13585 ( .A1(P3_U3151), .A2(n11061), .B1(n12306), .B2(n11060), 
        .C1(n11059), .C2(n12423), .ZN(P3_U3275) );
  XNOR2_X1 U13586 ( .A(n11063), .B(n11062), .ZN(n15166) );
  INV_X1 U13587 ( .A(n15166), .ZN(n11086) );
  NAND2_X1 U13588 ( .A1(n11065), .A2(n11064), .ZN(n12255) );
  INV_X1 U13589 ( .A(n11068), .ZN(n11069) );
  XNOR2_X1 U13590 ( .A(n11070), .B(n11071), .ZN(n11072) );
  NAND2_X1 U13591 ( .A1(n11072), .A2(n15098), .ZN(n11073) );
  AOI22_X1 U13592 ( .A1(n14812), .A2(n13961), .B1(n14979), .B2(n13963), .ZN(
        n11599) );
  NAND2_X1 U13593 ( .A1(n11073), .A2(n11599), .ZN(n11074) );
  AOI21_X1 U13594 ( .B1(n15166), .B2(n15102), .A(n11074), .ZN(n15168) );
  MUX2_X1 U13595 ( .A(n11075), .B(n15168), .S(n14804), .Z(n11085) );
  NAND2_X1 U13596 ( .A1(n15110), .A2(n11594), .ZN(n11076) );
  NAND2_X1 U13597 ( .A1(n11076), .A2(n15111), .ZN(n11077) );
  NOR2_X1 U13598 ( .A1(n15090), .A2(n11077), .ZN(n15164) );
  INV_X1 U13599 ( .A(n11078), .ZN(n11080) );
  NAND2_X1 U13600 ( .A1(n11080), .A2(n11079), .ZN(n11081) );
  INV_X1 U13601 ( .A(n11594), .ZN(n11082) );
  OAI22_X1 U13602 ( .A1(n15107), .A2(n11082), .B1(n11597), .B2(n14801), .ZN(
        n11083) );
  AOI21_X1 U13603 ( .B1(n15113), .B2(n15164), .A(n11083), .ZN(n11084) );
  OAI211_X1 U13604 ( .C1(n11086), .C2(n11765), .A(n11085), .B(n11084), .ZN(
        P1_U3287) );
  NOR3_X1 U13605 ( .A1(n15463), .A2(n14832), .A3(n12954), .ZN(n11097) );
  INV_X1 U13606 ( .A(n11087), .ZN(n11088) );
  NAND2_X1 U13607 ( .A1(n12954), .A2(n11088), .ZN(n11089) );
  MUX2_X1 U13608 ( .A(n11089), .B(n15454), .S(P3_IR_REG_0__SCAN_IN), .Z(n11095) );
  AOI22_X1 U13609 ( .A1(n15460), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11090) );
  OAI21_X1 U13610 ( .B1(n11091), .B2(n12949), .A(n11090), .ZN(n11092) );
  AOI21_X1 U13611 ( .B1(n14832), .B2(n11093), .A(n11092), .ZN(n11094) );
  OAI211_X1 U13612 ( .C1(n11097), .C2(n11096), .A(n11095), .B(n11094), .ZN(
        P3_U3182) );
  INV_X1 U13613 ( .A(n11098), .ZN(n11103) );
  OAI21_X1 U13614 ( .B1(n11100), .B2(n15342), .A(n11099), .ZN(n11102) );
  AOI211_X1 U13615 ( .C1(n9298), .C2(n11103), .A(n11102), .B(n11101), .ZN(
        n11203) );
  NAND2_X1 U13616 ( .A1(n15371), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11105) );
  OAI21_X1 U13617 ( .B1(n11203), .B2(n15371), .A(n11105), .ZN(P2_U3504) );
  INV_X1 U13618 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14623) );
  INV_X1 U13619 ( .A(n14964), .ZN(n13939) );
  NAND2_X1 U13620 ( .A1(n14921), .A2(n11150), .ZN(n11109) );
  OAI22_X1 U13621 ( .A1(n14910), .A2(n11106), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14623), .ZN(n11107) );
  INV_X1 U13622 ( .A(n11107), .ZN(n11108) );
  OAI211_X1 U13623 ( .C1(n11145), .C2(n14909), .A(n11109), .B(n11108), .ZN(
        n11114) );
  AOI211_X1 U13624 ( .C1(n11112), .C2(n11111), .A(n14916), .B(n11110), .ZN(
        n11113) );
  AOI211_X1 U13625 ( .C1(n14623), .C2(n13939), .A(n11114), .B(n11113), .ZN(
        n11115) );
  INV_X1 U13626 ( .A(n11115), .ZN(P1_U3218) );
  INV_X1 U13627 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11116) );
  OAI22_X1 U13628 ( .A1(n15105), .A2(n11117), .B1(n11116), .B2(n14801), .ZN(
        n11119) );
  NAND2_X1 U13629 ( .A1(n15113), .A2(n15111), .ZN(n12251) );
  AOI21_X1 U13630 ( .B1(n12251), .B2(n15107), .A(n14256), .ZN(n11118) );
  AOI211_X1 U13631 ( .C1(n14251), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11119), .B(
        n11118), .ZN(n11123) );
  OR2_X1 U13632 ( .A1(n15118), .A2(n15083), .ZN(n14233) );
  INV_X1 U13633 ( .A(n14233), .ZN(n14182) );
  OAI21_X1 U13634 ( .B1(n14182), .B2(n14809), .A(n11121), .ZN(n11122) );
  NAND2_X1 U13635 ( .A1(n11123), .A2(n11122), .ZN(P1_U3293) );
  INV_X1 U13636 ( .A(n11124), .ZN(n11125) );
  AOI21_X1 U13637 ( .B1(n11126), .B2(n11125), .A(n13417), .ZN(n11129) );
  NOR3_X1 U13638 ( .A1(n13408), .A2(n11127), .A3(n11130), .ZN(n11128) );
  OAI21_X1 U13639 ( .B1(n11129), .B2(n11128), .A(n11159), .ZN(n11134) );
  OAI22_X1 U13640 ( .A1(n13389), .A2(n11130), .B1(n11363), .B2(n13406), .ZN(
        n11131) );
  AOI211_X1 U13641 ( .C1(n13422), .C2(n13446), .A(n11132), .B(n11131), .ZN(
        n11133) );
  OAI211_X1 U13642 ( .C1(n7484), .C2(n13369), .A(n11134), .B(n11133), .ZN(
        P2_U3185) );
  INV_X1 U13643 ( .A(n13483), .ZN(n13476) );
  INV_X1 U13644 ( .A(n11135), .ZN(n11136) );
  OAI222_X1 U13645 ( .A1(P2_U3088), .A2(n13476), .B1(n13850), .B2(n11136), 
        .C1(n14648), .C2(n13844), .ZN(P2_U3311) );
  OAI222_X1 U13646 ( .A1(P1_U3086), .A2(n12060), .B1(n14383), .B2(n11136), 
        .C1(n14636), .C2(n14395), .ZN(P1_U3339) );
  OR2_X1 U13647 ( .A1(n11138), .A2(n11137), .ZN(n11139) );
  NAND2_X1 U13648 ( .A1(n11140), .A2(n11139), .ZN(n15139) );
  OAI21_X1 U13649 ( .B1(n11143), .B2(n11142), .A(n11141), .ZN(n11147) );
  NAND2_X1 U13650 ( .A1(n14979), .A2(n14267), .ZN(n11144) );
  OAI21_X1 U13651 ( .B1(n11145), .B2(n14220), .A(n11144), .ZN(n11146) );
  AOI21_X1 U13652 ( .B1(n11147), .B2(n15098), .A(n11146), .ZN(n11149) );
  NAND2_X1 U13653 ( .A1(n15139), .A2(n15102), .ZN(n11148) );
  NAND2_X1 U13654 ( .A1(n11149), .A2(n11148), .ZN(n15144) );
  MUX2_X1 U13655 ( .A(n15144), .B(P1_REG2_REG_3__SCAN_IN), .S(n15118), .Z(
        n11155) );
  NAND2_X1 U13656 ( .A1(n11185), .A2(n11150), .ZN(n11151) );
  NAND2_X1 U13657 ( .A1(n11151), .A2(n15111), .ZN(n11152) );
  NOR2_X1 U13658 ( .A1(n11171), .A2(n11152), .ZN(n15140) );
  INV_X1 U13659 ( .A(n14801), .ZN(n15103) );
  AOI22_X1 U13660 ( .A1(n15113), .A2(n15140), .B1(n15103), .B2(n14623), .ZN(
        n11153) );
  OAI21_X1 U13661 ( .B1(n6946), .B2(n15107), .A(n11153), .ZN(n11154) );
  AOI211_X1 U13662 ( .C1(n15114), .C2(n15139), .A(n11155), .B(n11154), .ZN(
        n11156) );
  INV_X1 U13663 ( .A(n11156), .ZN(P1_U3290) );
  NAND3_X1 U13664 ( .A1(n13415), .A2(n13447), .A3(n11157), .ZN(n11158) );
  OAI21_X1 U13665 ( .B1(n11159), .B2(n13417), .A(n11158), .ZN(n11162) );
  INV_X1 U13666 ( .A(n11160), .ZN(n11161) );
  NAND2_X1 U13667 ( .A1(n11162), .A2(n11161), .ZN(n11169) );
  OAI21_X1 U13668 ( .B1(n13389), .B2(n11164), .A(n11163), .ZN(n11167) );
  OAI22_X1 U13669 ( .A1(n13390), .A2(n11165), .B1(n13406), .B2(n11431), .ZN(
        n11166) );
  AOI211_X1 U13670 ( .C1(n11484), .C2(n13425), .A(n11167), .B(n11166), .ZN(
        n11168) );
  OAI211_X1 U13671 ( .C1(n11251), .C2(n13417), .A(n11169), .B(n11168), .ZN(
        P2_U3193) );
  XNOR2_X1 U13672 ( .A(n11170), .B(n11176), .ZN(n15146) );
  OAI211_X1 U13673 ( .C1(n11171), .C2(n15149), .A(n15111), .B(n15109), .ZN(
        n15148) );
  OAI22_X1 U13674 ( .A1(n14816), .A2(n15148), .B1(n11172), .B2(n14801), .ZN(
        n11173) );
  AOI21_X1 U13675 ( .B1(n14255), .B2(n11174), .A(n11173), .ZN(n11181) );
  XNOR2_X1 U13676 ( .A(n11175), .B(n11176), .ZN(n11177) );
  NAND2_X1 U13677 ( .A1(n11177), .A2(n15098), .ZN(n15150) );
  AOI22_X1 U13678 ( .A1(n14812), .A2(n13963), .B1(n14979), .B2(n13965), .ZN(
        n15147) );
  AND2_X1 U13679 ( .A1(n15150), .A2(n15147), .ZN(n11179) );
  MUX2_X1 U13680 ( .A(n11179), .B(n11178), .S(n14251), .Z(n11180) );
  OAI211_X1 U13681 ( .C1(n14210), .C2(n15146), .A(n11181), .B(n11180), .ZN(
        P1_U3289) );
  OAI21_X1 U13682 ( .B1(n11184), .B2(n11183), .A(n11182), .ZN(n15132) );
  INV_X1 U13683 ( .A(n15132), .ZN(n11202) );
  OAI211_X1 U13684 ( .C1(n14258), .C2(n15135), .A(n15111), .B(n11185), .ZN(
        n15133) );
  OAI22_X1 U13685 ( .A1(n14816), .A2(n15133), .B1(n11186), .B2(n14801), .ZN(
        n11187) );
  AOI21_X1 U13686 ( .B1(n14255), .B2(n11188), .A(n11187), .ZN(n11201) );
  OAI21_X1 U13687 ( .B1(n11191), .B2(n11190), .A(n11189), .ZN(n11195) );
  NAND2_X1 U13688 ( .A1(n14979), .A2(n13966), .ZN(n11192) );
  OAI21_X1 U13689 ( .B1(n11193), .B2(n14220), .A(n11192), .ZN(n11194) );
  AOI21_X1 U13690 ( .B1(n11195), .B2(n15098), .A(n11194), .ZN(n11197) );
  NAND2_X1 U13691 ( .A1(n15132), .A2(n15102), .ZN(n11196) );
  NAND2_X1 U13692 ( .A1(n11197), .A2(n11196), .ZN(n15137) );
  INV_X1 U13693 ( .A(n15137), .ZN(n11199) );
  MUX2_X1 U13694 ( .A(n11199), .B(n11198), .S(n14251), .Z(n11200) );
  OAI211_X1 U13695 ( .C1(n11202), .C2(n11765), .A(n11201), .B(n11200), .ZN(
        P1_U3291) );
  OR2_X1 U13696 ( .A1(n11203), .A2(n15362), .ZN(n11204) );
  OAI21_X1 U13697 ( .B1(n15364), .B2(n7834), .A(n11204), .ZN(P2_U3445) );
  INV_X1 U13698 ( .A(n11205), .ZN(n11207) );
  OAI222_X1 U13699 ( .A1(P3_U3151), .A2(n12651), .B1(n12306), .B2(n11207), 
        .C1(n11206), .C2(n12423), .ZN(P3_U3274) );
  NAND2_X1 U13700 ( .A1(n11219), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U13701 ( .A1(n11209), .A2(n11208), .ZN(n11212) );
  INV_X1 U13702 ( .A(n11212), .ZN(n11214) );
  MUX2_X1 U13703 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11210), .S(n11396), .Z(
        n11213) );
  MUX2_X1 U13704 ( .A(n11210), .B(P2_REG2_REG_11__SCAN_IN), .S(n11396), .Z(
        n11211) );
  OAI21_X1 U13705 ( .B1(n11214), .B2(n11213), .A(n11405), .ZN(n11224) );
  INV_X1 U13706 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n11217) );
  NOR2_X1 U13707 ( .A1(n11215), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11782) );
  AOI21_X1 U13708 ( .B1(n15281), .B2(n11396), .A(n11782), .ZN(n11216) );
  OAI21_X1 U13709 ( .B1(n15269), .B2(n11217), .A(n11216), .ZN(n11223) );
  MUX2_X1 U13710 ( .A(n11814), .B(P2_REG1_REG_11__SCAN_IN), .S(n11396), .Z(
        n11220) );
  AOI211_X1 U13711 ( .C1(n11221), .C2(n11220), .A(n15271), .B(n11395), .ZN(
        n11222) );
  AOI211_X1 U13712 ( .C1(n15277), .C2(n11224), .A(n11223), .B(n11222), .ZN(
        n11225) );
  INV_X1 U13713 ( .A(n11225), .ZN(P2_U3225) );
  INV_X1 U13714 ( .A(n14027), .ZN(n14023) );
  INV_X1 U13715 ( .A(n11226), .ZN(n11228) );
  OAI222_X1 U13716 ( .A1(P1_U3086), .A2(n14023), .B1(n14398), .B2(n11228), 
        .C1(n14610), .C2(n14395), .ZN(P1_U3338) );
  INV_X1 U13717 ( .A(n15280), .ZN(n13479) );
  OAI222_X1 U13718 ( .A1(P2_U3088), .A2(n13479), .B1(n13850), .B2(n11228), 
        .C1(n11227), .C2(n13844), .ZN(P2_U3310) );
  INV_X1 U13719 ( .A(n11229), .ZN(n11230) );
  NAND2_X1 U13720 ( .A1(n11230), .A2(n12825), .ZN(n11231) );
  INV_X1 U13721 ( .A(n12824), .ZN(n11552) );
  NAND2_X1 U13722 ( .A1(n11233), .A2(n11552), .ZN(n11453) );
  INV_X1 U13723 ( .A(n11233), .ZN(n11234) );
  NAND2_X1 U13724 ( .A1(n11234), .A2(n12824), .ZN(n11235) );
  OAI21_X1 U13725 ( .B1(n11237), .B2(n11236), .A(n11454), .ZN(n11238) );
  NAND2_X1 U13726 ( .A1(n11238), .A2(n12572), .ZN(n11244) );
  AOI21_X1 U13727 ( .B1(n12574), .B2(n11859), .A(n11239), .ZN(n11240) );
  OAI21_X1 U13728 ( .B1(n15488), .B2(n12576), .A(n11240), .ZN(n11241) );
  AOI21_X1 U13729 ( .B1(n12590), .B2(n11242), .A(n11241), .ZN(n11243) );
  OAI211_X1 U13730 ( .C1(n11857), .C2(n12588), .A(n11244), .B(n11243), .ZN(
        P3_U3170) );
  INV_X1 U13731 ( .A(n11245), .ZN(n11250) );
  NAND2_X1 U13732 ( .A1(n11246), .A2(n10187), .ZN(n11247) );
  OAI21_X1 U13733 ( .B1(n11248), .B2(n13408), .A(n11247), .ZN(n11249) );
  NAND3_X1 U13734 ( .A1(n11251), .A2(n11250), .A3(n11249), .ZN(n11257) );
  AOI21_X1 U13735 ( .B1(n13422), .B2(n13444), .A(n11252), .ZN(n11256) );
  INV_X1 U13736 ( .A(n11647), .ZN(n11253) );
  AOI22_X1 U13737 ( .A1(n11253), .A2(n13424), .B1(n13421), .B2(n13446), .ZN(
        n11255) );
  NAND2_X1 U13738 ( .A1(n15355), .A2(n13425), .ZN(n11254) );
  AND4_X1 U13739 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11258) );
  OAI21_X1 U13740 ( .B1(n11259), .B2(n13417), .A(n11258), .ZN(P2_U3203) );
  INV_X1 U13741 ( .A(n11260), .ZN(n11262) );
  OAI22_X1 U13742 ( .A1(n12810), .A2(P3_U3151), .B1(SI_22_), .B2(n12423), .ZN(
        n11261) );
  AOI21_X1 U13743 ( .B1(n11262), .B2(n13291), .A(n11261), .ZN(P3_U3273) );
  NOR2_X1 U13744 ( .A1(n15374), .A2(n6715), .ZN(n15373) );
  NOR2_X1 U13745 ( .A1(n11265), .A2(n15373), .ZN(n15390) );
  AOI22_X1 U13746 ( .A1(n11297), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n11296), 
        .B2(n15397), .ZN(n15389) );
  NOR2_X1 U13747 ( .A1(n15390), .A2(n15389), .ZN(n15388) );
  AOI21_X1 U13748 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n15397), .A(n15388), .ZN(
        n11266) );
  NOR2_X1 U13749 ( .A1(n11304), .A2(n11266), .ZN(n11267) );
  XNOR2_X1 U13750 ( .A(n11304), .B(n11266), .ZN(n15409) );
  NOR2_X1 U13751 ( .A1(n11303), .A2(n15409), .ZN(n15408) );
  AOI22_X1 U13752 ( .A1(n11311), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n11310), 
        .B2(n15435), .ZN(n15427) );
  INV_X1 U13753 ( .A(n11268), .ZN(n11270) );
  NAND2_X1 U13754 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11470), .ZN(n11271) );
  OAI21_X1 U13755 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11470), .A(n11271), 
        .ZN(n11272) );
  AOI21_X1 U13756 ( .B1(n6821), .B2(n11272), .A(n11463), .ZN(n11336) );
  AOI22_X1 U13757 ( .A1(n11323), .A2(n11322), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11470), .ZN(n11281) );
  AOI22_X1 U13758 ( .A1(n11311), .A2(n11309), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n15435), .ZN(n15440) );
  AOI22_X1 U13759 ( .A1(n11297), .A2(n11295), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n15397), .ZN(n15402) );
  OAI21_X1 U13760 ( .B1(n11288), .B2(n9598), .A(n11273), .ZN(n11274) );
  NAND2_X1 U13761 ( .A1(n11274), .A2(n7028), .ZN(n11275) );
  XNOR2_X1 U13762 ( .A(n11274), .B(n11293), .ZN(n15383) );
  NAND2_X1 U13763 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n15383), .ZN(n15382) );
  NAND2_X1 U13764 ( .A1(n15416), .A2(n11276), .ZN(n11277) );
  NAND2_X1 U13765 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15421), .ZN(n15420) );
  NAND2_X1 U13766 ( .A1(n11278), .A2(n15455), .ZN(n11279) );
  NAND2_X1 U13767 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15462), .ZN(n15461) );
  NAND2_X1 U13768 ( .A1(n11279), .A2(n15461), .ZN(n11280) );
  NAND2_X1 U13769 ( .A1(n11281), .A2(n11280), .ZN(n11471) );
  OAI21_X1 U13770 ( .B1(n11281), .B2(n11280), .A(n11471), .ZN(n11284) );
  AND2_X1 U13771 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11745) );
  AOI21_X1 U13772 ( .B1(n15460), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11745), 
        .ZN(n11282) );
  OAI21_X1 U13773 ( .B1(n15454), .B2(n11470), .A(n11282), .ZN(n11283) );
  AOI21_X1 U13774 ( .B1(n11284), .B2(n15463), .A(n11283), .ZN(n11335) );
  NAND2_X1 U13775 ( .A1(n11286), .A2(n11285), .ZN(n11291) );
  INV_X1 U13776 ( .A(n11287), .ZN(n11289) );
  NAND2_X1 U13777 ( .A1(n11289), .A2(n11288), .ZN(n11290) );
  NAND2_X1 U13778 ( .A1(n11291), .A2(n11290), .ZN(n15375) );
  MUX2_X1 U13779 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12913), .Z(n11292) );
  NAND2_X1 U13780 ( .A1(n11292), .A2(n7028), .ZN(n15376) );
  NAND2_X1 U13781 ( .A1(n15375), .A2(n15376), .ZN(n15395) );
  INV_X1 U13782 ( .A(n11292), .ZN(n11294) );
  NAND2_X1 U13783 ( .A1(n11294), .A2(n11293), .ZN(n15391) );
  NAND2_X1 U13784 ( .A1(n15395), .A2(n15391), .ZN(n11301) );
  MUX2_X1 U13785 ( .A(n11296), .B(n11295), .S(n12913), .Z(n11298) );
  NAND2_X1 U13786 ( .A1(n11298), .A2(n11297), .ZN(n15410) );
  INV_X1 U13787 ( .A(n11298), .ZN(n11299) );
  NAND2_X1 U13788 ( .A1(n11299), .A2(n15397), .ZN(n11300) );
  AND2_X1 U13789 ( .A1(n15410), .A2(n11300), .ZN(n15393) );
  NAND2_X1 U13790 ( .A1(n11301), .A2(n15393), .ZN(n15414) );
  NAND2_X1 U13791 ( .A1(n15414), .A2(n15410), .ZN(n11308) );
  MUX2_X1 U13792 ( .A(n11303), .B(n11302), .S(n12913), .Z(n11305) );
  NAND2_X1 U13793 ( .A1(n11305), .A2(n11304), .ZN(n15429) );
  INV_X1 U13794 ( .A(n11305), .ZN(n11306) );
  NAND2_X1 U13795 ( .A1(n11306), .A2(n15416), .ZN(n11307) );
  AND2_X1 U13796 ( .A1(n15429), .A2(n11307), .ZN(n15412) );
  NAND2_X1 U13797 ( .A1(n11308), .A2(n15412), .ZN(n15433) );
  NAND2_X1 U13798 ( .A1(n15433), .A2(n15429), .ZN(n11315) );
  MUX2_X1 U13799 ( .A(n11310), .B(n11309), .S(n12913), .Z(n11312) );
  NAND2_X1 U13800 ( .A1(n11312), .A2(n11311), .ZN(n15448) );
  INV_X1 U13801 ( .A(n11312), .ZN(n11313) );
  NAND2_X1 U13802 ( .A1(n11313), .A2(n15435), .ZN(n11314) );
  AND2_X1 U13803 ( .A1(n15448), .A2(n11314), .ZN(n15431) );
  NAND2_X1 U13804 ( .A1(n11315), .A2(n15431), .ZN(n15452) );
  NAND2_X1 U13805 ( .A1(n15452), .A2(n15448), .ZN(n11321) );
  MUX2_X1 U13806 ( .A(n11851), .B(n11316), .S(n12913), .Z(n11318) );
  NAND2_X1 U13807 ( .A1(n11318), .A2(n11317), .ZN(n11328) );
  INV_X1 U13808 ( .A(n11318), .ZN(n11319) );
  NAND2_X1 U13809 ( .A1(n11319), .A2(n15455), .ZN(n11320) );
  AND2_X1 U13810 ( .A1(n11328), .A2(n11320), .ZN(n15450) );
  NAND2_X1 U13811 ( .A1(n11321), .A2(n15450), .ZN(n11329) );
  INV_X1 U13812 ( .A(n11329), .ZN(n15451) );
  INV_X1 U13813 ( .A(n11328), .ZN(n11327) );
  MUX2_X1 U13814 ( .A(n11988), .B(n11322), .S(n12936), .Z(n11324) );
  NAND2_X1 U13815 ( .A1(n11324), .A2(n11323), .ZN(n11466) );
  INV_X1 U13816 ( .A(n11324), .ZN(n11325) );
  NAND2_X1 U13817 ( .A1(n11325), .A2(n11470), .ZN(n11326) );
  AND2_X1 U13818 ( .A1(n11466), .A2(n11326), .ZN(n11330) );
  NOR3_X1 U13819 ( .A1(n15451), .A2(n11327), .A3(n11330), .ZN(n11333) );
  NAND2_X1 U13820 ( .A1(n11329), .A2(n11328), .ZN(n11331) );
  NAND2_X1 U13821 ( .A1(n11331), .A2(n11330), .ZN(n11467) );
  INV_X1 U13822 ( .A(n11467), .ZN(n11332) );
  OAI21_X1 U13823 ( .B1(n11333), .B2(n11332), .A(n12954), .ZN(n11334) );
  OAI211_X1 U13824 ( .C1(n11336), .C2(n15467), .A(n11335), .B(n11334), .ZN(
        P3_U3192) );
  MUX2_X1 U13825 ( .A(n11922), .B(P1_REG1_REG_14__SCAN_IN), .S(n11343), .Z(
        n11339) );
  OAI21_X1 U13826 ( .B1(n14987), .B2(n11342), .A(n11337), .ZN(n11338) );
  AOI21_X1 U13827 ( .B1(n11339), .B2(n11338), .A(n11921), .ZN(n11351) );
  NAND2_X1 U13828 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14922)
         );
  INV_X1 U13829 ( .A(n14922), .ZN(n11341) );
  NOR2_X1 U13830 ( .A1(n15054), .A2(n11927), .ZN(n11340) );
  AOI211_X1 U13831 ( .C1(n15031), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n11341), 
        .B(n11340), .ZN(n11350) );
  NOR2_X1 U13832 ( .A1(n11342), .A2(n14803), .ZN(n11346) );
  MUX2_X1 U13833 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11344), .S(n11343), .Z(
        n11345) );
  OAI21_X1 U13834 ( .B1(n11347), .B2(n11346), .A(n11345), .ZN(n11926) );
  OR3_X1 U13835 ( .A1(n11347), .A2(n11346), .A3(n11345), .ZN(n11348) );
  NAND3_X1 U13836 ( .A1(n11926), .A2(n15044), .A3(n11348), .ZN(n11349) );
  OAI211_X1 U13837 ( .C1(n11351), .C2(n12065), .A(n11350), .B(n11349), .ZN(
        P1_U3257) );
  XNOR2_X1 U13838 ( .A(n11352), .B(n7042), .ZN(n15347) );
  INV_X1 U13839 ( .A(n11353), .ZN(n11354) );
  NAND2_X1 U13840 ( .A1(n11444), .A2(n11354), .ZN(n11356) );
  NAND2_X1 U13841 ( .A1(n11356), .A2(n11355), .ZN(n11358) );
  NAND3_X1 U13842 ( .A1(n11358), .A2(n13586), .A3(n11357), .ZN(n11360) );
  AOI22_X1 U13843 ( .A1(n13607), .A2(n13448), .B1(n13446), .B2(n13604), .ZN(
        n11359) );
  NAND2_X1 U13844 ( .A1(n11360), .A2(n11359), .ZN(n15353) );
  MUX2_X1 U13845 ( .A(n15353), .B(P2_REG2_REG_7__SCAN_IN), .S(n15301), .Z(
        n11361) );
  INV_X1 U13846 ( .A(n11361), .ZN(n11366) );
  XNOR2_X1 U13847 ( .A(n11438), .B(n7484), .ZN(n11362) );
  AND2_X1 U13848 ( .A1(n11362), .A2(n10146), .ZN(n15350) );
  OAI22_X1 U13849 ( .A1(n15292), .A2(n7484), .B1(n11363), .B2(n13683), .ZN(
        n11364) );
  AOI21_X1 U13850 ( .B1(n15297), .B2(n15350), .A(n11364), .ZN(n11365) );
  OAI211_X1 U13851 ( .C1(n15347), .C2(n15293), .A(n11366), .B(n11365), .ZN(
        P2_U3258) );
  XNOR2_X1 U13852 ( .A(n11367), .B(n11371), .ZN(n11368) );
  NAND2_X1 U13853 ( .A1(n11368), .A2(n15098), .ZN(n11369) );
  AOI22_X1 U13854 ( .A1(n14812), .A2(n14927), .B1(n14979), .B2(n13961), .ZN(
        n11875) );
  NAND2_X1 U13855 ( .A1(n11369), .A2(n11875), .ZN(n15180) );
  INV_X1 U13856 ( .A(n15180), .ZN(n11378) );
  XNOR2_X1 U13857 ( .A(n11370), .B(n11371), .ZN(n15182) );
  AOI21_X1 U13858 ( .B1(n15089), .B2(n15177), .A(n15125), .ZN(n11372) );
  NAND2_X1 U13859 ( .A1(n11372), .A2(n15074), .ZN(n15178) );
  NAND2_X1 U13860 ( .A1(n14255), .A2(n15177), .ZN(n11375) );
  NOR2_X1 U13861 ( .A1(n14801), .A2(n11876), .ZN(n11373) );
  AOI21_X1 U13862 ( .B1(n14251), .B2(P1_REG2_REG_8__SCAN_IN), .A(n11373), .ZN(
        n11374) );
  OAI211_X1 U13863 ( .C1(n15178), .C2(n14816), .A(n11375), .B(n11374), .ZN(
        n11376) );
  AOI21_X1 U13864 ( .B1(n15182), .B2(n14809), .A(n11376), .ZN(n11377) );
  OAI21_X1 U13865 ( .B1(n11378), .B2(n15118), .A(n11377), .ZN(P1_U3285) );
  XNOR2_X1 U13866 ( .A(n11379), .B(n11380), .ZN(n15532) );
  INV_X1 U13867 ( .A(n15532), .ZN(n11393) );
  AND2_X1 U13868 ( .A1(n12804), .A2(n11381), .ZN(n15498) );
  NAND2_X1 U13869 ( .A1(n15501), .A2(n15498), .ZN(n12290) );
  OAI22_X1 U13870 ( .A1(n15508), .A2(n15509), .B1(n11552), .B2(n15507), .ZN(
        n11387) );
  INV_X1 U13871 ( .A(n11382), .ZN(n11385) );
  AOI21_X1 U13872 ( .B1(n15492), .B2(n11383), .A(n12626), .ZN(n11384) );
  NOR3_X1 U13873 ( .A1(n11385), .A2(n11384), .A3(n15490), .ZN(n11386) );
  AOI211_X1 U13874 ( .C1(n15532), .C2(n15495), .A(n11387), .B(n11386), .ZN(
        n15529) );
  MUX2_X1 U13875 ( .A(n11388), .B(n15529), .S(n15501), .Z(n11392) );
  INV_X1 U13876 ( .A(n15482), .ZN(n14860) );
  NOR2_X1 U13877 ( .A1(n11389), .A2(n15545), .ZN(n15531) );
  AOI22_X1 U13878 ( .A1(n14860), .A2(n15531), .B1(n15517), .B2(n11390), .ZN(
        n11391) );
  OAI211_X1 U13879 ( .C1(n11393), .C2(n12290), .A(n11392), .B(n11391), .ZN(
        P3_U3230) );
  NAND2_X1 U13880 ( .A1(n12816), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11394) );
  OAI21_X1 U13881 ( .B1(n12473), .B2(n12816), .A(n11394), .ZN(P3_U3519) );
  MUX2_X1 U13882 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11397), .S(n11618), .Z(
        n11398) );
  NAND2_X1 U13883 ( .A1(n11399), .A2(n11398), .ZN(n11617) );
  OAI21_X1 U13884 ( .B1(n11399), .B2(n11398), .A(n11617), .ZN(n11410) );
  NAND2_X1 U13885 ( .A1(n11400), .A2(n11210), .ZN(n11403) );
  NAND2_X1 U13886 ( .A1(n11405), .A2(n11403), .ZN(n11401) );
  MUX2_X1 U13887 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11912), .S(n11618), .Z(
        n11402) );
  NAND2_X1 U13888 ( .A1(n11401), .A2(n11402), .ZN(n11623) );
  INV_X1 U13889 ( .A(n11402), .ZN(n11404) );
  NAND3_X1 U13890 ( .A1(n11405), .A2(n11404), .A3(n11403), .ZN(n11406) );
  AOI21_X1 U13891 ( .B1(n11623), .B2(n11406), .A(n13489), .ZN(n11409) );
  NAND2_X1 U13892 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11726)
         );
  NAND2_X1 U13893 ( .A1(n15281), .A2(n11618), .ZN(n11407) );
  OAI211_X1 U13894 ( .C1(n15269), .C2(n15008), .A(n11726), .B(n11407), .ZN(
        n11408) );
  AOI211_X1 U13895 ( .C1(n11410), .C2(n15231), .A(n11409), .B(n11408), .ZN(
        n11411) );
  INV_X1 U13896 ( .A(n11411), .ZN(P2_U3226) );
  NAND2_X1 U13897 ( .A1(n12816), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11412) );
  OAI21_X1 U13898 ( .B1(n12977), .B2(n12816), .A(n11412), .ZN(P3_U3520) );
  NAND2_X1 U13899 ( .A1(n11413), .A2(n13291), .ZN(n11414) );
  OAI211_X1 U13900 ( .C1(n11415), .C2(n12423), .A(n11414), .B(n12812), .ZN(
        P3_U3272) );
  NAND2_X1 U13901 ( .A1(n11416), .A2(n11421), .ZN(n11417) );
  NAND2_X1 U13902 ( .A1(n11418), .A2(n11417), .ZN(n11487) );
  OR2_X1 U13903 ( .A1(n11487), .A2(n10061), .ZN(n11420) );
  AOI22_X1 U13904 ( .A1(n13607), .A2(n13447), .B1(n13445), .B2(n13604), .ZN(
        n11419) );
  AND2_X1 U13905 ( .A1(n11420), .A2(n11419), .ZN(n11426) );
  INV_X1 U13906 ( .A(n11421), .ZN(n11422) );
  XNOR2_X1 U13907 ( .A(n11423), .B(n11422), .ZN(n11424) );
  NAND2_X1 U13908 ( .A1(n11424), .A2(n13705), .ZN(n11425) );
  NAND2_X1 U13909 ( .A1(n11426), .A2(n11425), .ZN(n11482) );
  MUX2_X1 U13910 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11482), .S(n13689), .Z(
        n11427) );
  INV_X1 U13911 ( .A(n11427), .ZN(n11435) );
  NAND2_X1 U13912 ( .A1(n11484), .A2(n11428), .ZN(n11429) );
  NAND2_X1 U13913 ( .A1(n11429), .A2(n10146), .ZN(n11430) );
  NOR2_X1 U13914 ( .A1(n11643), .A2(n11430), .ZN(n11483) );
  INV_X1 U13915 ( .A(n11484), .ZN(n11432) );
  OAI22_X1 U13916 ( .A1(n11432), .A2(n15292), .B1(n13683), .B2(n11431), .ZN(
        n11433) );
  AOI21_X1 U13917 ( .B1(n11483), .B2(n15297), .A(n11433), .ZN(n11434) );
  OAI211_X1 U13918 ( .C1(n11487), .C2(n13618), .A(n11435), .B(n11434), .ZN(
        P2_U3257) );
  XNOR2_X1 U13919 ( .A(n11437), .B(n11436), .ZN(n15340) );
  OAI211_X1 U13920 ( .C1(n11439), .C2(n15343), .A(n10146), .B(n11438), .ZN(
        n15341) );
  INV_X1 U13921 ( .A(n11440), .ZN(n11441) );
  AOI22_X1 U13922 ( .A1(n13685), .A2(n11442), .B1(n15288), .B2(n11441), .ZN(
        n11443) );
  OAI21_X1 U13923 ( .B1(n13519), .B2(n15341), .A(n11443), .ZN(n11451) );
  OAI21_X1 U13924 ( .B1(n11446), .B2(n11445), .A(n11444), .ZN(n11447) );
  NAND2_X1 U13925 ( .A1(n11447), .A2(n13705), .ZN(n11449) );
  AOI22_X1 U13926 ( .A1(n13607), .A2(n13449), .B1(n13447), .B2(n13604), .ZN(
        n11448) );
  NAND2_X1 U13927 ( .A1(n11449), .A2(n11448), .ZN(n15346) );
  MUX2_X1 U13928 ( .A(n15346), .B(P2_REG2_REG_6__SCAN_IN), .S(n15301), .Z(
        n11450) );
  AOI211_X1 U13929 ( .C1(n13652), .C2(n15340), .A(n11451), .B(n11450), .ZN(
        n11452) );
  INV_X1 U13930 ( .A(n11452), .ZN(P2_U3259) );
  XNOR2_X1 U13931 ( .A(n12466), .B(n11460), .ZN(n11579) );
  XNOR2_X1 U13932 ( .A(n11579), .B(n11859), .ZN(n11456) );
  NAND2_X1 U13933 ( .A1(n11454), .A2(n11453), .ZN(n11455) );
  NAND2_X1 U13934 ( .A1(n11455), .A2(n11456), .ZN(n11685) );
  OAI21_X1 U13935 ( .B1(n11456), .B2(n11455), .A(n11685), .ZN(n11457) );
  NAND2_X1 U13936 ( .A1(n11457), .A2(n12572), .ZN(n11462) );
  INV_X1 U13937 ( .A(n12823), .ZN(n15473) );
  INV_X1 U13938 ( .A(n12576), .ZN(n12586) );
  NOR2_X1 U13939 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14661), .ZN(n15381) );
  AOI21_X1 U13940 ( .B1(n12586), .B2(n12824), .A(n15381), .ZN(n11458) );
  OAI21_X1 U13941 ( .B1(n15473), .B2(n12584), .A(n11458), .ZN(n11459) );
  AOI21_X1 U13942 ( .B1(n12590), .B2(n11460), .A(n11459), .ZN(n11461) );
  OAI211_X1 U13943 ( .C1(n11559), .C2(n12588), .A(n11462), .B(n11461), .ZN(
        P3_U3167) );
  AOI21_X1 U13944 ( .B1(n11465), .B2(n9708), .A(n11653), .ZN(n11481) );
  NAND2_X1 U13945 ( .A1(n11467), .A2(n11466), .ZN(n11469) );
  MUX2_X1 U13946 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12913), .Z(n11666) );
  XNOR2_X1 U13947 ( .A(n11666), .B(n11667), .ZN(n11468) );
  NAND2_X1 U13948 ( .A1(n11469), .A2(n11468), .ZN(n11672) );
  OAI21_X1 U13949 ( .B1(n11469), .B2(n11468), .A(n11672), .ZN(n11479) );
  NAND2_X1 U13950 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11470), .ZN(n11472) );
  NAND2_X1 U13951 ( .A1(n11472), .A2(n11471), .ZN(n11659) );
  XNOR2_X1 U13952 ( .A(n11659), .B(n11667), .ZN(n11473) );
  NAND2_X1 U13953 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11473), .ZN(n11660) );
  OAI21_X1 U13954 ( .B1(n11473), .B2(P3_REG1_REG_11__SCAN_IN), .A(n11660), 
        .ZN(n11474) );
  NAND2_X1 U13955 ( .A1(n11474), .A2(n15463), .ZN(n11477) );
  INV_X1 U13956 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11475) );
  NOR2_X1 U13957 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11475), .ZN(n12002) );
  AOI21_X1 U13958 ( .B1(n15460), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12002), 
        .ZN(n11476) );
  OAI211_X1 U13959 ( .C1(n15454), .C2(n11658), .A(n11477), .B(n11476), .ZN(
        n11478) );
  AOI21_X1 U13960 ( .B1(n12954), .B2(n11479), .A(n11478), .ZN(n11480) );
  OAI21_X1 U13961 ( .B1(n11481), .B2(n15467), .A(n11480), .ZN(P3_U3193) );
  INV_X1 U13962 ( .A(n11482), .ZN(n11486) );
  AOI21_X1 U13963 ( .B1(n15356), .B2(n11484), .A(n11483), .ZN(n11485) );
  OAI211_X1 U13964 ( .C1(n13756), .C2(n11487), .A(n11486), .B(n11485), .ZN(
        n13814) );
  NAND2_X1 U13965 ( .A1(n13814), .A2(n15364), .ZN(n11488) );
  OAI21_X1 U13966 ( .B1(n15364), .B2(n7910), .A(n11488), .ZN(P2_U3454) );
  INV_X1 U13967 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n11491) );
  INV_X1 U13968 ( .A(n12616), .ZN(n11489) );
  NAND2_X1 U13969 ( .A1(n11489), .A2(P3_U3897), .ZN(n11490) );
  OAI21_X1 U13970 ( .B1(P3_U3897), .B2(n11491), .A(n11490), .ZN(P3_U3521) );
  XNOR2_X1 U13971 ( .A(n11492), .B(n11496), .ZN(n15197) );
  INV_X1 U13972 ( .A(n15197), .ZN(n11505) );
  INV_X1 U13973 ( .A(n11493), .ZN(n11494) );
  AOI211_X1 U13974 ( .C1(n11496), .C2(n11495), .A(n15083), .B(n11494), .ZN(
        n15195) );
  INV_X1 U13975 ( .A(n14925), .ZN(n11502) );
  AOI211_X1 U13976 ( .C1(n14925), .C2(n15075), .A(n15125), .B(n11541), .ZN(
        n15194) );
  NAND2_X1 U13977 ( .A1(n14812), .A2(n13959), .ZN(n14929) );
  INV_X1 U13978 ( .A(n14929), .ZN(n11497) );
  OAI21_X1 U13979 ( .B1(n15194), .B2(n11497), .A(n15113), .ZN(n11501) );
  NOR2_X1 U13980 ( .A1(n15105), .A2(n14265), .ZN(n14806) );
  OAI22_X1 U13981 ( .A1(n14804), .A2(n11498), .B1(n14937), .B2(n14801), .ZN(
        n11499) );
  AOI21_X1 U13982 ( .B1(n14806), .B2(n14927), .A(n11499), .ZN(n11500) );
  OAI211_X1 U13983 ( .C1(n11502), .C2(n15107), .A(n11501), .B(n11500), .ZN(
        n11503) );
  AOI21_X1 U13984 ( .B1(n15195), .B2(n14804), .A(n11503), .ZN(n11504) );
  OAI21_X1 U13985 ( .B1(n11505), .B2(n14210), .A(n11504), .ZN(P1_U3283) );
  INV_X1 U13986 ( .A(n15104), .ZN(n11526) );
  INV_X1 U13987 ( .A(n11506), .ZN(n11508) );
  AOI22_X1 U13988 ( .A1(n11519), .A2(n10208), .B1(n12409), .B2(n13963), .ZN(
        n11512) );
  XOR2_X1 U13989 ( .A(n10223), .B(n11512), .Z(n11515) );
  OAI22_X1 U13990 ( .A1(n6947), .A2(n12363), .B1(n11513), .B2(n10229), .ZN(
        n11514) );
  NOR2_X1 U13991 ( .A1(n11515), .A2(n11514), .ZN(n11589) );
  NAND2_X1 U13992 ( .A1(n11515), .A2(n11514), .ZN(n11588) );
  INV_X1 U13993 ( .A(n11588), .ZN(n11516) );
  NOR2_X1 U13994 ( .A1(n11589), .A2(n11516), .ZN(n11517) );
  XNOR2_X1 U13995 ( .A(n11590), .B(n11517), .ZN(n11518) );
  NAND2_X1 U13996 ( .A1(n11518), .A2(n14960), .ZN(n11525) );
  AND2_X1 U13997 ( .A1(n11519), .A2(n14980), .ZN(n15154) );
  NAND2_X1 U13998 ( .A1(n13964), .A2(n14979), .ZN(n11521) );
  NAND2_X1 U13999 ( .A1(n14812), .A2(n13962), .ZN(n11520) );
  AND2_X1 U14000 ( .A1(n11521), .A2(n11520), .ZN(n15157) );
  INV_X1 U14001 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n11522) );
  OAI22_X1 U14002 ( .A1(n13949), .A2(n15157), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11522), .ZN(n11523) );
  AOI21_X1 U14003 ( .B1(n14926), .B2(n15154), .A(n11523), .ZN(n11524) );
  OAI211_X1 U14004 ( .C1(n14964), .C2(n11526), .A(n11525), .B(n11524), .ZN(
        P1_U3227) );
  XNOR2_X1 U14005 ( .A(n11527), .B(n12625), .ZN(n15544) );
  INV_X1 U14006 ( .A(n15495), .ZN(n15514) );
  AOI22_X1 U14007 ( .A1(n14851), .A2(n11859), .B1(n12822), .B2(n14853), .ZN(
        n11532) );
  AND2_X1 U14008 ( .A1(n11555), .A2(n11528), .ZN(n11530) );
  OAI211_X1 U14009 ( .C1(n11530), .C2(n12625), .A(n11529), .B(n15511), .ZN(
        n11531) );
  OAI211_X1 U14010 ( .C1(n15544), .C2(n15514), .A(n11532), .B(n11531), .ZN(
        n15547) );
  NAND2_X1 U14011 ( .A1(n15547), .A2(n15501), .ZN(n11535) );
  OAI22_X1 U14012 ( .A1(n15501), .A2(n11296), .B1(n11587), .B2(n15479), .ZN(
        n11533) );
  AOI21_X1 U14013 ( .B1(n13148), .B2(n11584), .A(n11533), .ZN(n11534) );
  OAI211_X1 U14014 ( .C1(n15544), .C2(n12290), .A(n11535), .B(n11534), .ZN(
        P3_U3227) );
  XNOR2_X1 U14015 ( .A(n11537), .B(n11536), .ZN(n11538) );
  OAI222_X1 U14016 ( .A1(n14220), .A2(n12246), .B1(n11538), .B2(n15083), .C1(
        n14265), .C2(n12209), .ZN(n14989) );
  INV_X1 U14017 ( .A(n14989), .ZN(n11546) );
  XNOR2_X1 U14018 ( .A(n11539), .B(n11540), .ZN(n14991) );
  OAI21_X1 U14019 ( .B1(n6956), .B2(n11541), .A(n11759), .ZN(n14988) );
  OAI22_X1 U14020 ( .A1(n14804), .A2(n10739), .B1(n14949), .B2(n14801), .ZN(
        n11542) );
  AOI21_X1 U14021 ( .B1(n12216), .B2(n14255), .A(n11542), .ZN(n11543) );
  OAI21_X1 U14022 ( .B1(n14988), .B2(n12251), .A(n11543), .ZN(n11544) );
  AOI21_X1 U14023 ( .B1(n14991), .B2(n14809), .A(n11544), .ZN(n11545) );
  OAI21_X1 U14024 ( .B1(n11546), .B2(n14251), .A(n11545), .ZN(P1_U3282) );
  INV_X1 U14025 ( .A(n11547), .ZN(n11550) );
  INV_X1 U14026 ( .A(n13492), .ZN(n13496) );
  OAI222_X1 U14027 ( .A1(n13852), .A2(n11548), .B1(n13850), .B2(n11550), .C1(
        n13496), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U14028 ( .A(n14041), .ZN(n14035) );
  OAI222_X1 U14029 ( .A1(P1_U3086), .A2(n14035), .B1(n14398), .B2(n11550), 
        .C1(n11549), .C2(n14395), .ZN(P1_U3337) );
  XNOR2_X1 U14030 ( .A(n11551), .B(n12676), .ZN(n15542) );
  INV_X1 U14031 ( .A(n15542), .ZN(n11563) );
  OAI22_X1 U14032 ( .A1(n11552), .A2(n15509), .B1(n15473), .B2(n15507), .ZN(
        n11557) );
  NAND2_X1 U14033 ( .A1(n11553), .A2(n12676), .ZN(n11554) );
  AOI21_X1 U14034 ( .B1(n11555), .B2(n11554), .A(n15490), .ZN(n11556) );
  AOI211_X1 U14035 ( .C1(n15542), .C2(n15495), .A(n11557), .B(n11556), .ZN(
        n15539) );
  MUX2_X1 U14036 ( .A(n15374), .B(n15539), .S(n15501), .Z(n11562) );
  NOR2_X1 U14037 ( .A1(n11558), .A2(n15545), .ZN(n15541) );
  INV_X1 U14038 ( .A(n11559), .ZN(n11560) );
  AOI22_X1 U14039 ( .A1(n14860), .A2(n15541), .B1(n15517), .B2(n11560), .ZN(
        n11561) );
  OAI211_X1 U14040 ( .C1(n11563), .C2(n12290), .A(n11562), .B(n11561), .ZN(
        P3_U3228) );
  XNOR2_X1 U14041 ( .A(n11565), .B(n11564), .ZN(n11571) );
  OR2_X1 U14042 ( .A1(n11567), .A2(n11566), .ZN(n11568) );
  NAND2_X1 U14043 ( .A1(n11569), .A2(n11568), .ZN(n11734) );
  AOI22_X1 U14044 ( .A1(n13607), .A2(n13445), .B1(n13443), .B2(n13604), .ZN(
        n11794) );
  OAI21_X1 U14045 ( .B1(n11734), .B2(n10061), .A(n11794), .ZN(n11570) );
  AOI21_X1 U14046 ( .B1(n13705), .B2(n11571), .A(n11570), .ZN(n11733) );
  AOI211_X1 U14047 ( .C1(n11803), .C2(n11644), .A(n10861), .B(n6868), .ZN(
        n11731) );
  INV_X1 U14048 ( .A(n11803), .ZN(n11574) );
  INV_X1 U14049 ( .A(n11797), .ZN(n11572) );
  AOI22_X1 U14050 ( .A1(n15290), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11572), 
        .B2(n15288), .ZN(n11573) );
  OAI21_X1 U14051 ( .B1(n11574), .B2(n15292), .A(n11573), .ZN(n11576) );
  NOR2_X1 U14052 ( .A1(n11734), .A2(n13618), .ZN(n11575) );
  AOI211_X1 U14053 ( .C1(n11731), .C2(n15297), .A(n11576), .B(n11575), .ZN(
        n11577) );
  OAI21_X1 U14054 ( .B1(n15290), .B2(n11733), .A(n11577), .ZN(P2_U3255) );
  INV_X1 U14055 ( .A(n11859), .ZN(n11578) );
  NAND2_X1 U14056 ( .A1(n11579), .A2(n11578), .ZN(n11683) );
  AND2_X1 U14057 ( .A1(n11685), .A2(n11683), .ZN(n11581) );
  XNOR2_X1 U14058 ( .A(n12469), .B(n11584), .ZN(n11681) );
  XNOR2_X1 U14059 ( .A(n11681), .B(n12823), .ZN(n11580) );
  NAND2_X1 U14060 ( .A1(n11581), .A2(n11580), .ZN(n11608) );
  OAI211_X1 U14061 ( .C1(n11581), .C2(n11580), .A(n11608), .B(n12572), .ZN(
        n11586) );
  INV_X1 U14062 ( .A(n12822), .ZN(n11688) );
  AND2_X1 U14063 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n15400) );
  AOI21_X1 U14064 ( .B1(n12586), .B2(n11859), .A(n15400), .ZN(n11582) );
  OAI21_X1 U14065 ( .B1(n11688), .B2(n12584), .A(n11582), .ZN(n11583) );
  AOI21_X1 U14066 ( .B1(n12590), .B2(n11584), .A(n11583), .ZN(n11585) );
  OAI211_X1 U14067 ( .C1(n11587), .C2(n12588), .A(n11586), .B(n11585), .ZN(
        P3_U3179) );
  INV_X1 U14068 ( .A(n14926), .ZN(n11604) );
  NAND2_X1 U14069 ( .A1(n11594), .A2(n14980), .ZN(n15162) );
  NAND2_X1 U14070 ( .A1(n11594), .A2(n10208), .ZN(n11592) );
  NAND2_X1 U14071 ( .A1(n12409), .A2(n13962), .ZN(n11591) );
  NAND2_X1 U14072 ( .A1(n11592), .A2(n11591), .ZN(n11593) );
  XNOR2_X1 U14073 ( .A(n11593), .B(n10223), .ZN(n11766) );
  AOI22_X1 U14074 ( .A1(n11594), .A2(n12409), .B1(n12408), .B2(n13962), .ZN(
        n11767) );
  XNOR2_X1 U14075 ( .A(n11766), .B(n11767), .ZN(n11595) );
  NAND2_X1 U14076 ( .A1(n11596), .A2(n11595), .ZN(n11770) );
  OAI211_X1 U14077 ( .C1(n11596), .C2(n11595), .A(n11770), .B(n14960), .ZN(
        n11603) );
  INV_X1 U14078 ( .A(n11597), .ZN(n11601) );
  OAI21_X1 U14079 ( .B1(n13949), .B2(n11599), .A(n11598), .ZN(n11600) );
  AOI21_X1 U14080 ( .B1(n13939), .B2(n11601), .A(n11600), .ZN(n11602) );
  OAI211_X1 U14081 ( .C1(n11604), .C2(n15162), .A(n11603), .B(n11602), .ZN(
        P1_U3239) );
  INV_X1 U14082 ( .A(n8811), .ZN(n11606) );
  INV_X1 U14083 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11605) );
  OAI222_X1 U14084 ( .A1(P1_U3086), .A2(n14206), .B1(n14398), .B2(n11606), 
        .C1(n11605), .C2(n14395), .ZN(P1_U3336) );
  OAI222_X1 U14085 ( .A1(n13844), .A2(n14521), .B1(n13850), .B2(n11606), .C1(
        n13504), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U14086 ( .A(n11681), .ZN(n11607) );
  NAND2_X1 U14087 ( .A1(n11607), .A2(n12823), .ZN(n11686) );
  NAND2_X1 U14088 ( .A1(n11608), .A2(n11686), .ZN(n11818) );
  XNOR2_X1 U14089 ( .A(n15470), .B(n12452), .ZN(n11687) );
  XNOR2_X1 U14090 ( .A(n11818), .B(n11687), .ZN(n11615) );
  INV_X1 U14091 ( .A(n12572), .ZN(n12592) );
  INV_X1 U14092 ( .A(n12821), .ZN(n15472) );
  INV_X1 U14093 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11609) );
  NOR2_X1 U14094 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11609), .ZN(n15419) );
  AOI21_X1 U14095 ( .B1(n12586), .B2(n12823), .A(n15419), .ZN(n11610) );
  OAI21_X1 U14096 ( .B1(n15472), .B2(n12584), .A(n11610), .ZN(n11612) );
  NOR2_X1 U14097 ( .A1(n12588), .A2(n15480), .ZN(n11611) );
  AOI211_X1 U14098 ( .C1(n11613), .C2(n12590), .A(n11612), .B(n11611), .ZN(
        n11614) );
  OAI21_X1 U14099 ( .B1(n11615), .B2(n12592), .A(n11614), .ZN(P3_U3153) );
  MUX2_X1 U14100 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n11616), .S(n11629), .Z(
        n11620) );
  OAI21_X1 U14101 ( .B1(n11618), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11617), 
        .ZN(n11619) );
  NOR2_X1 U14102 ( .A1(n11619), .A2(n11620), .ZN(n11896) );
  AOI211_X1 U14103 ( .C1(n11620), .C2(n11619), .A(n15271), .B(n11896), .ZN(
        n11635) );
  NAND2_X1 U14104 ( .A1(n11621), .A2(n11912), .ZN(n11622) );
  NAND2_X1 U14105 ( .A1(n11623), .A2(n11622), .ZN(n11626) );
  INV_X1 U14106 ( .A(n11626), .ZN(n11628) );
  MUX2_X1 U14107 ( .A(n11624), .B(P2_REG2_REG_13__SCAN_IN), .S(n11629), .Z(
        n11627) );
  MUX2_X1 U14108 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11624), .S(n11629), .Z(
        n11625) );
  OAI211_X1 U14109 ( .C1(n11628), .C2(n11627), .A(n15277), .B(n11894), .ZN(
        n11633) );
  INV_X1 U14110 ( .A(n11629), .ZN(n11897) );
  NOR2_X1 U14111 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11630), .ZN(n11631) );
  AOI21_X1 U14112 ( .B1(n15281), .B2(n11897), .A(n11631), .ZN(n11632) );
  OAI211_X1 U14113 ( .C1(n15269), .C2(n7384), .A(n11633), .B(n11632), .ZN(
        n11634) );
  OR2_X1 U14114 ( .A1(n11635), .A2(n11634), .ZN(P2_U3227) );
  OAI21_X1 U14115 ( .B1(n11637), .B2(n11638), .A(n11636), .ZN(n15359) );
  OAI21_X1 U14116 ( .B1(n11640), .B2(n7527), .A(n11639), .ZN(n11641) );
  AOI222_X1 U14117 ( .A1(n13586), .A2(n11641), .B1(n13444), .B2(n13604), .C1(
        n13446), .C2(n13607), .ZN(n15358) );
  MUX2_X1 U14118 ( .A(n11642), .B(n15358), .S(n13689), .Z(n11651) );
  INV_X1 U14119 ( .A(n11643), .ZN(n11646) );
  INV_X1 U14120 ( .A(n11644), .ZN(n11645) );
  AOI211_X1 U14121 ( .C1(n15355), .C2(n11646), .A(n10861), .B(n11645), .ZN(
        n15354) );
  OAI22_X1 U14122 ( .A1(n11648), .A2(n15292), .B1(n11647), .B2(n13683), .ZN(
        n11649) );
  AOI21_X1 U14123 ( .B1(n15354), .B2(n15297), .A(n11649), .ZN(n11650) );
  OAI211_X1 U14124 ( .C1(n15293), .C2(n15359), .A(n11651), .B(n11650), .ZN(
        P2_U3256) );
  INV_X1 U14125 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11655) );
  NOR2_X1 U14126 ( .A1(n11665), .A2(n11655), .ZN(n11951) );
  INV_X1 U14127 ( .A(n11951), .ZN(n11656) );
  OAI21_X1 U14128 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n11958), .A(n11656), 
        .ZN(n11657) );
  AOI21_X1 U14129 ( .B1(n6814), .B2(n11657), .A(n11952), .ZN(n11679) );
  AOI22_X1 U14130 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11958), .B1(n11665), 
        .B2(n9731), .ZN(n11663) );
  NAND2_X1 U14131 ( .A1(n11659), .A2(n11658), .ZN(n11661) );
  NAND2_X1 U14132 ( .A1(n11661), .A2(n11660), .ZN(n11662) );
  NAND2_X1 U14133 ( .A1(n11663), .A2(n11662), .ZN(n11955) );
  OAI21_X1 U14134 ( .B1(n11663), .B2(n11662), .A(n11955), .ZN(n11677) );
  AND2_X1 U14135 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12052) );
  AOI21_X1 U14136 ( .B1(n15460), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12052), 
        .ZN(n11664) );
  OAI21_X1 U14137 ( .B1(n15454), .B2(n11958), .A(n11664), .ZN(n11676) );
  MUX2_X1 U14138 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12913), .Z(n11959) );
  XNOR2_X1 U14139 ( .A(n11959), .B(n11665), .ZN(n11670) );
  INV_X1 U14140 ( .A(n11666), .ZN(n11668) );
  NAND2_X1 U14141 ( .A1(n11668), .A2(n11667), .ZN(n11671) );
  AND2_X1 U14142 ( .A1(n11670), .A2(n11671), .ZN(n11669) );
  NAND2_X1 U14143 ( .A1(n11672), .A2(n11669), .ZN(n11963) );
  INV_X1 U14144 ( .A(n11963), .ZN(n11674) );
  AOI21_X1 U14145 ( .B1(n11672), .B2(n11671), .A(n11670), .ZN(n11673) );
  NOR3_X1 U14146 ( .A1(n11674), .A2(n11673), .A3(n15456), .ZN(n11675) );
  AOI211_X1 U14147 ( .C1(n15463), .C2(n11677), .A(n11676), .B(n11675), .ZN(
        n11678) );
  OAI21_X1 U14148 ( .B1(n11679), .B2(n15467), .A(n11678), .ZN(P3_U3194) );
  XNOR2_X1 U14149 ( .A(n12469), .B(n11703), .ZN(n11738) );
  XNOR2_X1 U14150 ( .A(n11738), .B(n12820), .ZN(n11698) );
  XNOR2_X1 U14151 ( .A(n12466), .B(n11680), .ZN(n11690) );
  XNOR2_X1 U14152 ( .A(n11690), .B(n12821), .ZN(n11819) );
  NAND2_X1 U14153 ( .A1(n11681), .A2(n15473), .ZN(n11682) );
  AND4_X1 U14154 ( .A1(n11819), .A2(n11687), .A3(n11683), .A4(n11682), .ZN(
        n11684) );
  NAND2_X1 U14155 ( .A1(n11685), .A2(n11684), .ZN(n11695) );
  INV_X1 U14156 ( .A(n11819), .ZN(n11689) );
  OAI21_X1 U14157 ( .B1(n11689), .B2(n11686), .A(n11687), .ZN(n11693) );
  INV_X1 U14158 ( .A(n11687), .ZN(n11817) );
  OAI21_X1 U14159 ( .B1(n11689), .B2(n11688), .A(n11817), .ZN(n11692) );
  INV_X1 U14160 ( .A(n11690), .ZN(n11691) );
  AOI22_X1 U14161 ( .A1(n11693), .A2(n11692), .B1(n11691), .B2(n12821), .ZN(
        n11694) );
  OR2_X2 U14162 ( .A1(n11697), .A2(n11698), .ZN(n11742) );
  INV_X1 U14163 ( .A(n11742), .ZN(n11696) );
  AOI21_X1 U14164 ( .B1(n11698), .B2(n11697), .A(n11696), .ZN(n11706) );
  INV_X1 U14165 ( .A(n11699), .ZN(n11849) );
  NOR2_X1 U14166 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11700), .ZN(n15459) );
  NOR2_X1 U14167 ( .A1(n12576), .A2(n15472), .ZN(n11701) );
  AOI211_X1 U14168 ( .C1(n12574), .C2(n14852), .A(n15459), .B(n11701), .ZN(
        n11702) );
  OAI21_X1 U14169 ( .B1(n12581), .B2(n11703), .A(n11702), .ZN(n11704) );
  AOI21_X1 U14170 ( .B1(n11849), .B2(n12578), .A(n11704), .ZN(n11705) );
  OAI21_X1 U14171 ( .B1(n11706), .B2(n12592), .A(n11705), .ZN(P3_U3171) );
  XNOR2_X1 U14172 ( .A(n11707), .B(n12690), .ZN(n15555) );
  NAND2_X1 U14173 ( .A1(n15555), .A2(n15495), .ZN(n11715) );
  NAND2_X1 U14174 ( .A1(n11708), .A2(n12690), .ZN(n11709) );
  NAND2_X1 U14175 ( .A1(n11841), .A2(n11709), .ZN(n11713) );
  NAND2_X1 U14176 ( .A1(n12822), .A2(n14851), .ZN(n11711) );
  NAND2_X1 U14177 ( .A1(n12820), .A2(n14853), .ZN(n11710) );
  NAND2_X1 U14178 ( .A1(n11711), .A2(n11710), .ZN(n11712) );
  AOI21_X1 U14179 ( .B1(n11713), .B2(n15511), .A(n11712), .ZN(n11714) );
  AND2_X1 U14180 ( .A1(n11715), .A2(n11714), .ZN(n15557) );
  INV_X1 U14181 ( .A(n12290), .ZN(n15518) );
  NOR2_X1 U14182 ( .A1(n11824), .A2(n15545), .ZN(n15554) );
  AOI22_X1 U14183 ( .A1(n14860), .A2(n15554), .B1(n15517), .B2(n11826), .ZN(
        n11716) );
  OAI21_X1 U14184 ( .B1(n11310), .B2(n15501), .A(n11716), .ZN(n11717) );
  AOI21_X1 U14185 ( .B1(n15555), .B2(n15518), .A(n11717), .ZN(n11718) );
  OAI21_X1 U14186 ( .B1(n15557), .B2(n13166), .A(n11718), .ZN(P3_U3225) );
  INV_X1 U14187 ( .A(n14759), .ZN(n11720) );
  OAI222_X1 U14188 ( .A1(n13844), .A2(n11721), .B1(n13850), .B2(n11720), .C1(
        n11719), .C2(P2_U3088), .ZN(P2_U3307) );
  NAND2_X1 U14189 ( .A1(n10115), .A2(n11723), .ZN(n11724) );
  XNOR2_X1 U14190 ( .A(n11725), .B(n11724), .ZN(n11730) );
  OAI21_X1 U14191 ( .B1(n13390), .B2(n12119), .A(n11726), .ZN(n11728) );
  OAI22_X1 U14192 ( .A1(n13389), .A2(n11907), .B1(n11911), .B2(n13406), .ZN(
        n11727) );
  AOI211_X1 U14193 ( .C1(n11917), .C2(n13425), .A(n11728), .B(n11727), .ZN(
        n11729) );
  OAI21_X1 U14194 ( .B1(n11730), .B2(n13417), .A(n11729), .ZN(P2_U3196) );
  INV_X2 U14195 ( .A(n15371), .ZN(n13815) );
  AOI21_X1 U14196 ( .B1(n15356), .B2(n11803), .A(n11731), .ZN(n11732) );
  OAI211_X1 U14197 ( .C1(n13756), .C2(n11734), .A(n11733), .B(n11732), .ZN(
        n11736) );
  NAND2_X1 U14198 ( .A1(n11736), .A2(n13815), .ZN(n11735) );
  OAI21_X1 U14199 ( .B1(n13815), .B2(n10867), .A(n11735), .ZN(P2_U3509) );
  NAND2_X1 U14200 ( .A1(n11736), .A2(n15364), .ZN(n11737) );
  OAI21_X1 U14201 ( .B1(n15364), .B2(n7953), .A(n11737), .ZN(P2_U3460) );
  INV_X1 U14202 ( .A(n11738), .ZN(n11739) );
  INV_X1 U14203 ( .A(n12820), .ZN(n11821) );
  NAND2_X1 U14204 ( .A1(n11739), .A2(n11821), .ZN(n11740) );
  AND2_X1 U14205 ( .A1(n11742), .A2(n11740), .ZN(n11744) );
  XNOR2_X1 U14206 ( .A(n12469), .B(n11748), .ZN(n11992) );
  XNOR2_X1 U14207 ( .A(n11992), .B(n14852), .ZN(n11743) );
  AND2_X1 U14208 ( .A1(n11743), .A2(n11740), .ZN(n11741) );
  NAND2_X2 U14209 ( .A1(n11742), .A2(n11741), .ZN(n11995) );
  OAI211_X1 U14210 ( .C1(n11744), .C2(n11743), .A(n12572), .B(n11995), .ZN(
        n11750) );
  AOI21_X1 U14211 ( .B1(n12574), .B2(n12819), .A(n11745), .ZN(n11746) );
  OAI21_X1 U14212 ( .B1(n11821), .B2(n12576), .A(n11746), .ZN(n11747) );
  AOI21_X1 U14213 ( .B1(n12590), .B2(n11748), .A(n11747), .ZN(n11749) );
  OAI211_X1 U14214 ( .C1(n11985), .C2(n12588), .A(n11750), .B(n11749), .ZN(
        P3_U3157) );
  XNOR2_X1 U14215 ( .A(n11752), .B(n11751), .ZN(n14792) );
  XNOR2_X1 U14216 ( .A(n11753), .B(n11754), .ZN(n11756) );
  OAI22_X1 U14217 ( .A1(n14911), .A2(n14220), .B1(n12230), .B2(n14265), .ZN(
        n11755) );
  AOI21_X1 U14218 ( .B1(n11756), .B2(n15098), .A(n11755), .ZN(n11757) );
  OAI21_X1 U14219 ( .B1(n14792), .B2(n11758), .A(n11757), .ZN(n14795) );
  NAND2_X1 U14220 ( .A1(n14795), .A2(n14804), .ZN(n11764) );
  OAI22_X1 U14221 ( .A1(n14804), .A2(n11023), .B1(n12231), .B2(n14801), .ZN(
        n11762) );
  INV_X1 U14222 ( .A(n11759), .ZN(n11760) );
  OAI211_X1 U14223 ( .C1(n11760), .C2(n14794), .A(n15111), .B(n14814), .ZN(
        n14793) );
  NOR2_X1 U14224 ( .A1(n14793), .A2(n14816), .ZN(n11761) );
  AOI211_X1 U14225 ( .C1(n14255), .C2(n12227), .A(n11762), .B(n11761), .ZN(
        n11763) );
  OAI211_X1 U14226 ( .C1(n14792), .C2(n11765), .A(n11764), .B(n11763), .ZN(
        P1_U3281) );
  NAND2_X1 U14227 ( .A1(n11766), .A2(n11768), .ZN(n11769) );
  NAND2_X1 U14228 ( .A1(n11770), .A2(n11769), .ZN(n11776) );
  NOR2_X1 U14229 ( .A1(n10229), .A2(n11771), .ZN(n11772) );
  AOI21_X1 U14230 ( .B1(n11773), .B2(n12404), .A(n11772), .ZN(n11868) );
  AOI22_X1 U14231 ( .A1(n11773), .A2(n10208), .B1(n12409), .B2(n13961), .ZN(
        n11774) );
  XNOR2_X1 U14232 ( .A(n11774), .B(n10223), .ZN(n11867) );
  XOR2_X1 U14233 ( .A(n11868), .B(n11867), .Z(n11775) );
  OAI211_X1 U14234 ( .C1(n11776), .C2(n11775), .A(n11872), .B(n14960), .ZN(
        n11780) );
  INV_X1 U14235 ( .A(n11777), .ZN(n15086) );
  AOI22_X1 U14236 ( .A1(n14812), .A2(n13960), .B1(n14979), .B2(n13962), .ZN(
        n15082) );
  OAI22_X1 U14237 ( .A1(n13949), .A2(n15082), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8658), .ZN(n11778) );
  AOI21_X1 U14238 ( .B1(n13939), .B2(n15086), .A(n11778), .ZN(n11779) );
  OAI211_X1 U14239 ( .C1(n15171), .C2(n14958), .A(n11780), .B(n11779), .ZN(
        P1_U3213) );
  INV_X1 U14240 ( .A(n13397), .ZN(n13361) );
  OAI22_X1 U14241 ( .A1(n11785), .A2(n13661), .B1(n11781), .B2(n13663), .ZN(
        n11808) );
  AOI21_X1 U14242 ( .B1(n13361), .B2(n11808), .A(n11782), .ZN(n11783) );
  OAI21_X1 U14243 ( .B1(n15287), .B2(n13406), .A(n11783), .ZN(n11791) );
  INV_X1 U14244 ( .A(n11784), .ZN(n11798) );
  NOR3_X1 U14245 ( .A1(n11786), .A2(n11785), .A3(n13408), .ZN(n11787) );
  AOI21_X1 U14246 ( .B1(n11798), .B2(n10187), .A(n11787), .ZN(n11789) );
  NOR2_X1 U14247 ( .A1(n11789), .A2(n11788), .ZN(n11790) );
  AOI211_X1 U14248 ( .C1(n15286), .C2(n13425), .A(n11791), .B(n11790), .ZN(
        n11792) );
  OAI21_X1 U14249 ( .B1(n11793), .B2(n13417), .A(n11792), .ZN(P2_U3208) );
  INV_X1 U14250 ( .A(n11794), .ZN(n11795) );
  AOI22_X1 U14251 ( .A1(n13361), .A2(n11795), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11796) );
  OAI21_X1 U14252 ( .B1(n11797), .B2(n13406), .A(n11796), .ZN(n11802) );
  AOI211_X1 U14253 ( .C1(n11800), .C2(n11799), .A(n13417), .B(n11798), .ZN(
        n11801) );
  AOI211_X1 U14254 ( .C1(n11803), .C2(n13425), .A(n11802), .B(n11801), .ZN(
        n11804) );
  INV_X1 U14255 ( .A(n11804), .ZN(P2_U3189) );
  INV_X1 U14256 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11814) );
  XOR2_X1 U14257 ( .A(n11807), .B(n11805), .Z(n15294) );
  XNOR2_X1 U14258 ( .A(n11806), .B(n11807), .ZN(n11809) );
  AOI21_X1 U14259 ( .B1(n11809), .B2(n13586), .A(n11808), .ZN(n15300) );
  INV_X1 U14260 ( .A(n11810), .ZN(n11914) );
  AOI211_X1 U14261 ( .C1(n15286), .C2(n11811), .A(n10861), .B(n11914), .ZN(
        n15298) );
  AOI21_X1 U14262 ( .B1(n15356), .B2(n15286), .A(n15298), .ZN(n11812) );
  OAI211_X1 U14263 ( .C1(n15294), .C2(n15360), .A(n15300), .B(n11812), .ZN(
        n11815) );
  NAND2_X1 U14264 ( .A1(n11815), .A2(n13815), .ZN(n11813) );
  OAI21_X1 U14265 ( .B1(n13815), .B2(n11814), .A(n11813), .ZN(P2_U3510) );
  NAND2_X1 U14266 ( .A1(n11815), .A2(n15364), .ZN(n11816) );
  OAI21_X1 U14267 ( .B1(n15364), .B2(n7980), .A(n11816), .ZN(P2_U3463) );
  MUX2_X1 U14268 ( .A(n11818), .B(n12822), .S(n11817), .Z(n11820) );
  XNOR2_X1 U14269 ( .A(n11820), .B(n11819), .ZN(n11828) );
  NOR2_X1 U14270 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9659), .ZN(n15438) );
  NOR2_X1 U14271 ( .A1(n12584), .A2(n11821), .ZN(n11822) );
  AOI211_X1 U14272 ( .C1(n12586), .C2(n12822), .A(n15438), .B(n11822), .ZN(
        n11823) );
  OAI21_X1 U14273 ( .B1(n11824), .B2(n12581), .A(n11823), .ZN(n11825) );
  AOI21_X1 U14274 ( .B1(n11826), .B2(n12578), .A(n11825), .ZN(n11827) );
  OAI21_X1 U14275 ( .B1(n11828), .B2(n12592), .A(n11827), .ZN(P3_U3161) );
  AOI222_X1 U14276 ( .A1(n11830), .A2(n13840), .B1(P1_DATAO_REG_22__SCAN_IN), 
        .B2(n12008), .C1(n11829), .C2(P2_STATE_REG_SCAN_IN), .ZN(n11831) );
  INV_X1 U14277 ( .A(n11831), .ZN(P2_U3305) );
  INV_X1 U14278 ( .A(n11832), .ZN(n11836) );
  INV_X1 U14279 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11833) );
  OAI222_X1 U14280 ( .A1(P1_U3086), .A2(n11834), .B1(n14398), .B2(n11836), 
        .C1(n11833), .C2(n14395), .ZN(P1_U3334) );
  OAI222_X1 U14281 ( .A1(n13852), .A2(n11837), .B1(n13850), .B2(n11836), .C1(
        n11835), .C2(P2_U3088), .ZN(P2_U3306) );
  XNOR2_X1 U14282 ( .A(n11838), .B(n12696), .ZN(n15560) );
  INV_X1 U14283 ( .A(n11839), .ZN(n11840) );
  NAND2_X1 U14284 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  NAND2_X1 U14285 ( .A1(n11842), .A2(n12696), .ZN(n11844) );
  NAND3_X1 U14286 ( .A1(n11844), .A2(n15511), .A3(n11843), .ZN(n11846) );
  AOI22_X1 U14287 ( .A1(n14851), .A2(n12821), .B1(n14852), .B2(n14853), .ZN(
        n11845) );
  NAND2_X1 U14288 ( .A1(n11846), .A2(n11845), .ZN(n11847) );
  AOI21_X1 U14289 ( .B1(n15560), .B2(n15495), .A(n11847), .ZN(n15562) );
  AND2_X1 U14290 ( .A1(n12698), .A2(n11848), .ZN(n15559) );
  AOI22_X1 U14291 ( .A1(n14860), .A2(n15559), .B1(n15517), .B2(n11849), .ZN(
        n11850) );
  OAI21_X1 U14292 ( .B1(n11851), .B2(n15501), .A(n11850), .ZN(n11852) );
  AOI21_X1 U14293 ( .B1(n15560), .B2(n15518), .A(n11852), .ZN(n11853) );
  OAI21_X1 U14294 ( .B1(n15562), .B2(n13166), .A(n11853), .ZN(P3_U3224) );
  OR2_X1 U14295 ( .A1(n11854), .A2(n12671), .ZN(n11855) );
  NAND2_X1 U14296 ( .A1(n11856), .A2(n11855), .ZN(n15537) );
  OAI22_X1 U14297 ( .A1(n13163), .A2(n15534), .B1(n11857), .B2(n15479), .ZN(
        n11864) );
  XNOR2_X1 U14298 ( .A(n11858), .B(n12630), .ZN(n11862) );
  NAND2_X1 U14299 ( .A1(n15537), .A2(n15495), .ZN(n11861) );
  AOI22_X1 U14300 ( .A1(n14851), .A2(n12825), .B1(n11859), .B2(n14853), .ZN(
        n11860) );
  OAI211_X1 U14301 ( .C1(n15490), .C2(n11862), .A(n11861), .B(n11860), .ZN(
        n15535) );
  MUX2_X1 U14302 ( .A(n15535), .B(P3_REG2_REG_4__SCAN_IN), .S(n13166), .Z(
        n11863) );
  AOI211_X1 U14303 ( .C1(n15518), .C2(n15537), .A(n11864), .B(n11863), .ZN(
        n11865) );
  INV_X1 U14304 ( .A(n11865), .ZN(P3_U3229) );
  AOI22_X1 U14305 ( .A1(n15177), .A2(n10208), .B1(n12409), .B2(n13960), .ZN(
        n11866) );
  XNOR2_X1 U14306 ( .A(n11866), .B(n10223), .ZN(n12023) );
  AOI22_X1 U14307 ( .A1(n15177), .A2(n12409), .B1(n12408), .B2(n13960), .ZN(
        n12022) );
  XNOR2_X1 U14308 ( .A(n12023), .B(n12022), .ZN(n11874) );
  INV_X1 U14309 ( .A(n11867), .ZN(n11870) );
  INV_X1 U14310 ( .A(n11868), .ZN(n11869) );
  AOI21_X1 U14311 ( .B1(n11874), .B2(n11873), .A(n6820), .ZN(n11880) );
  INV_X1 U14312 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n14004) );
  OAI22_X1 U14313 ( .A1(n13949), .A2(n11875), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14004), .ZN(n11878) );
  NOR2_X1 U14314 ( .A1(n14964), .A2(n11876), .ZN(n11877) );
  AOI211_X1 U14315 ( .C1(n14921), .C2(n15177), .A(n11878), .B(n11877), .ZN(
        n11879) );
  OAI21_X1 U14316 ( .B1(n11880), .B2(n14916), .A(n11879), .ZN(P1_U3221) );
  INV_X1 U14317 ( .A(n11881), .ZN(n11882) );
  OAI222_X1 U14318 ( .A1(n11883), .A2(P3_U3151), .B1(n12306), .B2(n11882), 
        .C1(n14664), .C2(n12423), .ZN(P3_U3270) );
  XNOR2_X1 U14319 ( .A(n11885), .B(n11884), .ZN(n11892) );
  INV_X1 U14320 ( .A(n12038), .ZN(n11889) );
  NAND2_X1 U14321 ( .A1(n13442), .A2(n13607), .ZN(n11887) );
  NAND2_X1 U14322 ( .A1(n13440), .A2(n13604), .ZN(n11886) );
  NAND2_X1 U14323 ( .A1(n11887), .A2(n11886), .ZN(n12044) );
  AOI22_X1 U14324 ( .A1(n13361), .A2(n12044), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11888) );
  OAI21_X1 U14325 ( .B1(n11889), .B2(n13406), .A(n11888), .ZN(n11890) );
  AOI21_X1 U14326 ( .B1(n12039), .B2(n13425), .A(n11890), .ZN(n11891) );
  OAI21_X1 U14327 ( .B1(n11892), .B2(n13417), .A(n11891), .ZN(P2_U3206) );
  NAND2_X1 U14328 ( .A1(n11897), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11893) );
  NAND2_X1 U14329 ( .A1(n11894), .A2(n11893), .ZN(n13452) );
  XNOR2_X1 U14330 ( .A(n13452), .B(n13467), .ZN(n13454) );
  XOR2_X1 U14331 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n13454), .Z(n11903) );
  AND2_X1 U14332 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n12019) );
  AOI21_X1 U14333 ( .B1(n15281), .B2(n13467), .A(n12019), .ZN(n11895) );
  INV_X1 U14334 ( .A(n11895), .ZN(n11901) );
  XNOR2_X1 U14335 ( .A(n13467), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11898) );
  AOI211_X1 U14336 ( .C1(n11899), .C2(n11898), .A(n15271), .B(n13466), .ZN(
        n11900) );
  AOI211_X1 U14337 ( .C1(n15275), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n11901), 
        .B(n11900), .ZN(n11902) );
  OAI21_X1 U14338 ( .B1(n11903), .B2(n13489), .A(n11902), .ZN(P2_U3228) );
  XNOR2_X1 U14339 ( .A(n11904), .B(n11906), .ZN(n14899) );
  XOR2_X1 U14340 ( .A(n11905), .B(n11906), .Z(n11909) );
  OAI22_X1 U14341 ( .A1(n11907), .A2(n13661), .B1(n12119), .B2(n13663), .ZN(
        n11908) );
  AOI21_X1 U14342 ( .B1(n11909), .B2(n13705), .A(n11908), .ZN(n11910) );
  OAI21_X1 U14343 ( .B1(n14899), .B2(n10061), .A(n11910), .ZN(n14902) );
  NAND2_X1 U14344 ( .A1(n14902), .A2(n13689), .ZN(n11919) );
  OAI22_X1 U14345 ( .A1(n13689), .A2(n11912), .B1(n11911), .B2(n13683), .ZN(
        n11916) );
  INV_X1 U14346 ( .A(n11917), .ZN(n14901) );
  INV_X1 U14347 ( .A(n12037), .ZN(n11913) );
  OAI211_X1 U14348 ( .C1(n14901), .C2(n11914), .A(n11913), .B(n10146), .ZN(
        n14900) );
  NOR2_X1 U14349 ( .A1(n14900), .A2(n13519), .ZN(n11915) );
  AOI211_X1 U14350 ( .C1(n13685), .C2(n11917), .A(n11916), .B(n11915), .ZN(
        n11918) );
  OAI211_X1 U14351 ( .C1(n14899), .C2(n13618), .A(n11919), .B(n11918), .ZN(
        P2_U3253) );
  INV_X1 U14352 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11920) );
  MUX2_X1 U14353 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n11920), .S(n12060), .Z(
        n11925) );
  AOI21_X1 U14354 ( .B1(n11922), .B2(n11927), .A(n11921), .ZN(n11923) );
  XOR2_X1 U14355 ( .A(n11928), .B(n11923), .Z(n15051) );
  INV_X1 U14356 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15050) );
  NAND2_X1 U14357 ( .A1(n15051), .A2(n15050), .ZN(n15049) );
  AOI211_X1 U14358 ( .C1(n11925), .C2(n11924), .A(n12065), .B(n12063), .ZN(
        n11936) );
  OAI21_X1 U14359 ( .B1(n11344), .B2(n11927), .A(n11926), .ZN(n11929) );
  NOR2_X1 U14360 ( .A1(n11929), .A2(n11928), .ZN(n11931) );
  XNOR2_X1 U14361 ( .A(n11929), .B(n11928), .ZN(n15053) );
  NOR2_X1 U14362 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15053), .ZN(n15052) );
  INV_X1 U14363 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12061) );
  MUX2_X1 U14364 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n12061), .S(n12060), .Z(
        n11930) );
  OAI21_X1 U14365 ( .B1(n11931), .B2(n15052), .A(n11930), .ZN(n11932) );
  AND3_X1 U14366 ( .A1(n11932), .A2(n15044), .A3(n12059), .ZN(n11935) );
  NAND2_X1 U14367 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13898)
         );
  NAND2_X1 U14368 ( .A1(n15031), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n11933) );
  OAI211_X1 U14369 ( .C1(n15054), .C2(n12060), .A(n13898), .B(n11933), .ZN(
        n11934) );
  OR3_X1 U14370 ( .A1(n11936), .A2(n11935), .A3(n11934), .ZN(P1_U3259) );
  OAI211_X1 U14371 ( .C1(n11938), .C2(n11944), .A(n11937), .B(n15098), .ZN(
        n11940) );
  AOI22_X1 U14372 ( .A1(n13957), .A2(n14812), .B1(n14979), .B2(n13958), .ZN(
        n11939) );
  NAND2_X1 U14373 ( .A1(n11940), .A2(n11939), .ZN(n14976) );
  AOI21_X1 U14374 ( .B1(n14971), .B2(n14815), .A(n15125), .ZN(n11941) );
  NAND2_X1 U14375 ( .A1(n11941), .A2(n12088), .ZN(n14974) );
  OR2_X1 U14376 ( .A1(n15118), .A2(n11942), .ZN(n14164) );
  NAND2_X1 U14377 ( .A1(n11943), .A2(n11944), .ZN(n14972) );
  NAND3_X1 U14378 ( .A1(n14973), .A2(n14972), .A3(n14809), .ZN(n11948) );
  NAND2_X1 U14379 ( .A1(n15105), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11945) );
  OAI21_X1 U14380 ( .B1(n14801), .B2(n14924), .A(n11945), .ZN(n11946) );
  AOI21_X1 U14381 ( .B1(n14971), .B2(n14255), .A(n11946), .ZN(n11947) );
  OAI211_X1 U14382 ( .C1(n14974), .C2(n14164), .A(n11948), .B(n11947), .ZN(
        n11949) );
  AOI21_X1 U14383 ( .B1(n14804), .B2(n14976), .A(n11949), .ZN(n11950) );
  INV_X1 U14384 ( .A(n11950), .ZN(P1_U3279) );
  AOI21_X1 U14385 ( .B1(n11954), .B2(n9759), .A(n12844), .ZN(n11972) );
  NAND2_X1 U14386 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11958), .ZN(n11956) );
  NAND2_X1 U14387 ( .A1(n11956), .A2(n11955), .ZN(n12837) );
  XNOR2_X1 U14388 ( .A(n12837), .B(n12828), .ZN(n11957) );
  NAND2_X1 U14389 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11957), .ZN(n12838) );
  OAI21_X1 U14390 ( .B1(n11957), .B2(P3_REG1_REG_13__SCAN_IN), .A(n12838), 
        .ZN(n11970) );
  MUX2_X1 U14391 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12913), .Z(n12827) );
  XNOR2_X1 U14392 ( .A(n12827), .B(n12828), .ZN(n11961) );
  NAND2_X1 U14393 ( .A1(n11959), .A2(n11958), .ZN(n11962) );
  AND2_X1 U14394 ( .A1(n11961), .A2(n11962), .ZN(n11960) );
  NAND2_X1 U14395 ( .A1(n11963), .A2(n11960), .ZN(n12835) );
  INV_X1 U14396 ( .A(n12835), .ZN(n11965) );
  AOI21_X1 U14397 ( .B1(n11963), .B2(n11962), .A(n11961), .ZN(n11964) );
  OAI21_X1 U14398 ( .B1(n11965), .B2(n11964), .A(n12954), .ZN(n11968) );
  NOR2_X1 U14399 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11966), .ZN(n12145) );
  AOI21_X1 U14400 ( .B1(n15460), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12145), 
        .ZN(n11967) );
  OAI211_X1 U14401 ( .C1(n15454), .C2(n12836), .A(n11968), .B(n11967), .ZN(
        n11969) );
  AOI21_X1 U14402 ( .B1(n11970), .B2(n15463), .A(n11969), .ZN(n11971) );
  OAI21_X1 U14403 ( .B1(n11972), .B2(n15467), .A(n11971), .ZN(P3_U3195) );
  INV_X1 U14404 ( .A(n11973), .ZN(n11974) );
  OAI222_X1 U14405 ( .A1(P3_U3151), .A2(n11976), .B1(n12423), .B2(n11975), 
        .C1(n12306), .C2(n11974), .ZN(P3_U3269) );
  XNOR2_X1 U14406 ( .A(n11977), .B(n12701), .ZN(n11983) );
  INV_X1 U14407 ( .A(n11978), .ZN(n11979) );
  AOI21_X1 U14408 ( .B1(n11980), .B2(n12701), .A(n11979), .ZN(n15567) );
  NAND2_X1 U14409 ( .A1(n15567), .A2(n15495), .ZN(n11982) );
  AOI22_X1 U14410 ( .A1(n14851), .A2(n12820), .B1(n12819), .B2(n14853), .ZN(
        n11981) );
  OAI211_X1 U14411 ( .C1(n15490), .C2(n11983), .A(n11982), .B(n11981), .ZN(
        n15564) );
  INV_X1 U14412 ( .A(n15564), .ZN(n11991) );
  NOR2_X1 U14413 ( .A1(n11984), .A2(n15545), .ZN(n15565) );
  INV_X1 U14414 ( .A(n11985), .ZN(n11986) );
  AOI22_X1 U14415 ( .A1(n14860), .A2(n15565), .B1(n15517), .B2(n11986), .ZN(
        n11987) );
  OAI21_X1 U14416 ( .B1(n11988), .B2(n15501), .A(n11987), .ZN(n11989) );
  AOI21_X1 U14417 ( .B1(n15567), .B2(n15518), .A(n11989), .ZN(n11990) );
  OAI21_X1 U14418 ( .B1(n11991), .B2(n13166), .A(n11990), .ZN(P3_U3223) );
  INV_X1 U14419 ( .A(n11992), .ZN(n11993) );
  NAND2_X1 U14420 ( .A1(n11993), .A2(n14852), .ZN(n11994) );
  XNOR2_X1 U14421 ( .A(n12466), .B(n11996), .ZN(n11997) );
  INV_X1 U14422 ( .A(n11997), .ZN(n11998) );
  INV_X1 U14423 ( .A(n12050), .ZN(n11999) );
  AOI21_X1 U14424 ( .B1(n12819), .B2(n12000), .A(n11999), .ZN(n12006) );
  INV_X1 U14425 ( .A(n14854), .ZN(n12143) );
  NOR2_X1 U14426 ( .A1(n12584), .A2(n12143), .ZN(n12001) );
  AOI211_X1 U14427 ( .C1(n12586), .C2(n14852), .A(n12002), .B(n12001), .ZN(
        n12003) );
  OAI21_X1 U14428 ( .B1(n12581), .B2(n14859), .A(n12003), .ZN(n12004) );
  AOI21_X1 U14429 ( .B1(n14856), .B2(n12578), .A(n12004), .ZN(n12005) );
  OAI21_X1 U14430 ( .B1(n12006), .B2(n12592), .A(n12005), .ZN(P3_U3176) );
  INV_X1 U14431 ( .A(n12007), .ZN(n12013) );
  NAND2_X1 U14432 ( .A1(n12008), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12010) );
  OAI211_X1 U14433 ( .C1(n12013), .C2(n13850), .A(n12010), .B(n12009), .ZN(
        P2_U3304) );
  NAND2_X1 U14434 ( .A1(n14756), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12012) );
  OAI211_X1 U14435 ( .C1(n12013), .C2(n14383), .A(n12012), .B(n12011), .ZN(
        P1_U3332) );
  INV_X1 U14436 ( .A(n13811), .ZN(n12125) );
  OAI21_X1 U14437 ( .B1(n12016), .B2(n12015), .A(n12014), .ZN(n12017) );
  NAND2_X1 U14438 ( .A1(n12017), .A2(n10187), .ZN(n12021) );
  OAI22_X1 U14439 ( .A1(n13389), .A2(n12119), .B1(n12121), .B2(n13406), .ZN(
        n12018) );
  AOI211_X1 U14440 ( .C1(n13422), .C2(n13439), .A(n12019), .B(n12018), .ZN(
        n12020) );
  OAI211_X1 U14441 ( .C1(n12125), .C2(n13369), .A(n12021), .B(n12020), .ZN(
        P2_U3187) );
  NAND2_X1 U14442 ( .A1(n12029), .A2(n10208), .ZN(n12025) );
  NAND2_X1 U14443 ( .A1(n12409), .A2(n14927), .ZN(n12024) );
  NAND2_X1 U14444 ( .A1(n12025), .A2(n12024), .ZN(n12026) );
  XNOR2_X1 U14445 ( .A(n12026), .B(n10223), .ZN(n12205) );
  NOR2_X1 U14446 ( .A1(n10229), .A2(n12027), .ZN(n12028) );
  AOI21_X1 U14447 ( .B1(n12029), .B2(n12404), .A(n12028), .ZN(n12206) );
  XNOR2_X1 U14448 ( .A(n12205), .B(n12206), .ZN(n12030) );
  NAND2_X1 U14449 ( .A1(n12031), .A2(n12030), .ZN(n12208) );
  OAI211_X1 U14450 ( .C1(n12031), .C2(n12030), .A(n12208), .B(n14960), .ZN(
        n12035) );
  INV_X1 U14451 ( .A(n12032), .ZN(n15071) );
  AOI22_X1 U14452 ( .A1(n14812), .A2(n14943), .B1(n14979), .B2(n13960), .ZN(
        n15068) );
  OAI22_X1 U14453 ( .A1(n13949), .A2(n15068), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8688), .ZN(n12033) );
  AOI21_X1 U14454 ( .B1(n13939), .B2(n15071), .A(n12033), .ZN(n12034) );
  OAI211_X1 U14455 ( .C1(n7364), .C2(n14958), .A(n12035), .B(n12034), .ZN(
        P1_U3231) );
  XNOR2_X1 U14456 ( .A(n12036), .B(n12043), .ZN(n14898) );
  OAI211_X1 U14457 ( .C1(n14896), .C2(n12037), .A(n10146), .B(n12120), .ZN(
        n14894) );
  AOI22_X1 U14458 ( .A1(n15290), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12038), 
        .B2(n15288), .ZN(n12041) );
  NAND2_X1 U14459 ( .A1(n12039), .A2(n13685), .ZN(n12040) );
  OAI211_X1 U14460 ( .C1(n14894), .C2(n13519), .A(n12041), .B(n12040), .ZN(
        n12047) );
  XOR2_X1 U14461 ( .A(n12043), .B(n12042), .Z(n12045) );
  AOI21_X1 U14462 ( .B1(n12045), .B2(n13705), .A(n12044), .ZN(n14895) );
  NOR2_X1 U14463 ( .A1(n14895), .A2(n15301), .ZN(n12046) );
  AOI211_X1 U14464 ( .C1(n14898), .C2(n13652), .A(n12047), .B(n12046), .ZN(
        n12048) );
  INV_X1 U14465 ( .A(n12048), .ZN(P2_U3252) );
  XNOR2_X1 U14466 ( .A(n12466), .B(n12056), .ZN(n12139) );
  XNOR2_X1 U14467 ( .A(n12139), .B(n12143), .ZN(n12051) );
  XNOR2_X1 U14468 ( .A(n12141), .B(n12051), .ZN(n12058) );
  AOI21_X1 U14469 ( .B1(n12574), .B2(n12818), .A(n12052), .ZN(n12053) );
  OAI21_X1 U14470 ( .B1(n7242), .B2(n12576), .A(n12053), .ZN(n12055) );
  NOR2_X1 U14471 ( .A1(n12588), .A2(n12080), .ZN(n12054) );
  AOI211_X1 U14472 ( .C1(n12056), .C2(n12590), .A(n12055), .B(n12054), .ZN(
        n12057) );
  OAI21_X1 U14473 ( .B1(n12058), .B2(n12592), .A(n12057), .ZN(P3_U3164) );
  OAI21_X1 U14474 ( .B1(n12061), .B2(n12060), .A(n12059), .ZN(n14021) );
  INV_X1 U14475 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14024) );
  MUX2_X1 U14476 ( .A(n14024), .B(P1_REG2_REG_17__SCAN_IN), .S(n14027), .Z(
        n14019) );
  XNOR2_X1 U14477 ( .A(n14021), .B(n14019), .ZN(n12070) );
  NAND2_X1 U14478 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13906)
         );
  NAND2_X1 U14479 ( .A1(n15031), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n12062) );
  OAI211_X1 U14480 ( .C1(n15054), .C2(n14023), .A(n13906), .B(n12062), .ZN(
        n12069) );
  AOI21_X1 U14481 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n12064), .A(n12063), 
        .ZN(n12067) );
  XNOR2_X1 U14482 ( .A(n14027), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n12066) );
  NOR2_X1 U14483 ( .A1(n12067), .A2(n12066), .ZN(n14026) );
  AOI211_X1 U14484 ( .C1(n12067), .C2(n12066), .A(n12065), .B(n14026), .ZN(
        n12068) );
  AOI211_X1 U14485 ( .C1(n15044), .C2(n12070), .A(n12069), .B(n12068), .ZN(
        n12071) );
  INV_X1 U14486 ( .A(n12071), .ZN(P1_U3260) );
  OAI211_X1 U14487 ( .C1(n12074), .C2(n12073), .A(n12072), .B(n15511), .ZN(
        n12076) );
  AOI22_X1 U14488 ( .A1(n14851), .A2(n12819), .B1(n12818), .B2(n14853), .ZN(
        n12075) );
  NAND2_X1 U14489 ( .A1(n12076), .A2(n12075), .ZN(n14876) );
  INV_X1 U14490 ( .A(n14876), .ZN(n12085) );
  XNOR2_X1 U14491 ( .A(n12077), .B(n7340), .ZN(n14878) );
  OR2_X1 U14492 ( .A1(n15495), .A2(n15498), .ZN(n12078) );
  NAND2_X1 U14493 ( .A1(n14878), .A2(n14861), .ZN(n12084) );
  NOR2_X1 U14494 ( .A1(n12079), .A2(n15545), .ZN(n14877) );
  INV_X1 U14495 ( .A(n14877), .ZN(n12081) );
  OAI22_X1 U14496 ( .A1(n15482), .A2(n12081), .B1(n12080), .B2(n15479), .ZN(
        n12082) );
  AOI21_X1 U14497 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n13166), .A(n12082), 
        .ZN(n12083) );
  OAI211_X1 U14498 ( .C1(n12085), .C2(n13166), .A(n12084), .B(n12083), .ZN(
        P3_U3221) );
  XNOR2_X1 U14499 ( .A(n12086), .B(n12092), .ZN(n12087) );
  AOI222_X1 U14500 ( .A1(n15098), .A2(n12087), .B1(n14953), .B2(n14812), .C1(
        n14955), .C2(n14979), .ZN(n14357) );
  AND2_X1 U14501 ( .A1(n14354), .A2(n12088), .ZN(n12089) );
  NOR2_X1 U14502 ( .A1(n6808), .A2(n12089), .ZN(n14355) );
  INV_X1 U14503 ( .A(n12251), .ZN(n14260) );
  INV_X1 U14504 ( .A(n14963), .ZN(n12090) );
  AOI22_X1 U14505 ( .A1(n15105), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n12090), 
        .B2(n15103), .ZN(n12091) );
  OAI21_X1 U14506 ( .B1(n6955), .B2(n15107), .A(n12091), .ZN(n12095) );
  XNOR2_X1 U14507 ( .A(n12093), .B(n12092), .ZN(n14358) );
  NOR2_X1 U14508 ( .A1(n14358), .A2(n14210), .ZN(n12094) );
  AOI211_X1 U14509 ( .C1(n14355), .C2(n14260), .A(n12095), .B(n12094), .ZN(
        n12096) );
  OAI21_X1 U14510 ( .B1(n14251), .B2(n14357), .A(n12096), .ZN(P1_U3278) );
  XNOR2_X1 U14511 ( .A(n12097), .B(n12098), .ZN(n14970) );
  INV_X1 U14512 ( .A(n14970), .ZN(n12109) );
  NAND2_X1 U14513 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  AOI21_X1 U14514 ( .B1(n12101), .B2(n12100), .A(n15083), .ZN(n14968) );
  AND2_X1 U14515 ( .A1(n13957), .A2(n14979), .ZN(n12102) );
  AOI21_X1 U14516 ( .B1(n14237), .B2(n14812), .A(n12102), .ZN(n14965) );
  INV_X1 U14517 ( .A(n14965), .ZN(n12103) );
  OAI21_X1 U14518 ( .B1(n14968), .B2(n12103), .A(n14804), .ZN(n12108) );
  OAI22_X1 U14519 ( .A1(n14804), .A2(n12061), .B1(n13899), .B2(n14801), .ZN(
        n12105) );
  OAI211_X1 U14520 ( .C1(n14967), .C2(n6808), .A(n15111), .B(n12131), .ZN(
        n14966) );
  NOR2_X1 U14521 ( .A1(n14966), .A2(n14816), .ZN(n12104) );
  AOI211_X1 U14522 ( .C1(n14255), .C2(n12106), .A(n12105), .B(n12104), .ZN(
        n12107) );
  OAI211_X1 U14523 ( .C1(n12109), .C2(n14210), .A(n12108), .B(n12107), .ZN(
        P1_U3277) );
  INV_X1 U14524 ( .A(n12110), .ZN(n12112) );
  OAI222_X1 U14525 ( .A1(n12306), .A2(n12112), .B1(n12423), .B2(n12111), .C1(
        P3_U3151), .C2(n9968), .ZN(P3_U3267) );
  XNOR2_X1 U14526 ( .A(n12113), .B(n12117), .ZN(n13813) );
  INV_X1 U14527 ( .A(n12114), .ZN(n12115) );
  AOI21_X1 U14528 ( .B1(n12117), .B2(n12116), .A(n12115), .ZN(n12118) );
  OAI222_X1 U14529 ( .A1(n13663), .A2(n13348), .B1(n13661), .B2(n12119), .C1(
        n13676), .C2(n12118), .ZN(n13809) );
  AOI211_X1 U14530 ( .C1(n13811), .C2(n12120), .A(n10861), .B(n7500), .ZN(
        n13810) );
  NAND2_X1 U14531 ( .A1(n13810), .A2(n15297), .ZN(n12124) );
  INV_X1 U14532 ( .A(n12121), .ZN(n12122) );
  AOI22_X1 U14533 ( .A1(n15290), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12122), 
        .B2(n15288), .ZN(n12123) );
  OAI211_X1 U14534 ( .C1(n12125), .C2(n15292), .A(n12124), .B(n12123), .ZN(
        n12126) );
  AOI21_X1 U14535 ( .B1(n13809), .B2(n13689), .A(n12126), .ZN(n12127) );
  OAI21_X1 U14536 ( .B1(n15293), .B2(n13813), .A(n12127), .ZN(P2_U3251) );
  XOR2_X1 U14537 ( .A(n12128), .B(n12129), .Z(n14353) );
  XNOR2_X1 U14538 ( .A(n12130), .B(n12129), .ZN(n14351) );
  INV_X1 U14539 ( .A(n12131), .ZN(n12132) );
  OAI211_X1 U14540 ( .C1(n14349), .C2(n12132), .A(n15111), .B(n14244), .ZN(
        n14348) );
  AOI22_X1 U14541 ( .A1(n14222), .A2(n14812), .B1(n14979), .B2(n14953), .ZN(
        n14347) );
  OAI21_X1 U14542 ( .B1(n13910), .B2(n14801), .A(n14347), .ZN(n12133) );
  MUX2_X1 U14543 ( .A(n12133), .B(P1_REG2_REG_17__SCAN_IN), .S(n14251), .Z(
        n12134) );
  AOI21_X1 U14544 ( .B1(n13912), .B2(n14255), .A(n12134), .ZN(n12135) );
  OAI21_X1 U14545 ( .B1(n14348), .B2(n14816), .A(n12135), .ZN(n12136) );
  AOI21_X1 U14546 ( .B1(n14351), .B2(n14182), .A(n12136), .ZN(n12137) );
  OAI21_X1 U14547 ( .B1(n14353), .B2(n14210), .A(n12137), .ZN(P1_U3276) );
  XNOR2_X1 U14548 ( .A(n14846), .B(n12469), .ZN(n12138) );
  OR2_X1 U14549 ( .A1(n12138), .A2(n13158), .ZN(n12180) );
  NAND2_X1 U14550 ( .A1(n12138), .A2(n13158), .ZN(n12178) );
  NAND2_X1 U14551 ( .A1(n12180), .A2(n12178), .ZN(n12142) );
  AND2_X1 U14552 ( .A1(n12139), .A2(n12143), .ZN(n12140) );
  XOR2_X1 U14553 ( .A(n12142), .B(n12179), .Z(n12150) );
  NOR2_X1 U14554 ( .A1(n12576), .A2(n12143), .ZN(n12144) );
  AOI211_X1 U14555 ( .C1(n12574), .C2(n14841), .A(n12145), .B(n12144), .ZN(
        n12146) );
  OAI21_X1 U14556 ( .B1(n12147), .B2(n12588), .A(n12146), .ZN(n12148) );
  AOI21_X1 U14557 ( .B1(n14846), .B2(n12590), .A(n12148), .ZN(n12149) );
  OAI21_X1 U14558 ( .B1(n12150), .B2(n12592), .A(n12149), .ZN(P3_U3174) );
  INV_X1 U14559 ( .A(n12151), .ZN(n12189) );
  AOI22_X1 U14560 ( .A1(n8978), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n14756), .ZN(n12152) );
  OAI21_X1 U14561 ( .B1(n12189), .B2(n14383), .A(n12152), .ZN(P1_U3331) );
  OAI211_X1 U14562 ( .C1(n12155), .C2(n12154), .A(n12153), .B(n13586), .ZN(
        n12157) );
  AOI22_X1 U14563 ( .A1(n13437), .A2(n13604), .B1(n13607), .B2(n13439), .ZN(
        n12156) );
  AND2_X1 U14564 ( .A1(n12157), .A2(n12156), .ZN(n13803) );
  AOI211_X1 U14565 ( .C1(n13798), .C2(n12171), .A(n10861), .B(n7498), .ZN(
        n13797) );
  INV_X1 U14566 ( .A(n13798), .ZN(n12158) );
  NOR2_X1 U14567 ( .A1(n12158), .A2(n15292), .ZN(n12160) );
  OAI22_X1 U14568 ( .A1(n13689), .A2(n13459), .B1(n13347), .B2(n13683), .ZN(
        n12159) );
  AOI211_X1 U14569 ( .C1(n13797), .C2(n15297), .A(n12160), .B(n12159), .ZN(
        n12164) );
  OR2_X1 U14570 ( .A1(n12162), .A2(n12161), .ZN(n13800) );
  NAND3_X1 U14571 ( .A1(n13800), .A2(n13799), .A3(n13652), .ZN(n12163) );
  OAI211_X1 U14572 ( .C1(n13803), .C2(n15301), .A(n12164), .B(n12163), .ZN(
        P2_U3249) );
  XNOR2_X1 U14573 ( .A(n12165), .B(n12167), .ZN(n13808) );
  OAI21_X1 U14574 ( .B1(n12168), .B2(n12167), .A(n12166), .ZN(n12169) );
  AOI222_X1 U14575 ( .A1(n13705), .A2(n12169), .B1(n13438), .B2(n13604), .C1(
        n13440), .C2(n13607), .ZN(n13807) );
  INV_X1 U14576 ( .A(n13807), .ZN(n12176) );
  AOI21_X1 U14577 ( .B1(n13805), .B2(n12170), .A(n10861), .ZN(n12172) );
  AND2_X1 U14578 ( .A1(n12172), .A2(n12171), .ZN(n13804) );
  NAND2_X1 U14579 ( .A1(n13804), .A2(n15297), .ZN(n12174) );
  AOI22_X1 U14580 ( .A1(n15290), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13423), 
        .B2(n15288), .ZN(n12173) );
  OAI211_X1 U14581 ( .C1(n7499), .C2(n15292), .A(n12174), .B(n12173), .ZN(
        n12175) );
  AOI21_X1 U14582 ( .B1(n12176), .B2(n13689), .A(n12175), .ZN(n12177) );
  OAI21_X1 U14583 ( .B1(n15293), .B2(n13808), .A(n12177), .ZN(P2_U3250) );
  XNOR2_X1 U14584 ( .A(n13284), .B(n12469), .ZN(n12428) );
  XNOR2_X1 U14585 ( .A(n12428), .B(n14841), .ZN(n12426) );
  XOR2_X1 U14586 ( .A(n12427), .B(n12426), .Z(n12186) );
  INV_X1 U14587 ( .A(n12181), .ZN(n13161) );
  NAND2_X1 U14588 ( .A1(n12586), .A2(n12818), .ZN(n12182) );
  NAND2_X1 U14589 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12850)
         );
  OAI211_X1 U14590 ( .C1(n13159), .C2(n12584), .A(n12182), .B(n12850), .ZN(
        n12184) );
  NOR2_X1 U14591 ( .A1(n12581), .A2(n13284), .ZN(n12183) );
  AOI211_X1 U14592 ( .C1(n13161), .C2(n12578), .A(n12184), .B(n12183), .ZN(
        n12185) );
  OAI21_X1 U14593 ( .B1(n12186), .B2(n12592), .A(n12185), .ZN(P3_U3155) );
  INV_X1 U14594 ( .A(n12187), .ZN(n12188) );
  OAI222_X1 U14595 ( .A1(n13852), .A2(n12190), .B1(n13850), .B2(n12189), .C1(
        n12188), .C2(P2_U3088), .ZN(P2_U3303) );
  XNOR2_X1 U14596 ( .A(n12192), .B(n12191), .ZN(n12195) );
  NAND2_X1 U14597 ( .A1(n13436), .A2(n13604), .ZN(n12194) );
  NAND2_X1 U14598 ( .A1(n13438), .A2(n13607), .ZN(n12193) );
  NAND2_X1 U14599 ( .A1(n12194), .A2(n12193), .ZN(n13360) );
  AOI21_X1 U14600 ( .B1(n12195), .B2(n13705), .A(n13360), .ZN(n13796) );
  XNOR2_X1 U14601 ( .A(n12197), .B(n12196), .ZN(n13794) );
  XNOR2_X1 U14602 ( .A(n12201), .B(n12198), .ZN(n12199) );
  OR2_X1 U14603 ( .A1(n12199), .A2(n10861), .ZN(n13791) );
  OAI22_X1 U14604 ( .A1(n13689), .A2(n13477), .B1(n13357), .B2(n13683), .ZN(
        n12200) );
  AOI21_X1 U14605 ( .B1(n12201), .B2(n13685), .A(n12200), .ZN(n12202) );
  OAI21_X1 U14606 ( .B1(n13791), .B2(n13519), .A(n12202), .ZN(n12203) );
  AOI21_X1 U14607 ( .B1(n13794), .B2(n13652), .A(n12203), .ZN(n12204) );
  OAI21_X1 U14608 ( .B1(n13796), .B2(n15301), .A(n12204), .ZN(P2_U3248) );
  INV_X1 U14609 ( .A(n12205), .ZN(n12207) );
  NOR2_X1 U14610 ( .A1(n10229), .A2(n12209), .ZN(n12210) );
  AOI21_X1 U14611 ( .B1(n14925), .B2(n12404), .A(n12210), .ZN(n12217) );
  AOI22_X1 U14612 ( .A1(n14925), .A2(n10208), .B1(n12409), .B2(n14943), .ZN(
        n12211) );
  XNOR2_X1 U14613 ( .A(n12211), .B(n10223), .ZN(n12218) );
  XOR2_X1 U14614 ( .A(n12217), .B(n12218), .Z(n14930) );
  NAND2_X1 U14615 ( .A1(n12216), .A2(n10208), .ZN(n12213) );
  NAND2_X1 U14616 ( .A1(n12409), .A2(n13959), .ZN(n12212) );
  NAND2_X1 U14617 ( .A1(n12213), .A2(n12212), .ZN(n12214) );
  XNOR2_X1 U14618 ( .A(n12214), .B(n10223), .ZN(n12220) );
  NOR2_X1 U14619 ( .A1(n10229), .A2(n12230), .ZN(n12215) );
  AOI21_X1 U14620 ( .B1(n12216), .B2(n12404), .A(n12215), .ZN(n12221) );
  XNOR2_X1 U14621 ( .A(n12220), .B(n12221), .ZN(n14938) );
  OR2_X1 U14622 ( .A1(n12218), .A2(n12217), .ZN(n14939) );
  AND2_X1 U14623 ( .A1(n14938), .A2(n14939), .ZN(n12219) );
  INV_X1 U14624 ( .A(n12220), .ZN(n12222) );
  NAND2_X1 U14625 ( .A1(n12227), .A2(n10208), .ZN(n12224) );
  NAND2_X1 U14626 ( .A1(n12409), .A2(n14978), .ZN(n12223) );
  NAND2_X1 U14627 ( .A1(n12224), .A2(n12223), .ZN(n12225) );
  XNOR2_X1 U14628 ( .A(n12225), .B(n10223), .ZN(n12236) );
  NOR2_X1 U14629 ( .A1(n10229), .A2(n12246), .ZN(n12226) );
  AOI21_X1 U14630 ( .B1(n12227), .B2(n12404), .A(n12226), .ZN(n12237) );
  XNOR2_X1 U14631 ( .A(n12236), .B(n12237), .ZN(n12228) );
  OAI211_X1 U14632 ( .C1(n12229), .C2(n12228), .A(n12240), .B(n14960), .ZN(
        n12235) );
  NAND2_X1 U14633 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n15046)
         );
  OAI21_X1 U14634 ( .B1(n14910), .B2(n12230), .A(n15046), .ZN(n12233) );
  NOR2_X1 U14635 ( .A1(n14964), .A2(n12231), .ZN(n12232) );
  AOI211_X1 U14636 ( .C1(n14954), .C2(n13958), .A(n12233), .B(n12232), .ZN(
        n12234) );
  OAI211_X1 U14637 ( .C1(n14794), .C2(n14958), .A(n12235), .B(n12234), .ZN(
        P1_U3224) );
  INV_X1 U14638 ( .A(n12237), .ZN(n12238) );
  NAND2_X1 U14639 ( .A1(n12236), .A2(n12238), .ZN(n12239) );
  NOR2_X1 U14640 ( .A1(n10229), .A2(n14911), .ZN(n12241) );
  AOI21_X1 U14641 ( .B1(n14981), .B2(n12404), .A(n12241), .ZN(n12312) );
  AOI22_X1 U14642 ( .A1(n14981), .A2(n10208), .B1(n12409), .B2(n13958), .ZN(
        n12242) );
  XNOR2_X1 U14643 ( .A(n12242), .B(n10223), .ZN(n12313) );
  XOR2_X1 U14644 ( .A(n12312), .B(n12313), .Z(n12243) );
  OAI211_X1 U14645 ( .C1(n12244), .C2(n12243), .A(n14914), .B(n14960), .ZN(
        n12250) );
  OAI22_X1 U14646 ( .A1(n14910), .A2(n12246), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12245), .ZN(n12248) );
  NOR2_X1 U14647 ( .A1(n14964), .A2(n14802), .ZN(n12247) );
  AOI211_X1 U14648 ( .C1(n14954), .C2(n14955), .A(n12248), .B(n12247), .ZN(
        n12249) );
  OAI211_X1 U14649 ( .C1(n7372), .C2(n14958), .A(n12250), .B(n12249), .ZN(
        P1_U3234) );
  NOR2_X1 U14650 ( .A1(n12252), .A2(n12251), .ZN(n12261) );
  OAI22_X1 U14651 ( .A1(n12255), .A2(n12254), .B1(n12253), .B2(n14801), .ZN(
        n12256) );
  AOI21_X1 U14652 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n15105), .A(n12256), 
        .ZN(n12258) );
  NAND2_X1 U14653 ( .A1(n14806), .A2(n14095), .ZN(n12257) );
  OAI211_X1 U14654 ( .C1(n12259), .C2(n15107), .A(n12258), .B(n12257), .ZN(
        n12260) );
  AOI211_X1 U14655 ( .C1(n12262), .C2(n14809), .A(n12261), .B(n12260), .ZN(
        n12263) );
  OAI21_X1 U14656 ( .B1(n12264), .B2(n14233), .A(n12263), .ZN(P1_U3356) );
  INV_X1 U14657 ( .A(n12265), .ZN(n12267) );
  OAI222_X1 U14658 ( .A1(n12268), .A2(P3_U3151), .B1(n12306), .B2(n12267), 
        .C1(n12266), .C2(n12423), .ZN(P3_U3271) );
  INV_X1 U14659 ( .A(n12269), .ZN(n14391) );
  OAI222_X1 U14660 ( .A1(n13844), .A2(n12271), .B1(n13850), .B2(n14391), .C1(
        n12270), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U14661 ( .A(n12272), .ZN(n14382) );
  OAI222_X1 U14662 ( .A1(n13852), .A2(n12422), .B1(P2_U3088), .B2(n12273), 
        .C1(n13850), .C2(n14382), .ZN(P2_U3297) );
  INV_X1 U14663 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12282) );
  AOI21_X1 U14664 ( .B1(n12275), .B2(n12783), .A(n12274), .ZN(n12291) );
  INV_X1 U14665 ( .A(n12291), .ZN(n12281) );
  AOI21_X1 U14666 ( .B1(n12645), .B2(n12277), .A(n12276), .ZN(n12280) );
  OAI22_X1 U14667 ( .A1(n12473), .A2(n15507), .B1(n9927), .B2(n15509), .ZN(
        n12278) );
  MUX2_X1 U14668 ( .A(n12282), .B(n13172), .S(n15570), .Z(n12283) );
  NAND2_X1 U14669 ( .A1(n12284), .A2(n15501), .ZN(n12289) );
  INV_X1 U14670 ( .A(n12475), .ZN(n12286) );
  OAI22_X1 U14671 ( .A1(n12286), .A2(n15479), .B1(n15501), .B2(n12285), .ZN(
        n12287) );
  AOI21_X1 U14672 ( .B1(n12470), .B2(n13148), .A(n12287), .ZN(n12288) );
  OAI211_X1 U14673 ( .C1(n12291), .C2(n12290), .A(n12289), .B(n12288), .ZN(
        P3_U3206) );
  INV_X1 U14674 ( .A(n12292), .ZN(n14385) );
  OAI222_X1 U14675 ( .A1(n13844), .A2(n12294), .B1(P2_U3088), .B2(n12293), 
        .C1(n13850), .C2(n14385), .ZN(P2_U3298) );
  INV_X1 U14676 ( .A(n12295), .ZN(n12296) );
  OAI222_X1 U14677 ( .A1(P3_U3151), .A2(n9459), .B1(n12423), .B2(n12297), .C1(
        n12306), .C2(n12296), .ZN(P3_U3266) );
  INV_X1 U14678 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n12298) );
  MUX2_X1 U14679 ( .A(n12298), .B(n12300), .S(n15570), .Z(n12299) );
  OAI21_X1 U14680 ( .B1(n10790), .B2(n13285), .A(n12299), .ZN(P3_U3390) );
  MUX2_X1 U14681 ( .A(n12301), .B(n12300), .S(n15585), .Z(n12302) );
  OAI21_X1 U14682 ( .B1(n10790), .B2(n13232), .A(n12302), .ZN(P3_U3459) );
  INV_X1 U14683 ( .A(n12303), .ZN(n12305) );
  OAI222_X1 U14684 ( .A1(n12306), .A2(n12305), .B1(n12423), .B2(n12304), .C1(
        P3_U3151), .C2(n12936), .ZN(P3_U3268) );
  NAND2_X1 U14685 ( .A1(n14971), .A2(n10208), .ZN(n12308) );
  NAND2_X1 U14686 ( .A1(n12404), .A2(n14955), .ZN(n12307) );
  NAND2_X1 U14687 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  XNOR2_X1 U14688 ( .A(n12309), .B(n10223), .ZN(n12317) );
  NOR2_X1 U14689 ( .A1(n10229), .A2(n12310), .ZN(n12311) );
  AOI21_X1 U14690 ( .B1(n14971), .B2(n12404), .A(n12311), .ZN(n12315) );
  XNOR2_X1 U14691 ( .A(n12317), .B(n12315), .ZN(n14912) );
  OR2_X1 U14692 ( .A1(n12313), .A2(n12312), .ZN(n14913) );
  INV_X1 U14693 ( .A(n12315), .ZN(n12316) );
  OR2_X1 U14694 ( .A1(n12317), .A2(n12316), .ZN(n12318) );
  NAND2_X1 U14695 ( .A1(n14354), .A2(n10208), .ZN(n12320) );
  NAND2_X1 U14696 ( .A1(n12409), .A2(n13957), .ZN(n12319) );
  NAND2_X1 U14697 ( .A1(n12320), .A2(n12319), .ZN(n12321) );
  XNOR2_X1 U14698 ( .A(n12321), .B(n10223), .ZN(n12323) );
  XNOR2_X1 U14699 ( .A(n12322), .B(n12323), .ZN(n14951) );
  AOI22_X1 U14700 ( .A1(n14354), .A2(n12404), .B1(n12408), .B2(n13957), .ZN(
        n14952) );
  NAND2_X1 U14701 ( .A1(n14951), .A2(n14952), .ZN(n14950) );
  INV_X1 U14702 ( .A(n12322), .ZN(n12324) );
  OR2_X1 U14703 ( .A1(n14967), .A2(n12363), .ZN(n12327) );
  NAND2_X1 U14704 ( .A1(n12408), .A2(n14953), .ZN(n12326) );
  NAND2_X1 U14705 ( .A1(n12327), .A2(n12326), .ZN(n12331) );
  OAI22_X1 U14706 ( .A1(n14967), .A2(n12353), .B1(n12328), .B2(n12363), .ZN(
        n12329) );
  XNOR2_X1 U14707 ( .A(n12329), .B(n10223), .ZN(n12330) );
  XOR2_X1 U14708 ( .A(n12331), .B(n12330), .Z(n13896) );
  INV_X1 U14709 ( .A(n12330), .ZN(n12333) );
  INV_X1 U14710 ( .A(n12331), .ZN(n12332) );
  NAND2_X1 U14711 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  OAI22_X1 U14712 ( .A1(n14349), .A2(n12363), .B1(n13943), .B2(n10229), .ZN(
        n12339) );
  NAND2_X1 U14713 ( .A1(n13912), .A2(n10208), .ZN(n12336) );
  NAND2_X1 U14714 ( .A1(n14237), .A2(n12409), .ZN(n12335) );
  NAND2_X1 U14715 ( .A1(n12336), .A2(n12335), .ZN(n12337) );
  XNOR2_X1 U14716 ( .A(n12337), .B(n10223), .ZN(n12338) );
  XOR2_X1 U14717 ( .A(n12339), .B(n12338), .Z(n13904) );
  INV_X1 U14718 ( .A(n12338), .ZN(n12341) );
  INV_X1 U14719 ( .A(n12339), .ZN(n12340) );
  NAND2_X1 U14720 ( .A1(n14342), .A2(n10208), .ZN(n12343) );
  NAND2_X1 U14721 ( .A1(n14222), .A2(n12409), .ZN(n12342) );
  NAND2_X1 U14722 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  XNOR2_X1 U14723 ( .A(n12344), .B(n10223), .ZN(n12347) );
  AOI22_X1 U14724 ( .A1(n14342), .A2(n12409), .B1(n12408), .B2(n14222), .ZN(
        n12345) );
  XNOR2_X1 U14725 ( .A(n12347), .B(n12345), .ZN(n13938) );
  INV_X1 U14726 ( .A(n12345), .ZN(n12346) );
  NOR2_X1 U14727 ( .A1(n12347), .A2(n12346), .ZN(n12348) );
  OAI22_X1 U14728 ( .A1(n14335), .A2(n12363), .B1(n14199), .B2(n10229), .ZN(
        n12350) );
  OAI22_X1 U14729 ( .A1(n14335), .A2(n12353), .B1(n14199), .B2(n12363), .ZN(
        n12349) );
  XNOR2_X1 U14730 ( .A(n12349), .B(n10223), .ZN(n12351) );
  XOR2_X1 U14731 ( .A(n12350), .B(n12351), .Z(n13870) );
  NAND2_X1 U14732 ( .A1(n12351), .A2(n12350), .ZN(n12352) );
  NAND2_X1 U14733 ( .A1(n13869), .A2(n12352), .ZN(n13924) );
  OAI22_X1 U14734 ( .A1(n14212), .A2(n12363), .B1(n14221), .B2(n10229), .ZN(
        n12355) );
  OAI22_X1 U14735 ( .A1(n14212), .A2(n12353), .B1(n14221), .B2(n12363), .ZN(
        n12354) );
  XNOR2_X1 U14736 ( .A(n12354), .B(n10223), .ZN(n12356) );
  XOR2_X1 U14737 ( .A(n12355), .B(n12356), .Z(n13923) );
  NAND2_X1 U14738 ( .A1(n12356), .A2(n12355), .ZN(n12357) );
  AOI22_X1 U14739 ( .A1(n14324), .A2(n10208), .B1(n12409), .B2(n14175), .ZN(
        n12358) );
  XNOR2_X1 U14740 ( .A(n12358), .B(n10223), .ZN(n12361) );
  AOI22_X1 U14741 ( .A1(n14324), .A2(n12409), .B1(n12408), .B2(n14175), .ZN(
        n12360) );
  XNOR2_X1 U14742 ( .A(n12361), .B(n12360), .ZN(n13880) );
  NAND2_X1 U14743 ( .A1(n12361), .A2(n12360), .ZN(n12362) );
  OAI22_X1 U14744 ( .A1(n7369), .A2(n12363), .B1(n13881), .B2(n10229), .ZN(
        n12369) );
  NAND2_X1 U14745 ( .A1(n12364), .A2(n10208), .ZN(n12366) );
  NAND2_X1 U14746 ( .A1(n14156), .A2(n12409), .ZN(n12365) );
  NAND2_X1 U14747 ( .A1(n12366), .A2(n12365), .ZN(n12367) );
  XNOR2_X1 U14748 ( .A(n12367), .B(n10223), .ZN(n12368) );
  XOR2_X1 U14749 ( .A(n12369), .B(n12368), .Z(n13931) );
  INV_X1 U14750 ( .A(n12368), .ZN(n12371) );
  INV_X1 U14751 ( .A(n12369), .ZN(n12370) );
  NAND2_X1 U14752 ( .A1(n14313), .A2(n10208), .ZN(n12373) );
  NAND2_X1 U14753 ( .A1(n12409), .A2(n14174), .ZN(n12372) );
  NAND2_X1 U14754 ( .A1(n12373), .A2(n12372), .ZN(n12374) );
  XNOR2_X1 U14755 ( .A(n12374), .B(n10223), .ZN(n12375) );
  AOI22_X1 U14756 ( .A1(n14313), .A2(n12409), .B1(n12408), .B2(n14174), .ZN(
        n12376) );
  XNOR2_X1 U14757 ( .A(n12375), .B(n12376), .ZN(n13863) );
  INV_X1 U14758 ( .A(n12375), .ZN(n12377) );
  NAND2_X1 U14759 ( .A1(n12377), .A2(n12376), .ZN(n12378) );
  NAND2_X1 U14760 ( .A1(n14308), .A2(n10208), .ZN(n12381) );
  NAND2_X1 U14761 ( .A1(n12409), .A2(n14157), .ZN(n12380) );
  NAND2_X1 U14762 ( .A1(n12381), .A2(n12380), .ZN(n12382) );
  XNOR2_X1 U14763 ( .A(n12382), .B(n10223), .ZN(n12383) );
  AOI22_X1 U14764 ( .A1(n14308), .A2(n12409), .B1(n12408), .B2(n14157), .ZN(
        n12384) );
  XNOR2_X1 U14765 ( .A(n12383), .B(n12384), .ZN(n13916) );
  NAND2_X1 U14766 ( .A1(n13915), .A2(n13916), .ZN(n12387) );
  INV_X1 U14767 ( .A(n12383), .ZN(n12385) );
  NAND2_X1 U14768 ( .A1(n12385), .A2(n12384), .ZN(n12386) );
  NAND2_X1 U14769 ( .A1(n14131), .A2(n10208), .ZN(n12389) );
  NAND2_X1 U14770 ( .A1(n12409), .A2(n13955), .ZN(n12388) );
  NAND2_X1 U14771 ( .A1(n12389), .A2(n12388), .ZN(n12390) );
  XNOR2_X1 U14772 ( .A(n12390), .B(n10223), .ZN(n12391) );
  AOI22_X1 U14773 ( .A1(n14131), .A2(n12409), .B1(n12408), .B2(n13955), .ZN(
        n12392) );
  XNOR2_X1 U14774 ( .A(n12391), .B(n12392), .ZN(n13887) );
  INV_X1 U14775 ( .A(n12391), .ZN(n12393) );
  NAND2_X1 U14776 ( .A1(n12393), .A2(n12392), .ZN(n12394) );
  NAND2_X1 U14777 ( .A1(n14112), .A2(n10208), .ZN(n12396) );
  NAND2_X1 U14778 ( .A1(n12409), .A2(n14094), .ZN(n12395) );
  NAND2_X1 U14779 ( .A1(n12396), .A2(n12395), .ZN(n12397) );
  XNOR2_X1 U14780 ( .A(n12397), .B(n10223), .ZN(n12398) );
  AOI22_X1 U14781 ( .A1(n14112), .A2(n12409), .B1(n12408), .B2(n14094), .ZN(
        n12399) );
  XNOR2_X1 U14782 ( .A(n12398), .B(n12399), .ZN(n13948) );
  INV_X1 U14783 ( .A(n12398), .ZN(n12400) );
  NAND2_X1 U14784 ( .A1(n14285), .A2(n10208), .ZN(n12402) );
  NAND2_X1 U14785 ( .A1(n12409), .A2(n14069), .ZN(n12401) );
  NAND2_X1 U14786 ( .A1(n12402), .A2(n12401), .ZN(n12403) );
  XNOR2_X1 U14787 ( .A(n12403), .B(n10223), .ZN(n12405) );
  AOI22_X1 U14788 ( .A1(n14285), .A2(n12404), .B1(n12408), .B2(n14069), .ZN(
        n12406) );
  XNOR2_X1 U14789 ( .A(n12405), .B(n12406), .ZN(n13855) );
  INV_X1 U14790 ( .A(n12405), .ZN(n12407) );
  AOI22_X1 U14791 ( .A1(n14279), .A2(n10208), .B1(n12409), .B2(n14095), .ZN(
        n12412) );
  AOI22_X1 U14792 ( .A1(n14279), .A2(n12409), .B1(n12408), .B2(n14095), .ZN(
        n12410) );
  XNOR2_X1 U14793 ( .A(n12410), .B(n10223), .ZN(n12411) );
  XOR2_X1 U14794 ( .A(n12412), .B(n12411), .Z(n12413) );
  NOR2_X1 U14795 ( .A1(n14964), .A2(n14081), .ZN(n12417) );
  AOI22_X1 U14796 ( .A1(n14954), .A2(n14070), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12414) );
  OAI21_X1 U14797 ( .B1(n12415), .B2(n14910), .A(n12414), .ZN(n12416) );
  AOI211_X1 U14798 ( .C1(n14279), .C2(n14921), .A(n12417), .B(n12416), .ZN(
        n12418) );
  OAI21_X1 U14799 ( .B1(n12419), .B2(n14916), .A(n12418), .ZN(P1_U3220) );
  INV_X1 U14800 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14381) );
  OAI22_X1 U14801 ( .A1(n14381), .A2(n12422), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12594) );
  XOR2_X1 U14802 ( .A(n12595), .B(n12594), .Z(n12601) );
  INV_X1 U14803 ( .A(SI_30_), .ZN(n12604) );
  INV_X1 U14804 ( .A(n12428), .ZN(n12430) );
  NAND2_X1 U14805 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  XNOR2_X1 U14806 ( .A(n13278), .B(n12469), .ZN(n12433) );
  XNOR2_X1 U14807 ( .A(n12433), .B(n12817), .ZN(n12582) );
  NAND2_X1 U14808 ( .A1(n12583), .A2(n12582), .ZN(n12435) );
  NAND2_X1 U14809 ( .A1(n12433), .A2(n13159), .ZN(n12434) );
  NAND2_X1 U14810 ( .A1(n12435), .A2(n12434), .ZN(n12517) );
  XNOR2_X1 U14811 ( .A(n12515), .B(n12466), .ZN(n12436) );
  XNOR2_X1 U14812 ( .A(n12436), .B(n13142), .ZN(n12516) );
  OR2_X2 U14813 ( .A1(n12517), .A2(n12516), .ZN(n12518) );
  INV_X1 U14814 ( .A(n12436), .ZN(n12437) );
  NAND2_X1 U14815 ( .A1(n12437), .A2(n12531), .ZN(n12438) );
  XNOR2_X1 U14816 ( .A(n13271), .B(n12466), .ZN(n12439) );
  XNOR2_X1 U14817 ( .A(n12439), .B(n13130), .ZN(n12526) );
  INV_X1 U14818 ( .A(n12439), .ZN(n12440) );
  NAND2_X1 U14819 ( .A1(n12440), .A2(n13130), .ZN(n12441) );
  XNOR2_X1 U14820 ( .A(n13267), .B(n12469), .ZN(n12561) );
  AND2_X1 U14821 ( .A1(n12561), .A2(n13118), .ZN(n12442) );
  XNOR2_X1 U14822 ( .A(n13264), .B(n12469), .ZN(n12443) );
  XNOR2_X1 U14823 ( .A(n12443), .B(n12549), .ZN(n12483) );
  NAND2_X1 U14824 ( .A1(n12482), .A2(n12483), .ZN(n12445) );
  NAND2_X1 U14825 ( .A1(n12443), .A2(n13100), .ZN(n12444) );
  XNOR2_X1 U14826 ( .A(n13076), .B(n12452), .ZN(n12545) );
  AND2_X1 U14827 ( .A1(n12545), .A2(n13085), .ZN(n12446) );
  INV_X1 U14828 ( .A(n12545), .ZN(n12447) );
  NAND2_X1 U14829 ( .A1(n12447), .A2(n13058), .ZN(n12448) );
  XNOR2_X1 U14830 ( .A(n13258), .B(n12469), .ZN(n12449) );
  XNOR2_X1 U14831 ( .A(n12449), .B(n13070), .ZN(n12500) );
  NAND2_X1 U14832 ( .A1(n12449), .A2(n13042), .ZN(n12450) );
  XNOR2_X1 U14833 ( .A(n12453), .B(n12452), .ZN(n12454) );
  INV_X1 U14834 ( .A(n12454), .ZN(n12455) );
  AND2_X1 U14835 ( .A1(n12456), .A2(n12455), .ZN(n12457) );
  AOI21_X2 U14836 ( .B1(n12555), .B2(n12554), .A(n12457), .ZN(n12535) );
  XNOR2_X1 U14837 ( .A(n12458), .B(n12466), .ZN(n12537) );
  XNOR2_X1 U14838 ( .A(n12767), .B(n12466), .ZN(n12460) );
  OAI22_X1 U14839 ( .A1(n12537), .A2(n12511), .B1(n13043), .B2(n12460), .ZN(
        n12463) );
  INV_X1 U14840 ( .A(n12460), .ZN(n12534) );
  INV_X1 U14841 ( .A(n13043), .ZN(n12815) );
  NOR2_X1 U14842 ( .A1(n12534), .A2(n12815), .ZN(n12459) );
  OAI21_X1 U14843 ( .B1(n12511), .B2(n12459), .A(n12537), .ZN(n12462) );
  NAND3_X1 U14844 ( .A1(n12460), .A2(n12511), .A3(n13043), .ZN(n12461) );
  XNOR2_X1 U14845 ( .A(n13243), .B(n12469), .ZN(n12464) );
  XNOR2_X1 U14846 ( .A(n12464), .B(n13013), .ZN(n12507) );
  INV_X1 U14847 ( .A(n12464), .ZN(n12465) );
  XNOR2_X1 U14848 ( .A(n12467), .B(n12466), .ZN(n12468) );
  XNOR2_X1 U14849 ( .A(n12468), .B(n9927), .ZN(n12570) );
  XNOR2_X1 U14850 ( .A(n12470), .B(n12469), .ZN(n12489) );
  XNOR2_X1 U14851 ( .A(n12489), .B(n9945), .ZN(n12490) );
  XNOR2_X1 U14852 ( .A(n12491), .B(n12490), .ZN(n12471) );
  AOI22_X1 U14853 ( .A1(n12996), .A2(n12586), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12472) );
  OAI21_X1 U14854 ( .B1(n12473), .B2(n12584), .A(n12472), .ZN(n12474) );
  AOI21_X1 U14855 ( .B1(n12475), .B2(n12578), .A(n12474), .ZN(n12476) );
  XNOR2_X1 U14856 ( .A(n12535), .B(n12534), .ZN(n12536) );
  XNOR2_X1 U14857 ( .A(n12536), .B(n12815), .ZN(n12477) );
  NAND2_X1 U14858 ( .A1(n12477), .A2(n12572), .ZN(n12481) );
  AOI22_X1 U14859 ( .A1(n9912), .A2(n12574), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12478) );
  OAI21_X1 U14860 ( .B1(n12554), .B2(n12576), .A(n12478), .ZN(n12479) );
  AOI21_X1 U14861 ( .B1(n13036), .B2(n12578), .A(n12479), .ZN(n12480) );
  OAI211_X1 U14862 ( .C1(n13251), .C2(n12581), .A(n12481), .B(n12480), .ZN(
        P3_U3156) );
  XOR2_X1 U14863 ( .A(n12483), .B(n12482), .Z(n12484) );
  NAND2_X1 U14864 ( .A1(n12484), .A2(n12572), .ZN(n12488) );
  NAND2_X1 U14865 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12941)
         );
  OAI21_X1 U14866 ( .B1(n12584), .B2(n13058), .A(n12941), .ZN(n12486) );
  NOR2_X1 U14867 ( .A1(n12588), .A2(n13089), .ZN(n12485) );
  AOI211_X1 U14868 ( .C1(n12586), .C2(n13086), .A(n12486), .B(n12485), .ZN(
        n12487) );
  OAI211_X1 U14869 ( .C1(n12581), .C2(n13264), .A(n12488), .B(n12487), .ZN(
        P3_U3159) );
  XNOR2_X1 U14870 ( .A(n12974), .B(n12466), .ZN(n12492) );
  NAND2_X1 U14871 ( .A1(n12493), .A2(n12572), .ZN(n12498) );
  INV_X1 U14872 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12494) );
  OAI22_X1 U14873 ( .A1(n12986), .A2(n12576), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12494), .ZN(n12496) );
  NOR2_X1 U14874 ( .A1(n12977), .A2(n12584), .ZN(n12495) );
  AOI211_X1 U14875 ( .C1(n12979), .C2(n12578), .A(n12496), .B(n12495), .ZN(
        n12497) );
  OAI211_X1 U14876 ( .C1(n13236), .C2(n12581), .A(n12498), .B(n12497), .ZN(
        P3_U3160) );
  XOR2_X1 U14877 ( .A(n12499), .B(n12500), .Z(n12506) );
  OAI22_X1 U14878 ( .A1(n12576), .A2(n13058), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12501), .ZN(n12503) );
  NOR2_X1 U14879 ( .A1(n12554), .A2(n12584), .ZN(n12502) );
  AOI211_X1 U14880 ( .C1(n12578), .C2(n13061), .A(n12503), .B(n12502), .ZN(
        n12505) );
  NAND2_X1 U14881 ( .A1(n13258), .A2(n12590), .ZN(n12504) );
  OAI211_X1 U14882 ( .C1(n12506), .C2(n12592), .A(n12505), .B(n12504), .ZN(
        P3_U3163) );
  XNOR2_X1 U14883 ( .A(n12508), .B(n12507), .ZN(n12509) );
  NAND2_X1 U14884 ( .A1(n12509), .A2(n12572), .ZN(n12514) );
  AOI22_X1 U14885 ( .A1(n12996), .A2(n12574), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12510) );
  OAI21_X1 U14886 ( .B1(n12511), .B2(n12576), .A(n12510), .ZN(n12512) );
  AOI21_X1 U14887 ( .B1(n13003), .B2(n12578), .A(n12512), .ZN(n12513) );
  OAI211_X1 U14888 ( .C1(n13243), .C2(n12581), .A(n12514), .B(n12513), .ZN(
        P3_U3165) );
  INV_X1 U14889 ( .A(n12515), .ZN(n13275) );
  AOI21_X1 U14890 ( .B1(n12517), .B2(n12516), .A(n12592), .ZN(n12519) );
  NAND2_X1 U14891 ( .A1(n12519), .A2(n12518), .ZN(n12523) );
  NAND2_X1 U14892 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12890)
         );
  OAI21_X1 U14893 ( .B1(n12584), .B2(n13130), .A(n12890), .ZN(n12521) );
  NOR2_X1 U14894 ( .A1(n12588), .A2(n13131), .ZN(n12520) );
  AOI211_X1 U14895 ( .C1(n12586), .C2(n12817), .A(n12521), .B(n12520), .ZN(
        n12522) );
  OAI211_X1 U14896 ( .C1(n13275), .C2(n12581), .A(n12523), .B(n12522), .ZN(
        P3_U3166) );
  OAI21_X1 U14897 ( .B1(n12526), .B2(n12525), .A(n12524), .ZN(n12527) );
  NAND2_X1 U14898 ( .A1(n12527), .A2(n12572), .ZN(n12533) );
  OAI22_X1 U14899 ( .A1(n12584), .A2(n13118), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12528), .ZN(n12530) );
  NOR2_X1 U14900 ( .A1(n12588), .A2(n13119), .ZN(n12529) );
  AOI211_X1 U14901 ( .C1(n12586), .C2(n12531), .A(n12530), .B(n12529), .ZN(
        n12532) );
  OAI211_X1 U14902 ( .C1(n12581), .C2(n13271), .A(n12533), .B(n12532), .ZN(
        P3_U3168) );
  OAI22_X1 U14903 ( .A1(n12536), .A2(n12815), .B1(n12535), .B2(n12534), .ZN(
        n12539) );
  XNOR2_X1 U14904 ( .A(n12537), .B(n9912), .ZN(n12538) );
  XNOR2_X1 U14905 ( .A(n12539), .B(n12538), .ZN(n12540) );
  NAND2_X1 U14906 ( .A1(n12540), .A2(n12572), .ZN(n12544) );
  INV_X1 U14907 ( .A(n13013), .ZN(n12814) );
  AOI22_X1 U14908 ( .A1(n12814), .A2(n12574), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12541) );
  OAI21_X1 U14909 ( .B1(n13043), .B2(n12576), .A(n12541), .ZN(n12542) );
  AOI21_X1 U14910 ( .B1(n13021), .B2(n12578), .A(n12542), .ZN(n12543) );
  OAI211_X1 U14911 ( .C1(n13247), .C2(n12581), .A(n12544), .B(n12543), .ZN(
        P3_U3169) );
  INV_X1 U14912 ( .A(n13076), .ZN(n13203) );
  XNOR2_X1 U14913 ( .A(n12545), .B(n13085), .ZN(n12546) );
  XNOR2_X1 U14914 ( .A(n12547), .B(n12546), .ZN(n12548) );
  NAND2_X1 U14915 ( .A1(n12548), .A2(n12572), .ZN(n12553) );
  NOR2_X1 U14916 ( .A1(n12576), .A2(n12549), .ZN(n12551) );
  INV_X1 U14917 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n14571) );
  OAI22_X1 U14918 ( .A1(n12584), .A2(n13042), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14571), .ZN(n12550) );
  AOI211_X1 U14919 ( .C1(n12578), .C2(n13072), .A(n12551), .B(n12550), .ZN(
        n12552) );
  OAI211_X1 U14920 ( .C1(n13203), .C2(n12581), .A(n12553), .B(n12552), .ZN(
        P3_U3173) );
  XNOR2_X1 U14921 ( .A(n12555), .B(n12554), .ZN(n12556) );
  NAND2_X1 U14922 ( .A1(n12556), .A2(n12572), .ZN(n12560) );
  AOI22_X1 U14923 ( .A1(n12586), .A2(n13070), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12557) );
  OAI21_X1 U14924 ( .B1(n13043), .B2(n12584), .A(n12557), .ZN(n12558) );
  AOI21_X1 U14925 ( .B1(n13048), .B2(n12578), .A(n12558), .ZN(n12559) );
  OAI211_X1 U14926 ( .C1(n13255), .C2(n12581), .A(n12560), .B(n12559), .ZN(
        P3_U3175) );
  XNOR2_X1 U14927 ( .A(n12561), .B(n13118), .ZN(n12562) );
  XNOR2_X1 U14928 ( .A(n12563), .B(n12562), .ZN(n12569) );
  NOR2_X1 U14929 ( .A1(n12564), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12922) );
  NOR2_X1 U14930 ( .A1(n12576), .A2(n13130), .ZN(n12565) );
  AOI211_X1 U14931 ( .C1(n12574), .C2(n13100), .A(n12922), .B(n12565), .ZN(
        n12566) );
  OAI21_X1 U14932 ( .B1(n12588), .B2(n13104), .A(n12566), .ZN(n12567) );
  AOI21_X1 U14933 ( .B1(n13267), .B2(n12590), .A(n12567), .ZN(n12568) );
  OAI21_X1 U14934 ( .B1(n12569), .B2(n12592), .A(n12568), .ZN(P3_U3178) );
  XNOR2_X1 U14935 ( .A(n12571), .B(n12570), .ZN(n12573) );
  NAND2_X1 U14936 ( .A1(n12573), .A2(n12572), .ZN(n12580) );
  AOI22_X1 U14937 ( .A1(n9945), .A2(n12574), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12575) );
  OAI21_X1 U14938 ( .B1(n13013), .B2(n12576), .A(n12575), .ZN(n12577) );
  AOI21_X1 U14939 ( .B1(n12989), .B2(n12578), .A(n12577), .ZN(n12579) );
  OAI211_X1 U14940 ( .C1(n9928), .C2(n12581), .A(n12580), .B(n12579), .ZN(
        P3_U3180) );
  XOR2_X1 U14941 ( .A(n12583), .B(n12582), .Z(n12593) );
  NAND2_X1 U14942 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12867)
         );
  OAI21_X1 U14943 ( .B1(n12584), .B2(n13142), .A(n12867), .ZN(n12585) );
  AOI21_X1 U14944 ( .B1(n12586), .B2(n14841), .A(n12585), .ZN(n12587) );
  OAI21_X1 U14945 ( .B1(n12588), .B2(n13145), .A(n12587), .ZN(n12589) );
  AOI21_X1 U14946 ( .B1(n13278), .B2(n12590), .A(n12589), .ZN(n12591) );
  OAI21_X1 U14947 ( .B1(n12593), .B2(n12592), .A(n12591), .ZN(P3_U3181) );
  OAI21_X1 U14948 ( .B1(n14381), .B2(P1_DATAO_REG_30__SCAN_IN), .A(n12596), 
        .ZN(n12599) );
  INV_X1 U14949 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U14950 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n13836), .B2(n12597), .ZN(n12598) );
  XOR2_X1 U14951 ( .A(n12599), .B(n12598), .Z(n13292) );
  INV_X1 U14952 ( .A(SI_31_), .ZN(n13288) );
  NOR2_X1 U14953 ( .A1(n6687), .A2(n13288), .ZN(n12600) );
  AOI21_X1 U14954 ( .B1(n13292), .B2(n12602), .A(n12600), .ZN(n14864) );
  INV_X1 U14955 ( .A(n14864), .ZN(n12621) );
  INV_X1 U14956 ( .A(n12601), .ZN(n12603) );
  OR2_X1 U14957 ( .A1(n12618), .A2(n12616), .ZN(n12615) );
  INV_X1 U14958 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14866) );
  NAND2_X1 U14959 ( .A1(n6688), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12608) );
  INV_X1 U14960 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12606) );
  OR2_X1 U14961 ( .A1(n6683), .A2(n12606), .ZN(n12607) );
  OAI211_X1 U14962 ( .C1(n6667), .C2(n14866), .A(n12608), .B(n12607), .ZN(
        n12610) );
  INV_X1 U14963 ( .A(n12610), .ZN(n12611) );
  NAND2_X1 U14964 ( .A1(n12612), .A2(n12611), .ZN(n12959) );
  INV_X1 U14965 ( .A(n12959), .ZN(n12613) );
  NAND2_X1 U14966 ( .A1(n12621), .A2(n12613), .ZN(n12614) );
  NAND2_X1 U14967 ( .A1(n12615), .A2(n12614), .ZN(n12800) );
  NAND2_X1 U14968 ( .A1(n12623), .A2(n12617), .ZN(n12796) );
  NAND2_X1 U14969 ( .A1(n14864), .A2(n12959), .ZN(n12799) );
  OAI21_X1 U14970 ( .B1(n14867), .B2(n12959), .A(n12799), .ZN(n12619) );
  INV_X1 U14971 ( .A(n12622), .ZN(n12806) );
  INV_X1 U14972 ( .A(n12623), .ZN(n12647) );
  INV_X1 U14973 ( .A(n12624), .ZN(n12781) );
  NAND2_X1 U14974 ( .A1(n12756), .A2(n12757), .ZN(n13046) );
  INV_X1 U14975 ( .A(n13052), .ZN(n13065) );
  NOR2_X1 U14976 ( .A1(n12626), .A2(n12625), .ZN(n12629) );
  INV_X1 U14977 ( .A(n11008), .ZN(n12628) );
  NAND4_X1 U14978 ( .A1(n12629), .A2(n12628), .A3(n12627), .A4(n12696), .ZN(
        n12631) );
  NOR2_X1 U14979 ( .A1(n12631), .A2(n12630), .ZN(n12635) );
  NAND4_X1 U14980 ( .A1(n12676), .A2(n6673), .A3(n12690), .A4(n12632), .ZN(
        n12633) );
  NOR2_X1 U14981 ( .A1(n12633), .A2(n12701), .ZN(n12634) );
  NAND4_X1 U14982 ( .A1(n12635), .A2(n9987), .A3(n7340), .A4(n12634), .ZN(
        n12638) );
  INV_X1 U14983 ( .A(n12636), .ZN(n12718) );
  INV_X1 U14984 ( .A(n14844), .ZN(n12637) );
  NOR3_X1 U14985 ( .A1(n12638), .A2(n13156), .A3(n12637), .ZN(n12639) );
  NAND3_X1 U14986 ( .A1(n13125), .A2(n13149), .A3(n12639), .ZN(n12640) );
  NOR2_X1 U14987 ( .A1(n12640), .A2(n13115), .ZN(n12641) );
  NAND3_X1 U14988 ( .A1(n13083), .A2(n13095), .A3(n12641), .ZN(n12642) );
  OR3_X1 U14989 ( .A1(n12761), .A2(n13031), .A3(n12642), .ZN(n12643) );
  NOR2_X1 U14990 ( .A1(n12998), .A2(n12643), .ZN(n12644) );
  NAND4_X1 U14991 ( .A1(n12645), .A2(n12987), .A3(n12644), .A4(n13008), .ZN(
        n12646) );
  NAND2_X1 U14992 ( .A1(n10789), .A2(n12651), .ZN(n12652) );
  NAND2_X1 U14993 ( .A1(n12652), .A2(n12653), .ZN(n12655) );
  AND2_X1 U14994 ( .A1(n12657), .A2(n12653), .ZN(n12654) );
  MUX2_X1 U14995 ( .A(n12655), .B(n12654), .S(n12780), .Z(n12656) );
  NAND2_X1 U14996 ( .A1(n12656), .A2(n12663), .ZN(n12662) );
  NOR2_X1 U14997 ( .A1(n12657), .A2(n12780), .ZN(n12658) );
  NOR2_X1 U14998 ( .A1(n12658), .A2(n9979), .ZN(n12661) );
  NAND2_X1 U14999 ( .A1(n12669), .A2(n12659), .ZN(n12660) );
  AOI21_X1 U15000 ( .B1(n12662), .B2(n12661), .A(n12660), .ZN(n12667) );
  AOI21_X1 U15001 ( .B1(n12627), .B2(n12663), .A(n12794), .ZN(n12666) );
  AND2_X1 U15002 ( .A1(n12668), .A2(n12664), .ZN(n12665) );
  OAI22_X1 U15003 ( .A1(n12667), .A2(n12666), .B1(n12665), .B2(n12794), .ZN(
        n12672) );
  MUX2_X1 U15004 ( .A(n12669), .B(n12668), .S(n12794), .Z(n12670) );
  NAND3_X1 U15005 ( .A1(n12672), .A2(n12671), .A3(n12670), .ZN(n12677) );
  OR2_X1 U15006 ( .A1(n15534), .A2(n12780), .ZN(n12674) );
  NAND2_X1 U15007 ( .A1(n15534), .A2(n12780), .ZN(n12673) );
  MUX2_X1 U15008 ( .A(n12674), .B(n12673), .S(n12824), .Z(n12675) );
  NAND3_X1 U15009 ( .A1(n12677), .A2(n12676), .A3(n12675), .ZN(n12681) );
  NAND2_X1 U15010 ( .A1(n12686), .A2(n12678), .ZN(n12679) );
  NAND2_X1 U15011 ( .A1(n12679), .A2(n12780), .ZN(n12680) );
  NAND2_X1 U15012 ( .A1(n12681), .A2(n12680), .ZN(n12685) );
  AOI21_X1 U15013 ( .B1(n12684), .B2(n12682), .A(n12780), .ZN(n12683) );
  AOI21_X1 U15014 ( .B1(n12685), .B2(n12684), .A(n12683), .ZN(n12692) );
  OAI21_X1 U15015 ( .B1(n12780), .B2(n12686), .A(n6673), .ZN(n12691) );
  MUX2_X1 U15016 ( .A(n12688), .B(n12687), .S(n12794), .Z(n12689) );
  OAI211_X1 U15017 ( .C1(n12692), .C2(n12691), .A(n12690), .B(n12689), .ZN(
        n12697) );
  MUX2_X1 U15018 ( .A(n12694), .B(n12693), .S(n12780), .Z(n12695) );
  NAND3_X1 U15019 ( .A1(n12697), .A2(n12696), .A3(n12695), .ZN(n12707) );
  AND2_X1 U15020 ( .A1(n12820), .A2(n12794), .ZN(n12700) );
  NOR2_X1 U15021 ( .A1(n12820), .A2(n12794), .ZN(n12699) );
  MUX2_X1 U15022 ( .A(n12700), .B(n12699), .S(n12698), .Z(n12702) );
  NOR3_X1 U15023 ( .A1(n12702), .A2(n12711), .A3(n12701), .ZN(n12706) );
  OAI211_X1 U15024 ( .C1(n12711), .C2(n12704), .A(n12717), .B(n12703), .ZN(
        n12705) );
  AOI22_X1 U15025 ( .A1(n12707), .A2(n12706), .B1(n12794), .B2(n12705), .ZN(
        n12715) );
  INV_X1 U15026 ( .A(n12709), .ZN(n12714) );
  NAND2_X1 U15027 ( .A1(n12819), .A2(n14859), .ZN(n12708) );
  OAI211_X1 U15028 ( .C1(n12711), .C2(n12710), .A(n12709), .B(n12708), .ZN(
        n12712) );
  NAND2_X1 U15029 ( .A1(n12712), .A2(n12780), .ZN(n12713) );
  OAI21_X1 U15030 ( .B1(n12715), .B2(n12714), .A(n12713), .ZN(n12716) );
  OAI211_X1 U15031 ( .C1(n12794), .C2(n12717), .A(n12716), .B(n14844), .ZN(
        n12721) );
  MUX2_X1 U15032 ( .A(n12719), .B(n12718), .S(n12794), .Z(n12720) );
  NAND3_X1 U15033 ( .A1(n12721), .A2(n7465), .A3(n12720), .ZN(n12725) );
  MUX2_X1 U15034 ( .A(n12723), .B(n12722), .S(n12780), .Z(n12724) );
  NAND2_X1 U15035 ( .A1(n12725), .A2(n12724), .ZN(n12726) );
  NAND2_X1 U15036 ( .A1(n12726), .A2(n13149), .ZN(n12730) );
  NAND2_X1 U15037 ( .A1(n12733), .A2(n12727), .ZN(n12728) );
  NAND2_X1 U15038 ( .A1(n12728), .A2(n12794), .ZN(n12729) );
  AOI21_X1 U15039 ( .B1(n12730), .B2(n12729), .A(n7470), .ZN(n12735) );
  AOI21_X1 U15040 ( .B1(n12732), .B2(n12731), .A(n12794), .ZN(n12734) );
  OAI22_X1 U15041 ( .A1(n12735), .A2(n12734), .B1(n12733), .B2(n12794), .ZN(
        n12742) );
  INV_X1 U15042 ( .A(n12736), .ZN(n12741) );
  INV_X1 U15043 ( .A(n12737), .ZN(n12738) );
  NAND2_X1 U15044 ( .A1(n12743), .A2(n12738), .ZN(n12739) );
  NAND4_X1 U15045 ( .A1(n12759), .A2(n12780), .A3(n12740), .A4(n12739), .ZN(
        n12745) );
  AOI22_X1 U15046 ( .A1(n12742), .A2(n13114), .B1(n12741), .B2(n12745), .ZN(
        n12748) );
  INV_X1 U15047 ( .A(n12761), .ZN(n12747) );
  NAND3_X1 U15048 ( .A1(n12758), .A2(n12743), .A3(n12794), .ZN(n12744) );
  NAND2_X1 U15049 ( .A1(n12745), .A2(n12744), .ZN(n12746) );
  OAI211_X1 U15050 ( .C1(n12748), .C2(n13107), .A(n12747), .B(n12746), .ZN(
        n12765) );
  INV_X1 U15051 ( .A(n13046), .ZN(n12755) );
  MUX2_X1 U15052 ( .A(n12750), .B(n12749), .S(n12780), .Z(n12754) );
  MUX2_X1 U15053 ( .A(n12794), .B(n13058), .S(n13076), .Z(n12751) );
  OAI21_X1 U15054 ( .B1(n12780), .B2(n13085), .A(n12751), .ZN(n12752) );
  NAND2_X1 U15055 ( .A1(n13052), .A2(n12752), .ZN(n12753) );
  NAND3_X1 U15056 ( .A1(n12755), .A2(n12754), .A3(n12753), .ZN(n12764) );
  MUX2_X1 U15057 ( .A(n12757), .B(n12756), .S(n12794), .Z(n12763) );
  MUX2_X1 U15058 ( .A(n12759), .B(n12758), .S(n12780), .Z(n12760) );
  OR2_X1 U15059 ( .A1(n12761), .A2(n12760), .ZN(n12762) );
  NAND4_X1 U15060 ( .A1(n12765), .A2(n12764), .A3(n12763), .A4(n12762), .ZN(
        n12766) );
  NAND2_X1 U15061 ( .A1(n12766), .A2(n13026), .ZN(n12769) );
  NAND3_X1 U15062 ( .A1(n12767), .A2(n13043), .A3(n12780), .ZN(n12768) );
  NAND2_X1 U15063 ( .A1(n12769), .A2(n12768), .ZN(n12770) );
  NAND2_X1 U15064 ( .A1(n12770), .A2(n13008), .ZN(n12775) );
  INV_X1 U15065 ( .A(n12998), .ZN(n12994) );
  XNOR2_X1 U15066 ( .A(n12771), .B(n12780), .ZN(n12772) );
  NAND2_X1 U15067 ( .A1(n12773), .A2(n12772), .ZN(n12774) );
  NAND3_X1 U15068 ( .A1(n12775), .A2(n12994), .A3(n12774), .ZN(n12779) );
  MUX2_X1 U15069 ( .A(n12777), .B(n12776), .S(n12780), .Z(n12778) );
  NAND3_X1 U15070 ( .A1(n12987), .A2(n12779), .A3(n12778), .ZN(n12785) );
  MUX2_X1 U15071 ( .A(n12782), .B(n12781), .S(n12780), .Z(n12784) );
  OAI211_X1 U15072 ( .C1(n12788), .C2(n12794), .A(n12787), .B(n12786), .ZN(
        n12789) );
  NAND3_X1 U15073 ( .A1(n12791), .A2(n12790), .A3(n12789), .ZN(n12798) );
  INV_X1 U15074 ( .A(n12792), .ZN(n12793) );
  AOI21_X1 U15075 ( .B1(n12795), .B2(n12794), .A(n12793), .ZN(n12797) );
  AOI21_X1 U15076 ( .B1(n12798), .B2(n12797), .A(n12796), .ZN(n12801) );
  MUX2_X1 U15077 ( .A(n12804), .B(n12803), .S(n12802), .Z(n12805) );
  NAND3_X1 U15078 ( .A1(n12808), .A2(n12807), .A3(n12913), .ZN(n12809) );
  OAI211_X1 U15079 ( .C1(n12810), .C2(n12812), .A(n12809), .B(P3_B_REG_SCAN_IN), .ZN(n12811) );
  OAI21_X1 U15080 ( .B1(n12813), .B2(n12812), .A(n12811), .ZN(P3_U3296) );
  MUX2_X1 U15081 ( .A(n12959), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12816), .Z(
        P3_U3522) );
  MUX2_X1 U15082 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n9945), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15083 ( .A(n12996), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12816), .Z(
        P3_U3517) );
  MUX2_X1 U15084 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12814), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15085 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n9912), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15086 ( .A(n12815), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12816), .Z(
        P3_U3514) );
  MUX2_X1 U15087 ( .A(n13056), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12816), .Z(
        P3_U3513) );
  MUX2_X1 U15088 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13070), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15089 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13085), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15090 ( .A(n13100), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12816), .Z(
        P3_U3510) );
  MUX2_X1 U15091 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13086), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15092 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13101), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15093 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12817), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15094 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n14841), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15095 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12818), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15096 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n14854), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15097 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12819), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15098 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n14852), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15099 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12820), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15100 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12821), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15101 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12822), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15102 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12823), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15103 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12824), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15104 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12825), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15105 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12826), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15106 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n10788), .S(P3_U3897), .Z(
        P3_U3492) );
  INV_X1 U15107 ( .A(n12827), .ZN(n12829) );
  NAND2_X1 U15108 ( .A1(n12829), .A2(n12828), .ZN(n12834) );
  NAND2_X1 U15109 ( .A1(n14781), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12870) );
  OR2_X1 U15110 ( .A1(n14781), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12830) );
  NAND2_X1 U15111 ( .A1(n12870), .A2(n12830), .ZN(n12845) );
  INV_X1 U15112 ( .A(n12845), .ZN(n12832) );
  NAND2_X1 U15113 ( .A1(n14781), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12865) );
  OR2_X1 U15114 ( .A1(n14781), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12831) );
  AND2_X1 U15115 ( .A1(n12865), .A2(n12831), .ZN(n12841) );
  MUX2_X1 U15116 ( .A(n12832), .B(n12841), .S(n12913), .Z(n12833) );
  NAND3_X1 U15117 ( .A1(n12835), .A2(n12834), .A3(n12833), .ZN(n12861) );
  NAND2_X1 U15118 ( .A1(n12861), .A2(n12954), .ZN(n12859) );
  AOI21_X1 U15119 ( .B1(n12835), .B2(n12834), .A(n12833), .ZN(n12858) );
  INV_X1 U15120 ( .A(n14781), .ZN(n12856) );
  NAND2_X1 U15121 ( .A1(n12837), .A2(n12836), .ZN(n12839) );
  NAND2_X1 U15122 ( .A1(n12839), .A2(n12838), .ZN(n12840) );
  NAND2_X1 U15123 ( .A1(n12841), .A2(n12840), .ZN(n12864) );
  OAI21_X1 U15124 ( .B1(n12841), .B2(n12840), .A(n12864), .ZN(n12842) );
  INV_X1 U15125 ( .A(n12842), .ZN(n12854) );
  NAND2_X1 U15126 ( .A1(n12845), .A2(n12846), .ZN(n12848) );
  NOR2_X1 U15127 ( .A1(n12846), .A2(n12845), .ZN(n12847) );
  NAND2_X1 U15128 ( .A1(n12848), .A2(n12869), .ZN(n12849) );
  NAND2_X1 U15129 ( .A1(n14832), .A2(n12849), .ZN(n12853) );
  INV_X1 U15130 ( .A(n12850), .ZN(n12851) );
  AOI21_X1 U15131 ( .B1(n15460), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12851), 
        .ZN(n12852) );
  OAI211_X1 U15132 ( .C1(n12854), .C2(n12949), .A(n12853), .B(n12852), .ZN(
        n12855) );
  AOI21_X1 U15133 ( .B1(n14825), .B2(n12856), .A(n12855), .ZN(n12857) );
  OAI21_X1 U15134 ( .B1(n12859), .B2(n12858), .A(n12857), .ZN(P3_U3196) );
  MUX2_X1 U15135 ( .A(n12870), .B(n12865), .S(n12913), .Z(n12860) );
  NAND2_X1 U15136 ( .A1(n12861), .A2(n12860), .ZN(n12896) );
  XOR2_X1 U15137 ( .A(n12898), .B(n12896), .Z(n12863) );
  MUX2_X1 U15138 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12913), .Z(n12862) );
  NOR2_X1 U15139 ( .A1(n12863), .A2(n12862), .ZN(n12897) );
  AOI21_X1 U15140 ( .B1(n12863), .B2(n12862), .A(n12897), .ZN(n12879) );
  NAND2_X1 U15141 ( .A1(n12865), .A2(n12864), .ZN(n12883) );
  XNOR2_X1 U15142 ( .A(n12898), .B(n12883), .ZN(n12866) );
  NAND2_X1 U15143 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12866), .ZN(n12885) );
  OAI21_X1 U15144 ( .B1(n12866), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12885), 
        .ZN(n12876) );
  NAND2_X1 U15145 ( .A1(n15460), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n12868) );
  NAND2_X1 U15146 ( .A1(n12868), .A2(n12867), .ZN(n12875) );
  AOI21_X1 U15147 ( .B1(n12872), .B2(n13146), .A(n12881), .ZN(n12873) );
  NOR2_X1 U15148 ( .A1(n15467), .A2(n12873), .ZN(n12874) );
  AOI211_X1 U15149 ( .C1(n15463), .C2(n12876), .A(n12875), .B(n12874), .ZN(
        n12878) );
  NAND2_X1 U15150 ( .A1(n14825), .A2(n12898), .ZN(n12877) );
  OAI211_X1 U15151 ( .C1(n12879), .C2(n15456), .A(n12878), .B(n12877), .ZN(
        P3_U3197) );
  AOI22_X1 U15152 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12912), .B1(n12889), 
        .B2(n13132), .ZN(n12882) );
  AOI21_X1 U15153 ( .B1(n6798), .B2(n12882), .A(n12908), .ZN(n12906) );
  AOI22_X1 U15154 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12889), .B1(n12912), 
        .B2(n13220), .ZN(n12888) );
  NAND2_X1 U15155 ( .A1(n12884), .A2(n12883), .ZN(n12886) );
  NAND2_X1 U15156 ( .A1(n12886), .A2(n12885), .ZN(n12887) );
  NAND2_X1 U15157 ( .A1(n12888), .A2(n12887), .ZN(n12911) );
  OAI21_X1 U15158 ( .B1(n12888), .B2(n12887), .A(n12911), .ZN(n12895) );
  NOR2_X1 U15159 ( .A1(n15454), .A2(n12889), .ZN(n12894) );
  OAI21_X1 U15160 ( .B1(n12892), .B2(n12891), .A(n12890), .ZN(n12893) );
  AOI211_X1 U15161 ( .C1(n12895), .C2(n15463), .A(n12894), .B(n12893), .ZN(
        n12905) );
  INV_X1 U15162 ( .A(n12896), .ZN(n12899) );
  AOI21_X1 U15163 ( .B1(n12899), .B2(n12898), .A(n12897), .ZN(n12916) );
  MUX2_X1 U15164 ( .A(n13132), .B(n13220), .S(n12913), .Z(n12900) );
  NOR2_X1 U15165 ( .A1(n12900), .A2(n12912), .ZN(n12915) );
  INV_X1 U15166 ( .A(n12915), .ZN(n12901) );
  NAND2_X1 U15167 ( .A1(n12900), .A2(n12912), .ZN(n12914) );
  NAND2_X1 U15168 ( .A1(n12901), .A2(n12914), .ZN(n12902) );
  XNOR2_X1 U15169 ( .A(n12916), .B(n12902), .ZN(n12903) );
  NAND2_X1 U15170 ( .A1(n12903), .A2(n12954), .ZN(n12904) );
  OAI211_X1 U15171 ( .C1(n12906), .C2(n15467), .A(n12905), .B(n12904), .ZN(
        P3_U3198) );
  NOR2_X1 U15172 ( .A1(n12912), .A2(n13132), .ZN(n12907) );
  NAND2_X1 U15173 ( .A1(n12920), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12929) );
  OAI21_X1 U15174 ( .B1(n12920), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12929), 
        .ZN(n12910) );
  AOI21_X1 U15175 ( .B1(n6804), .B2(n12910), .A(n12931), .ZN(n12928) );
  XOR2_X1 U15176 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12944), .Z(n12945) );
  XNOR2_X1 U15177 ( .A(n12946), .B(n12945), .ZN(n12926) );
  MUX2_X1 U15178 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12936), .Z(n12919) );
  MUX2_X1 U15179 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12913), .Z(n12917) );
  OAI21_X1 U15180 ( .B1(n12916), .B2(n12915), .A(n12914), .ZN(n14828) );
  XNOR2_X1 U15181 ( .A(n12917), .B(n14824), .ZN(n14829) );
  NOR2_X1 U15182 ( .A1(n14828), .A2(n14829), .ZN(n14827) );
  AOI21_X1 U15183 ( .B1(n12917), .B2(n14824), .A(n14827), .ZN(n12934) );
  XNOR2_X1 U15184 ( .A(n12934), .B(n12944), .ZN(n12918) );
  NOR2_X1 U15185 ( .A1(n12918), .A2(n12919), .ZN(n12933) );
  AOI21_X1 U15186 ( .B1(n12919), .B2(n12918), .A(n12933), .ZN(n12924) );
  NOR2_X1 U15187 ( .A1(n15454), .A2(n12920), .ZN(n12921) );
  AOI211_X1 U15188 ( .C1(n15460), .C2(P3_ADDR_REG_18__SCAN_IN), .A(n12922), 
        .B(n12921), .ZN(n12923) );
  OAI21_X1 U15189 ( .B1(n12924), .B2(n15456), .A(n12923), .ZN(n12925) );
  AOI21_X1 U15190 ( .B1(n15463), .B2(n12926), .A(n12925), .ZN(n12927) );
  OAI21_X1 U15191 ( .B1(n12928), .B2(n15467), .A(n12927), .ZN(P3_U3200) );
  INV_X1 U15192 ( .A(n12929), .ZN(n12930) );
  XNOR2_X1 U15193 ( .A(n12942), .B(n13090), .ZN(n12935) );
  XNOR2_X1 U15194 ( .A(n12932), .B(n12935), .ZN(n12956) );
  AOI21_X1 U15195 ( .B1(n12934), .B2(n12944), .A(n12933), .ZN(n12939) );
  INV_X1 U15196 ( .A(n12935), .ZN(n12937) );
  XNOR2_X1 U15197 ( .A(n12942), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12947) );
  MUX2_X1 U15198 ( .A(n12937), .B(n12947), .S(n12936), .Z(n12938) );
  XNOR2_X1 U15199 ( .A(n12939), .B(n12938), .ZN(n12953) );
  NAND2_X1 U15200 ( .A1(n15460), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12940) );
  OAI211_X1 U15201 ( .C1(n15454), .C2(n12942), .A(n12941), .B(n12940), .ZN(
        n12952) );
  XNOR2_X1 U15202 ( .A(n12948), .B(n12947), .ZN(n12950) );
  NOR2_X1 U15203 ( .A1(n12950), .A2(n12949), .ZN(n12951) );
  OAI21_X1 U15204 ( .B1(n12956), .B2(n15467), .A(n12955), .ZN(P3_U3201) );
  INV_X1 U15205 ( .A(n12957), .ZN(n12958) );
  NAND2_X1 U15206 ( .A1(n12959), .A2(n12958), .ZN(n14868) );
  NAND2_X1 U15207 ( .A1(n12960), .A2(n15517), .ZN(n12965) );
  OAI21_X1 U15208 ( .B1(n13166), .B2(n14868), .A(n12965), .ZN(n12962) );
  AOI21_X1 U15209 ( .B1(n13166), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12962), 
        .ZN(n12961) );
  OAI21_X1 U15210 ( .B1(n14864), .B2(n13163), .A(n12961), .ZN(P3_U3202) );
  AOI21_X1 U15211 ( .B1(n13166), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12962), 
        .ZN(n12963) );
  OAI21_X1 U15212 ( .B1(n14867), .B2(n13163), .A(n12963), .ZN(P3_U3203) );
  INV_X1 U15213 ( .A(n12964), .ZN(n12972) );
  OAI21_X1 U15214 ( .B1(n15501), .B2(n12966), .A(n12965), .ZN(n12967) );
  AOI21_X1 U15215 ( .B1(n12968), .B2(n13148), .A(n12967), .ZN(n12971) );
  NAND2_X1 U15216 ( .A1(n12969), .A2(n15501), .ZN(n12970) );
  OAI211_X1 U15217 ( .C1(n12972), .C2(n13137), .A(n12971), .B(n12970), .ZN(
        P3_U3204) );
  XNOR2_X1 U15218 ( .A(n12973), .B(n12974), .ZN(n13169) );
  INV_X1 U15219 ( .A(n13169), .ZN(n12983) );
  NAND2_X1 U15220 ( .A1(n9945), .A2(n14851), .ZN(n12978) );
  AOI22_X1 U15221 ( .A1(n12979), .A2(n15517), .B1(n13166), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12980) );
  OAI21_X1 U15222 ( .B1(n13236), .B2(n13163), .A(n12980), .ZN(n12981) );
  AOI21_X1 U15223 ( .B1(n13168), .B2(n15501), .A(n12981), .ZN(n12982) );
  OAI21_X1 U15224 ( .B1(n12983), .B2(n13137), .A(n12982), .ZN(P3_U3205) );
  XOR2_X1 U15225 ( .A(n12987), .B(n12984), .Z(n12985) );
  OAI222_X1 U15226 ( .A1(n15507), .A2(n12986), .B1(n15509), .B2(n13013), .C1(
        n12985), .C2(n15490), .ZN(n13175) );
  INV_X1 U15227 ( .A(n13175), .ZN(n12993) );
  XNOR2_X1 U15228 ( .A(n12988), .B(n12987), .ZN(n13176) );
  AOI22_X1 U15229 ( .A1(n15517), .A2(n12989), .B1(n13166), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12990) );
  OAI21_X1 U15230 ( .B1(n9928), .B2(n13163), .A(n12990), .ZN(n12991) );
  AOI21_X1 U15231 ( .B1(n13176), .B2(n14861), .A(n12991), .ZN(n12992) );
  OAI21_X1 U15232 ( .B1(n12993), .B2(n13166), .A(n12992), .ZN(P3_U3207) );
  XNOR2_X1 U15233 ( .A(n12995), .B(n12994), .ZN(n13002) );
  AOI22_X1 U15234 ( .A1(n12996), .A2(n14853), .B1(n9912), .B2(n14851), .ZN(
        n13001) );
  OAI211_X1 U15235 ( .C1(n12999), .C2(n12998), .A(n12997), .B(n15511), .ZN(
        n13000) );
  OAI211_X1 U15236 ( .C1(n13002), .C2(n15514), .A(n13001), .B(n13000), .ZN(
        n13179) );
  INV_X1 U15237 ( .A(n13179), .ZN(n13007) );
  INV_X1 U15238 ( .A(n13002), .ZN(n13180) );
  AOI22_X1 U15239 ( .A1(n13166), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n13003), 
        .B2(n15517), .ZN(n13004) );
  OAI21_X1 U15240 ( .B1(n13243), .B2(n13163), .A(n13004), .ZN(n13005) );
  AOI21_X1 U15241 ( .B1(n13180), .B2(n15518), .A(n13005), .ZN(n13006) );
  OAI21_X1 U15242 ( .B1(n13007), .B2(n13166), .A(n13006), .ZN(P3_U3208) );
  INV_X1 U15243 ( .A(n13029), .ZN(n13010) );
  AOI21_X1 U15244 ( .B1(n13010), .B2(n13009), .A(n13008), .ZN(n13012) );
  NOR2_X1 U15245 ( .A1(n13012), .A2(n13011), .ZN(n13020) );
  OAI22_X1 U15246 ( .A1(n13013), .A2(n15507), .B1(n13043), .B2(n15509), .ZN(
        n13014) );
  INV_X1 U15247 ( .A(n13014), .ZN(n13019) );
  OAI211_X1 U15248 ( .C1(n13017), .C2(n13016), .A(n13015), .B(n15511), .ZN(
        n13018) );
  OAI211_X1 U15249 ( .C1(n13020), .C2(n15514), .A(n13019), .B(n13018), .ZN(
        n13183) );
  INV_X1 U15250 ( .A(n13183), .ZN(n13025) );
  INV_X1 U15251 ( .A(n13020), .ZN(n13184) );
  AOI22_X1 U15252 ( .A1(n13166), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15517), 
        .B2(n13021), .ZN(n13022) );
  OAI21_X1 U15253 ( .B1(n13247), .B2(n13163), .A(n13022), .ZN(n13023) );
  AOI21_X1 U15254 ( .B1(n13184), .B2(n15518), .A(n13023), .ZN(n13024) );
  OAI21_X1 U15255 ( .B1(n13025), .B2(n13166), .A(n13024), .ZN(P3_U3209) );
  NOR2_X1 U15256 ( .A1(n13027), .A2(n13026), .ZN(n13028) );
  AOI22_X1 U15257 ( .A1(n9912), .A2(n14853), .B1(n14851), .B2(n13056), .ZN(
        n13034) );
  OAI211_X1 U15258 ( .C1(n13032), .C2(n13031), .A(n13030), .B(n15511), .ZN(
        n13033) );
  OAI211_X1 U15259 ( .C1(n13035), .C2(n15514), .A(n13034), .B(n13033), .ZN(
        n13187) );
  INV_X1 U15260 ( .A(n13187), .ZN(n13040) );
  AOI22_X1 U15261 ( .A1(n13166), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15517), 
        .B2(n13036), .ZN(n13037) );
  OAI21_X1 U15262 ( .B1(n13251), .B2(n13163), .A(n13037), .ZN(n13038) );
  AOI21_X1 U15263 ( .B1(n13188), .B2(n15518), .A(n13038), .ZN(n13039) );
  OAI21_X1 U15264 ( .B1(n13040), .B2(n13166), .A(n13039), .ZN(P3_U3210) );
  XNOR2_X1 U15265 ( .A(n13041), .B(n13046), .ZN(n13045) );
  OAI22_X1 U15266 ( .A1(n13043), .A2(n15507), .B1(n13042), .B2(n15509), .ZN(
        n13044) );
  AOI21_X1 U15267 ( .B1(n13045), .B2(n15511), .A(n13044), .ZN(n13191) );
  XNOR2_X1 U15268 ( .A(n13047), .B(n13046), .ZN(n13190) );
  AOI22_X1 U15269 ( .A1(n13166), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15517), 
        .B2(n13048), .ZN(n13049) );
  OAI21_X1 U15270 ( .B1(n13255), .B2(n13163), .A(n13049), .ZN(n13050) );
  AOI21_X1 U15271 ( .B1(n13190), .B2(n14861), .A(n13050), .ZN(n13051) );
  OAI21_X1 U15272 ( .B1(n13166), .B2(n13191), .A(n13051), .ZN(P3_U3211) );
  OR2_X1 U15273 ( .A1(n13053), .A2(n13052), .ZN(n13055) );
  NAND2_X1 U15274 ( .A1(n13053), .A2(n13052), .ZN(n13054) );
  NAND2_X1 U15275 ( .A1(n13055), .A2(n13054), .ZN(n13060) );
  NAND2_X1 U15276 ( .A1(n13056), .A2(n14853), .ZN(n13057) );
  OAI21_X1 U15277 ( .B1(n13058), .B2(n15509), .A(n13057), .ZN(n13059) );
  AOI21_X1 U15278 ( .B1(n13060), .B2(n15511), .A(n13059), .ZN(n13196) );
  INV_X1 U15279 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13063) );
  INV_X1 U15280 ( .A(n13061), .ZN(n13062) );
  OAI22_X1 U15281 ( .A1(n15501), .A2(n13063), .B1(n13062), .B2(n15479), .ZN(
        n13064) );
  AOI21_X1 U15282 ( .B1(n13258), .B2(n13148), .A(n13064), .ZN(n13068) );
  XNOR2_X1 U15283 ( .A(n13066), .B(n13065), .ZN(n13195) );
  NAND2_X1 U15284 ( .A1(n13195), .A2(n14861), .ZN(n13067) );
  OAI211_X1 U15285 ( .C1(n13196), .C2(n13166), .A(n13068), .B(n13067), .ZN(
        P3_U3212) );
  XOR2_X1 U15286 ( .A(n13069), .B(n13079), .Z(n13071) );
  AOI222_X1 U15287 ( .A1(n15511), .A2(n13071), .B1(n13070), .B2(n14853), .C1(
        n13100), .C2(n14851), .ZN(n13202) );
  INV_X1 U15288 ( .A(n13072), .ZN(n13073) );
  OAI22_X1 U15289 ( .A1(n15501), .A2(n13074), .B1(n13073), .B2(n15479), .ZN(
        n13075) );
  AOI21_X1 U15290 ( .B1(n13076), .B2(n13148), .A(n13075), .ZN(n13081) );
  NAND2_X1 U15291 ( .A1(n13078), .A2(n13079), .ZN(n13200) );
  NAND3_X1 U15292 ( .A1(n13077), .A2(n13200), .A3(n14861), .ZN(n13080) );
  OAI211_X1 U15293 ( .C1(n13202), .C2(n13166), .A(n13081), .B(n13080), .ZN(
        P3_U3213) );
  XOR2_X1 U15294 ( .A(n13082), .B(n13083), .Z(n13205) );
  INV_X1 U15295 ( .A(n13205), .ZN(n13094) );
  OAI211_X1 U15296 ( .C1(n6815), .C2(n7356), .A(n15511), .B(n13084), .ZN(
        n13088) );
  AOI22_X1 U15297 ( .A1(n14851), .A2(n13086), .B1(n13085), .B2(n14853), .ZN(
        n13087) );
  NAND2_X1 U15298 ( .A1(n13088), .A2(n13087), .ZN(n13204) );
  NOR2_X1 U15299 ( .A1(n13264), .A2(n13163), .ZN(n13092) );
  OAI22_X1 U15300 ( .A1(n15501), .A2(n13090), .B1(n13089), .B2(n15479), .ZN(
        n13091) );
  AOI211_X1 U15301 ( .C1(n13204), .C2(n15501), .A(n13092), .B(n13091), .ZN(
        n13093) );
  OAI21_X1 U15302 ( .B1(n13094), .B2(n13137), .A(n13093), .ZN(P3_U3214) );
  NAND2_X1 U15303 ( .A1(n13096), .A2(n13095), .ZN(n13097) );
  NAND2_X1 U15304 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  NAND2_X1 U15305 ( .A1(n13099), .A2(n15511), .ZN(n13103) );
  AOI22_X1 U15306 ( .A1(n14851), .A2(n13101), .B1(n13100), .B2(n14853), .ZN(
        n13102) );
  OAI22_X1 U15307 ( .A1(n15501), .A2(n13105), .B1(n13104), .B2(n15479), .ZN(
        n13111) );
  NAND2_X1 U15308 ( .A1(n13106), .A2(n13107), .ZN(n13108) );
  NAND2_X1 U15309 ( .A1(n13109), .A2(n13108), .ZN(n13209) );
  NOR2_X1 U15310 ( .A1(n13209), .A2(n13137), .ZN(n13110) );
  AOI211_X1 U15311 ( .C1(n13148), .C2(n13267), .A(n13111), .B(n13110), .ZN(
        n13112) );
  OAI21_X1 U15312 ( .B1(n13166), .B2(n13210), .A(n13112), .ZN(P3_U3215) );
  XNOR2_X1 U15313 ( .A(n13113), .B(n13114), .ZN(n13215) );
  INV_X1 U15314 ( .A(n13215), .ZN(n13124) );
  XNOR2_X1 U15315 ( .A(n13116), .B(n13115), .ZN(n13117) );
  OAI222_X1 U15316 ( .A1(n15507), .A2(n13118), .B1(n15509), .B2(n13142), .C1(
        n13117), .C2(n15490), .ZN(n13214) );
  INV_X1 U15317 ( .A(n13119), .ZN(n13120) );
  AOI22_X1 U15318 ( .A1(n13166), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15517), 
        .B2(n13120), .ZN(n13121) );
  OAI21_X1 U15319 ( .B1(n13271), .B2(n13163), .A(n13121), .ZN(n13122) );
  AOI21_X1 U15320 ( .B1(n13214), .B2(n15501), .A(n13122), .ZN(n13123) );
  OAI21_X1 U15321 ( .B1(n13137), .B2(n13124), .A(n13123), .ZN(P3_U3216) );
  XNOR2_X1 U15322 ( .A(n13126), .B(n13125), .ZN(n13219) );
  INV_X1 U15323 ( .A(n13219), .ZN(n13136) );
  XNOR2_X1 U15324 ( .A(n13127), .B(n13128), .ZN(n13129) );
  OAI222_X1 U15325 ( .A1(n15507), .A2(n13130), .B1(n15509), .B2(n13159), .C1(
        n13129), .C2(n15490), .ZN(n13218) );
  NOR2_X1 U15326 ( .A1(n13275), .A2(n13163), .ZN(n13134) );
  OAI22_X1 U15327 ( .A1(n15501), .A2(n13132), .B1(n13131), .B2(n15479), .ZN(
        n13133) );
  AOI211_X1 U15328 ( .C1(n13218), .C2(n15501), .A(n13134), .B(n13133), .ZN(
        n13135) );
  OAI21_X1 U15329 ( .B1(n13137), .B2(n13136), .A(n13135), .ZN(P3_U3217) );
  NAND2_X1 U15330 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  XNOR2_X1 U15331 ( .A(n13140), .B(n13149), .ZN(n13144) );
  NAND2_X1 U15332 ( .A1(n14841), .A2(n14851), .ZN(n13141) );
  OAI21_X1 U15333 ( .B1(n13142), .B2(n15507), .A(n13141), .ZN(n13143) );
  AOI21_X1 U15334 ( .B1(n13144), .B2(n15511), .A(n13143), .ZN(n13224) );
  OAI22_X1 U15335 ( .A1(n15501), .A2(n13146), .B1(n13145), .B2(n15479), .ZN(
        n13147) );
  AOI21_X1 U15336 ( .B1(n13148), .B2(n13278), .A(n13147), .ZN(n13154) );
  OR2_X1 U15337 ( .A1(n13150), .A2(n13149), .ZN(n13151) );
  NAND2_X1 U15338 ( .A1(n13152), .A2(n13151), .ZN(n13222) );
  NAND2_X1 U15339 ( .A1(n13222), .A2(n14861), .ZN(n13153) );
  OAI211_X1 U15340 ( .C1(n13224), .C2(n13166), .A(n13154), .B(n13153), .ZN(
        P3_U3218) );
  XNOR2_X1 U15341 ( .A(n13155), .B(n13156), .ZN(n13157) );
  OAI222_X1 U15342 ( .A1(n15507), .A2(n13159), .B1(n15509), .B2(n13158), .C1(
        n13157), .C2(n15490), .ZN(n13228) );
  INV_X1 U15343 ( .A(n13228), .ZN(n13167) );
  OAI21_X1 U15344 ( .B1(n6810), .B2(n7465), .A(n13160), .ZN(n13229) );
  AOI22_X1 U15345 ( .A1(n13166), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15517), 
        .B2(n13161), .ZN(n13162) );
  OAI21_X1 U15346 ( .B1(n13163), .B2(n13284), .A(n13162), .ZN(n13164) );
  AOI21_X1 U15347 ( .B1(n13229), .B2(n14861), .A(n13164), .ZN(n13165) );
  OAI21_X1 U15348 ( .B1(n13167), .B2(n13166), .A(n13165), .ZN(P3_U3219) );
  INV_X1 U15349 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13170) );
  AOI21_X1 U15350 ( .B1(n13169), .B2(n14883), .A(n13168), .ZN(n13233) );
  MUX2_X1 U15351 ( .A(n13170), .B(n13233), .S(n15585), .Z(n13171) );
  MUX2_X1 U15352 ( .A(n14580), .B(n13172), .S(n15585), .Z(n13173) );
  INV_X1 U15353 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13177) );
  AOI21_X1 U15354 ( .B1(n13176), .B2(n14883), .A(n13175), .ZN(n13237) );
  OAI21_X1 U15355 ( .B1(n9928), .B2(n13232), .A(n13178), .ZN(P3_U3485) );
  INV_X1 U15356 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13181) );
  AOI21_X1 U15357 ( .B1(n15566), .B2(n13180), .A(n13179), .ZN(n13240) );
  MUX2_X1 U15358 ( .A(n13181), .B(n13240), .S(n15585), .Z(n13182) );
  OAI21_X1 U15359 ( .B1(n13243), .B2(n13232), .A(n13182), .ZN(P3_U3484) );
  INV_X1 U15360 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13185) );
  AOI21_X1 U15361 ( .B1(n15566), .B2(n13184), .A(n13183), .ZN(n13244) );
  MUX2_X1 U15362 ( .A(n13185), .B(n13244), .S(n15585), .Z(n13186) );
  OAI21_X1 U15363 ( .B1(n13247), .B2(n13232), .A(n13186), .ZN(P3_U3483) );
  INV_X1 U15364 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n14626) );
  AOI21_X1 U15365 ( .B1(n15566), .B2(n13188), .A(n13187), .ZN(n13248) );
  MUX2_X1 U15366 ( .A(n14626), .B(n13248), .S(n15585), .Z(n13189) );
  OAI21_X1 U15367 ( .B1(n13251), .B2(n13232), .A(n13189), .ZN(P3_U3482) );
  NAND2_X1 U15368 ( .A1(n13190), .A2(n14883), .ZN(n13192) );
  NAND2_X1 U15369 ( .A1(n13192), .A2(n13191), .ZN(n13252) );
  MUX2_X1 U15370 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n13252), .S(n15585), .Z(
        n13193) );
  INV_X1 U15371 ( .A(n13193), .ZN(n13194) );
  OAI21_X1 U15372 ( .B1(n13255), .B2(n13232), .A(n13194), .ZN(P3_U3481) );
  INV_X1 U15373 ( .A(n13232), .ZN(n13226) );
  NAND2_X1 U15374 ( .A1(n13195), .A2(n14883), .ZN(n13197) );
  NAND2_X1 U15375 ( .A1(n13197), .A2(n13196), .ZN(n13256) );
  MUX2_X1 U15376 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n13256), .S(n15585), .Z(
        n13198) );
  AOI21_X1 U15377 ( .B1(n13226), .B2(n13258), .A(n13198), .ZN(n13199) );
  INV_X1 U15378 ( .A(n13199), .ZN(P3_U3480) );
  NAND3_X1 U15379 ( .A1(n13077), .A2(n14883), .A3(n13200), .ZN(n13201) );
  OAI211_X1 U15380 ( .C1(n13203), .C2(n15545), .A(n13202), .B(n13201), .ZN(
        n13260) );
  MUX2_X1 U15381 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13260), .S(n15585), .Z(
        P3_U3479) );
  AOI21_X1 U15382 ( .B1(n13205), .B2(n14883), .A(n13204), .ZN(n13261) );
  MUX2_X1 U15383 ( .A(n13206), .B(n13261), .S(n15585), .Z(n13207) );
  OAI21_X1 U15384 ( .B1(n13232), .B2(n13264), .A(n13207), .ZN(P3_U3478) );
  INV_X1 U15385 ( .A(n14883), .ZN(n13208) );
  OR2_X1 U15386 ( .A1(n13209), .A2(n13208), .ZN(n13211) );
  NAND2_X1 U15387 ( .A1(n13211), .A2(n13210), .ZN(n13265) );
  MUX2_X1 U15388 ( .A(n13265), .B(P3_REG1_REG_18__SCAN_IN), .S(n15583), .Z(
        n13212) );
  AOI21_X1 U15389 ( .B1(n13226), .B2(n13267), .A(n13212), .ZN(n13213) );
  INV_X1 U15390 ( .A(n13213), .ZN(P3_U3477) );
  INV_X1 U15391 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13216) );
  AOI21_X1 U15392 ( .B1(n13215), .B2(n14883), .A(n13214), .ZN(n13269) );
  MUX2_X1 U15393 ( .A(n13216), .B(n13269), .S(n15585), .Z(n13217) );
  OAI21_X1 U15394 ( .B1(n13232), .B2(n13271), .A(n13217), .ZN(P3_U3476) );
  AOI21_X1 U15395 ( .B1(n13219), .B2(n14883), .A(n13218), .ZN(n13272) );
  MUX2_X1 U15396 ( .A(n13220), .B(n13272), .S(n15585), .Z(n13221) );
  OAI21_X1 U15397 ( .B1(n13275), .B2(n13232), .A(n13221), .ZN(P3_U3475) );
  NAND2_X1 U15398 ( .A1(n13222), .A2(n14883), .ZN(n13223) );
  NAND2_X1 U15399 ( .A1(n13224), .A2(n13223), .ZN(n13276) );
  MUX2_X1 U15400 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13276), .S(n15585), .Z(
        n13225) );
  AOI21_X1 U15401 ( .B1(n13226), .B2(n13278), .A(n13225), .ZN(n13227) );
  INV_X1 U15402 ( .A(n13227), .ZN(P3_U3474) );
  AOI21_X1 U15403 ( .B1(n14883), .B2(n13229), .A(n13228), .ZN(n13281) );
  MUX2_X1 U15404 ( .A(n13230), .B(n13281), .S(n15585), .Z(n13231) );
  OAI21_X1 U15405 ( .B1(n13232), .B2(n13284), .A(n13231), .ZN(P3_U3473) );
  OAI21_X1 U15406 ( .B1(n9928), .B2(n13285), .A(n13239), .ZN(P3_U3453) );
  MUX2_X1 U15407 ( .A(n13241), .B(n13240), .S(n15570), .Z(n13242) );
  OAI21_X1 U15408 ( .B1(n13243), .B2(n13285), .A(n13242), .ZN(P3_U3452) );
  MUX2_X1 U15409 ( .A(n13245), .B(n13244), .S(n15570), .Z(n13246) );
  OAI21_X1 U15410 ( .B1(n13247), .B2(n13285), .A(n13246), .ZN(P3_U3451) );
  INV_X1 U15411 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13249) );
  MUX2_X1 U15412 ( .A(n13249), .B(n13248), .S(n15570), .Z(n13250) );
  OAI21_X1 U15413 ( .B1(n13251), .B2(n13285), .A(n13250), .ZN(P3_U3450) );
  MUX2_X1 U15414 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n13252), .S(n15570), .Z(
        n13253) );
  INV_X1 U15415 ( .A(n13253), .ZN(n13254) );
  OAI21_X1 U15416 ( .B1(n13255), .B2(n13285), .A(n13254), .ZN(P3_U3449) );
  INV_X1 U15417 ( .A(n13285), .ZN(n13279) );
  MUX2_X1 U15418 ( .A(n13256), .B(P3_REG0_REG_21__SCAN_IN), .S(n15568), .Z(
        n13257) );
  AOI21_X1 U15419 ( .B1(n13279), .B2(n13258), .A(n13257), .ZN(n13259) );
  INV_X1 U15420 ( .A(n13259), .ZN(P3_U3448) );
  MUX2_X1 U15421 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13260), .S(n15570), .Z(
        P3_U3447) );
  INV_X1 U15422 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13262) );
  MUX2_X1 U15423 ( .A(n13262), .B(n13261), .S(n15570), .Z(n13263) );
  OAI21_X1 U15424 ( .B1(n13285), .B2(n13264), .A(n13263), .ZN(P3_U3446) );
  MUX2_X1 U15425 ( .A(n13265), .B(P3_REG0_REG_18__SCAN_IN), .S(n15568), .Z(
        n13266) );
  AOI21_X1 U15426 ( .B1(n13279), .B2(n13267), .A(n13266), .ZN(n13268) );
  INV_X1 U15427 ( .A(n13268), .ZN(P3_U3444) );
  MUX2_X1 U15428 ( .A(n14567), .B(n13269), .S(n15570), .Z(n13270) );
  OAI21_X1 U15429 ( .B1(n13285), .B2(n13271), .A(n13270), .ZN(P3_U3441) );
  INV_X1 U15430 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13273) );
  MUX2_X1 U15431 ( .A(n13273), .B(n13272), .S(n15570), .Z(n13274) );
  OAI21_X1 U15432 ( .B1(n13275), .B2(n13285), .A(n13274), .ZN(P3_U3438) );
  MUX2_X1 U15433 ( .A(n13276), .B(P3_REG0_REG_15__SCAN_IN), .S(n15568), .Z(
        n13277) );
  AOI21_X1 U15434 ( .B1(n13279), .B2(n13278), .A(n13277), .ZN(n13280) );
  INV_X1 U15435 ( .A(n13280), .ZN(P3_U3435) );
  INV_X1 U15436 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13282) );
  MUX2_X1 U15437 ( .A(n13282), .B(n13281), .S(n15570), .Z(n13283) );
  OAI21_X1 U15438 ( .B1(n13285), .B2(n13284), .A(n13283), .ZN(P3_U3432) );
  NAND3_X1 U15439 ( .A1(n13287), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13289) );
  OAI22_X1 U15440 ( .A1(n13286), .A2(n13289), .B1(n13288), .B2(n12423), .ZN(
        n13290) );
  AOI21_X1 U15441 ( .B1(n13292), .B2(n13291), .A(n13290), .ZN(n13293) );
  INV_X1 U15442 ( .A(n13293), .ZN(P3_U3264) );
  INV_X1 U15443 ( .A(n13294), .ZN(n13295) );
  AOI22_X1 U15444 ( .A1(n13295), .A2(n10187), .B1(n13415), .B2(n13606), .ZN(
        n13300) );
  INV_X1 U15445 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13296) );
  OAI22_X1 U15446 ( .A1(n13390), .A2(n13629), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13296), .ZN(n13298) );
  OAI22_X1 U15447 ( .A1(n13389), .A2(n13662), .B1(n13406), .B2(n13631), .ZN(
        n13297) );
  AOI211_X1 U15448 ( .C1(n13759), .C2(n13425), .A(n13298), .B(n13297), .ZN(
        n13299) );
  OAI21_X1 U15449 ( .B1(n13301), .B2(n13300), .A(n13299), .ZN(P2_U3188) );
  XNOR2_X1 U15450 ( .A(n6990), .B(n13303), .ZN(n13304) );
  XNOR2_X1 U15451 ( .A(n13373), .B(n13304), .ZN(n13311) );
  NAND2_X1 U15452 ( .A1(n13434), .A2(n13604), .ZN(n13306) );
  NAND2_X1 U15453 ( .A1(n13436), .A2(n13607), .ZN(n13305) );
  NAND2_X1 U15454 ( .A1(n13306), .A2(n13305), .ZN(n13781) );
  INV_X1 U15455 ( .A(n13781), .ZN(n13308) );
  NAND2_X1 U15456 ( .A1(n13424), .A2(n13698), .ZN(n13307) );
  NAND2_X1 U15457 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13506)
         );
  OAI211_X1 U15458 ( .C1(n13308), .C2(n13397), .A(n13307), .B(n13506), .ZN(
        n13309) );
  AOI21_X1 U15459 ( .B1(n13782), .B2(n13425), .A(n13309), .ZN(n13310) );
  OAI21_X1 U15460 ( .B1(n13311), .B2(n13417), .A(n13310), .ZN(P2_U3191) );
  INV_X1 U15461 ( .A(n13312), .ZN(n13313) );
  NAND2_X1 U15462 ( .A1(n13551), .A2(n10861), .ZN(n13315) );
  XOR2_X1 U15463 ( .A(n13316), .B(n13315), .Z(n13317) );
  XNOR2_X1 U15464 ( .A(n13729), .B(n13317), .ZN(n13318) );
  NOR2_X1 U15465 ( .A1(n13406), .A2(n13538), .ZN(n13323) );
  NAND2_X1 U15466 ( .A1(n13431), .A2(n13604), .ZN(n13320) );
  NAND2_X1 U15467 ( .A1(n13575), .A2(n13607), .ZN(n13319) );
  AND2_X1 U15468 ( .A1(n13320), .A2(n13319), .ZN(n13536) );
  OAI22_X1 U15469 ( .A1(n13397), .A2(n13536), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13321), .ZN(n13322) );
  AOI211_X1 U15470 ( .C1(n13729), .C2(n13425), .A(n13323), .B(n13322), .ZN(
        n13324) );
  AOI22_X1 U15471 ( .A1(n13422), .A2(n13432), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13329) );
  AOI22_X1 U15472 ( .A1(n13666), .A2(n13424), .B1(n13421), .B2(n13434), .ZN(
        n13328) );
  NAND2_X1 U15473 ( .A1(n13772), .A2(n13425), .ZN(n13327) );
  NAND4_X1 U15474 ( .A1(n13330), .A2(n13329), .A3(n13328), .A4(n13327), .ZN(
        P2_U3195) );
  INV_X1 U15475 ( .A(n13403), .ZN(n13341) );
  OR2_X1 U15476 ( .A1(n13364), .A2(n13331), .ZN(n13334) );
  NOR2_X1 U15477 ( .A1(n13408), .A2(n13629), .ZN(n13333) );
  AOI22_X1 U15478 ( .A1(n13334), .A2(n10187), .B1(n13333), .B2(n13332), .ZN(
        n13340) );
  OAI22_X1 U15479 ( .A1(n13390), .A2(n13336), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13335), .ZN(n13338) );
  OAI22_X1 U15480 ( .A1(n13389), .A2(n13629), .B1(n13588), .B2(n13406), .ZN(
        n13337) );
  AOI211_X1 U15481 ( .C1(n13747), .C2(n13425), .A(n13338), .B(n13337), .ZN(
        n13339) );
  OAI21_X1 U15482 ( .B1(n13341), .B2(n13340), .A(n13339), .ZN(P2_U3197) );
  INV_X1 U15483 ( .A(n13342), .ZN(n13343) );
  AOI21_X1 U15484 ( .B1(n13345), .B2(n13344), .A(n13343), .ZN(n13352) );
  INV_X1 U15485 ( .A(n13437), .ZN(n13346) );
  NAND2_X1 U15486 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n13462)
         );
  OAI21_X1 U15487 ( .B1(n13390), .B2(n13346), .A(n13462), .ZN(n13350) );
  OAI22_X1 U15488 ( .A1(n13389), .A2(n13348), .B1(n13347), .B2(n13406), .ZN(
        n13349) );
  AOI211_X1 U15489 ( .C1(n13798), .C2(n13425), .A(n13350), .B(n13349), .ZN(
        n13351) );
  OAI21_X1 U15490 ( .B1(n13352), .B2(n13417), .A(n13351), .ZN(P2_U3198) );
  OAI21_X1 U15491 ( .B1(n13355), .B2(n13354), .A(n13353), .ZN(n13356) );
  NAND2_X1 U15492 ( .A1(n13356), .A2(n10187), .ZN(n13363) );
  NAND2_X1 U15493 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15284)
         );
  INV_X1 U15494 ( .A(n15284), .ZN(n13359) );
  NOR2_X1 U15495 ( .A1(n13406), .A2(n13357), .ZN(n13358) );
  AOI211_X1 U15496 ( .C1(n13361), .C2(n13360), .A(n13359), .B(n13358), .ZN(
        n13362) );
  OAI211_X1 U15497 ( .C1(n13792), .C2(n13369), .A(n13363), .B(n13362), .ZN(
        P2_U3200) );
  AOI211_X1 U15498 ( .C1(n6738), .C2(n13365), .A(n13417), .B(n13364), .ZN(
        n13371) );
  AOI22_X1 U15499 ( .A1(n13422), .A2(n13605), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13368) );
  INV_X1 U15500 ( .A(n13366), .ZN(n13614) );
  AOI22_X1 U15501 ( .A1(n13424), .A2(n13614), .B1(n13421), .B2(n13606), .ZN(
        n13367) );
  OAI211_X1 U15502 ( .C1(n13616), .C2(n13369), .A(n13368), .B(n13367), .ZN(
        n13370) );
  OR2_X1 U15503 ( .A1(n13371), .A2(n13370), .ZN(P2_U3201) );
  INV_X1 U15504 ( .A(n13372), .ZN(n13376) );
  INV_X1 U15505 ( .A(n13373), .ZN(n13374) );
  OAI33_X1 U15506 ( .A1(n13408), .A2(n13376), .A3(n13375), .B1(n13417), .B2(
        n6990), .B3(n13374), .ZN(n13378) );
  NAND2_X1 U15507 ( .A1(n13378), .A2(n13377), .ZN(n13383) );
  NOR2_X1 U15508 ( .A1(n13406), .A2(n13682), .ZN(n13381) );
  AOI22_X1 U15509 ( .A1(n13433), .A2(n13604), .B1(n13607), .B2(n13435), .ZN(
        n13675) );
  OAI22_X1 U15510 ( .A1(n13675), .A2(n13397), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13379), .ZN(n13380) );
  AOI211_X1 U15511 ( .C1(n13777), .C2(n13425), .A(n13381), .B(n13380), .ZN(
        n13382) );
  OAI211_X1 U15512 ( .C1(n13417), .C2(n13384), .A(n13383), .B(n13382), .ZN(
        P2_U3205) );
  NAND2_X1 U15513 ( .A1(n13415), .A2(n13432), .ZN(n13388) );
  NAND2_X1 U15514 ( .A1(n13385), .A2(n10187), .ZN(n13387) );
  MUX2_X1 U15515 ( .A(n13388), .B(n13387), .S(n13386), .Z(n13394) );
  OAI22_X1 U15516 ( .A1(n13389), .A2(n13641), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14574), .ZN(n13392) );
  OAI22_X1 U15517 ( .A1(n13390), .A2(n13640), .B1(n13644), .B2(n13406), .ZN(
        n13391) );
  AOI211_X1 U15518 ( .C1(n13765), .C2(n13425), .A(n13392), .B(n13391), .ZN(
        n13393) );
  NAND2_X1 U15519 ( .A1(n13394), .A2(n13393), .ZN(P2_U3207) );
  XNOR2_X1 U15520 ( .A(n13396), .B(n13395), .ZN(n13401) );
  NOR2_X1 U15521 ( .A1(n13406), .A2(n13712), .ZN(n13399) );
  AOI22_X1 U15522 ( .A1(n13435), .A2(n13604), .B1(n13607), .B2(n13437), .ZN(
        n13710) );
  NAND2_X1 U15523 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13481)
         );
  OAI21_X1 U15524 ( .B1(n13710), .B2(n13397), .A(n13481), .ZN(n13398) );
  AOI211_X1 U15525 ( .C1(n13787), .C2(n13425), .A(n13399), .B(n13398), .ZN(
        n13400) );
  OAI21_X1 U15526 ( .B1(n13401), .B2(n13417), .A(n13400), .ZN(P2_U3210) );
  OAI21_X1 U15527 ( .B1(n13410), .B2(n13403), .A(n13402), .ZN(n13404) );
  INV_X1 U15528 ( .A(n13404), .ZN(n13414) );
  AOI22_X1 U15529 ( .A1(n13422), .A2(n13575), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13405) );
  OAI21_X1 U15530 ( .B1(n13568), .B2(n13406), .A(n13405), .ZN(n13407) );
  AOI21_X1 U15531 ( .B1(n13742), .B2(n13425), .A(n13407), .ZN(n13413) );
  NOR3_X1 U15532 ( .A1(n13410), .A2(n13409), .A3(n13408), .ZN(n13411) );
  OAI21_X1 U15533 ( .B1(n13411), .B2(n13421), .A(n13605), .ZN(n13412) );
  OAI211_X1 U15534 ( .C1(n13414), .C2(n13417), .A(n13413), .B(n13412), .ZN(
        P2_U3212) );
  NAND2_X1 U15535 ( .A1(n13415), .A2(n13439), .ZN(n13420) );
  OR2_X1 U15536 ( .A1(n13417), .A2(n13416), .ZN(n13419) );
  MUX2_X1 U15537 ( .A(n13420), .B(n13419), .S(n13418), .Z(n13429) );
  AOI22_X1 U15538 ( .A1(n13421), .A2(n13440), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13428) );
  AOI22_X1 U15539 ( .A1(n13424), .A2(n13423), .B1(n13422), .B2(n13438), .ZN(
        n13427) );
  NAND2_X1 U15540 ( .A1(n13805), .A2(n13425), .ZN(n13426) );
  NAND4_X1 U15541 ( .A1(n13429), .A2(n13428), .A3(n13427), .A4(n13426), .ZN(
        P2_U3213) );
  MUX2_X1 U15542 ( .A(n13510), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13451), .Z(
        P2_U3562) );
  MUX2_X1 U15543 ( .A(n13430), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13451), .Z(
        P2_U3561) );
  MUX2_X1 U15544 ( .A(n13431), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13451), .Z(
        P2_U3560) );
  MUX2_X1 U15545 ( .A(n13551), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13451), .Z(
        P2_U3559) );
  MUX2_X1 U15546 ( .A(n13575), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13451), .Z(
        P2_U3558) );
  MUX2_X1 U15547 ( .A(n13583), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13451), .Z(
        P2_U3557) );
  MUX2_X1 U15548 ( .A(n13605), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13451), .Z(
        P2_U3556) );
  MUX2_X1 U15549 ( .A(n13584), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13451), .Z(
        P2_U3555) );
  MUX2_X1 U15550 ( .A(n13606), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13451), .Z(
        P2_U3554) );
  MUX2_X1 U15551 ( .A(n13432), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13451), .Z(
        P2_U3553) );
  MUX2_X1 U15552 ( .A(n13433), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13451), .Z(
        P2_U3552) );
  MUX2_X1 U15553 ( .A(n13434), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13451), .Z(
        P2_U3551) );
  MUX2_X1 U15554 ( .A(n13435), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13451), .Z(
        P2_U3550) );
  MUX2_X1 U15555 ( .A(n13436), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13451), .Z(
        P2_U3549) );
  MUX2_X1 U15556 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13437), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U15557 ( .A(n13438), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13451), .Z(
        P2_U3547) );
  MUX2_X1 U15558 ( .A(n13439), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13451), .Z(
        P2_U3546) );
  MUX2_X1 U15559 ( .A(n13440), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13451), .Z(
        P2_U3545) );
  MUX2_X1 U15560 ( .A(n13441), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13451), .Z(
        P2_U3544) );
  MUX2_X1 U15561 ( .A(n13442), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13451), .Z(
        P2_U3543) );
  MUX2_X1 U15562 ( .A(n13443), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13451), .Z(
        P2_U3542) );
  MUX2_X1 U15563 ( .A(n13444), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13451), .Z(
        P2_U3541) );
  MUX2_X1 U15564 ( .A(n13445), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13451), .Z(
        P2_U3540) );
  MUX2_X1 U15565 ( .A(n13446), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13451), .Z(
        P2_U3539) );
  MUX2_X1 U15566 ( .A(n13447), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13451), .Z(
        P2_U3538) );
  MUX2_X1 U15567 ( .A(n13448), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13451), .Z(
        P2_U3537) );
  MUX2_X1 U15568 ( .A(n13449), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13451), .Z(
        P2_U3536) );
  MUX2_X1 U15569 ( .A(n13450), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13451), .Z(
        P2_U3535) );
  MUX2_X1 U15570 ( .A(n8479), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13451), .Z(
        P2_U3534) );
  MUX2_X1 U15571 ( .A(n8475), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13451), .Z(
        P2_U3533) );
  MUX2_X1 U15572 ( .A(n10062), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13451), .Z(
        P2_U3532) );
  MUX2_X1 U15573 ( .A(n8473), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13451), .Z(
        P2_U3531) );
  NAND2_X1 U15574 ( .A1(n13467), .A2(n13452), .ZN(n13456) );
  OR2_X1 U15575 ( .A1(n13454), .A2(n13453), .ZN(n13455) );
  NAND2_X1 U15576 ( .A1(n13456), .A2(n13455), .ZN(n13457) );
  NAND2_X1 U15577 ( .A1(n15263), .A2(n13457), .ZN(n13458) );
  XNOR2_X1 U15578 ( .A(n13468), .B(n13457), .ZN(n15265) );
  NAND2_X1 U15579 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15265), .ZN(n15264) );
  NAND2_X1 U15580 ( .A1(n13458), .A2(n15264), .ZN(n13461) );
  MUX2_X1 U15581 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n13459), .S(n13483), .Z(
        n13460) );
  NAND2_X1 U15582 ( .A1(n13460), .A2(n13461), .ZN(n13475) );
  OAI211_X1 U15583 ( .C1(n13461), .C2(n13460), .A(n15277), .B(n13475), .ZN(
        n13465) );
  INV_X1 U15584 ( .A(n13462), .ZN(n13463) );
  AOI21_X1 U15585 ( .B1(n15281), .B2(n13483), .A(n13463), .ZN(n13464) );
  OAI211_X1 U15586 ( .C1(n15269), .C2(n7375), .A(n13465), .B(n13464), .ZN(
        n13474) );
  NOR2_X1 U15587 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  NOR2_X1 U15588 ( .A1(n15259), .A2(n15260), .ZN(n15258) );
  NOR2_X1 U15589 ( .A1(n13470), .A2(n15258), .ZN(n13472) );
  XNOR2_X1 U15590 ( .A(n13483), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13471) );
  NOR2_X1 U15591 ( .A1(n13472), .A2(n13471), .ZN(n13482) );
  AOI211_X1 U15592 ( .C1(n13472), .C2(n13471), .A(n13482), .B(n15271), .ZN(
        n13473) );
  OR2_X1 U15593 ( .A1(n13474), .A2(n13473), .ZN(P2_U3230) );
  OAI21_X1 U15594 ( .B1(n13476), .B2(n13459), .A(n13475), .ZN(n15278) );
  NOR2_X1 U15595 ( .A1(n13479), .A2(n13477), .ZN(n13478) );
  AOI21_X1 U15596 ( .B1(n13477), .B2(n13479), .A(n13478), .ZN(n15279) );
  NAND2_X1 U15597 ( .A1(n15278), .A2(n15279), .ZN(n15276) );
  OAI21_X1 U15598 ( .B1(n13477), .B2(n13479), .A(n15276), .ZN(n13491) );
  XNOR2_X1 U15599 ( .A(n13491), .B(n13492), .ZN(n13480) );
  NOR2_X1 U15600 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13480), .ZN(n13493) );
  AOI21_X1 U15601 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13480), .A(n13493), 
        .ZN(n13490) );
  OAI21_X1 U15602 ( .B1(n15236), .B2(n13496), .A(n13481), .ZN(n13487) );
  XNOR2_X1 U15603 ( .A(n15280), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15272) );
  INV_X1 U15604 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13484) );
  NOR2_X1 U15605 ( .A1(n13484), .A2(n13485), .ZN(n13499) );
  AOI211_X1 U15606 ( .C1(n13485), .C2(n13484), .A(n13499), .B(n15271), .ZN(
        n13486) );
  AOI211_X1 U15607 ( .C1(n15275), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13487), 
        .B(n13486), .ZN(n13488) );
  OAI21_X1 U15608 ( .B1(n13490), .B2(n13489), .A(n13488), .ZN(P2_U3232) );
  NOR2_X1 U15609 ( .A1(n13492), .A2(n13491), .ZN(n13494) );
  NOR2_X1 U15610 ( .A1(n13494), .A2(n13493), .ZN(n13495) );
  XOR2_X1 U15611 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13495), .Z(n13503) );
  INV_X1 U15612 ( .A(n13503), .ZN(n13501) );
  NOR2_X1 U15613 ( .A1(n13497), .A2(n13496), .ZN(n13498) );
  NOR2_X1 U15614 ( .A1(n13499), .A2(n13498), .ZN(n13500) );
  XNOR2_X1 U15615 ( .A(n13500), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13502) );
  AOI22_X1 U15616 ( .A1(n13503), .A2(n15277), .B1(n15231), .B2(n13502), .ZN(
        n13505) );
  INV_X1 U15617 ( .A(n13508), .ZN(n13509) );
  NAND2_X1 U15618 ( .A1(n13510), .A2(n13509), .ZN(n13724) );
  NOR2_X1 U15619 ( .A1(n15301), .A2(n13724), .ZN(n13517) );
  NOR2_X1 U15620 ( .A1(n7487), .A2(n15292), .ZN(n13512) );
  AOI211_X1 U15621 ( .C1(n15290), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13517), 
        .B(n13512), .ZN(n13513) );
  OAI21_X1 U15622 ( .B1(n13723), .B2(n13519), .A(n13513), .ZN(P2_U3234) );
  OAI211_X1 U15623 ( .C1(n13726), .C2(n13515), .A(n10146), .B(n13514), .ZN(
        n13725) );
  NOR2_X1 U15624 ( .A1(n13726), .A2(n15292), .ZN(n13516) );
  AOI211_X1 U15625 ( .C1(n15290), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13517), 
        .B(n13516), .ZN(n13518) );
  OAI21_X1 U15626 ( .B1(n13519), .B2(n13725), .A(n13518), .ZN(P2_U3235) );
  INV_X1 U15627 ( .A(n13521), .ZN(n13522) );
  NOR2_X1 U15628 ( .A1(n13522), .A2(n15292), .ZN(n13526) );
  OAI22_X1 U15629 ( .A1(n13689), .A2(n13524), .B1(n13523), .B2(n13683), .ZN(
        n13525) );
  AOI211_X1 U15630 ( .C1(n13527), .C2(n15297), .A(n13526), .B(n13525), .ZN(
        n13530) );
  NAND2_X1 U15631 ( .A1(n13528), .A2(n13652), .ZN(n13529) );
  OAI211_X1 U15632 ( .C1(n13520), .C2(n15301), .A(n13530), .B(n13529), .ZN(
        P2_U3236) );
  OAI211_X1 U15633 ( .C1(n13535), .C2(n13534), .A(n13533), .B(n13586), .ZN(
        n13537) );
  INV_X1 U15634 ( .A(n13731), .ZN(n13540) );
  OAI22_X1 U15635 ( .A1(n13732), .A2(n10061), .B1(n13538), .B2(n13683), .ZN(
        n13539) );
  OAI21_X1 U15636 ( .B1(n13540), .B2(n13539), .A(n13689), .ZN(n13548) );
  INV_X1 U15637 ( .A(n13555), .ZN(n13543) );
  INV_X1 U15638 ( .A(n13541), .ZN(n13542) );
  AOI211_X1 U15639 ( .C1(n13729), .C2(n13543), .A(n10861), .B(n13542), .ZN(
        n13728) );
  OAI22_X1 U15640 ( .A1(n13545), .A2(n15292), .B1(n13544), .B2(n13689), .ZN(
        n13546) );
  AOI21_X1 U15641 ( .B1(n13728), .B2(n15297), .A(n13546), .ZN(n13547) );
  OAI211_X1 U15642 ( .C1(n13732), .C2(n13618), .A(n13548), .B(n13547), .ZN(
        P2_U3237) );
  NAND2_X1 U15643 ( .A1(n13551), .A2(n13604), .ZN(n13553) );
  NAND2_X1 U15644 ( .A1(n13583), .A2(n13607), .ZN(n13552) );
  AOI211_X1 U15645 ( .C1(n13734), .C2(n13565), .A(n10861), .B(n13555), .ZN(
        n13733) );
  AOI22_X1 U15646 ( .A1(n15290), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13556), 
        .B2(n15288), .ZN(n13557) );
  OAI21_X1 U15647 ( .B1(n13558), .B2(n15292), .A(n13557), .ZN(n13559) );
  AOI21_X1 U15648 ( .B1(n13733), .B2(n15297), .A(n13559), .ZN(n13563) );
  NAND2_X1 U15649 ( .A1(n13561), .A2(n13560), .ZN(n13735) );
  NAND3_X1 U15650 ( .A1(n13736), .A2(n13735), .A3(n13652), .ZN(n13562) );
  OAI211_X1 U15651 ( .C1(n13740), .C2(n15301), .A(n13563), .B(n13562), .ZN(
        P2_U3238) );
  XNOR2_X1 U15652 ( .A(n13564), .B(n13574), .ZN(n13745) );
  INV_X1 U15653 ( .A(n13587), .ZN(n13567) );
  INV_X1 U15654 ( .A(n13565), .ZN(n13566) );
  AOI211_X1 U15655 ( .C1(n13742), .C2(n13567), .A(n10861), .B(n13566), .ZN(
        n13741) );
  INV_X1 U15656 ( .A(n13568), .ZN(n13569) );
  AOI22_X1 U15657 ( .A1(n15290), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13569), 
        .B2(n15288), .ZN(n13570) );
  OAI21_X1 U15658 ( .B1(n13571), .B2(n15292), .A(n13570), .ZN(n13578) );
  AOI222_X1 U15659 ( .A1(n13705), .A2(n13576), .B1(n13575), .B2(n13604), .C1(
        n13605), .C2(n13607), .ZN(n13744) );
  OAI21_X1 U15660 ( .B1(n13745), .B2(n15293), .A(n13579), .ZN(P2_U3239) );
  OR3_X1 U15661 ( .A1(n13601), .A2(n13594), .A3(n13580), .ZN(n13581) );
  NAND2_X1 U15662 ( .A1(n13582), .A2(n13581), .ZN(n13585) );
  AOI222_X1 U15663 ( .A1(n13586), .A2(n13585), .B1(n13584), .B2(n13607), .C1(
        n13583), .C2(n13604), .ZN(n13749) );
  AOI211_X1 U15664 ( .C1(n13747), .C2(n13612), .A(n10861), .B(n13587), .ZN(
        n13746) );
  INV_X1 U15665 ( .A(n13588), .ZN(n13589) );
  AOI22_X1 U15666 ( .A1(n15290), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13589), 
        .B2(n15288), .ZN(n13590) );
  OAI21_X1 U15667 ( .B1(n7492), .B2(n15292), .A(n13590), .ZN(n13596) );
  INV_X1 U15668 ( .A(n13591), .ZN(n13592) );
  AOI21_X1 U15669 ( .B1(n13594), .B2(n13593), .A(n13592), .ZN(n13750) );
  NOR2_X1 U15670 ( .A1(n13750), .A2(n15293), .ZN(n13595) );
  AOI211_X1 U15671 ( .C1(n13746), .C2(n15297), .A(n13596), .B(n13595), .ZN(
        n13597) );
  OAI21_X1 U15672 ( .B1(n6682), .B2(n15301), .A(n13597), .ZN(P2_U3240) );
  OR2_X1 U15673 ( .A1(n13598), .A2(n13602), .ZN(n13599) );
  AND2_X1 U15674 ( .A1(n13600), .A2(n13599), .ZN(n13617) );
  AOI21_X1 U15675 ( .B1(n13603), .B2(n13602), .A(n13601), .ZN(n13609) );
  AOI22_X1 U15676 ( .A1(n13607), .A2(n13606), .B1(n13605), .B2(n13604), .ZN(
        n13608) );
  OAI21_X1 U15677 ( .B1(n13609), .B2(n13676), .A(n13608), .ZN(n13610) );
  AOI21_X1 U15678 ( .B1(n13611), .B2(n13617), .A(n13610), .ZN(n13754) );
  INV_X1 U15679 ( .A(n13630), .ZN(n13613) );
  AOI211_X1 U15680 ( .C1(n13752), .C2(n13613), .A(n10861), .B(n7489), .ZN(
        n13751) );
  AOI22_X1 U15681 ( .A1(n15290), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13614), 
        .B2(n15288), .ZN(n13615) );
  OAI21_X1 U15682 ( .B1(n13616), .B2(n15292), .A(n13615), .ZN(n13620) );
  NOR2_X1 U15683 ( .A1(n13755), .A2(n13618), .ZN(n13619) );
  AOI211_X1 U15684 ( .C1(n13751), .C2(n15297), .A(n13620), .B(n13619), .ZN(
        n13621) );
  OAI21_X1 U15685 ( .B1(n13754), .B2(n15301), .A(n13621), .ZN(P2_U3241) );
  OR2_X1 U15686 ( .A1(n13622), .A2(n13626), .ZN(n13623) );
  NAND2_X1 U15687 ( .A1(n13624), .A2(n13623), .ZN(n13762) );
  AOI21_X1 U15688 ( .B1(n13627), .B2(n13626), .A(n13625), .ZN(n13628) );
  OAI222_X1 U15689 ( .A1(n13661), .A2(n13662), .B1(n13663), .B2(n13629), .C1(
        n13676), .C2(n13628), .ZN(n13757) );
  NAND2_X1 U15690 ( .A1(n13757), .A2(n13689), .ZN(n13636) );
  AOI211_X1 U15691 ( .C1(n13759), .C2(n13642), .A(n10861), .B(n13630), .ZN(
        n13758) );
  NOR2_X1 U15692 ( .A1(n7491), .A2(n15292), .ZN(n13634) );
  OAI22_X1 U15693 ( .A1(n13689), .A2(n13632), .B1(n13631), .B2(n13683), .ZN(
        n13633) );
  AOI211_X1 U15694 ( .C1(n13758), .C2(n15297), .A(n13634), .B(n13633), .ZN(
        n13635) );
  OAI211_X1 U15695 ( .C1(n13762), .C2(n15293), .A(n13636), .B(n13635), .ZN(
        P2_U3242) );
  AOI21_X1 U15696 ( .B1(n7541), .B2(n13638), .A(n13637), .ZN(n13639) );
  OAI222_X1 U15697 ( .A1(n13661), .A2(n13641), .B1(n13663), .B2(n13640), .C1(
        n13676), .C2(n13639), .ZN(n13763) );
  INV_X1 U15698 ( .A(n13765), .ZN(n13648) );
  AOI21_X1 U15699 ( .B1(n13665), .B2(n13765), .A(n10861), .ZN(n13643) );
  AND2_X1 U15700 ( .A1(n13643), .A2(n13642), .ZN(n13764) );
  NAND2_X1 U15701 ( .A1(n13764), .A2(n15297), .ZN(n13647) );
  INV_X1 U15702 ( .A(n13644), .ZN(n13645) );
  AOI22_X1 U15703 ( .A1(n13645), .A2(n15288), .B1(n15290), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n13646) );
  OAI211_X1 U15704 ( .C1(n13648), .C2(n15292), .A(n13647), .B(n13646), .ZN(
        n13649) );
  AOI21_X1 U15705 ( .B1(n13763), .B2(n13689), .A(n13649), .ZN(n13654) );
  NAND2_X1 U15706 ( .A1(n13651), .A2(n13650), .ZN(n13766) );
  NAND3_X1 U15707 ( .A1(n13767), .A2(n13766), .A3(n13652), .ZN(n13653) );
  NAND2_X1 U15708 ( .A1(n13654), .A2(n13653), .ZN(P2_U3243) );
  XNOR2_X1 U15709 ( .A(n13656), .B(n13655), .ZN(n13774) );
  XNOR2_X1 U15710 ( .A(n13658), .B(n13657), .ZN(n13659) );
  OAI222_X1 U15711 ( .A1(n13663), .A2(n13662), .B1(n13661), .B2(n13660), .C1(
        n13676), .C2(n13659), .ZN(n13770) );
  OR2_X1 U15712 ( .A1(n13680), .A2(n13669), .ZN(n13664) );
  AND3_X1 U15713 ( .A1(n13665), .A2(n10146), .A3(n13664), .ZN(n13771) );
  NAND2_X1 U15714 ( .A1(n13771), .A2(n15297), .ZN(n13668) );
  AOI22_X1 U15715 ( .A1(n15290), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13666), 
        .B2(n15288), .ZN(n13667) );
  OAI211_X1 U15716 ( .C1(n13669), .C2(n15292), .A(n13668), .B(n13667), .ZN(
        n13670) );
  AOI21_X1 U15717 ( .B1(n13770), .B2(n13689), .A(n13670), .ZN(n13671) );
  OAI21_X1 U15718 ( .B1(n15293), .B2(n13774), .A(n13671), .ZN(P2_U3244) );
  XNOR2_X1 U15719 ( .A(n13672), .B(n13674), .ZN(n13779) );
  XOR2_X1 U15720 ( .A(n13673), .B(n13674), .Z(n13677) );
  OAI21_X1 U15721 ( .B1(n13677), .B2(n13676), .A(n13675), .ZN(n13775) );
  NAND2_X1 U15722 ( .A1(n13696), .A2(n13777), .ZN(n13678) );
  NAND2_X1 U15723 ( .A1(n13678), .A2(n10146), .ZN(n13679) );
  NOR2_X1 U15724 ( .A1(n13680), .A2(n13679), .ZN(n13776) );
  NAND2_X1 U15725 ( .A1(n13776), .A2(n15297), .ZN(n13687) );
  NAND2_X1 U15726 ( .A1(n15290), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n13681) );
  OAI21_X1 U15727 ( .B1(n13683), .B2(n13682), .A(n13681), .ZN(n13684) );
  AOI21_X1 U15728 ( .B1(n13777), .B2(n13685), .A(n13684), .ZN(n13686) );
  NAND2_X1 U15729 ( .A1(n13687), .A2(n13686), .ZN(n13688) );
  AOI21_X1 U15730 ( .B1(n13775), .B2(n13689), .A(n13688), .ZN(n13690) );
  OAI21_X1 U15731 ( .B1(n13779), .B2(n15293), .A(n13690), .ZN(P2_U3245) );
  XOR2_X1 U15732 ( .A(n13692), .B(n13691), .Z(n13785) );
  XNOR2_X1 U15733 ( .A(n13693), .B(n13692), .ZN(n13694) );
  NAND2_X1 U15734 ( .A1(n13694), .A2(n13705), .ZN(n13783) );
  INV_X1 U15735 ( .A(n13783), .ZN(n13695) );
  OAI21_X1 U15736 ( .B1(n13695), .B2(n13781), .A(n13689), .ZN(n13703) );
  INV_X1 U15737 ( .A(n13696), .ZN(n13697) );
  AOI211_X1 U15738 ( .C1(n13782), .C2(n13708), .A(n10861), .B(n13697), .ZN(
        n13780) );
  AOI22_X1 U15739 ( .A1(n15290), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13698), 
        .B2(n15288), .ZN(n13699) );
  OAI21_X1 U15740 ( .B1(n13700), .B2(n15292), .A(n13699), .ZN(n13701) );
  AOI21_X1 U15741 ( .B1(n13780), .B2(n15297), .A(n13701), .ZN(n13702) );
  OAI211_X1 U15742 ( .C1(n13785), .C2(n15293), .A(n13703), .B(n13702), .ZN(
        P2_U3246) );
  XNOR2_X1 U15743 ( .A(n13704), .B(n13719), .ZN(n13706) );
  NAND2_X1 U15744 ( .A1(n13706), .A2(n13705), .ZN(n13788) );
  INV_X1 U15745 ( .A(n13707), .ZN(n13709) );
  OAI211_X1 U15746 ( .C1(n13715), .C2(n13709), .A(n10146), .B(n13708), .ZN(
        n13711) );
  NAND2_X1 U15747 ( .A1(n13711), .A2(n13710), .ZN(n13786) );
  INV_X1 U15748 ( .A(n13712), .ZN(n13713) );
  AOI22_X1 U15749 ( .A1(n15290), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13713), 
        .B2(n15288), .ZN(n13714) );
  OAI21_X1 U15750 ( .B1(n13715), .B2(n15292), .A(n13714), .ZN(n13721) );
  INV_X1 U15751 ( .A(n13716), .ZN(n13717) );
  AOI21_X1 U15752 ( .B1(n13719), .B2(n13718), .A(n13717), .ZN(n13790) );
  NOR2_X1 U15753 ( .A1(n13790), .A2(n15293), .ZN(n13720) );
  AOI211_X1 U15754 ( .C1(n15297), .C2(n13786), .A(n13721), .B(n13720), .ZN(
        n13722) );
  OAI21_X1 U15755 ( .B1(n15290), .B2(n13788), .A(n13722), .ZN(P2_U3247) );
  OAI211_X1 U15756 ( .C1(n7487), .C2(n15342), .A(n13723), .B(n13724), .ZN(
        n13817) );
  MUX2_X1 U15757 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13817), .S(n13815), .Z(
        P2_U3530) );
  OAI211_X1 U15758 ( .C1(n13726), .C2(n15342), .A(n13725), .B(n13724), .ZN(
        n13818) );
  MUX2_X1 U15759 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13818), .S(n13815), .Z(
        P2_U3529) );
  AOI21_X1 U15760 ( .B1(n15356), .B2(n13729), .A(n13728), .ZN(n13730) );
  OAI211_X1 U15761 ( .C1(n15360), .C2(n13732), .A(n13731), .B(n13730), .ZN(
        n13819) );
  MUX2_X1 U15762 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13819), .S(n13815), .Z(
        P2_U3527) );
  AOI21_X1 U15763 ( .B1(n15356), .B2(n13734), .A(n13733), .ZN(n13738) );
  NAND3_X1 U15764 ( .A1(n13736), .A2(n13735), .A3(n15339), .ZN(n13737) );
  MUX2_X1 U15765 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13820), .S(n13815), .Z(
        P2_U3526) );
  AOI21_X1 U15766 ( .B1(n15356), .B2(n13742), .A(n13741), .ZN(n13743) );
  OAI211_X1 U15767 ( .C1(n15360), .C2(n13745), .A(n13744), .B(n13743), .ZN(
        n13821) );
  MUX2_X1 U15768 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13821), .S(n13815), .Z(
        P2_U3525) );
  AOI21_X1 U15769 ( .B1(n15356), .B2(n13747), .A(n13746), .ZN(n13748) );
  OAI211_X1 U15770 ( .C1(n15360), .C2(n13750), .A(n6682), .B(n13748), .ZN(
        n13822) );
  MUX2_X1 U15771 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13822), .S(n13815), .Z(
        P2_U3524) );
  AOI21_X1 U15772 ( .B1(n15356), .B2(n13752), .A(n13751), .ZN(n13753) );
  OAI211_X1 U15773 ( .C1(n13756), .C2(n13755), .A(n13754), .B(n13753), .ZN(
        n13823) );
  MUX2_X1 U15774 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13823), .S(n13815), .Z(
        P2_U3523) );
  INV_X1 U15775 ( .A(n13757), .ZN(n13761) );
  AOI21_X1 U15776 ( .B1(n15356), .B2(n13759), .A(n13758), .ZN(n13760) );
  OAI211_X1 U15777 ( .C1(n15360), .C2(n13762), .A(n13761), .B(n13760), .ZN(
        n13824) );
  MUX2_X1 U15778 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13824), .S(n13815), .Z(
        P2_U3522) );
  AOI211_X1 U15779 ( .C1(n15356), .C2(n13765), .A(n13764), .B(n13763), .ZN(
        n13769) );
  NAND3_X1 U15780 ( .A1(n13767), .A2(n13766), .A3(n15339), .ZN(n13768) );
  NAND2_X1 U15781 ( .A1(n13769), .A2(n13768), .ZN(n13825) );
  MUX2_X1 U15782 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13825), .S(n13815), .Z(
        P2_U3521) );
  AOI211_X1 U15783 ( .C1(n15356), .C2(n13772), .A(n13771), .B(n13770), .ZN(
        n13773) );
  OAI21_X1 U15784 ( .B1(n15360), .B2(n13774), .A(n13773), .ZN(n13826) );
  MUX2_X1 U15785 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13826), .S(n13815), .Z(
        P2_U3520) );
  AOI211_X1 U15786 ( .C1(n15356), .C2(n13777), .A(n13776), .B(n13775), .ZN(
        n13778) );
  OAI21_X1 U15787 ( .B1(n15360), .B2(n13779), .A(n13778), .ZN(n13827) );
  MUX2_X1 U15788 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13827), .S(n13815), .Z(
        P2_U3519) );
  AOI211_X1 U15789 ( .C1(n15356), .C2(n13782), .A(n13781), .B(n13780), .ZN(
        n13784) );
  OAI211_X1 U15790 ( .C1(n15360), .C2(n13785), .A(n13784), .B(n13783), .ZN(
        n13828) );
  MUX2_X1 U15791 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13828), .S(n13815), .Z(
        P2_U3518) );
  AOI21_X1 U15792 ( .B1(n15356), .B2(n13787), .A(n13786), .ZN(n13789) );
  OAI211_X1 U15793 ( .C1(n13790), .C2(n15360), .A(n13789), .B(n13788), .ZN(
        n13829) );
  MUX2_X1 U15794 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13829), .S(n13815), .Z(
        P2_U3517) );
  OAI21_X1 U15795 ( .B1(n13792), .B2(n15342), .A(n13791), .ZN(n13793) );
  AOI21_X1 U15796 ( .B1(n13794), .B2(n15339), .A(n13793), .ZN(n13795) );
  NAND2_X1 U15797 ( .A1(n13796), .A2(n13795), .ZN(n13830) );
  MUX2_X1 U15798 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13830), .S(n13815), .Z(
        P2_U3516) );
  AOI21_X1 U15799 ( .B1(n15356), .B2(n13798), .A(n13797), .ZN(n13802) );
  NAND3_X1 U15800 ( .A1(n13800), .A2(n13799), .A3(n15339), .ZN(n13801) );
  NAND3_X1 U15801 ( .A1(n13803), .A2(n13802), .A3(n13801), .ZN(n13831) );
  MUX2_X1 U15802 ( .A(n13831), .B(P2_REG1_REG_16__SCAN_IN), .S(n15371), .Z(
        P2_U3515) );
  AOI21_X1 U15803 ( .B1(n15356), .B2(n13805), .A(n13804), .ZN(n13806) );
  OAI211_X1 U15804 ( .C1(n15360), .C2(n13808), .A(n13807), .B(n13806), .ZN(
        n13832) );
  MUX2_X1 U15805 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13832), .S(n13815), .Z(
        P2_U3514) );
  AOI211_X1 U15806 ( .C1(n15356), .C2(n13811), .A(n13810), .B(n13809), .ZN(
        n13812) );
  OAI21_X1 U15807 ( .B1(n15360), .B2(n13813), .A(n13812), .ZN(n13833) );
  MUX2_X1 U15808 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13833), .S(n13815), .Z(
        P2_U3513) );
  MUX2_X1 U15809 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n13814), .S(n13815), .Z(
        P2_U3507) );
  MUX2_X1 U15810 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n13816), .S(n13815), .Z(
        P2_U3499) );
  MUX2_X1 U15811 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13817), .S(n15364), .Z(
        P2_U3498) );
  MUX2_X1 U15812 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13818), .S(n15364), .Z(
        P2_U3497) );
  MUX2_X1 U15813 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13819), .S(n15364), .Z(
        P2_U3495) );
  MUX2_X1 U15814 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13820), .S(n15364), .Z(
        P2_U3494) );
  MUX2_X1 U15815 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13821), .S(n15364), .Z(
        P2_U3493) );
  MUX2_X1 U15816 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13822), .S(n15364), .Z(
        P2_U3492) );
  MUX2_X1 U15817 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13823), .S(n15364), .Z(
        P2_U3491) );
  MUX2_X1 U15818 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13824), .S(n15364), .Z(
        P2_U3490) );
  MUX2_X1 U15819 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13825), .S(n15364), .Z(
        P2_U3489) );
  MUX2_X1 U15820 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13826), .S(n15364), .Z(
        P2_U3488) );
  MUX2_X1 U15821 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13827), .S(n15364), .Z(
        P2_U3487) );
  MUX2_X1 U15822 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13828), .S(n15364), .Z(
        P2_U3486) );
  MUX2_X1 U15823 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13829), .S(n15364), .Z(
        P2_U3484) );
  MUX2_X1 U15824 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13830), .S(n15364), .Z(
        P2_U3481) );
  MUX2_X1 U15825 ( .A(n13831), .B(P2_REG0_REG_16__SCAN_IN), .S(n15362), .Z(
        P2_U3478) );
  MUX2_X1 U15826 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13832), .S(n15364), .Z(
        P2_U3475) );
  MUX2_X1 U15827 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13833), .S(n15364), .Z(
        P2_U3472) );
  NAND3_X1 U15828 ( .A1(n13835), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13837) );
  OAI22_X1 U15829 ( .A1(n13834), .A2(n13837), .B1(n13836), .B2(n13844), .ZN(
        n13838) );
  AOI21_X1 U15830 ( .B1(n14376), .B2(n13840), .A(n13838), .ZN(n13839) );
  INV_X1 U15831 ( .A(n13839), .ZN(P2_U3296) );
  NAND2_X1 U15832 ( .A1(n14387), .A2(n13840), .ZN(n13842) );
  OAI211_X1 U15833 ( .C1(n13844), .C2(n14552), .A(n13842), .B(n13841), .ZN(
        P2_U3299) );
  INV_X1 U15834 ( .A(n13843), .ZN(n14393) );
  OAI222_X1 U15835 ( .A1(n13846), .A2(P2_U3088), .B1(n13850), .B2(n14393), 
        .C1(n13845), .C2(n13844), .ZN(P2_U3301) );
  INV_X1 U15836 ( .A(n13847), .ZN(n14397) );
  OAI222_X1 U15837 ( .A1(n13852), .A2(n13851), .B1(n13850), .B2(n14397), .C1(
        n13849), .C2(P2_U3088), .ZN(P2_U3302) );
  MUX2_X1 U15838 ( .A(n13853), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15839 ( .A(n13855), .B(n13854), .Z(n13861) );
  NOR2_X1 U15840 ( .A1(n14964), .A2(n14101), .ZN(n13859) );
  AOI22_X1 U15841 ( .A1(n14954), .A2(n14095), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13856) );
  OAI21_X1 U15842 ( .B1(n13857), .B2(n14910), .A(n13856), .ZN(n13858) );
  AOI211_X1 U15843 ( .C1(n14285), .C2(n14921), .A(n13859), .B(n13858), .ZN(
        n13860) );
  OAI21_X1 U15844 ( .B1(n13861), .B2(n14916), .A(n13860), .ZN(P1_U3214) );
  XOR2_X1 U15845 ( .A(n13863), .B(n13862), .Z(n13868) );
  NOR2_X1 U15846 ( .A1(n14964), .A2(n14160), .ZN(n13866) );
  AOI22_X1 U15847 ( .A1(n14954), .A2(n14157), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13864) );
  OAI21_X1 U15848 ( .B1(n13881), .B2(n14910), .A(n13864), .ZN(n13865) );
  AOI211_X1 U15849 ( .C1(n14313), .C2(n14921), .A(n13866), .B(n13865), .ZN(
        n13867) );
  OAI21_X1 U15850 ( .B1(n13868), .B2(n14916), .A(n13867), .ZN(P1_U3216) );
  OAI211_X1 U15851 ( .C1(n13871), .C2(n13870), .A(n13869), .B(n14960), .ZN(
        n13876) );
  NOR2_X1 U15852 ( .A1(n13872), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14051) );
  AOI21_X1 U15853 ( .B1(n14956), .B2(n14222), .A(n14051), .ZN(n13873) );
  OAI21_X1 U15854 ( .B1(n14221), .B2(n14909), .A(n13873), .ZN(n13874) );
  AOI21_X1 U15855 ( .B1(n14225), .B2(n13939), .A(n13874), .ZN(n13875) );
  OAI211_X1 U15856 ( .C1(n14335), .C2(n14958), .A(n13876), .B(n13875), .ZN(
        P1_U3219) );
  INV_X1 U15857 ( .A(n13877), .ZN(n13878) );
  AOI21_X1 U15858 ( .B1(n13880), .B2(n13879), .A(n13878), .ZN(n13885) );
  OAI22_X1 U15859 ( .A1(n13881), .A2(n14220), .B1(n14221), .B2(n14265), .ZN(
        n14186) );
  INV_X1 U15860 ( .A(n13949), .ZN(n14934) );
  AOI22_X1 U15861 ( .A1(n14186), .A2(n14934), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13882) );
  OAI21_X1 U15862 ( .B1(n14964), .B2(n14188), .A(n13882), .ZN(n13883) );
  AOI21_X1 U15863 ( .B1(n14324), .B2(n14921), .A(n13883), .ZN(n13884) );
  OAI21_X1 U15864 ( .B1(n13885), .B2(n14916), .A(n13884), .ZN(P1_U3223) );
  XOR2_X1 U15865 ( .A(n13887), .B(n13886), .Z(n13893) );
  NAND2_X1 U15866 ( .A1(n14812), .A2(n14094), .ZN(n13889) );
  NAND2_X1 U15867 ( .A1(n14979), .A2(n14157), .ZN(n13888) );
  NAND2_X1 U15868 ( .A1(n13889), .A2(n13888), .ZN(n14125) );
  AOI22_X1 U15869 ( .A1(n14934), .A2(n14125), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13890) );
  OAI21_X1 U15870 ( .B1(n14964), .B2(n14126), .A(n13890), .ZN(n13891) );
  AOI21_X1 U15871 ( .B1(n14131), .B2(n14921), .A(n13891), .ZN(n13892) );
  OAI21_X1 U15872 ( .B1(n13893), .B2(n14916), .A(n13892), .ZN(P1_U3225) );
  OAI21_X1 U15873 ( .B1(n13896), .B2(n13895), .A(n13894), .ZN(n13897) );
  NAND2_X1 U15874 ( .A1(n13897), .A2(n14960), .ZN(n13903) );
  OAI21_X1 U15875 ( .B1(n14910), .B2(n14908), .A(n13898), .ZN(n13901) );
  NOR2_X1 U15876 ( .A1(n14964), .A2(n13899), .ZN(n13900) );
  AOI211_X1 U15877 ( .C1(n14954), .C2(n14237), .A(n13901), .B(n13900), .ZN(
        n13902) );
  OAI211_X1 U15878 ( .C1(n14967), .C2(n14958), .A(n13903), .B(n13902), .ZN(
        P1_U3226) );
  XOR2_X1 U15879 ( .A(n13905), .B(n13904), .Z(n13914) );
  OAI21_X1 U15880 ( .B1(n14909), .B2(n13907), .A(n13906), .ZN(n13908) );
  AOI21_X1 U15881 ( .B1(n14956), .B2(n14953), .A(n13908), .ZN(n13909) );
  OAI21_X1 U15882 ( .B1(n14964), .B2(n13910), .A(n13909), .ZN(n13911) );
  AOI21_X1 U15883 ( .B1(n13912), .B2(n14921), .A(n13911), .ZN(n13913) );
  OAI21_X1 U15884 ( .B1(n13914), .B2(n14916), .A(n13913), .ZN(P1_U3228) );
  XOR2_X1 U15885 ( .A(n13916), .B(n13915), .Z(n13921) );
  NOR2_X1 U15886 ( .A1(n14964), .A2(n14146), .ZN(n13919) );
  AOI22_X1 U15887 ( .A1(n14954), .A2(n13955), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13917) );
  OAI21_X1 U15888 ( .B1(n14137), .B2(n14910), .A(n13917), .ZN(n13918) );
  AOI211_X1 U15889 ( .C1(n14308), .C2(n14921), .A(n13919), .B(n13918), .ZN(
        n13920) );
  OAI21_X1 U15890 ( .B1(n13921), .B2(n14916), .A(n13920), .ZN(P1_U3229) );
  OAI211_X1 U15891 ( .C1(n13924), .C2(n13923), .A(n13922), .B(n14960), .ZN(
        n13928) );
  AOI22_X1 U15892 ( .A1(n14956), .A2(n14238), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13925) );
  OAI21_X1 U15893 ( .B1(n14200), .B2(n14909), .A(n13925), .ZN(n13926) );
  AOI21_X1 U15894 ( .B1(n14205), .B2(n13939), .A(n13926), .ZN(n13927) );
  OAI211_X1 U15895 ( .C1(n14212), .C2(n14958), .A(n13928), .B(n13927), .ZN(
        P1_U3233) );
  OAI21_X1 U15896 ( .B1(n13931), .B2(n13930), .A(n13929), .ZN(n13932) );
  NAND2_X1 U15897 ( .A1(n13932), .A2(n14960), .ZN(n13936) );
  AOI22_X1 U15898 ( .A1(n14956), .A2(n14175), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13933) );
  OAI21_X1 U15899 ( .B1(n14137), .B2(n14909), .A(n13933), .ZN(n13934) );
  AOI21_X1 U15900 ( .B1(n14176), .B2(n13939), .A(n13934), .ZN(n13935) );
  OAI211_X1 U15901 ( .C1(n14958), .C2(n7369), .A(n13936), .B(n13935), .ZN(
        P1_U3235) );
  XOR2_X1 U15902 ( .A(n13938), .B(n13937), .Z(n13946) );
  NAND2_X1 U15903 ( .A1(n13939), .A2(n14245), .ZN(n13942) );
  NOR2_X1 U15904 ( .A1(n13940), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14018) );
  AOI21_X1 U15905 ( .B1(n14954), .B2(n14238), .A(n14018), .ZN(n13941) );
  OAI211_X1 U15906 ( .C1(n13943), .C2(n14910), .A(n13942), .B(n13941), .ZN(
        n13944) );
  AOI21_X1 U15907 ( .B1(n14342), .B2(n14921), .A(n13944), .ZN(n13945) );
  OAI21_X1 U15908 ( .B1(n13946), .B2(n14916), .A(n13945), .ZN(P1_U3238) );
  XOR2_X1 U15909 ( .A(n13948), .B(n13947), .Z(n13953) );
  NOR2_X1 U15910 ( .A1(n14964), .A2(n14113), .ZN(n13951) );
  AOI22_X1 U15911 ( .A1(n14812), .A2(n14069), .B1(n14979), .B2(n13955), .ZN(
        n14292) );
  OAI22_X1 U15912 ( .A1(n13949), .A2(n14292), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14599), .ZN(n13950) );
  AOI211_X1 U15913 ( .C1(n14112), .C2(n14921), .A(n13951), .B(n13950), .ZN(
        n13952) );
  OAI21_X1 U15914 ( .B1(n13953), .B2(n14916), .A(n13952), .ZN(P1_U3240) );
  MUX2_X1 U15915 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14056), .S(n13967), .Z(
        P1_U3591) );
  MUX2_X1 U15916 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13954), .S(n13967), .Z(
        P1_U3590) );
  MUX2_X1 U15917 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14070), .S(n13967), .Z(
        P1_U3589) );
  MUX2_X1 U15918 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14095), .S(n13967), .Z(
        P1_U3588) );
  MUX2_X1 U15919 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14069), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15920 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14094), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15921 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13955), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15922 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14157), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15923 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14174), .S(n13967), .Z(
        P1_U3583) );
  MUX2_X1 U15924 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14156), .S(n13967), .Z(
        P1_U3582) );
  MUX2_X1 U15925 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14175), .S(n13967), .Z(
        P1_U3581) );
  MUX2_X1 U15926 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13956), .S(n13967), .Z(
        P1_U3580) );
  MUX2_X1 U15927 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14238), .S(n13967), .Z(
        P1_U3579) );
  MUX2_X1 U15928 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14222), .S(n13967), .Z(
        P1_U3578) );
  MUX2_X1 U15929 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14237), .S(n13967), .Z(
        P1_U3577) );
  MUX2_X1 U15930 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14953), .S(n13967), .Z(
        P1_U3576) );
  MUX2_X1 U15931 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13957), .S(n13967), .Z(
        P1_U3575) );
  MUX2_X1 U15932 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14955), .S(n13967), .Z(
        P1_U3574) );
  MUX2_X1 U15933 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13958), .S(n13967), .Z(
        P1_U3573) );
  MUX2_X1 U15934 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14978), .S(n13967), .Z(
        P1_U3572) );
  MUX2_X1 U15935 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13959), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15936 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14943), .S(n13967), .Z(
        P1_U3570) );
  MUX2_X1 U15937 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14927), .S(n13967), .Z(
        P1_U3569) );
  MUX2_X1 U15938 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13960), .S(n13967), .Z(
        P1_U3568) );
  MUX2_X1 U15939 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13961), .S(n13967), .Z(
        P1_U3567) );
  MUX2_X1 U15940 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13962), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15941 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13963), .S(n13967), .Z(
        P1_U3565) );
  MUX2_X1 U15942 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13964), .S(n13967), .Z(
        P1_U3564) );
  MUX2_X1 U15943 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13965), .S(n13967), .Z(
        P1_U3563) );
  MUX2_X1 U15944 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14267), .S(n13967), .Z(
        P1_U3562) );
  MUX2_X1 U15945 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13966), .S(n13967), .Z(
        P1_U3561) );
  MUX2_X1 U15946 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14262), .S(n13967), .Z(
        P1_U3560) );
  NOR2_X1 U15947 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14623), .ZN(n13970) );
  NOR2_X1 U15948 ( .A1(n15054), .A2(n13968), .ZN(n13969) );
  AOI211_X1 U15949 ( .C1(n15031), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n13970), .B(
        n13969), .ZN(n13981) );
  OAI211_X1 U15950 ( .C1(n13973), .C2(n13972), .A(n15059), .B(n13971), .ZN(
        n13980) );
  INV_X1 U15951 ( .A(n13986), .ZN(n13978) );
  NAND3_X1 U15952 ( .A1(n13976), .A2(n13975), .A3(n13974), .ZN(n13977) );
  NAND3_X1 U15953 ( .A1(n15044), .A2(n13978), .A3(n13977), .ZN(n13979) );
  NAND3_X1 U15954 ( .A1(n13981), .A2(n13980), .A3(n13979), .ZN(P1_U3246) );
  INV_X1 U15955 ( .A(n13982), .ZN(n13990) );
  INV_X1 U15956 ( .A(n13983), .ZN(n13988) );
  NOR3_X1 U15957 ( .A1(n13986), .A2(n13985), .A3(n13984), .ZN(n13987) );
  NOR3_X1 U15958 ( .A1(n15056), .A2(n13988), .A3(n13987), .ZN(n13989) );
  AOI211_X1 U15959 ( .C1(n15031), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n13990), .B(
        n13989), .ZN(n13998) );
  NAND2_X1 U15960 ( .A1(n15042), .A2(n13991), .ZN(n13997) );
  INV_X1 U15961 ( .A(n13992), .ZN(n13993) );
  OAI211_X1 U15962 ( .C1(n13995), .C2(n13994), .A(n15059), .B(n13993), .ZN(
        n13996) );
  NAND4_X1 U15963 ( .A1(n13999), .A2(n13998), .A3(n13997), .A4(n13996), .ZN(
        P1_U3247) );
  OAI21_X1 U15964 ( .B1(n14002), .B2(n14001), .A(n14000), .ZN(n14003) );
  NAND2_X1 U15965 ( .A1(n14003), .A2(n15059), .ZN(n14016) );
  NOR2_X1 U15966 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14004), .ZN(n14005) );
  AOI21_X1 U15967 ( .B1(n15031), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n14005), .ZN(
        n14015) );
  INV_X1 U15968 ( .A(n14006), .ZN(n14008) );
  MUX2_X1 U15969 ( .A(n10524), .B(P1_REG2_REG_8__SCAN_IN), .S(n14012), .Z(
        n14007) );
  NAND3_X1 U15970 ( .A1(n14009), .A2(n14008), .A3(n14007), .ZN(n14010) );
  NAND3_X1 U15971 ( .A1(n15044), .A2(n14011), .A3(n14010), .ZN(n14014) );
  NAND2_X1 U15972 ( .A1(n15042), .A2(n14012), .ZN(n14013) );
  NAND4_X1 U15973 ( .A1(n14016), .A2(n14015), .A3(n14014), .A4(n14013), .ZN(
        P1_U3251) );
  NOR2_X1 U15974 ( .A1(n15054), .A2(n14035), .ZN(n14017) );
  AOI211_X1 U15975 ( .C1(n15031), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n14018), 
        .B(n14017), .ZN(n14034) );
  INV_X1 U15976 ( .A(n14019), .ZN(n14020) );
  NAND2_X1 U15977 ( .A1(n14021), .A2(n14020), .ZN(n14022) );
  OAI21_X1 U15978 ( .B1(n14024), .B2(n14023), .A(n14022), .ZN(n14040) );
  XNOR2_X1 U15979 ( .A(n14035), .B(n14040), .ZN(n14025) );
  NAND2_X1 U15980 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14025), .ZN(n14043) );
  OAI211_X1 U15981 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14025), .A(n15044), 
        .B(n14043), .ZN(n14033) );
  XNOR2_X1 U15982 ( .A(n14035), .B(n14036), .ZN(n14028) );
  INV_X1 U15983 ( .A(n14028), .ZN(n14031) );
  NOR2_X1 U15984 ( .A1(n14029), .A2(n14028), .ZN(n14038) );
  INV_X1 U15985 ( .A(n14038), .ZN(n14030) );
  OAI211_X1 U15986 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14031), .A(n15059), 
        .B(n14030), .ZN(n14032) );
  NAND3_X1 U15987 ( .A1(n14034), .A2(n14033), .A3(n14032), .ZN(P1_U3261) );
  NOR2_X1 U15988 ( .A1(n14036), .A2(n14035), .ZN(n14037) );
  NOR2_X1 U15989 ( .A1(n14038), .A2(n14037), .ZN(n14039) );
  XNOR2_X1 U15990 ( .A(n14039), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14048) );
  INV_X1 U15991 ( .A(n14048), .ZN(n14046) );
  NAND2_X1 U15992 ( .A1(n14041), .A2(n14040), .ZN(n14042) );
  NAND2_X1 U15993 ( .A1(n14043), .A2(n14042), .ZN(n14044) );
  XOR2_X1 U15994 ( .A(n14044), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14047) );
  OAI21_X1 U15995 ( .B1(n14047), .B2(n15056), .A(n15054), .ZN(n14045) );
  AOI21_X1 U15996 ( .B1(n14046), .B2(n15059), .A(n14045), .ZN(n14050) );
  AOI22_X1 U15997 ( .A1(n14048), .A2(n15059), .B1(n15044), .B2(n14047), .ZN(
        n14049) );
  MUX2_X1 U15998 ( .A(n14050), .B(n14049), .S(n14206), .Z(n14053) );
  AOI21_X1 U15999 ( .B1(n15031), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n14051), 
        .ZN(n14052) );
  NAND2_X1 U16000 ( .A1(n14053), .A2(n14052), .ZN(P1_U3262) );
  NOR2_X1 U16001 ( .A1(n14054), .A2(n14060), .ZN(n14061) );
  XOR2_X1 U16002 ( .A(n6685), .B(n14061), .Z(n14055) );
  NAND2_X1 U16003 ( .A1(n14055), .A2(n15111), .ZN(n14273) );
  NAND2_X1 U16004 ( .A1(n14057), .A2(n14056), .ZN(n14275) );
  NOR2_X1 U16005 ( .A1(n14251), .A2(n14275), .ZN(n14064) );
  NOR2_X1 U16006 ( .A1(n6685), .A2(n15107), .ZN(n14058) );
  AOI211_X1 U16007 ( .C1(n14251), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14064), 
        .B(n14058), .ZN(n14059) );
  OAI21_X1 U16008 ( .B1(n14273), .B2(n14816), .A(n14059), .ZN(P1_U3263) );
  INV_X1 U16009 ( .A(n14060), .ZN(n14063) );
  INV_X1 U16010 ( .A(n14061), .ZN(n14062) );
  OAI211_X1 U16011 ( .C1(n14277), .C2(n14063), .A(n14062), .B(n15111), .ZN(
        n14276) );
  NAND2_X1 U16012 ( .A1(n15105), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14066) );
  INV_X1 U16013 ( .A(n14064), .ZN(n14065) );
  OAI211_X1 U16014 ( .C1(n14277), .C2(n15107), .A(n14066), .B(n14065), .ZN(
        n14067) );
  INV_X1 U16015 ( .A(n14067), .ZN(n14068) );
  OAI21_X1 U16016 ( .B1(n14276), .B2(n14816), .A(n14068), .ZN(P1_U3264) );
  OAI21_X1 U16017 ( .B1(n14077), .B2(n14072), .A(n14071), .ZN(n14073) );
  AOI21_X1 U16018 ( .B1(n14077), .B2(n14076), .A(n14075), .ZN(n14278) );
  AND2_X1 U16019 ( .A1(n14279), .A2(n14099), .ZN(n14078) );
  NAND2_X1 U16020 ( .A1(n15105), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14080) );
  OAI21_X1 U16021 ( .B1(n14801), .B2(n14081), .A(n14080), .ZN(n14082) );
  AOI21_X1 U16022 ( .B1(n14279), .B2(n14255), .A(n14082), .ZN(n14083) );
  OAI21_X1 U16023 ( .B1(n14281), .B2(n14816), .A(n14083), .ZN(n14084) );
  AOI21_X1 U16024 ( .B1(n14278), .B2(n14809), .A(n14084), .ZN(n14085) );
  OAI21_X1 U16025 ( .B1(n14284), .B2(n15105), .A(n14085), .ZN(P1_U3265) );
  OR2_X1 U16026 ( .A1(n14090), .A2(n14086), .ZN(n14087) );
  NAND2_X1 U16027 ( .A1(n14088), .A2(n14087), .ZN(n14289) );
  NAND2_X1 U16028 ( .A1(n14289), .A2(n15102), .ZN(n14098) );
  NAND2_X1 U16029 ( .A1(n14090), .A2(n14089), .ZN(n14091) );
  NAND2_X1 U16030 ( .A1(n14092), .A2(n14091), .ZN(n14093) );
  NAND2_X1 U16031 ( .A1(n14093), .A2(n15098), .ZN(n14097) );
  AOI22_X1 U16032 ( .A1(n14812), .A2(n14095), .B1(n14979), .B2(n14094), .ZN(
        n14096) );
  AOI21_X1 U16033 ( .B1(n14285), .B2(n14111), .A(n15125), .ZN(n14100) );
  NAND2_X1 U16034 ( .A1(n14100), .A2(n14099), .ZN(n14287) );
  INV_X1 U16035 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14102) );
  OAI22_X1 U16036 ( .A1(n14804), .A2(n14102), .B1(n14101), .B2(n14801), .ZN(
        n14103) );
  AOI21_X1 U16037 ( .B1(n14285), .B2(n14255), .A(n14103), .ZN(n14104) );
  OAI21_X1 U16038 ( .B1(n14287), .B2(n14164), .A(n14104), .ZN(n14105) );
  AOI21_X1 U16039 ( .B1(n15114), .B2(n14289), .A(n14105), .ZN(n14106) );
  OAI21_X1 U16040 ( .B1(n14291), .B2(n14251), .A(n14106), .ZN(P1_U3266) );
  XNOR2_X1 U16041 ( .A(n14108), .B(n14107), .ZN(n14298) );
  OAI21_X1 U16042 ( .B1(n7276), .B2(n14110), .A(n14109), .ZN(n14296) );
  INV_X1 U16043 ( .A(n14112), .ZN(n14293) );
  AOI211_X1 U16044 ( .C1(n14112), .C2(n14124), .A(n15125), .B(n7367), .ZN(
        n14294) );
  NAND2_X1 U16045 ( .A1(n14294), .A2(n15113), .ZN(n14116) );
  OAI22_X1 U16046 ( .A1(n15105), .A2(n14292), .B1(n14113), .B2(n14801), .ZN(
        n14114) );
  AOI21_X1 U16047 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n15105), .A(n14114), 
        .ZN(n14115) );
  OAI211_X1 U16048 ( .C1(n14293), .C2(n15107), .A(n14116), .B(n14115), .ZN(
        n14117) );
  AOI21_X1 U16049 ( .B1(n14182), .B2(n14296), .A(n14117), .ZN(n14118) );
  OAI21_X1 U16050 ( .B1(n14298), .B2(n14210), .A(n14118), .ZN(P1_U3267) );
  XNOR2_X1 U16051 ( .A(n14119), .B(n14123), .ZN(n14305) );
  INV_X1 U16052 ( .A(n14120), .ZN(n14121) );
  AOI21_X1 U16053 ( .B1(n14123), .B2(n14122), .A(n14121), .ZN(n14303) );
  OAI211_X1 U16054 ( .C1(n14301), .C2(n14145), .A(n15111), .B(n14124), .ZN(
        n14300) );
  INV_X1 U16055 ( .A(n14125), .ZN(n14299) );
  OAI21_X1 U16056 ( .B1(n14801), .B2(n14126), .A(n14299), .ZN(n14127) );
  INV_X1 U16057 ( .A(n14127), .ZN(n14129) );
  NAND2_X1 U16058 ( .A1(n15105), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14128) );
  OAI21_X1 U16059 ( .B1(n14251), .B2(n14129), .A(n14128), .ZN(n14130) );
  AOI21_X1 U16060 ( .B1(n14131), .B2(n14255), .A(n14130), .ZN(n14132) );
  OAI21_X1 U16061 ( .B1(n14300), .B2(n14816), .A(n14132), .ZN(n14133) );
  AOI21_X1 U16062 ( .B1(n14303), .B2(n14809), .A(n14133), .ZN(n14134) );
  OAI21_X1 U16063 ( .B1(n14233), .B2(n14305), .A(n14134), .ZN(P1_U3268) );
  OAI21_X1 U16064 ( .B1(n14136), .B2(n14142), .A(n14135), .ZN(n14306) );
  OAI22_X1 U16065 ( .A1(n14138), .A2(n14220), .B1(n14137), .B2(n14265), .ZN(
        n14144) );
  INV_X1 U16066 ( .A(n6854), .ZN(n14140) );
  AOI211_X1 U16067 ( .C1(n14142), .C2(n14141), .A(n15083), .B(n14140), .ZN(
        n14143) );
  AOI211_X1 U16068 ( .C1(n15102), .C2(n14306), .A(n14144), .B(n14143), .ZN(
        n14310) );
  AOI211_X1 U16069 ( .C1(n14308), .C2(n14163), .A(n15125), .B(n14145), .ZN(
        n14307) );
  NAND2_X1 U16070 ( .A1(n14307), .A2(n15113), .ZN(n14149) );
  INV_X1 U16071 ( .A(n14146), .ZN(n14147) );
  AOI22_X1 U16072 ( .A1(n15105), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14147), 
        .B2(n15103), .ZN(n14148) );
  OAI211_X1 U16073 ( .C1(n6943), .C2(n15107), .A(n14149), .B(n14148), .ZN(
        n14150) );
  AOI21_X1 U16074 ( .B1(n15114), .B2(n14306), .A(n14150), .ZN(n14151) );
  OAI21_X1 U16075 ( .B1(n14310), .B2(n15105), .A(n14151), .ZN(P1_U3269) );
  XNOR2_X1 U16076 ( .A(n14152), .B(n14154), .ZN(n14316) );
  OAI21_X1 U16077 ( .B1(n14155), .B2(n14154), .A(n14153), .ZN(n14158) );
  AOI222_X1 U16078 ( .A1(n15098), .A2(n14158), .B1(n14157), .B2(n14812), .C1(
        n14156), .C2(n14979), .ZN(n14315) );
  NAND2_X1 U16079 ( .A1(n15105), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14159) );
  OAI21_X1 U16080 ( .B1(n14801), .B2(n14160), .A(n14159), .ZN(n14161) );
  AOI21_X1 U16081 ( .B1(n14313), .B2(n14255), .A(n14161), .ZN(n14167) );
  AOI21_X1 U16082 ( .B1(n14313), .B2(n6691), .A(n15125), .ZN(n14162) );
  AND2_X1 U16083 ( .A1(n14163), .A2(n14162), .ZN(n14312) );
  INV_X1 U16084 ( .A(n14164), .ZN(n14165) );
  NAND2_X1 U16085 ( .A1(n14312), .A2(n14165), .ZN(n14166) );
  OAI211_X1 U16086 ( .C1(n14315), .C2(n14251), .A(n14167), .B(n14166), .ZN(
        n14168) );
  INV_X1 U16087 ( .A(n14168), .ZN(n14169) );
  OAI21_X1 U16088 ( .B1(n14210), .B2(n14316), .A(n14169), .ZN(P1_U3270) );
  XNOR2_X1 U16089 ( .A(n14171), .B(n14170), .ZN(n14322) );
  XNOR2_X1 U16090 ( .A(n14173), .B(n14172), .ZN(n14320) );
  OAI211_X1 U16091 ( .C1(n6713), .C2(n7369), .A(n15111), .B(n6691), .ZN(n14318) );
  AOI22_X1 U16092 ( .A1(n14175), .A2(n14979), .B1(n14812), .B2(n14174), .ZN(
        n14317) );
  INV_X1 U16093 ( .A(n14176), .ZN(n14177) );
  OAI22_X1 U16094 ( .A1(n14317), .A2(n15105), .B1(n14177), .B2(n14801), .ZN(
        n14179) );
  NOR2_X1 U16095 ( .A1(n7369), .A2(n15107), .ZN(n14178) );
  AOI211_X1 U16096 ( .C1(n14251), .C2(P1_REG2_REG_22__SCAN_IN), .A(n14179), 
        .B(n14178), .ZN(n14180) );
  OAI21_X1 U16097 ( .B1(n14816), .B2(n14318), .A(n14180), .ZN(n14181) );
  AOI21_X1 U16098 ( .B1(n14320), .B2(n14182), .A(n14181), .ZN(n14183) );
  OAI21_X1 U16099 ( .B1(n14322), .B2(n14210), .A(n14183), .ZN(P1_U3271) );
  XNOR2_X1 U16100 ( .A(n14185), .B(n14184), .ZN(n14187) );
  AOI21_X1 U16101 ( .B1(n14187), .B2(n15098), .A(n14186), .ZN(n14326) );
  AOI211_X1 U16102 ( .C1(n14324), .C2(n6813), .A(n15125), .B(n6713), .ZN(
        n14323) );
  INV_X1 U16103 ( .A(n14188), .ZN(n14189) );
  AOI22_X1 U16104 ( .A1(n15105), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14189), 
        .B2(n15103), .ZN(n14190) );
  OAI21_X1 U16105 ( .B1(n6950), .B2(n15107), .A(n14190), .ZN(n14196) );
  INV_X1 U16106 ( .A(n14191), .ZN(n14192) );
  AOI21_X1 U16107 ( .B1(n14194), .B2(n14193), .A(n14192), .ZN(n14327) );
  NOR2_X1 U16108 ( .A1(n14327), .A2(n14210), .ZN(n14195) );
  AOI211_X1 U16109 ( .C1(n14323), .C2(n15113), .A(n14196), .B(n14195), .ZN(
        n14197) );
  OAI21_X1 U16110 ( .B1(n14251), .B2(n14326), .A(n14197), .ZN(P1_U3272) );
  AOI21_X1 U16111 ( .B1(n14198), .B2(n14209), .A(n15083), .ZN(n14203) );
  OAI22_X1 U16112 ( .A1(n14200), .A2(n14220), .B1(n14199), .B2(n14265), .ZN(
        n14201) );
  AOI21_X1 U16113 ( .B1(n14203), .B2(n14202), .A(n14201), .ZN(n14331) );
  AOI21_X1 U16114 ( .B1(n14329), .B2(n6807), .A(n15125), .ZN(n14204) );
  AND2_X1 U16115 ( .A1(n14204), .A2(n6813), .ZN(n14328) );
  AOI22_X1 U16116 ( .A1(n14328), .A2(n14206), .B1(n15103), .B2(n14205), .ZN(
        n14207) );
  AOI21_X1 U16117 ( .B1(n14331), .B2(n14207), .A(n15105), .ZN(n14215) );
  OAI21_X1 U16118 ( .B1(n6818), .B2(n14209), .A(n14208), .ZN(n14332) );
  NOR2_X1 U16119 ( .A1(n14332), .A2(n14210), .ZN(n14214) );
  INV_X1 U16120 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14211) );
  OAI22_X1 U16121 ( .A1(n14212), .A2(n15107), .B1(n14804), .B2(n14211), .ZN(
        n14213) );
  OR3_X1 U16122 ( .A1(n14215), .A2(n14214), .A3(n14213), .ZN(P1_U3273) );
  XOR2_X1 U16123 ( .A(n14216), .B(n14217), .Z(n14339) );
  XNOR2_X1 U16124 ( .A(n14218), .B(n14217), .ZN(n14337) );
  NAND2_X1 U16125 ( .A1(n14229), .A2(n14242), .ZN(n14219) );
  NAND3_X1 U16126 ( .A1(n6807), .A2(n15111), .A3(n14219), .ZN(n14334) );
  OR2_X1 U16127 ( .A1(n14221), .A2(n14220), .ZN(n14224) );
  NAND2_X1 U16128 ( .A1(n14222), .A2(n14979), .ZN(n14223) );
  AND2_X1 U16129 ( .A1(n14224), .A2(n14223), .ZN(n14333) );
  NAND2_X1 U16130 ( .A1(n14225), .A2(n15103), .ZN(n14227) );
  NAND2_X1 U16131 ( .A1(n15105), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n14226) );
  OAI211_X1 U16132 ( .C1(n14333), .C2(n15105), .A(n14227), .B(n14226), .ZN(
        n14228) );
  AOI21_X1 U16133 ( .B1(n14229), .B2(n14255), .A(n14228), .ZN(n14230) );
  OAI21_X1 U16134 ( .B1(n14334), .B2(n14816), .A(n14230), .ZN(n14231) );
  AOI21_X1 U16135 ( .B1(n14337), .B2(n14809), .A(n14231), .ZN(n14232) );
  OAI21_X1 U16136 ( .B1(n14339), .B2(n14233), .A(n14232), .ZN(P1_U3274) );
  XNOR2_X1 U16137 ( .A(n14234), .B(n14235), .ZN(n14340) );
  XNOR2_X1 U16138 ( .A(n14236), .B(n14235), .ZN(n14240) );
  AOI22_X1 U16139 ( .A1(n14238), .A2(n14812), .B1(n14979), .B2(n14237), .ZN(
        n14239) );
  OAI21_X1 U16140 ( .B1(n14240), .B2(n15083), .A(n14239), .ZN(n14241) );
  AOI21_X1 U16141 ( .B1(n15102), .B2(n14340), .A(n14241), .ZN(n14343) );
  INV_X1 U16142 ( .A(n14342), .ZN(n14248) );
  INV_X1 U16143 ( .A(n14242), .ZN(n14243) );
  AOI211_X1 U16144 ( .C1(n14342), .C2(n14244), .A(n15125), .B(n14243), .ZN(
        n14341) );
  NAND2_X1 U16145 ( .A1(n14341), .A2(n15113), .ZN(n14247) );
  AOI22_X1 U16146 ( .A1(n15118), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14245), 
        .B2(n15103), .ZN(n14246) );
  OAI211_X1 U16147 ( .C1(n14248), .C2(n15107), .A(n14247), .B(n14246), .ZN(
        n14249) );
  AOI21_X1 U16148 ( .B1(n15114), .B2(n14340), .A(n14249), .ZN(n14250) );
  OAI21_X1 U16149 ( .B1(n14251), .B2(n14343), .A(n14250), .ZN(P1_U3275) );
  OAI21_X1 U16150 ( .B1(n14264), .B2(n14253), .A(n14252), .ZN(n15130) );
  AOI22_X1 U16151 ( .A1(n15114), .A2(n15130), .B1(n14255), .B2(n14254), .ZN(
        n14272) );
  NOR2_X1 U16152 ( .A1(n15124), .A2(n14256), .ZN(n14257) );
  OR2_X1 U16153 ( .A1(n14258), .A2(n14257), .ZN(n15126) );
  INV_X1 U16154 ( .A(n15126), .ZN(n14259) );
  AOI22_X1 U16155 ( .A1(n14260), .A2(n14259), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n15103), .ZN(n14271) );
  XNOR2_X1 U16156 ( .A(n15126), .B(n14261), .ZN(n14263) );
  OAI21_X1 U16157 ( .B1(n14263), .B2(n15083), .A(n10210), .ZN(n14269) );
  OAI21_X1 U16158 ( .B1(n14264), .B2(n10210), .A(n15098), .ZN(n14266) );
  NAND2_X1 U16159 ( .A1(n14266), .A2(n14265), .ZN(n14268) );
  AOI222_X1 U16160 ( .A1(n14269), .A2(n14268), .B1(n14267), .B2(n14812), .C1(
        n15130), .C2(n15102), .ZN(n15127) );
  MUX2_X1 U16161 ( .A(n15127), .B(n10586), .S(n15118), .Z(n14270) );
  NAND3_X1 U16162 ( .A1(n14272), .A2(n14271), .A3(n14270), .ZN(P1_U3292) );
  OAI211_X1 U16163 ( .C1(n6685), .C2(n15185), .A(n14273), .B(n14275), .ZN(
        n14361) );
  MUX2_X1 U16164 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14361), .S(n15215), .Z(
        P1_U3559) );
  OAI211_X1 U16165 ( .C1(n14277), .C2(n15185), .A(n14276), .B(n14275), .ZN(
        n14362) );
  MUX2_X1 U16166 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14362), .S(n15215), .Z(
        P1_U3558) );
  NAND2_X1 U16167 ( .A1(n14279), .A2(n14980), .ZN(n14280) );
  MUX2_X1 U16168 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14363), .S(n15215), .Z(
        P1_U3556) );
  INV_X1 U16169 ( .A(n14345), .ZN(n15190) );
  NAND2_X1 U16170 ( .A1(n14285), .A2(n14980), .ZN(n14286) );
  NAND2_X1 U16171 ( .A1(n14287), .A2(n14286), .ZN(n14288) );
  AOI21_X1 U16172 ( .B1(n14289), .B2(n15190), .A(n14288), .ZN(n14290) );
  NAND2_X1 U16173 ( .A1(n14291), .A2(n14290), .ZN(n14364) );
  MUX2_X1 U16174 ( .A(n14364), .B(P1_REG1_REG_27__SCAN_IN), .S(n15213), .Z(
        P1_U3555) );
  OAI21_X1 U16175 ( .B1(n14293), .B2(n15185), .A(n14292), .ZN(n14295) );
  AOI211_X1 U16176 ( .C1(n15098), .C2(n14296), .A(n14295), .B(n14294), .ZN(
        n14297) );
  OAI21_X1 U16177 ( .B1(n14359), .B2(n14298), .A(n14297), .ZN(n14365) );
  MUX2_X1 U16178 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14365), .S(n15215), .Z(
        P1_U3554) );
  OAI211_X1 U16179 ( .C1(n14301), .C2(n15185), .A(n14300), .B(n14299), .ZN(
        n14302) );
  AOI21_X1 U16180 ( .B1(n14303), .B2(n15198), .A(n14302), .ZN(n14304) );
  OAI21_X1 U16181 ( .B1(n15083), .B2(n14305), .A(n14304), .ZN(n14366) );
  MUX2_X1 U16182 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14366), .S(n15215), .Z(
        P1_U3553) );
  INV_X1 U16183 ( .A(n14306), .ZN(n14311) );
  AOI21_X1 U16184 ( .B1(n14980), .B2(n14308), .A(n14307), .ZN(n14309) );
  OAI211_X1 U16185 ( .C1(n14311), .C2(n14345), .A(n14310), .B(n14309), .ZN(
        n14367) );
  MUX2_X1 U16186 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14367), .S(n15215), .Z(
        P1_U3552) );
  AOI21_X1 U16187 ( .B1(n14980), .B2(n14313), .A(n14312), .ZN(n14314) );
  OAI211_X1 U16188 ( .C1(n14359), .C2(n14316), .A(n14315), .B(n14314), .ZN(
        n14368) );
  MUX2_X1 U16189 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14368), .S(n15215), .Z(
        P1_U3551) );
  OAI211_X1 U16190 ( .C1(n15185), .C2(n7369), .A(n14318), .B(n14317), .ZN(
        n14319) );
  AOI21_X1 U16191 ( .B1(n14320), .B2(n15098), .A(n14319), .ZN(n14321) );
  OAI21_X1 U16192 ( .B1(n14322), .B2(n14359), .A(n14321), .ZN(n14369) );
  MUX2_X1 U16193 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14369), .S(n15215), .Z(
        P1_U3550) );
  AOI21_X1 U16194 ( .B1(n14980), .B2(n14324), .A(n14323), .ZN(n14325) );
  OAI211_X1 U16195 ( .C1(n14327), .C2(n14359), .A(n14326), .B(n14325), .ZN(
        n14370) );
  MUX2_X1 U16196 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14370), .S(n15215), .Z(
        P1_U3549) );
  AOI21_X1 U16197 ( .B1(n14980), .B2(n14329), .A(n14328), .ZN(n14330) );
  OAI211_X1 U16198 ( .C1(n14332), .C2(n14359), .A(n14331), .B(n14330), .ZN(
        n14371) );
  MUX2_X1 U16199 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14371), .S(n15215), .Z(
        P1_U3548) );
  OAI211_X1 U16200 ( .C1(n14335), .C2(n15185), .A(n14334), .B(n14333), .ZN(
        n14336) );
  AOI21_X1 U16201 ( .B1(n14337), .B2(n15198), .A(n14336), .ZN(n14338) );
  OAI21_X1 U16202 ( .B1(n14339), .B2(n15083), .A(n14338), .ZN(n14372) );
  MUX2_X1 U16203 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14372), .S(n15215), .Z(
        P1_U3547) );
  INV_X1 U16204 ( .A(n14340), .ZN(n14346) );
  AOI21_X1 U16205 ( .B1(n14980), .B2(n14342), .A(n14341), .ZN(n14344) );
  OAI211_X1 U16206 ( .C1(n14346), .C2(n14345), .A(n14344), .B(n14343), .ZN(
        n14373) );
  MUX2_X1 U16207 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14373), .S(n15215), .Z(
        P1_U3546) );
  OAI211_X1 U16208 ( .C1(n14349), .C2(n15185), .A(n14348), .B(n14347), .ZN(
        n14350) );
  AOI21_X1 U16209 ( .B1(n14351), .B2(n15098), .A(n14350), .ZN(n14352) );
  OAI21_X1 U16210 ( .B1(n14353), .B2(n14359), .A(n14352), .ZN(n14374) );
  MUX2_X1 U16211 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14374), .S(n15215), .Z(
        P1_U3545) );
  AOI22_X1 U16212 ( .A1(n14355), .A2(n15111), .B1(n14980), .B2(n14354), .ZN(
        n14356) );
  OAI211_X1 U16213 ( .C1(n14359), .C2(n14358), .A(n14357), .B(n14356), .ZN(
        n14375) );
  MUX2_X1 U16214 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14375), .S(n15215), .Z(
        P1_U3543) );
  MUX2_X1 U16215 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14360), .S(n15215), .Z(
        P1_U3528) );
  MUX2_X1 U16216 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14361), .S(n15201), .Z(
        P1_U3527) );
  MUX2_X1 U16217 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14362), .S(n15201), .Z(
        P1_U3526) );
  MUX2_X1 U16218 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14363), .S(n15201), .Z(
        P1_U3524) );
  MUX2_X1 U16219 ( .A(n14364), .B(P1_REG0_REG_27__SCAN_IN), .S(n15199), .Z(
        P1_U3523) );
  MUX2_X1 U16220 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14365), .S(n15201), .Z(
        P1_U3522) );
  MUX2_X1 U16221 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14366), .S(n15201), .Z(
        P1_U3521) );
  MUX2_X1 U16222 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14367), .S(n15201), .Z(
        P1_U3520) );
  MUX2_X1 U16223 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14368), .S(n15201), .Z(
        P1_U3519) );
  MUX2_X1 U16224 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14369), .S(n15201), .Z(
        P1_U3518) );
  MUX2_X1 U16225 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14370), .S(n15201), .Z(
        P1_U3517) );
  MUX2_X1 U16226 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14371), .S(n15201), .Z(
        P1_U3516) );
  MUX2_X1 U16227 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14372), .S(n15201), .Z(
        P1_U3515) );
  MUX2_X1 U16228 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14373), .S(n15201), .Z(
        P1_U3513) );
  MUX2_X1 U16229 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14374), .S(n15201), .Z(
        P1_U3510) );
  MUX2_X1 U16230 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14375), .S(n15201), .Z(
        P1_U3504) );
  INV_X1 U16231 ( .A(n14376), .ZN(n14380) );
  NOR4_X1 U16232 ( .A1(n14377), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n8787), .ZN(n14378) );
  AOI21_X1 U16233 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14756), .A(n14378), 
        .ZN(n14379) );
  OAI21_X1 U16234 ( .B1(n14380), .B2(n14383), .A(n14379), .ZN(P1_U3324) );
  INV_X1 U16235 ( .A(n14387), .ZN(n14388) );
  OAI222_X1 U16236 ( .A1(n6661), .A2(P1_U3086), .B1(n14398), .B2(n14388), .C1(
        n7129), .C2(n14395), .ZN(P1_U3327) );
  OAI222_X1 U16237 ( .A1(n15026), .A2(P1_U3086), .B1(n14398), .B2(n14391), 
        .C1(n14390), .C2(n14395), .ZN(P1_U3328) );
  OAI222_X1 U16238 ( .A1(n14394), .A2(P1_U3086), .B1(n14398), .B2(n14393), 
        .C1(n14392), .C2(n14395), .ZN(P1_U3329) );
  OAI222_X1 U16239 ( .A1(P1_U3086), .A2(n8976), .B1(n14398), .B2(n14397), .C1(
        n14396), .C2(n14395), .ZN(P1_U3330) );
  MUX2_X1 U16240 ( .A(n14400), .B(n14399), .S(P1_U3086), .Z(P1_U3333) );
  OAI22_X1 U16241 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(keyinput150), .B1(
        P1_REG3_REG_27__SCAN_IN), .B2(keyinput223), .ZN(n14401) );
  AOI221_X1 U16242 ( .B1(P2_IR_REG_21__SCAN_IN), .B2(keyinput150), .C1(
        keyinput223), .C2(P1_REG3_REG_27__SCAN_IN), .A(n14401), .ZN(n14408) );
  OAI22_X1 U16243 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(keyinput251), .B1(
        keyinput243), .B2(P1_D_REG_17__SCAN_IN), .ZN(n14402) );
  AOI221_X1 U16244 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(keyinput251), .C1(
        P1_D_REG_17__SCAN_IN), .C2(keyinput243), .A(n14402), .ZN(n14407) );
  OAI22_X1 U16245 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(keyinput170), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput132), .ZN(n14403) );
  AOI221_X1 U16246 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(keyinput170), .C1(
        keyinput132), .C2(P1_IR_REG_18__SCAN_IN), .A(n14403), .ZN(n14406) );
  OAI22_X1 U16247 ( .A1(P3_REG2_REG_5__SCAN_IN), .A2(keyinput157), .B1(
        P2_REG0_REG_12__SCAN_IN), .B2(keyinput158), .ZN(n14404) );
  AOI221_X1 U16248 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(keyinput157), .C1(
        keyinput158), .C2(P2_REG0_REG_12__SCAN_IN), .A(n14404), .ZN(n14405) );
  NAND4_X1 U16249 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        n14436) );
  OAI22_X1 U16250 ( .A1(P3_REG1_REG_1__SCAN_IN), .A2(keyinput244), .B1(
        P2_IR_REG_16__SCAN_IN), .B2(keyinput129), .ZN(n14409) );
  AOI221_X1 U16251 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(keyinput244), .C1(
        keyinput129), .C2(P2_IR_REG_16__SCAN_IN), .A(n14409), .ZN(n14416) );
  OAI22_X1 U16252 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(keyinput198), .B1(
        keyinput253), .B2(P2_REG2_REG_22__SCAN_IN), .ZN(n14410) );
  AOI221_X1 U16253 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(keyinput198), .C1(
        P2_REG2_REG_22__SCAN_IN), .C2(keyinput253), .A(n14410), .ZN(n14415) );
  OAI22_X1 U16254 ( .A1(P3_B_REG_SCAN_IN), .A2(keyinput186), .B1(keyinput187), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n14411) );
  AOI221_X1 U16255 ( .B1(P3_B_REG_SCAN_IN), .B2(keyinput186), .C1(
        P3_DATAO_REG_0__SCAN_IN), .C2(keyinput187), .A(n14411), .ZN(n14414) );
  OAI22_X1 U16256 ( .A1(P3_D_REG_14__SCAN_IN), .A2(keyinput255), .B1(
        P3_DATAO_REG_5__SCAN_IN), .B2(keyinput221), .ZN(n14412) );
  AOI221_X1 U16257 ( .B1(P3_D_REG_14__SCAN_IN), .B2(keyinput255), .C1(
        keyinput221), .C2(P3_DATAO_REG_5__SCAN_IN), .A(n14412), .ZN(n14413) );
  NAND4_X1 U16258 ( .A1(n14416), .A2(n14415), .A3(n14414), .A4(n14413), .ZN(
        n14435) );
  OAI22_X1 U16259 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(keyinput240), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput211), .ZN(n14417) );
  AOI221_X1 U16260 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(keyinput240), .C1(
        keyinput211), .C2(P2_REG3_REG_6__SCAN_IN), .A(n14417), .ZN(n14424) );
  OAI22_X1 U16261 ( .A1(P3_REG0_REG_17__SCAN_IN), .A2(keyinput181), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(keyinput200), .ZN(n14418) );
  AOI221_X1 U16262 ( .B1(P3_REG0_REG_17__SCAN_IN), .B2(keyinput181), .C1(
        keyinput200), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n14418), .ZN(n14423) );
  OAI22_X1 U16263 ( .A1(P2_D_REG_16__SCAN_IN), .A2(keyinput202), .B1(
        keyinput228), .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n14419) );
  AOI221_X1 U16264 ( .B1(P2_D_REG_16__SCAN_IN), .B2(keyinput202), .C1(
        P3_DATAO_REG_30__SCAN_IN), .C2(keyinput228), .A(n14419), .ZN(n14422)
         );
  OAI22_X1 U16265 ( .A1(P3_D_REG_19__SCAN_IN), .A2(keyinput188), .B1(
        P3_ADDR_REG_18__SCAN_IN), .B2(keyinput216), .ZN(n14420) );
  AOI221_X1 U16266 ( .B1(P3_D_REG_19__SCAN_IN), .B2(keyinput188), .C1(
        keyinput216), .C2(P3_ADDR_REG_18__SCAN_IN), .A(n14420), .ZN(n14421) );
  NAND4_X1 U16267 ( .A1(n14424), .A2(n14423), .A3(n14422), .A4(n14421), .ZN(
        n14434) );
  OAI22_X1 U16268 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput167), .B1(
        keyinput165), .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n14425) );
  AOI221_X1 U16269 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput167), .C1(
        P3_DATAO_REG_16__SCAN_IN), .C2(keyinput165), .A(n14425), .ZN(n14432)
         );
  OAI22_X1 U16270 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput183), .B1(
        P2_REG0_REG_27__SCAN_IN), .B2(keyinput217), .ZN(n14426) );
  AOI221_X1 U16271 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput183), .C1(
        keyinput217), .C2(P2_REG0_REG_27__SCAN_IN), .A(n14426), .ZN(n14431) );
  OAI22_X1 U16272 ( .A1(SI_14_), .A2(keyinput215), .B1(P1_REG3_REG_23__SCAN_IN), .B2(keyinput138), .ZN(n14427) );
  AOI221_X1 U16273 ( .B1(SI_14_), .B2(keyinput215), .C1(keyinput138), .C2(
        P1_REG3_REG_23__SCAN_IN), .A(n14427), .ZN(n14430) );
  OAI22_X1 U16274 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(keyinput252), .B1(
        keyinput220), .B2(P3_ADDR_REG_10__SCAN_IN), .ZN(n14428) );
  AOI221_X1 U16275 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(keyinput252), .C1(
        P3_ADDR_REG_10__SCAN_IN), .C2(keyinput220), .A(n14428), .ZN(n14429) );
  NAND4_X1 U16276 ( .A1(n14432), .A2(n14431), .A3(n14430), .A4(n14429), .ZN(
        n14433) );
  NOR4_X1 U16277 ( .A1(n14436), .A2(n14435), .A3(n14434), .A4(n14433), .ZN(
        n14515) );
  OAI22_X1 U16278 ( .A1(P2_D_REG_20__SCAN_IN), .A2(keyinput173), .B1(
        keyinput192), .B2(P1_REG0_REG_19__SCAN_IN), .ZN(n14437) );
  AOI221_X1 U16279 ( .B1(P2_D_REG_20__SCAN_IN), .B2(keyinput173), .C1(
        P1_REG0_REG_19__SCAN_IN), .C2(keyinput192), .A(n14437), .ZN(n14444) );
  OAI22_X1 U16280 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(keyinput159), .B1(
        P2_ADDR_REG_10__SCAN_IN), .B2(keyinput133), .ZN(n14438) );
  AOI221_X1 U16281 ( .B1(P2_REG1_REG_27__SCAN_IN), .B2(keyinput159), .C1(
        keyinput133), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n14438), .ZN(n14443) );
  OAI22_X1 U16282 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput134), .B1(
        P2_REG2_REG_23__SCAN_IN), .B2(keyinput254), .ZN(n14439) );
  AOI221_X1 U16283 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput134), .C1(
        keyinput254), .C2(P2_REG2_REG_23__SCAN_IN), .A(n14439), .ZN(n14442) );
  OAI22_X1 U16284 ( .A1(P3_D_REG_0__SCAN_IN), .A2(keyinput197), .B1(
        P1_REG3_REG_14__SCAN_IN), .B2(keyinput176), .ZN(n14440) );
  AOI221_X1 U16285 ( .B1(P3_D_REG_0__SCAN_IN), .B2(keyinput197), .C1(
        keyinput176), .C2(P1_REG3_REG_14__SCAN_IN), .A(n14440), .ZN(n14441) );
  NAND4_X1 U16286 ( .A1(n14444), .A2(n14443), .A3(n14442), .A4(n14441), .ZN(
        n14472) );
  OAI22_X1 U16287 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(keyinput201), .B1(SI_17_), 
        .B2(keyinput235), .ZN(n14445) );
  AOI221_X1 U16288 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(keyinput201), .C1(
        keyinput235), .C2(SI_17_), .A(n14445), .ZN(n14452) );
  OAI22_X1 U16289 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput242), .B1(
        keyinput199), .B2(P3_ADDR_REG_13__SCAN_IN), .ZN(n14446) );
  AOI221_X1 U16290 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput242), .C1(
        P3_ADDR_REG_13__SCAN_IN), .C2(keyinput199), .A(n14446), .ZN(n14451) );
  OAI22_X1 U16291 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(keyinput152), .B1(
        P2_REG2_REG_31__SCAN_IN), .B2(keyinput208), .ZN(n14447) );
  AOI221_X1 U16292 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(keyinput152), .C1(
        keyinput208), .C2(P2_REG2_REG_31__SCAN_IN), .A(n14447), .ZN(n14450) );
  OAI22_X1 U16293 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput190), .B1(
        P2_REG1_REG_13__SCAN_IN), .B2(keyinput227), .ZN(n14448) );
  AOI221_X1 U16294 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput190), .C1(
        keyinput227), .C2(P2_REG1_REG_13__SCAN_IN), .A(n14448), .ZN(n14449) );
  NAND4_X1 U16295 ( .A1(n14452), .A2(n14451), .A3(n14450), .A4(n14449), .ZN(
        n14471) );
  OAI22_X1 U16296 ( .A1(SI_18_), .A2(keyinput214), .B1(keyinput177), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14453) );
  AOI221_X1 U16297 ( .B1(SI_18_), .B2(keyinput214), .C1(
        P3_ADDR_REG_17__SCAN_IN), .C2(keyinput177), .A(n14453), .ZN(n14460) );
  OAI22_X1 U16298 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput213), .B1(
        keyinput191), .B2(P1_REG3_REG_6__SCAN_IN), .ZN(n14454) );
  AOI221_X1 U16299 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput213), .C1(
        P1_REG3_REG_6__SCAN_IN), .C2(keyinput191), .A(n14454), .ZN(n14459) );
  OAI22_X1 U16300 ( .A1(P3_D_REG_17__SCAN_IN), .A2(keyinput141), .B1(
        keyinput225), .B2(P3_REG1_REG_23__SCAN_IN), .ZN(n14455) );
  AOI221_X1 U16301 ( .B1(P3_D_REG_17__SCAN_IN), .B2(keyinput141), .C1(
        P3_REG1_REG_23__SCAN_IN), .C2(keyinput225), .A(n14455), .ZN(n14458) );
  OAI22_X1 U16302 ( .A1(SI_27_), .A2(keyinput239), .B1(SI_25_), .B2(
        keyinput247), .ZN(n14456) );
  AOI221_X1 U16303 ( .B1(SI_27_), .B2(keyinput239), .C1(keyinput247), .C2(
        SI_25_), .A(n14456), .ZN(n14457) );
  NAND4_X1 U16304 ( .A1(n14460), .A2(n14459), .A3(n14458), .A4(n14457), .ZN(
        n14470) );
  OAI22_X1 U16305 ( .A1(P3_REG0_REG_24__SCAN_IN), .A2(keyinput203), .B1(
        keyinput146), .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n14461) );
  AOI221_X1 U16306 ( .B1(P3_REG0_REG_24__SCAN_IN), .B2(keyinput203), .C1(
        P2_REG0_REG_18__SCAN_IN), .C2(keyinput146), .A(n14461), .ZN(n14468) );
  OAI22_X1 U16307 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(keyinput156), .B1(
        keyinput135), .B2(P1_ADDR_REG_9__SCAN_IN), .ZN(n14462) );
  AOI221_X1 U16308 ( .B1(P1_DATAO_REG_16__SCAN_IN), .B2(keyinput156), .C1(
        P1_ADDR_REG_9__SCAN_IN), .C2(keyinput135), .A(n14462), .ZN(n14467) );
  OAI22_X1 U16309 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput248), .B1(
        P2_ADDR_REG_3__SCAN_IN), .B2(keyinput182), .ZN(n14463) );
  AOI221_X1 U16310 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput248), .C1(
        keyinput182), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n14463), .ZN(n14466) );
  OAI22_X1 U16311 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput219), .B1(
        keyinput153), .B2(P1_REG0_REG_12__SCAN_IN), .ZN(n14464) );
  AOI221_X1 U16312 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput219), .C1(
        P1_REG0_REG_12__SCAN_IN), .C2(keyinput153), .A(n14464), .ZN(n14465) );
  NAND4_X1 U16313 ( .A1(n14468), .A2(n14467), .A3(n14466), .A4(n14465), .ZN(
        n14469) );
  NOR4_X1 U16314 ( .A1(n14472), .A2(n14471), .A3(n14470), .A4(n14469), .ZN(
        n14514) );
  INV_X1 U16315 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U16316 ( .A1(n11310), .A2(keyinput162), .B1(keyinput236), .B2(
        n15120), .ZN(n14473) );
  OAI221_X1 U16317 ( .B1(n11310), .B2(keyinput162), .C1(n15120), .C2(
        keyinput236), .A(n14473), .ZN(n14481) );
  INV_X1 U16318 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15145) );
  AOI22_X1 U16319 ( .A1(n15145), .A2(keyinput234), .B1(n15257), .B2(
        keyinput205), .ZN(n14474) );
  OAI221_X1 U16320 ( .B1(n15145), .B2(keyinput234), .C1(n15257), .C2(
        keyinput205), .A(n14474), .ZN(n14480) );
  INV_X1 U16321 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15119) );
  XNOR2_X1 U16322 ( .A(n15119), .B(keyinput207), .ZN(n14479) );
  XNOR2_X1 U16323 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput195), .ZN(n14477) );
  XNOR2_X1 U16324 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput180), .ZN(n14476) );
  XNOR2_X1 U16325 ( .A(P3_IR_REG_22__SCAN_IN), .B(keyinput142), .ZN(n14475) );
  NAND3_X1 U16326 ( .A1(n14477), .A2(n14476), .A3(n14475), .ZN(n14478) );
  NOR4_X1 U16327 ( .A1(n14481), .A2(n14480), .A3(n14479), .A4(n14478), .ZN(
        n14513) );
  OAI22_X1 U16328 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput229), .B1(
        P2_REG0_REG_8__SCAN_IN), .B2(keyinput148), .ZN(n14482) );
  AOI221_X1 U16329 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput229), .C1(
        keyinput148), .C2(P2_REG0_REG_8__SCAN_IN), .A(n14482), .ZN(n14489) );
  OAI22_X1 U16330 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput143), .B1(
        keyinput163), .B2(P1_REG1_REG_20__SCAN_IN), .ZN(n14483) );
  AOI221_X1 U16331 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput143), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput163), .A(n14483), .ZN(n14488) );
  OAI22_X1 U16332 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(keyinput168), .B1(
        keyinput139), .B2(P2_D_REG_30__SCAN_IN), .ZN(n14484) );
  AOI221_X1 U16333 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput168), .C1(
        P2_D_REG_30__SCAN_IN), .C2(keyinput139), .A(n14484), .ZN(n14487) );
  OAI22_X1 U16334 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(keyinput194), .B1(
        keyinput184), .B2(P1_REG0_REG_24__SCAN_IN), .ZN(n14485) );
  AOI221_X1 U16335 ( .B1(P1_REG0_REG_29__SCAN_IN), .B2(keyinput194), .C1(
        P1_REG0_REG_24__SCAN_IN), .C2(keyinput184), .A(n14485), .ZN(n14486) );
  NAND4_X1 U16336 ( .A1(n14489), .A2(n14488), .A3(n14487), .A4(n14486), .ZN(
        n14511) );
  OAI22_X1 U16337 ( .A1(n12966), .A2(keyinput238), .B1(n10379), .B2(
        keyinput149), .ZN(n14490) );
  AOI221_X1 U16338 ( .B1(n12966), .B2(keyinput238), .C1(keyinput149), .C2(
        n10379), .A(n14490), .ZN(n14498) );
  OAI22_X1 U16339 ( .A1(n14661), .A2(keyinput175), .B1(n15204), .B2(
        keyinput166), .ZN(n14491) );
  AOI221_X1 U16340 ( .B1(n14661), .B2(keyinput175), .C1(keyinput166), .C2(
        n15204), .A(n14491), .ZN(n14497) );
  OAI22_X1 U16341 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput155), .B1(
        keyinput209), .B2(P2_REG1_REG_7__SCAN_IN), .ZN(n14492) );
  AOI221_X1 U16342 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput155), .C1(
        P2_REG1_REG_7__SCAN_IN), .C2(keyinput209), .A(n14492), .ZN(n14496) );
  XOR2_X1 U16343 ( .A(SI_9_), .B(keyinput147), .Z(n14494) );
  XNOR2_X1 U16344 ( .A(keyinput250), .B(n8309), .ZN(n14493) );
  NOR2_X1 U16345 ( .A1(n14494), .A2(n14493), .ZN(n14495) );
  NAND4_X1 U16346 ( .A1(n14498), .A2(n14497), .A3(n14496), .A4(n14495), .ZN(
        n14510) );
  OAI22_X1 U16347 ( .A1(n14500), .A2(keyinput172), .B1(n15306), .B2(
        keyinput193), .ZN(n14499) );
  AOI221_X1 U16348 ( .B1(n14500), .B2(keyinput172), .C1(keyinput193), .C2(
        n15306), .A(n14499), .ZN(n14508) );
  OAI22_X1 U16349 ( .A1(n14588), .A2(keyinput128), .B1(n14599), .B2(
        keyinput164), .ZN(n14501) );
  AOI221_X1 U16350 ( .B1(n14588), .B2(keyinput128), .C1(keyinput164), .C2(
        n14599), .A(n14501), .ZN(n14507) );
  XNOR2_X1 U16351 ( .A(SI_4_), .B(keyinput137), .ZN(n14505) );
  XNOR2_X1 U16352 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput249), .ZN(n14504)
         );
  INV_X1 U16353 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n14583) );
  XNOR2_X1 U16354 ( .A(keyinput178), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14503) );
  XNOR2_X1 U16355 ( .A(keyinput174), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n14502)
         );
  AND4_X1 U16356 ( .A1(n14505), .A2(n14504), .A3(n14503), .A4(n14502), .ZN(
        n14506) );
  NAND3_X1 U16357 ( .A1(n14508), .A2(n14507), .A3(n14506), .ZN(n14509) );
  NOR3_X1 U16358 ( .A1(n14511), .A2(n14510), .A3(n14509), .ZN(n14512) );
  NAND4_X1 U16359 ( .A1(n14515), .A2(n14514), .A3(n14513), .A4(n14512), .ZN(
        n14755) );
  AOI22_X1 U16360 ( .A1(n14517), .A2(keyinput233), .B1(n9628), .B2(keyinput169), .ZN(n14516) );
  OAI221_X1 U16361 ( .B1(n14517), .B2(keyinput233), .C1(n9628), .C2(
        keyinput169), .A(n14516), .ZN(n14527) );
  INV_X1 U16362 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n14519) );
  AOI22_X1 U16363 ( .A1(n14102), .A2(keyinput171), .B1(n14519), .B2(
        keyinput206), .ZN(n14518) );
  OAI221_X1 U16364 ( .B1(n14102), .B2(keyinput171), .C1(n14519), .C2(
        keyinput206), .A(n14518), .ZN(n14526) );
  AOI22_X1 U16365 ( .A1(n14521), .A2(keyinput231), .B1(keyinput154), .B2(
        n14663), .ZN(n14520) );
  OAI221_X1 U16366 ( .B1(n14521), .B2(keyinput231), .C1(n14663), .C2(
        keyinput154), .A(n14520), .ZN(n14525) );
  XOR2_X1 U16367 ( .A(n8906), .B(keyinput136), .Z(n14523) );
  XNOR2_X1 U16368 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput210), .ZN(n14522) );
  NAND2_X1 U16369 ( .A1(n14523), .A2(n14522), .ZN(n14524) );
  NOR4_X1 U16370 ( .A1(n14527), .A2(n14526), .A3(n14525), .A4(n14524), .ZN(
        n14564) );
  AOI22_X1 U16371 ( .A1(n9897), .A2(keyinput224), .B1(n14580), .B2(keyinput218), .ZN(n14528) );
  OAI221_X1 U16372 ( .B1(n9897), .B2(keyinput224), .C1(n14580), .C2(
        keyinput218), .A(n14528), .ZN(n14539) );
  AOI22_X1 U16373 ( .A1(n14530), .A2(keyinput204), .B1(n12285), .B2(
        keyinput212), .ZN(n14529) );
  OAI221_X1 U16374 ( .B1(n14530), .B2(keyinput204), .C1(n12285), .C2(
        keyinput212), .A(n14529), .ZN(n14538) );
  INV_X1 U16375 ( .A(n6829), .ZN(n14533) );
  INV_X1 U16376 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n14532) );
  AOI22_X1 U16377 ( .A1(n14533), .A2(keyinput241), .B1(keyinput226), .B2(
        n14532), .ZN(n14531) );
  OAI221_X1 U16378 ( .B1(n14533), .B2(keyinput241), .C1(n14532), .C2(
        keyinput226), .A(n14531), .ZN(n14537) );
  XNOR2_X1 U16379 ( .A(P3_IR_REG_20__SCAN_IN), .B(keyinput179), .ZN(n14535) );
  XNOR2_X1 U16380 ( .A(SI_6_), .B(keyinput131), .ZN(n14534) );
  NAND2_X1 U16381 ( .A1(n14535), .A2(n14534), .ZN(n14536) );
  NOR4_X1 U16382 ( .A1(n14539), .A2(n14538), .A3(n14537), .A4(n14536), .ZN(
        n14563) );
  AOI22_X1 U16383 ( .A1(n14694), .A2(keyinput222), .B1(keyinput144), .B2(
        n14541), .ZN(n14540) );
  OAI221_X1 U16384 ( .B1(n14694), .B2(keyinput222), .C1(n14541), .C2(
        keyinput144), .A(n14540), .ZN(n14550) );
  AOI22_X1 U16385 ( .A1(n14572), .A2(keyinput161), .B1(n10875), .B2(
        keyinput185), .ZN(n14542) );
  OAI221_X1 U16386 ( .B1(n14572), .B2(keyinput161), .C1(n10875), .C2(
        keyinput185), .A(n14542), .ZN(n14549) );
  INV_X1 U16387 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14544) );
  AOI22_X1 U16388 ( .A1(n14544), .A2(keyinput145), .B1(keyinput230), .B2(
        n14623), .ZN(n14543) );
  OAI221_X1 U16389 ( .B1(n14544), .B2(keyinput145), .C1(n14623), .C2(
        keyinput230), .A(n14543), .ZN(n14548) );
  AOI22_X1 U16390 ( .A1(n14597), .A2(keyinput237), .B1(keyinput160), .B2(
        n14546), .ZN(n14545) );
  OAI221_X1 U16391 ( .B1(n14597), .B2(keyinput237), .C1(n14546), .C2(
        keyinput160), .A(n14545), .ZN(n14547) );
  NOR4_X1 U16392 ( .A1(n14550), .A2(n14549), .A3(n14548), .A4(n14547), .ZN(
        n14562) );
  AOI22_X1 U16393 ( .A1(n14552), .A2(keyinput151), .B1(n14608), .B2(
        keyinput232), .ZN(n14551) );
  OAI221_X1 U16394 ( .B1(n14552), .B2(keyinput151), .C1(n14608), .C2(
        keyinput232), .A(n14551), .ZN(n14560) );
  AOI22_X1 U16395 ( .A1(n10867), .A2(keyinput245), .B1(n14657), .B2(
        keyinput189), .ZN(n14553) );
  OAI221_X1 U16396 ( .B1(n10867), .B2(keyinput245), .C1(n14657), .C2(
        keyinput189), .A(n14553), .ZN(n14559) );
  XNOR2_X1 U16397 ( .A(SI_1_), .B(keyinput196), .ZN(n14557) );
  XNOR2_X1 U16398 ( .A(P2_REG0_REG_14__SCAN_IN), .B(keyinput140), .ZN(n14556)
         );
  XNOR2_X1 U16399 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput246), .ZN(n14555) );
  XNOR2_X1 U16400 ( .A(P1_REG3_REG_28__SCAN_IN), .B(keyinput130), .ZN(n14554)
         );
  NAND4_X1 U16401 ( .A1(n14557), .A2(n14556), .A3(n14555), .A4(n14554), .ZN(
        n14558) );
  NOR3_X1 U16402 ( .A1(n14560), .A2(n14559), .A3(n14558), .ZN(n14561) );
  NAND4_X1 U16403 ( .A1(n14564), .A2(n14563), .A3(n14562), .A4(n14561), .ZN(
        n14754) );
  AOI22_X1 U16404 ( .A1(n14567), .A2(keyinput53), .B1(keyinput72), .B2(n14566), 
        .ZN(n14565) );
  OAI221_X1 U16405 ( .B1(n14567), .B2(keyinput53), .C1(n14566), .C2(keyinput72), .A(n14565), .ZN(n14578) );
  AOI22_X1 U16406 ( .A1(n10676), .A2(keyinput114), .B1(keyinput37), .B2(n14569), .ZN(n14568) );
  OAI221_X1 U16407 ( .B1(n10676), .B2(keyinput114), .C1(n14569), .C2(
        keyinput37), .A(n14568), .ZN(n14577) );
  AOI22_X1 U16408 ( .A1(n14572), .A2(keyinput33), .B1(n14571), .B2(keyinput40), 
        .ZN(n14570) );
  OAI221_X1 U16409 ( .B1(n14572), .B2(keyinput33), .C1(n14571), .C2(keyinput40), .A(n14570), .ZN(n14576) );
  INV_X1 U16410 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14798) );
  AOI22_X1 U16411 ( .A1(n14574), .A2(keyinput15), .B1(keyinput25), .B2(n14798), 
        .ZN(n14573) );
  OAI221_X1 U16412 ( .B1(n14574), .B2(keyinput15), .C1(n14798), .C2(keyinput25), .A(n14573), .ZN(n14575) );
  NOR4_X1 U16413 ( .A1(n14578), .A2(n14577), .A3(n14576), .A4(n14575), .ZN(
        n14621) );
  AOI22_X1 U16414 ( .A1(n14581), .A2(keyinput89), .B1(n14580), .B2(keyinput90), 
        .ZN(n14579) );
  OAI221_X1 U16415 ( .B1(n14581), .B2(keyinput89), .C1(n14580), .C2(keyinput90), .A(n14579), .ZN(n14592) );
  AOI22_X1 U16416 ( .A1(n14583), .A2(keyinput50), .B1(n9659), .B2(keyinput101), 
        .ZN(n14582) );
  OAI221_X1 U16417 ( .B1(n14583), .B2(keyinput50), .C1(n9659), .C2(keyinput101), .A(n14582), .ZN(n14591) );
  AOI22_X1 U16418 ( .A1(n11851), .A2(keyinput42), .B1(n14585), .B2(keyinput127), .ZN(n14584) );
  OAI221_X1 U16419 ( .B1(n11851), .B2(keyinput42), .C1(n14585), .C2(
        keyinput127), .A(n14584), .ZN(n14590) );
  INV_X1 U16420 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14587) );
  AOI22_X1 U16421 ( .A1(n14588), .A2(keyinput0), .B1(keyinput18), .B2(n14587), 
        .ZN(n14586) );
  OAI221_X1 U16422 ( .B1(n14588), .B2(keyinput0), .C1(n14587), .C2(keyinput18), 
        .A(n14586), .ZN(n14589) );
  NOR4_X1 U16423 ( .A1(n14592), .A2(n14591), .A3(n14590), .A4(n14589), .ZN(
        n14620) );
  INV_X1 U16424 ( .A(P3_B_REG_SCAN_IN), .ZN(n14594) );
  AOI22_X1 U16425 ( .A1(n14594), .A2(keyinput58), .B1(keyinput95), .B2(n8568), 
        .ZN(n14593) );
  OAI221_X1 U16426 ( .B1(n14594), .B2(keyinput58), .C1(n8568), .C2(keyinput95), 
        .A(n14593), .ZN(n14606) );
  INV_X1 U16427 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n14596) );
  AOI22_X1 U16428 ( .A1(n14597), .A2(keyinput109), .B1(n14596), .B2(keyinput62), .ZN(n14595) );
  OAI221_X1 U16429 ( .B1(n14597), .B2(keyinput109), .C1(n14596), .C2(
        keyinput62), .A(n14595), .ZN(n14605) );
  AOI22_X1 U16430 ( .A1(n14600), .A2(keyinput35), .B1(n14599), .B2(keyinput36), 
        .ZN(n14598) );
  OAI221_X1 U16431 ( .B1(n14600), .B2(keyinput35), .C1(n14599), .C2(keyinput36), .A(n14598), .ZN(n14604) );
  XNOR2_X1 U16432 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput112), .ZN(n14602)
         );
  XNOR2_X1 U16433 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput44), .ZN(n14601)
         );
  NAND2_X1 U16434 ( .A1(n14602), .A2(n14601), .ZN(n14603) );
  NOR4_X1 U16435 ( .A1(n14606), .A2(n14605), .A3(n14604), .A4(n14603), .ZN(
        n14619) );
  INV_X1 U16436 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15599) );
  AOI22_X1 U16437 ( .A1(n14608), .A2(keyinput104), .B1(keyinput54), .B2(n15599), .ZN(n14607) );
  OAI221_X1 U16438 ( .B1(n14608), .B2(keyinput104), .C1(n15599), .C2(
        keyinput54), .A(n14607), .ZN(n14617) );
  AOI22_X1 U16439 ( .A1(n14610), .A2(keyinput91), .B1(keyinput81), .B2(n10451), 
        .ZN(n14609) );
  OAI221_X1 U16440 ( .B1(n14610), .B2(keyinput91), .C1(n10451), .C2(keyinput81), .A(n14609), .ZN(n14616) );
  INV_X1 U16441 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15121) );
  AOI22_X1 U16442 ( .A1(n10898), .A2(keyinput116), .B1(keyinput115), .B2(
        n15121), .ZN(n14611) );
  OAI221_X1 U16443 ( .B1(n10898), .B2(keyinput116), .C1(n15121), .C2(
        keyinput115), .A(n14611), .ZN(n14615) );
  XNOR2_X1 U16444 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput121), .ZN(n14613)
         );
  XNOR2_X1 U16445 ( .A(keyinput99), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14612)
         );
  NAND2_X1 U16446 ( .A1(n14613), .A2(n14612), .ZN(n14614) );
  NOR4_X1 U16447 ( .A1(n14617), .A2(n14616), .A3(n14615), .A4(n14614), .ZN(
        n14618) );
  NAND4_X1 U16448 ( .A1(n14621), .A2(n14620), .A3(n14619), .A4(n14618), .ZN(
        n14752) );
  AOI22_X1 U16449 ( .A1(n14623), .A2(keyinput102), .B1(keyinput124), .B2(
        n10524), .ZN(n14622) );
  OAI221_X1 U16450 ( .B1(n14623), .B2(keyinput102), .C1(n10524), .C2(
        keyinput124), .A(n14622), .ZN(n14633) );
  AOI22_X1 U16451 ( .A1(n7910), .A2(keyinput20), .B1(n13132), .B2(keyinput70), 
        .ZN(n14624) );
  OAI221_X1 U16452 ( .B1(n7910), .B2(keyinput20), .C1(n13132), .C2(keyinput70), 
        .A(n14624), .ZN(n14632) );
  INV_X1 U16453 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14906) );
  AOI22_X1 U16454 ( .A1(n14906), .A2(keyinput30), .B1(n14626), .B2(keyinput97), 
        .ZN(n14625) );
  OAI221_X1 U16455 ( .B1(n14906), .B2(keyinput30), .C1(n14626), .C2(keyinput97), .A(n14625), .ZN(n14631) );
  XOR2_X1 U16456 ( .A(n14627), .B(keyinput88), .Z(n14629) );
  XNOR2_X1 U16457 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput55), .ZN(n14628)
         );
  NAND2_X1 U16458 ( .A1(n14629), .A2(n14628), .ZN(n14630) );
  NOR4_X1 U16459 ( .A1(n14633), .A2(n14632), .A3(n14631), .A4(n14630), .ZN(
        n14674) );
  AOI22_X1 U16460 ( .A1(n14636), .A2(keyinput39), .B1(keyinput64), .B2(n14635), 
        .ZN(n14634) );
  OAI221_X1 U16461 ( .B1(n14636), .B2(keyinput39), .C1(n14635), .C2(keyinput64), .A(n14634), .ZN(n14644) );
  AOI22_X1 U16462 ( .A1(n15303), .A2(keyinput11), .B1(n10379), .B2(keyinput21), 
        .ZN(n14637) );
  OAI221_X1 U16463 ( .B1(n15303), .B2(keyinput11), .C1(n10379), .C2(keyinput21), .A(n14637), .ZN(n14643) );
  AOI22_X1 U16464 ( .A1(n9564), .A2(keyinput24), .B1(keyinput56), .B2(n14639), 
        .ZN(n14638) );
  OAI221_X1 U16465 ( .B1(n9564), .B2(keyinput24), .C1(n14639), .C2(keyinput56), 
        .A(n14638), .ZN(n14642) );
  AOI22_X1 U16466 ( .A1(n9897), .A2(keyinput96), .B1(keyinput43), .B2(n14102), 
        .ZN(n14640) );
  OAI221_X1 U16467 ( .B1(n9897), .B2(keyinput96), .C1(n14102), .C2(keyinput43), 
        .A(n14640), .ZN(n14641) );
  NOR4_X1 U16468 ( .A1(n14644), .A2(n14643), .A3(n14642), .A4(n14641), .ZN(
        n14673) );
  AOI22_X1 U16469 ( .A1(n15306), .A2(keyinput65), .B1(keyinput93), .B2(n14646), 
        .ZN(n14645) );
  OAI221_X1 U16470 ( .B1(n15306), .B2(keyinput65), .C1(n14646), .C2(keyinput93), .A(n14645), .ZN(n14655) );
  AOI22_X1 U16471 ( .A1(n10867), .A2(keyinput117), .B1(n14648), .B2(keyinput28), .ZN(n14647) );
  OAI221_X1 U16472 ( .B1(n10867), .B2(keyinput117), .C1(n14648), .C2(
        keyinput28), .A(n14647), .ZN(n14654) );
  XNOR2_X1 U16473 ( .A(SI_27_), .B(keyinput111), .ZN(n14652) );
  XNOR2_X1 U16474 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput52), .ZN(n14651) );
  XNOR2_X1 U16475 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput85), .ZN(n14650)
         );
  XNOR2_X1 U16476 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput83), .ZN(n14649) );
  NAND4_X1 U16477 ( .A1(n14652), .A2(n14651), .A3(n14650), .A4(n14649), .ZN(
        n14653) );
  NOR3_X1 U16478 ( .A1(n14655), .A2(n14654), .A3(n14653), .ZN(n14672) );
  AOI22_X1 U16479 ( .A1(n14658), .A2(keyinput13), .B1(keyinput61), .B2(n14657), 
        .ZN(n14656) );
  OAI221_X1 U16480 ( .B1(n14658), .B2(keyinput13), .C1(n14657), .C2(keyinput61), .A(n14656), .ZN(n14670) );
  AOI22_X1 U16481 ( .A1(n14661), .A2(keyinput47), .B1(keyinput10), .B2(n14660), 
        .ZN(n14659) );
  OAI221_X1 U16482 ( .B1(n14661), .B2(keyinput47), .C1(n14660), .C2(keyinput10), .A(n14659), .ZN(n14669) );
  AOI22_X1 U16483 ( .A1(n14664), .A2(keyinput119), .B1(keyinput26), .B2(n14663), .ZN(n14662) );
  OAI221_X1 U16484 ( .B1(n14664), .B2(keyinput119), .C1(n14663), .C2(
        keyinput26), .A(n14662), .ZN(n14668) );
  XOR2_X1 U16485 ( .A(n13632), .B(keyinput126), .Z(n14666) );
  XNOR2_X1 U16486 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput118), .ZN(n14665) );
  NAND2_X1 U16487 ( .A1(n14666), .A2(n14665), .ZN(n14667) );
  NOR4_X1 U16488 ( .A1(n14670), .A2(n14669), .A3(n14668), .A4(n14667), .ZN(
        n14671) );
  NAND4_X1 U16489 ( .A1(n14674), .A2(n14673), .A3(n14672), .A4(n14671), .ZN(
        n14751) );
  AOI22_X1 U16490 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput17), .B1(
        P2_IR_REG_16__SCAN_IN), .B2(keyinput1), .ZN(n14675) );
  OAI221_X1 U16491 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput17), .C1(
        P2_IR_REG_16__SCAN_IN), .C2(keyinput1), .A(n14675), .ZN(n14682) );
  AOI22_X1 U16492 ( .A1(P3_REG0_REG_24__SCAN_IN), .A2(keyinput75), .B1(
        P3_D_REG_0__SCAN_IN), .B2(keyinput69), .ZN(n14676) );
  OAI221_X1 U16493 ( .B1(P3_REG0_REG_24__SCAN_IN), .B2(keyinput75), .C1(
        P3_D_REG_0__SCAN_IN), .C2(keyinput69), .A(n14676), .ZN(n14681) );
  AOI22_X1 U16494 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(keyinput31), .B1(SI_1_), 
        .B2(keyinput68), .ZN(n14677) );
  OAI221_X1 U16495 ( .B1(P2_REG1_REG_27__SCAN_IN), .B2(keyinput31), .C1(SI_1_), 
        .C2(keyinput68), .A(n14677), .ZN(n14680) );
  AOI22_X1 U16496 ( .A1(P1_REG1_REG_31__SCAN_IN), .A2(keyinput32), .B1(
        P3_REG1_REG_5__SCAN_IN), .B2(keyinput73), .ZN(n14678) );
  OAI221_X1 U16497 ( .B1(P1_REG1_REG_31__SCAN_IN), .B2(keyinput32), .C1(
        P3_REG1_REG_5__SCAN_IN), .C2(keyinput73), .A(n14678), .ZN(n14679) );
  NOR4_X1 U16498 ( .A1(n14682), .A2(n14681), .A3(n14680), .A4(n14679), .ZN(
        n14712) );
  AOI22_X1 U16499 ( .A1(SI_6_), .A2(keyinput3), .B1(P3_IR_REG_22__SCAN_IN), 
        .B2(keyinput14), .ZN(n14683) );
  OAI221_X1 U16500 ( .B1(SI_6_), .B2(keyinput3), .C1(P3_IR_REG_22__SCAN_IN), 
        .C2(keyinput14), .A(n14683), .ZN(n14690) );
  AOI22_X1 U16501 ( .A1(P1_REG0_REG_3__SCAN_IN), .A2(keyinput106), .B1(
        P1_D_REG_31__SCAN_IN), .B2(keyinput79), .ZN(n14684) );
  OAI221_X1 U16502 ( .B1(P1_REG0_REG_3__SCAN_IN), .B2(keyinput106), .C1(
        P1_D_REG_31__SCAN_IN), .C2(keyinput79), .A(n14684), .ZN(n14689) );
  AOI22_X1 U16503 ( .A1(P3_REG0_REG_6__SCAN_IN), .A2(keyinput41), .B1(
        P3_REG2_REG_27__SCAN_IN), .B2(keyinput84), .ZN(n14685) );
  OAI221_X1 U16504 ( .B1(P3_REG0_REG_6__SCAN_IN), .B2(keyinput41), .C1(
        P3_REG2_REG_27__SCAN_IN), .C2(keyinput84), .A(n14685), .ZN(n14688) );
  AOI22_X1 U16505 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(keyinput66), .B1(
        P3_IR_REG_20__SCAN_IN), .B2(keyinput51), .ZN(n14686) );
  OAI221_X1 U16506 ( .B1(P1_REG0_REG_29__SCAN_IN), .B2(keyinput66), .C1(
        P3_IR_REG_20__SCAN_IN), .C2(keyinput51), .A(n14686), .ZN(n14687) );
  NOR4_X1 U16507 ( .A1(n14690), .A2(n14689), .A3(n14688), .A4(n14687), .ZN(
        n14711) );
  AOI22_X1 U16508 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(keyinput48), .B1(
        P2_IR_REG_21__SCAN_IN), .B2(keyinput22), .ZN(n14691) );
  OAI221_X1 U16509 ( .B1(P1_REG3_REG_14__SCAN_IN), .B2(keyinput48), .C1(
        P2_IR_REG_21__SCAN_IN), .C2(keyinput22), .A(n14691), .ZN(n14700) );
  AOI22_X1 U16510 ( .A1(P1_D_REG_18__SCAN_IN), .A2(keyinput108), .B1(
        P3_REG2_REG_29__SCAN_IN), .B2(keyinput110), .ZN(n14692) );
  OAI221_X1 U16511 ( .B1(P1_D_REG_18__SCAN_IN), .B2(keyinput108), .C1(
        P3_REG2_REG_29__SCAN_IN), .C2(keyinput110), .A(n14692), .ZN(n14699) );
  AOI22_X1 U16512 ( .A1(n7751), .A2(keyinput123), .B1(n14694), .B2(keyinput94), 
        .ZN(n14693) );
  OAI221_X1 U16513 ( .B1(n7751), .B2(keyinput123), .C1(n14694), .C2(keyinput94), .A(n14693), .ZN(n14698) );
  AOI22_X1 U16514 ( .A1(n8246), .A2(keyinput125), .B1(keyinput7), .B2(n14696), 
        .ZN(n14695) );
  OAI221_X1 U16515 ( .B1(n8246), .B2(keyinput125), .C1(n14696), .C2(keyinput7), 
        .A(n14695), .ZN(n14697) );
  NOR4_X1 U16516 ( .A1(n14700), .A2(n14699), .A3(n14698), .A4(n14697), .ZN(
        n14710) );
  AOI22_X1 U16517 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(keyinput76), .B1(SI_4_), 
        .B2(keyinput9), .ZN(n14701) );
  OAI221_X1 U16518 ( .B1(P1_REG1_REG_24__SCAN_IN), .B2(keyinput76), .C1(SI_4_), 
        .C2(keyinput9), .A(n14701), .ZN(n14708) );
  AOI22_X1 U16519 ( .A1(P2_REG1_REG_21__SCAN_IN), .A2(keyinput16), .B1(SI_9_), 
        .B2(keyinput19), .ZN(n14702) );
  OAI221_X1 U16520 ( .B1(P2_REG1_REG_21__SCAN_IN), .B2(keyinput16), .C1(SI_9_), 
        .C2(keyinput19), .A(n14702), .ZN(n14707) );
  AOI22_X1 U16521 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(keyinput2), .B1(SI_18_), 
        .B2(keyinput86), .ZN(n14703) );
  OAI221_X1 U16522 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(keyinput2), .C1(SI_18_), 
        .C2(keyinput86), .A(n14703), .ZN(n14706) );
  AOI22_X1 U16523 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput4), .B1(n6829), 
        .B2(keyinput113), .ZN(n14704) );
  OAI221_X1 U16524 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput4), .C1(n6829), 
        .C2(keyinput113), .A(n14704), .ZN(n14705) );
  NOR4_X1 U16525 ( .A1(n14708), .A2(n14707), .A3(n14706), .A4(n14705), .ZN(
        n14709) );
  NAND4_X1 U16526 ( .A1(n14712), .A2(n14711), .A3(n14710), .A4(n14709), .ZN(
        n14750) );
  AOI22_X1 U16527 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(keyinput105), .B1(
        P3_IR_REG_7__SCAN_IN), .B2(keyinput67), .ZN(n14713) );
  OAI221_X1 U16528 ( .B1(P1_REG1_REG_28__SCAN_IN), .B2(keyinput105), .C1(
        P3_IR_REG_7__SCAN_IN), .C2(keyinput67), .A(n14713), .ZN(n14720) );
  AOI22_X1 U16529 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput8), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput6), .ZN(n14714) );
  OAI221_X1 U16530 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput8), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput6), .A(n14714), .ZN(n14719) );
  AOI22_X1 U16531 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput120), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(keyinput46), .ZN(n14715) );
  OAI221_X1 U16532 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput120), .C1(
        P1_REG2_REG_1__SCAN_IN), .C2(keyinput46), .A(n14715), .ZN(n14718) );
  AOI22_X1 U16533 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(keyinput63), .B1(SI_14_), 
        .B2(keyinput87), .ZN(n14716) );
  OAI221_X1 U16534 ( .B1(P1_REG3_REG_6__SCAN_IN), .B2(keyinput63), .C1(SI_14_), 
        .C2(keyinput87), .A(n14716), .ZN(n14717) );
  NOR4_X1 U16535 ( .A1(n14720), .A2(n14719), .A3(n14718), .A4(n14717), .ZN(
        n14748) );
  AOI22_X1 U16536 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(keyinput122), .B1(
        P2_REG2_REG_31__SCAN_IN), .B2(keyinput80), .ZN(n14721) );
  OAI221_X1 U16537 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(keyinput122), .C1(
        P2_REG2_REG_31__SCAN_IN), .C2(keyinput80), .A(n14721), .ZN(n14728) );
  AOI22_X1 U16538 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(keyinput92), .B1(
        P2_D_REG_20__SCAN_IN), .B2(keyinput45), .ZN(n14722) );
  OAI221_X1 U16539 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(keyinput92), .C1(
        P2_D_REG_20__SCAN_IN), .C2(keyinput45), .A(n14722), .ZN(n14727) );
  AOI22_X1 U16540 ( .A1(P3_D_REG_19__SCAN_IN), .A2(keyinput60), .B1(
        P3_REG3_REG_9__SCAN_IN), .B2(keyinput27), .ZN(n14723) );
  OAI221_X1 U16541 ( .B1(P3_D_REG_19__SCAN_IN), .B2(keyinput60), .C1(
        P3_REG3_REG_9__SCAN_IN), .C2(keyinput27), .A(n14723), .ZN(n14726) );
  AOI22_X1 U16542 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(keyinput59), .B1(SI_17_), 
        .B2(keyinput107), .ZN(n14724) );
  OAI221_X1 U16543 ( .B1(P3_DATAO_REG_0__SCAN_IN), .B2(keyinput59), .C1(SI_17_), .C2(keyinput107), .A(n14724), .ZN(n14725) );
  NOR4_X1 U16544 ( .A1(n14728), .A2(n14727), .A3(n14726), .A4(n14725), .ZN(
        n14747) );
  AOI22_X1 U16545 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput82), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput98), .ZN(n14729) );
  OAI221_X1 U16546 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput82), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput98), .A(n14729), .ZN(n14736) );
  AOI22_X1 U16547 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(keyinput100), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput103), .ZN(n14730) );
  OAI221_X1 U16548 ( .B1(P3_DATAO_REG_30__SCAN_IN), .B2(keyinput100), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput103), .A(n14730), .ZN(n14735)
         );
  AOI22_X1 U16549 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(keyinput71), .B1(
        P2_D_REG_16__SCAN_IN), .B2(keyinput74), .ZN(n14731) );
  OAI221_X1 U16550 ( .B1(P3_ADDR_REG_13__SCAN_IN), .B2(keyinput71), .C1(
        P2_D_REG_16__SCAN_IN), .C2(keyinput74), .A(n14731), .ZN(n14734) );
  AOI22_X1 U16551 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(keyinput23), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput78), .ZN(n14732) );
  OAI221_X1 U16552 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(keyinput23), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput78), .A(n14732), .ZN(n14733) );
  NOR4_X1 U16553 ( .A1(n14736), .A2(n14735), .A3(n14734), .A4(n14733), .ZN(
        n14746) );
  AOI22_X1 U16554 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(keyinput5), .B1(
        P3_ADDR_REG_17__SCAN_IN), .B2(keyinput49), .ZN(n14737) );
  OAI221_X1 U16555 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(keyinput5), .C1(
        P3_ADDR_REG_17__SCAN_IN), .C2(keyinput49), .A(n14737), .ZN(n14744) );
  AOI22_X1 U16556 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(keyinput38), .B1(
        P3_REG2_REG_5__SCAN_IN), .B2(keyinput29), .ZN(n14738) );
  OAI221_X1 U16557 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(keyinput38), .C1(
        P3_REG2_REG_5__SCAN_IN), .C2(keyinput29), .A(n14738), .ZN(n14743) );
  AOI22_X1 U16558 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(keyinput57), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput77), .ZN(n14739) );
  OAI221_X1 U16559 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(keyinput57), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput77), .A(n14739), .ZN(n14742) );
  AOI22_X1 U16560 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(keyinput12), .B1(
        P3_REG2_REG_8__SCAN_IN), .B2(keyinput34), .ZN(n14740) );
  OAI221_X1 U16561 ( .B1(P2_REG0_REG_14__SCAN_IN), .B2(keyinput12), .C1(
        P3_REG2_REG_8__SCAN_IN), .C2(keyinput34), .A(n14740), .ZN(n14741) );
  NOR4_X1 U16562 ( .A1(n14744), .A2(n14743), .A3(n14742), .A4(n14741), .ZN(
        n14745) );
  NAND4_X1 U16563 ( .A1(n14748), .A2(n14747), .A3(n14746), .A4(n14745), .ZN(
        n14749) );
  NOR4_X1 U16564 ( .A1(n14752), .A2(n14751), .A3(n14750), .A4(n14749), .ZN(
        n14753) );
  OAI21_X1 U16565 ( .B1(n14755), .B2(n14754), .A(n14753), .ZN(n14761) );
  XOR2_X1 U16566 ( .A(n14761), .B(n14760), .Z(P1_U3335) );
  INV_X1 U16567 ( .A(n14762), .ZN(n14763) );
  MUX2_X1 U16568 ( .A(n14763), .B(n6664), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  OAI21_X1 U16569 ( .B1(n14766), .B2(n14765), .A(n14764), .ZN(n14767) );
  XNOR2_X1 U16570 ( .A(n14767), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16571 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14768) );
  OAI21_X1 U16572 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14768), 
        .ZN(U28) );
  AOI21_X1 U16573 ( .B1(n6842), .B2(n6829), .A(P3_RD_REG_SCAN_IN), .ZN(n14769)
         );
  OAI21_X1 U16574 ( .B1(n6842), .B2(n6829), .A(n14769), .ZN(U29) );
  OAI21_X1 U16575 ( .B1(n14772), .B2(n14771), .A(n14770), .ZN(n14773) );
  XNOR2_X1 U16576 ( .A(n14773), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16577 ( .B1(n14776), .B2(n14775), .A(n14774), .ZN(SUB_1596_U57) );
  OAI22_X1 U16578 ( .A1(n14778), .A2(n12306), .B1(n14777), .B2(n12423), .ZN(
        n14779) );
  INV_X1 U16579 ( .A(n14779), .ZN(n14780) );
  OAI21_X1 U16580 ( .B1(P3_U3151), .B2(n14781), .A(n14780), .ZN(P3_U3281) );
  OAI21_X1 U16581 ( .B1(n14784), .B2(n14783), .A(n14782), .ZN(SUB_1596_U55) );
  AOI21_X1 U16582 ( .B1(n14787), .B2(n14786), .A(n14785), .ZN(SUB_1596_U54) );
  AOI21_X1 U16583 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n14791) );
  XOR2_X1 U16584 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14791), .Z(SUB_1596_U70)
         );
  INV_X1 U16585 ( .A(n14792), .ZN(n14797) );
  OAI21_X1 U16586 ( .B1(n14794), .B2(n15185), .A(n14793), .ZN(n14796) );
  AOI211_X1 U16587 ( .C1(n15190), .C2(n14797), .A(n14796), .B(n14795), .ZN(
        n14799) );
  AOI22_X1 U16588 ( .A1(n15201), .A2(n14799), .B1(n14798), .B2(n15199), .ZN(
        P1_U3495) );
  AOI22_X1 U16589 ( .A1(n15215), .A2(n14799), .B1(n11018), .B2(n15213), .ZN(
        P1_U3540) );
  XNOR2_X1 U16590 ( .A(n14800), .B(n14811), .ZN(n14986) );
  OAI22_X1 U16591 ( .A1(n14804), .A2(n14803), .B1(n14802), .B2(n14801), .ZN(
        n14805) );
  AOI21_X1 U16592 ( .B1(n14806), .B2(n14978), .A(n14805), .ZN(n14807) );
  OAI21_X1 U16593 ( .B1(n7372), .B2(n15107), .A(n14807), .ZN(n14808) );
  AOI21_X1 U16594 ( .B1(n14986), .B2(n14809), .A(n14808), .ZN(n14819) );
  XNOR2_X1 U16595 ( .A(n14810), .B(n14811), .ZN(n14813) );
  AOI22_X1 U16596 ( .A1(n14813), .A2(n15098), .B1(n14812), .B2(n14955), .ZN(
        n14984) );
  OAI211_X1 U16597 ( .C1(n7372), .C2(n7373), .A(n15111), .B(n14815), .ZN(
        n14982) );
  OAI22_X1 U16598 ( .A1(n14984), .A2(n15118), .B1(n14982), .B2(n14816), .ZN(
        n14817) );
  INV_X1 U16599 ( .A(n14817), .ZN(n14818) );
  NAND2_X1 U16600 ( .A1(n14819), .A2(n14818), .ZN(P1_U3280) );
  OAI21_X1 U16601 ( .B1(n14822), .B2(n14821), .A(n14820), .ZN(n14823) );
  XNOR2_X1 U16602 ( .A(n14823), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  AOI22_X1 U16603 ( .A1(n14825), .A2(n7036), .B1(n15460), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14839) );
  XNOR2_X1 U16604 ( .A(n14826), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n14831) );
  AOI211_X1 U16605 ( .C1(n14829), .C2(n14828), .A(n15456), .B(n14827), .ZN(
        n14830) );
  AOI21_X1 U16606 ( .B1(n14831), .B2(n15463), .A(n14830), .ZN(n14838) );
  NAND2_X1 U16607 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14837)
         );
  OAI221_X1 U16608 ( .B1(n14835), .B2(n14834), .C1(n14835), .C2(n14833), .A(
        n14832), .ZN(n14836) );
  NAND4_X1 U16609 ( .A1(n14839), .A2(n14838), .A3(n14837), .A4(n14836), .ZN(
        P3_U3199) );
  XNOR2_X1 U16610 ( .A(n14840), .B(n14844), .ZN(n14842) );
  AOI222_X1 U16611 ( .A1(n15511), .A2(n14842), .B1(n14841), .B2(n14853), .C1(
        n14854), .C2(n14851), .ZN(n14871) );
  AOI22_X1 U16612 ( .A1(n15517), .A2(n14843), .B1(n13166), .B2(
        P3_REG2_REG_13__SCAN_IN), .ZN(n14849) );
  XNOR2_X1 U16613 ( .A(n14845), .B(n14844), .ZN(n14874) );
  INV_X1 U16614 ( .A(n14846), .ZN(n14847) );
  NOR2_X1 U16615 ( .A1(n14847), .A2(n15545), .ZN(n14873) );
  AOI22_X1 U16616 ( .A1(n14874), .A2(n14861), .B1(n14860), .B2(n14873), .ZN(
        n14848) );
  OAI211_X1 U16617 ( .C1(n13166), .C2(n14871), .A(n14849), .B(n14848), .ZN(
        P3_U3220) );
  XNOR2_X1 U16618 ( .A(n14850), .B(n9987), .ZN(n14855) );
  AOI222_X1 U16619 ( .A1(n15511), .A2(n14855), .B1(n14854), .B2(n14853), .C1(
        n14852), .C2(n14851), .ZN(n14879) );
  AOI22_X1 U16620 ( .A1(n15517), .A2(n14856), .B1(n13166), .B2(
        P3_REG2_REG_11__SCAN_IN), .ZN(n14863) );
  OAI21_X1 U16621 ( .B1(n14858), .B2(n9987), .A(n14857), .ZN(n14882) );
  NOR2_X1 U16622 ( .A1(n14859), .A2(n15545), .ZN(n14881) );
  AOI22_X1 U16623 ( .A1(n14882), .A2(n14861), .B1(n14860), .B2(n14881), .ZN(
        n14862) );
  OAI211_X1 U16624 ( .C1(n13166), .C2(n14879), .A(n14863), .B(n14862), .ZN(
        P3_U3222) );
  OR2_X1 U16625 ( .A1(n14864), .A2(n15545), .ZN(n14865) );
  AOI22_X1 U16626 ( .A1(n15585), .A2(n14885), .B1(n14866), .B2(n15583), .ZN(
        P3_U3490) );
  OR2_X1 U16627 ( .A1(n14867), .A2(n15545), .ZN(n14869) );
  AOI22_X1 U16628 ( .A1(n15585), .A2(n14886), .B1(n14870), .B2(n15583), .ZN(
        P3_U3489) );
  INV_X1 U16629 ( .A(n14871), .ZN(n14872) );
  AOI211_X1 U16630 ( .C1(n14874), .C2(n14883), .A(n14873), .B(n14872), .ZN(
        n14890) );
  INV_X1 U16631 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14875) );
  AOI22_X1 U16632 ( .A1(n15585), .A2(n14890), .B1(n14875), .B2(n15583), .ZN(
        P3_U3472) );
  AOI211_X1 U16633 ( .C1(n14878), .C2(n14883), .A(n14877), .B(n14876), .ZN(
        n14891) );
  AOI22_X1 U16634 ( .A1(n15585), .A2(n14891), .B1(n9731), .B2(n15583), .ZN(
        P3_U3471) );
  INV_X1 U16635 ( .A(n14879), .ZN(n14880) );
  AOI211_X1 U16636 ( .C1(n14883), .C2(n14882), .A(n14881), .B(n14880), .ZN(
        n14893) );
  AOI22_X1 U16637 ( .A1(n15585), .A2(n14893), .B1(n9707), .B2(n15583), .ZN(
        P3_U3470) );
  INV_X1 U16638 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14884) );
  AOI22_X1 U16639 ( .A1(n15570), .A2(n14885), .B1(n14884), .B2(n15568), .ZN(
        P3_U3458) );
  INV_X1 U16640 ( .A(n14886), .ZN(n14887) );
  OAI22_X1 U16641 ( .A1(n15568), .A2(n14887), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n15570), .ZN(n14888) );
  INV_X1 U16642 ( .A(n14888), .ZN(P3_U3457) );
  INV_X1 U16643 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14889) );
  AOI22_X1 U16644 ( .A1(n15570), .A2(n14890), .B1(n14889), .B2(n15568), .ZN(
        P3_U3429) );
  AOI22_X1 U16645 ( .A1(n15570), .A2(n14891), .B1(n9733), .B2(n15568), .ZN(
        P3_U3426) );
  INV_X1 U16646 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14892) );
  AOI22_X1 U16647 ( .A1(n15570), .A2(n14893), .B1(n14892), .B2(n15568), .ZN(
        P3_U3423) );
  OAI211_X1 U16648 ( .C1(n14896), .C2(n15342), .A(n14895), .B(n14894), .ZN(
        n14897) );
  AOI21_X1 U16649 ( .B1(n14898), .B2(n15339), .A(n14897), .ZN(n14905) );
  AOI22_X1 U16650 ( .A1(n13815), .A2(n14905), .B1(n11616), .B2(n15371), .ZN(
        P2_U3512) );
  INV_X1 U16651 ( .A(n14899), .ZN(n14904) );
  OAI21_X1 U16652 ( .B1(n14901), .B2(n15342), .A(n14900), .ZN(n14903) );
  AOI211_X1 U16653 ( .C1(n9298), .C2(n14904), .A(n14903), .B(n14902), .ZN(
        n14907) );
  AOI22_X1 U16654 ( .A1(n13815), .A2(n14907), .B1(n11397), .B2(n15371), .ZN(
        P2_U3511) );
  AOI22_X1 U16655 ( .A1(n15364), .A2(n14905), .B1(n8041), .B2(n15362), .ZN(
        P2_U3469) );
  AOI22_X1 U16656 ( .A1(n15364), .A2(n14907), .B1(n14906), .B2(n15362), .ZN(
        P2_U3466) );
  OAI22_X1 U16657 ( .A1(n14911), .A2(n14910), .B1(n14909), .B2(n14908), .ZN(
        n14920) );
  AOI21_X1 U16658 ( .B1(n14914), .B2(n14913), .A(n14912), .ZN(n14915) );
  INV_X1 U16659 ( .A(n14915), .ZN(n14918) );
  AOI21_X1 U16660 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(n14919) );
  AOI211_X1 U16661 ( .C1(n14921), .C2(n14971), .A(n14920), .B(n14919), .ZN(
        n14923) );
  OAI211_X1 U16662 ( .C1(n14964), .C2(n14924), .A(n14923), .B(n14922), .ZN(
        P1_U3215) );
  AND2_X1 U16663 ( .A1(n14925), .A2(n14980), .ZN(n15193) );
  AOI22_X1 U16664 ( .A1(n15193), .A2(n14926), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14936) );
  NAND2_X1 U16665 ( .A1(n14979), .A2(n14927), .ZN(n14928) );
  NAND2_X1 U16666 ( .A1(n14929), .A2(n14928), .ZN(n15192) );
  OAI211_X1 U16667 ( .C1(n14931), .C2(n14930), .A(n14940), .B(n14960), .ZN(
        n14932) );
  INV_X1 U16668 ( .A(n14932), .ZN(n14933) );
  AOI21_X1 U16669 ( .B1(n14934), .B2(n15192), .A(n14933), .ZN(n14935) );
  OAI211_X1 U16670 ( .C1(n14937), .C2(n14964), .A(n14936), .B(n14935), .ZN(
        P1_U3217) );
  AOI21_X1 U16671 ( .B1(n14940), .B2(n14939), .A(n14938), .ZN(n14941) );
  OAI21_X1 U16672 ( .B1(n14942), .B2(n14941), .A(n14960), .ZN(n14945) );
  AOI22_X1 U16673 ( .A1(n14956), .A2(n14943), .B1(n14954), .B2(n14978), .ZN(
        n14944) );
  OAI211_X1 U16674 ( .C1(n6956), .C2(n14958), .A(n14945), .B(n14944), .ZN(
        n14946) );
  INV_X1 U16675 ( .A(n14946), .ZN(n14948) );
  OAI211_X1 U16676 ( .C1(n14964), .C2(n14949), .A(n14948), .B(n14947), .ZN(
        P1_U3236) );
  OAI21_X1 U16677 ( .B1(n14952), .B2(n14951), .A(n14950), .ZN(n14961) );
  AOI22_X1 U16678 ( .A1(n14956), .A2(n14955), .B1(n14954), .B2(n14953), .ZN(
        n14957) );
  OAI21_X1 U16679 ( .B1(n6955), .B2(n14958), .A(n14957), .ZN(n14959) );
  AOI21_X1 U16680 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n14962) );
  NAND2_X1 U16681 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15061)
         );
  OAI211_X1 U16682 ( .C1(n14964), .C2(n14963), .A(n14962), .B(n15061), .ZN(
        P1_U3241) );
  OAI211_X1 U16683 ( .C1(n14967), .C2(n15185), .A(n14966), .B(n14965), .ZN(
        n14969) );
  AOI211_X1 U16684 ( .C1(n15198), .C2(n14970), .A(n14969), .B(n14968), .ZN(
        n14993) );
  AOI22_X1 U16685 ( .A1(n15215), .A2(n14993), .B1(n11920), .B2(n15213), .ZN(
        P1_U3544) );
  NAND3_X1 U16686 ( .A1(n14973), .A2(n14972), .A3(n15198), .ZN(n14975) );
  OAI211_X1 U16687 ( .C1(n7370), .C2(n15185), .A(n14975), .B(n14974), .ZN(
        n14977) );
  NOR2_X1 U16688 ( .A1(n14977), .A2(n14976), .ZN(n14995) );
  AOI22_X1 U16689 ( .A1(n15215), .A2(n14995), .B1(n11922), .B2(n15213), .ZN(
        P1_U3542) );
  AOI22_X1 U16690 ( .A1(n14981), .A2(n14980), .B1(n14979), .B2(n14978), .ZN(
        n14983) );
  NAND3_X1 U16691 ( .A1(n14984), .A2(n14983), .A3(n14982), .ZN(n14985) );
  AOI21_X1 U16692 ( .B1(n14986), .B2(n15198), .A(n14985), .ZN(n14997) );
  AOI22_X1 U16693 ( .A1(n15215), .A2(n14997), .B1(n14987), .B2(n15213), .ZN(
        P1_U3541) );
  OAI22_X1 U16694 ( .A1(n14988), .A2(n15125), .B1(n6956), .B2(n15185), .ZN(
        n14990) );
  AOI211_X1 U16695 ( .C1(n14991), .C2(n15198), .A(n14990), .B(n14989), .ZN(
        n14999) );
  AOI22_X1 U16696 ( .A1(n15215), .A2(n14999), .B1(n11015), .B2(n15213), .ZN(
        P1_U3539) );
  INV_X1 U16697 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U16698 ( .A1(n15201), .A2(n14993), .B1(n14992), .B2(n15199), .ZN(
        P1_U3507) );
  INV_X1 U16699 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14994) );
  AOI22_X1 U16700 ( .A1(n15201), .A2(n14995), .B1(n14994), .B2(n15199), .ZN(
        P1_U3501) );
  INV_X1 U16701 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14996) );
  AOI22_X1 U16702 ( .A1(n15201), .A2(n14997), .B1(n14996), .B2(n15199), .ZN(
        P1_U3498) );
  INV_X1 U16703 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14998) );
  AOI22_X1 U16704 ( .A1(n15201), .A2(n14999), .B1(n14998), .B2(n15199), .ZN(
        P1_U3492) );
  AOI21_X1 U16705 ( .B1(n15002), .B2(n15001), .A(n15000), .ZN(n15003) );
  XOR2_X1 U16706 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15003), .Z(SUB_1596_U69)
         );
  OAI222_X1 U16707 ( .A1(n15008), .A2(n15007), .B1(n15008), .B2(n15006), .C1(
        n15005), .C2(n15004), .ZN(SUB_1596_U68) );
  AOI21_X1 U16708 ( .B1(n15010), .B2(n15009), .A(n6816), .ZN(n15011) );
  XOR2_X1 U16709 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n15011), .Z(SUB_1596_U67)
         );
  OAI21_X1 U16710 ( .B1(n15014), .B2(n15013), .A(n15012), .ZN(n15015) );
  XNOR2_X1 U16711 ( .A(n15015), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16712 ( .A1(n15268), .A2(n15019), .B1(n15268), .B2(n15018), .C1(
        n15017), .C2(n15016), .ZN(SUB_1596_U65) );
  OAI21_X1 U16713 ( .B1(n15022), .B2(n15021), .A(n15020), .ZN(n15023) );
  XNOR2_X1 U16714 ( .A(n15023), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  INV_X1 U16715 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15025) );
  AOI21_X1 U16716 ( .B1(n15026), .B2(n15025), .A(n15024), .ZN(n15027) );
  XNOR2_X1 U16717 ( .A(n15027), .B(n6664), .ZN(n15030) );
  AOI22_X1 U16718 ( .A1(n15031), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15028) );
  OAI21_X1 U16719 ( .B1(n15030), .B2(n15029), .A(n15028), .ZN(P1_U3243) );
  INV_X1 U16720 ( .A(n15031), .ZN(n15063) );
  OAI21_X1 U16721 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15045) );
  INV_X1 U16722 ( .A(n15035), .ZN(n15040) );
  NAND3_X1 U16723 ( .A1(n15038), .A2(n15037), .A3(n15036), .ZN(n15039) );
  NAND2_X1 U16724 ( .A1(n15040), .A2(n15039), .ZN(n15041) );
  AOI222_X1 U16725 ( .A1(n15045), .A2(n15044), .B1(n15043), .B2(n15042), .C1(
        n15041), .C2(n15059), .ZN(n15047) );
  OAI211_X1 U16726 ( .C1(n15048), .C2(n15063), .A(n15047), .B(n15046), .ZN(
        P1_U3255) );
  OAI21_X1 U16727 ( .B1(n15051), .B2(n15050), .A(n15049), .ZN(n15060) );
  AOI21_X1 U16728 ( .B1(n15053), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15052), 
        .ZN(n15057) );
  OAI22_X1 U16729 ( .A1(n15057), .A2(n15056), .B1(n15055), .B2(n15054), .ZN(
        n15058) );
  AOI21_X1 U16730 ( .B1(n15060), .B2(n15059), .A(n15058), .ZN(n15062) );
  OAI211_X1 U16731 ( .C1(n15064), .C2(n15063), .A(n15062), .B(n15061), .ZN(
        P1_U3258) );
  XNOR2_X1 U16732 ( .A(n15065), .B(n15067), .ZN(n15189) );
  XNOR2_X1 U16733 ( .A(n15066), .B(n15067), .ZN(n15069) );
  OAI21_X1 U16734 ( .B1(n15069), .B2(n15083), .A(n15068), .ZN(n15070) );
  AOI21_X1 U16735 ( .B1(n15102), .B2(n15189), .A(n15070), .ZN(n15186) );
  AOI22_X1 U16736 ( .A1(n15105), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n15071), 
        .B2(n15103), .ZN(n15072) );
  OAI21_X1 U16737 ( .B1(n7364), .B2(n15107), .A(n15072), .ZN(n15073) );
  INV_X1 U16738 ( .A(n15073), .ZN(n15078) );
  OAI211_X1 U16739 ( .C1(n7364), .C2(n7365), .A(n15111), .B(n15075), .ZN(
        n15184) );
  INV_X1 U16740 ( .A(n15184), .ZN(n15076) );
  AOI22_X1 U16741 ( .A1(n15189), .A2(n15114), .B1(n15113), .B2(n15076), .ZN(
        n15077) );
  OAI211_X1 U16742 ( .C1(n15118), .C2(n15186), .A(n15078), .B(n15077), .ZN(
        P1_U3284) );
  XNOR2_X1 U16743 ( .A(n15079), .B(n15081), .ZN(n15175) );
  XNOR2_X1 U16744 ( .A(n15080), .B(n15081), .ZN(n15084) );
  OAI21_X1 U16745 ( .B1(n15084), .B2(n15083), .A(n15082), .ZN(n15085) );
  AOI21_X1 U16746 ( .B1(n15102), .B2(n15175), .A(n15085), .ZN(n15172) );
  AOI22_X1 U16747 ( .A1(n15105), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n15086), 
        .B2(n15103), .ZN(n15087) );
  OAI21_X1 U16748 ( .B1(n15107), .B2(n15171), .A(n15087), .ZN(n15088) );
  INV_X1 U16749 ( .A(n15088), .ZN(n15093) );
  OAI211_X1 U16750 ( .C1(n15171), .C2(n15090), .A(n15111), .B(n15089), .ZN(
        n15170) );
  INV_X1 U16751 ( .A(n15170), .ZN(n15091) );
  AOI22_X1 U16752 ( .A1(n15175), .A2(n15114), .B1(n15113), .B2(n15091), .ZN(
        n15092) );
  OAI211_X1 U16753 ( .C1(n15118), .C2(n15172), .A(n15093), .B(n15092), .ZN(
        P1_U3286) );
  XNOR2_X1 U16754 ( .A(n15095), .B(n15094), .ZN(n15160) );
  INV_X1 U16755 ( .A(n15157), .ZN(n15101) );
  XNOR2_X1 U16756 ( .A(n15096), .B(n15097), .ZN(n15099) );
  NAND2_X1 U16757 ( .A1(n15099), .A2(n15098), .ZN(n15158) );
  INV_X1 U16758 ( .A(n15158), .ZN(n15100) );
  AOI211_X1 U16759 ( .C1(n15102), .C2(n15160), .A(n15101), .B(n15100), .ZN(
        n15117) );
  AOI22_X1 U16760 ( .A1(n15105), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n15104), 
        .B2(n15103), .ZN(n15106) );
  OAI21_X1 U16761 ( .B1(n15107), .B2(n6947), .A(n15106), .ZN(n15108) );
  INV_X1 U16762 ( .A(n15108), .ZN(n15116) );
  OAI211_X1 U16763 ( .C1(n6948), .C2(n6947), .A(n15111), .B(n15110), .ZN(
        n15155) );
  INV_X1 U16764 ( .A(n15155), .ZN(n15112) );
  AOI22_X1 U16765 ( .A1(n15160), .A2(n15114), .B1(n15113), .B2(n15112), .ZN(
        n15115) );
  OAI211_X1 U16766 ( .C1(n15118), .C2(n15117), .A(n15116), .B(n15115), .ZN(
        P1_U3288) );
  INV_X1 U16767 ( .A(n15123), .ZN(n15122) );
  NOR2_X1 U16768 ( .A1(n15122), .A2(n15119), .ZN(P1_U3294) );
  AND2_X1 U16769 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15123), .ZN(P1_U3295) );
  AND2_X1 U16770 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15123), .ZN(P1_U3296) );
  AND2_X1 U16771 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15123), .ZN(P1_U3297) );
  AND2_X1 U16772 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15123), .ZN(P1_U3298) );
  AND2_X1 U16773 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15123), .ZN(P1_U3299) );
  AND2_X1 U16774 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15123), .ZN(P1_U3300) );
  AND2_X1 U16775 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15123), .ZN(P1_U3301) );
  AND2_X1 U16776 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15123), .ZN(P1_U3302) );
  AND2_X1 U16777 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15123), .ZN(P1_U3303) );
  AND2_X1 U16778 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15123), .ZN(P1_U3304) );
  AND2_X1 U16779 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15123), .ZN(P1_U3305) );
  AND2_X1 U16780 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15123), .ZN(P1_U3306) );
  NOR2_X1 U16781 ( .A1(n15122), .A2(n15120), .ZN(P1_U3307) );
  NOR2_X1 U16782 ( .A1(n15122), .A2(n15121), .ZN(P1_U3308) );
  AND2_X1 U16783 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15123), .ZN(P1_U3309) );
  AND2_X1 U16784 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15123), .ZN(P1_U3310) );
  AND2_X1 U16785 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15123), .ZN(P1_U3311) );
  AND2_X1 U16786 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15123), .ZN(P1_U3312) );
  AND2_X1 U16787 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15123), .ZN(P1_U3313) );
  AND2_X1 U16788 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15123), .ZN(P1_U3314) );
  AND2_X1 U16789 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15123), .ZN(P1_U3315) );
  AND2_X1 U16790 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15123), .ZN(P1_U3316) );
  AND2_X1 U16791 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15123), .ZN(P1_U3317) );
  AND2_X1 U16792 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15123), .ZN(P1_U3318) );
  AND2_X1 U16793 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15123), .ZN(P1_U3319) );
  AND2_X1 U16794 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15123), .ZN(P1_U3320) );
  AND2_X1 U16795 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15123), .ZN(P1_U3321) );
  AND2_X1 U16796 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15123), .ZN(P1_U3322) );
  AND2_X1 U16797 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15123), .ZN(P1_U3323) );
  OAI22_X1 U16798 ( .A1(n15126), .A2(n15125), .B1(n15124), .B2(n15185), .ZN(
        n15129) );
  INV_X1 U16799 ( .A(n15127), .ZN(n15128) );
  AOI211_X1 U16800 ( .C1(n15190), .C2(n15130), .A(n15129), .B(n15128), .ZN(
        n15203) );
  INV_X1 U16801 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15131) );
  AOI22_X1 U16802 ( .A1(n15201), .A2(n15203), .B1(n15131), .B2(n15199), .ZN(
        P1_U3462) );
  NAND2_X1 U16803 ( .A1(n15132), .A2(n15190), .ZN(n15134) );
  OAI211_X1 U16804 ( .C1(n15135), .C2(n15185), .A(n15134), .B(n15133), .ZN(
        n15136) );
  NOR2_X1 U16805 ( .A1(n15137), .A2(n15136), .ZN(n15205) );
  INV_X1 U16806 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U16807 ( .A1(n15201), .A2(n15205), .B1(n15138), .B2(n15199), .ZN(
        P1_U3465) );
  NAND2_X1 U16808 ( .A1(n15139), .A2(n15190), .ZN(n15142) );
  INV_X1 U16809 ( .A(n15140), .ZN(n15141) );
  OAI211_X1 U16810 ( .C1(n6946), .C2(n15185), .A(n15142), .B(n15141), .ZN(
        n15143) );
  NOR2_X1 U16811 ( .A1(n15144), .A2(n15143), .ZN(n15206) );
  AOI22_X1 U16812 ( .A1(n15201), .A2(n15206), .B1(n15145), .B2(n15199), .ZN(
        P1_U3468) );
  INV_X1 U16813 ( .A(n15146), .ZN(n15153) );
  OAI211_X1 U16814 ( .C1(n15149), .C2(n15185), .A(n15148), .B(n15147), .ZN(
        n15152) );
  INV_X1 U16815 ( .A(n15150), .ZN(n15151) );
  AOI211_X1 U16816 ( .C1(n15153), .C2(n15198), .A(n15152), .B(n15151), .ZN(
        n15207) );
  AOI22_X1 U16817 ( .A1(n15201), .A2(n15207), .B1(n8614), .B2(n15199), .ZN(
        P1_U3471) );
  INV_X1 U16818 ( .A(n15154), .ZN(n15156) );
  NAND4_X1 U16819 ( .A1(n15158), .A2(n15157), .A3(n15156), .A4(n15155), .ZN(
        n15159) );
  AOI21_X1 U16820 ( .B1(n15160), .B2(n15198), .A(n15159), .ZN(n15208) );
  INV_X1 U16821 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15161) );
  AOI22_X1 U16822 ( .A1(n15201), .A2(n15208), .B1(n15161), .B2(n15199), .ZN(
        P1_U3474) );
  INV_X1 U16823 ( .A(n15162), .ZN(n15163) );
  OR2_X1 U16824 ( .A1(n15164), .A2(n15163), .ZN(n15165) );
  AOI21_X1 U16825 ( .B1(n15166), .B2(n15190), .A(n15165), .ZN(n15167) );
  AND2_X1 U16826 ( .A1(n15168), .A2(n15167), .ZN(n15209) );
  INV_X1 U16827 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U16828 ( .A1(n15201), .A2(n15209), .B1(n15169), .B2(n15199), .ZN(
        P1_U3477) );
  OAI21_X1 U16829 ( .B1(n15171), .B2(n15185), .A(n15170), .ZN(n15174) );
  INV_X1 U16830 ( .A(n15172), .ZN(n15173) );
  AOI211_X1 U16831 ( .C1(n15190), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        n15210) );
  INV_X1 U16832 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15176) );
  AOI22_X1 U16833 ( .A1(n15201), .A2(n15210), .B1(n15176), .B2(n15199), .ZN(
        P1_U3480) );
  INV_X1 U16834 ( .A(n15177), .ZN(n15179) );
  OAI21_X1 U16835 ( .B1(n15179), .B2(n15185), .A(n15178), .ZN(n15181) );
  AOI211_X1 U16836 ( .C1(n15182), .C2(n15198), .A(n15181), .B(n15180), .ZN(
        n15211) );
  INV_X1 U16837 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15183) );
  AOI22_X1 U16838 ( .A1(n15201), .A2(n15211), .B1(n15183), .B2(n15199), .ZN(
        P1_U3483) );
  OAI21_X1 U16839 ( .B1(n7364), .B2(n15185), .A(n15184), .ZN(n15188) );
  INV_X1 U16840 ( .A(n15186), .ZN(n15187) );
  AOI211_X1 U16841 ( .C1(n15190), .C2(n15189), .A(n15188), .B(n15187), .ZN(
        n15212) );
  INV_X1 U16842 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U16843 ( .A1(n15201), .A2(n15212), .B1(n15191), .B2(n15199), .ZN(
        P1_U3486) );
  OR4_X1 U16844 ( .A1(n15195), .A2(n15194), .A3(n15193), .A4(n15192), .ZN(
        n15196) );
  AOI21_X1 U16845 ( .B1(n15198), .B2(n15197), .A(n15196), .ZN(n15214) );
  INV_X1 U16846 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15200) );
  AOI22_X1 U16847 ( .A1(n15201), .A2(n15214), .B1(n15200), .B2(n15199), .ZN(
        P1_U3489) );
  AOI22_X1 U16848 ( .A1(n15215), .A2(n15203), .B1(n15202), .B2(n15213), .ZN(
        P1_U3529) );
  AOI22_X1 U16849 ( .A1(n15215), .A2(n15205), .B1(n15204), .B2(n15213), .ZN(
        P1_U3530) );
  AOI22_X1 U16850 ( .A1(n15215), .A2(n15206), .B1(n10502), .B2(n15213), .ZN(
        P1_U3531) );
  AOI22_X1 U16851 ( .A1(n15215), .A2(n15207), .B1(n10504), .B2(n15213), .ZN(
        P1_U3532) );
  AOI22_X1 U16852 ( .A1(n15215), .A2(n15208), .B1(n10505), .B2(n15213), .ZN(
        P1_U3533) );
  AOI22_X1 U16853 ( .A1(n15215), .A2(n15209), .B1(n10532), .B2(n15213), .ZN(
        P1_U3534) );
  AOI22_X1 U16854 ( .A1(n15215), .A2(n15210), .B1(n10534), .B2(n15213), .ZN(
        P1_U3535) );
  AOI22_X1 U16855 ( .A1(n15215), .A2(n15211), .B1(n10536), .B2(n15213), .ZN(
        P1_U3536) );
  AOI22_X1 U16856 ( .A1(n15215), .A2(n15212), .B1(n10529), .B2(n15213), .ZN(
        P1_U3537) );
  AOI22_X1 U16857 ( .A1(n15215), .A2(n15214), .B1(n10632), .B2(n15213), .ZN(
        P1_U3538) );
  NOR2_X1 U16858 ( .A1(n15275), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16859 ( .A1(n15275), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15229) );
  OAI21_X1 U16860 ( .B1(n15218), .B2(n15217), .A(n15216), .ZN(n15222) );
  NAND2_X1 U16861 ( .A1(n8517), .A2(n15219), .ZN(n15220) );
  OAI22_X1 U16862 ( .A1(n15271), .A2(n15222), .B1(n15221), .B2(n15220), .ZN(
        n15223) );
  INV_X1 U16863 ( .A(n15223), .ZN(n15228) );
  OAI211_X1 U16864 ( .C1(n15226), .C2(n15225), .A(n15277), .B(n15224), .ZN(
        n15227) );
  NAND3_X1 U16865 ( .A1(n15229), .A2(n15228), .A3(n15227), .ZN(P2_U3215) );
  OAI211_X1 U16866 ( .C1(n15233), .C2(n15232), .A(n15231), .B(n15230), .ZN(
        n15234) );
  INV_X1 U16867 ( .A(n15234), .ZN(n15238) );
  OAI22_X1 U16868 ( .A1(n15236), .A2(n15235), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10676), .ZN(n15237) );
  AOI211_X1 U16869 ( .C1(n15275), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n15238), .B(
        n15237), .ZN(n15243) );
  OAI211_X1 U16870 ( .C1(n15241), .C2(n15240), .A(n15277), .B(n15239), .ZN(
        n15242) );
  NAND2_X1 U16871 ( .A1(n15243), .A2(n15242), .ZN(P2_U3216) );
  NOR2_X1 U16872 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15244), .ZN(n15250) );
  NOR2_X1 U16873 ( .A1(n15246), .A2(n15245), .ZN(n15247) );
  NOR3_X1 U16874 ( .A1(n15271), .A2(n15248), .A3(n15247), .ZN(n15249) );
  AOI211_X1 U16875 ( .C1(n15281), .C2(n15251), .A(n15250), .B(n15249), .ZN(
        n15256) );
  OAI211_X1 U16876 ( .C1(n15254), .C2(n15253), .A(n15277), .B(n15252), .ZN(
        n15255) );
  OAI211_X1 U16877 ( .C1(n15269), .C2(n15599), .A(n15256), .B(n15255), .ZN(
        P2_U3217) );
  NOR2_X1 U16878 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15257), .ZN(n15262) );
  AOI211_X1 U16879 ( .C1(n15260), .C2(n15259), .A(n15258), .B(n15271), .ZN(
        n15261) );
  AOI211_X1 U16880 ( .C1(n15281), .C2(n15263), .A(n15262), .B(n15261), .ZN(
        n15267) );
  OAI211_X1 U16881 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15265), .A(n15277), 
        .B(n15264), .ZN(n15266) );
  OAI211_X1 U16882 ( .C1(n15269), .C2(n15268), .A(n15267), .B(n15266), .ZN(
        P2_U3229) );
  AOI211_X1 U16883 ( .C1(n15273), .C2(n15272), .A(n15271), .B(n15270), .ZN(
        n15274) );
  AOI21_X1 U16884 ( .B1(n15275), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n15274), 
        .ZN(n15285) );
  OAI211_X1 U16885 ( .C1(n15279), .C2(n15278), .A(n15277), .B(n15276), .ZN(
        n15283) );
  NAND2_X1 U16886 ( .A1(n15281), .A2(n15280), .ZN(n15282) );
  NAND4_X1 U16887 ( .A1(n15285), .A2(n15284), .A3(n15283), .A4(n15282), .ZN(
        P2_U3231) );
  INV_X1 U16888 ( .A(n15287), .ZN(n15289) );
  AOI22_X1 U16889 ( .A1(n15290), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n15289), 
        .B2(n15288), .ZN(n15291) );
  OAI21_X1 U16890 ( .B1(n6867), .B2(n15292), .A(n15291), .ZN(n15296) );
  NOR2_X1 U16891 ( .A1(n15294), .A2(n15293), .ZN(n15295) );
  AOI211_X1 U16892 ( .C1(n15298), .C2(n15297), .A(n15296), .B(n15295), .ZN(
        n15299) );
  OAI21_X1 U16893 ( .B1(n15301), .B2(n15300), .A(n15299), .ZN(P2_U3254) );
  AND2_X1 U16894 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15308), .ZN(P2_U3266) );
  NOR2_X1 U16895 ( .A1(n15307), .A2(n15303), .ZN(P2_U3267) );
  AND2_X1 U16896 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15308), .ZN(P2_U3268) );
  AND2_X1 U16897 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15308), .ZN(P2_U3269) );
  AND2_X1 U16898 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15308), .ZN(P2_U3270) );
  AND2_X1 U16899 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15308), .ZN(P2_U3271) );
  AND2_X1 U16900 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15308), .ZN(P2_U3272) );
  AND2_X1 U16901 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15308), .ZN(P2_U3273) );
  AND2_X1 U16902 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15308), .ZN(P2_U3274) );
  AND2_X1 U16903 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15308), .ZN(P2_U3275) );
  AND2_X1 U16904 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15308), .ZN(P2_U3276) );
  NOR2_X1 U16905 ( .A1(n15307), .A2(n15304), .ZN(P2_U3277) );
  AND2_X1 U16906 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15308), .ZN(P2_U3278) );
  AND2_X1 U16907 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15308), .ZN(P2_U3279) );
  AND2_X1 U16908 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15308), .ZN(P2_U3280) );
  NOR2_X1 U16909 ( .A1(n15307), .A2(n15305), .ZN(P2_U3281) );
  AND2_X1 U16910 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15308), .ZN(P2_U3282) );
  NOR2_X1 U16911 ( .A1(n15307), .A2(n15306), .ZN(P2_U3283) );
  AND2_X1 U16912 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15308), .ZN(P2_U3284) );
  AND2_X1 U16913 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15308), .ZN(P2_U3285) );
  AND2_X1 U16914 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15308), .ZN(P2_U3286) );
  AND2_X1 U16915 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15308), .ZN(P2_U3287) );
  AND2_X1 U16916 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15308), .ZN(P2_U3288) );
  AND2_X1 U16917 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15308), .ZN(P2_U3289) );
  AND2_X1 U16918 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15308), .ZN(P2_U3290) );
  AND2_X1 U16919 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15308), .ZN(P2_U3291) );
  AND2_X1 U16920 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15308), .ZN(P2_U3292) );
  AND2_X1 U16921 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15308), .ZN(P2_U3293) );
  AND2_X1 U16922 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15308), .ZN(P2_U3294) );
  AND2_X1 U16923 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15308), .ZN(P2_U3295) );
  INV_X1 U16924 ( .A(n15311), .ZN(n15314) );
  AOI22_X1 U16925 ( .A1(n15314), .A2(n15310), .B1(n15309), .B2(n15311), .ZN(
        P2_U3416) );
  AOI22_X1 U16926 ( .A1(n15314), .A2(n15313), .B1(n15312), .B2(n15311), .ZN(
        P2_U3417) );
  OAI21_X1 U16927 ( .B1(n15316), .B2(n15342), .A(n15315), .ZN(n15318) );
  AOI211_X1 U16928 ( .C1(n9298), .C2(n15319), .A(n15318), .B(n15317), .ZN(
        n15365) );
  INV_X1 U16929 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15320) );
  AOI22_X1 U16930 ( .A1(n15364), .A2(n15365), .B1(n15320), .B2(n15362), .ZN(
        P2_U3433) );
  OAI21_X1 U16931 ( .B1(n8476), .B2(n15342), .A(n15321), .ZN(n15323) );
  AOI211_X1 U16932 ( .C1(n9298), .C2(n15324), .A(n15323), .B(n15322), .ZN(
        n15366) );
  INV_X1 U16933 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15325) );
  AOI22_X1 U16934 ( .A1(n15364), .A2(n15366), .B1(n15325), .B2(n15362), .ZN(
        P2_U3436) );
  INV_X1 U16935 ( .A(n15326), .ZN(n15331) );
  OAI21_X1 U16936 ( .B1(n15328), .B2(n15342), .A(n15327), .ZN(n15330) );
  AOI211_X1 U16937 ( .C1(n9298), .C2(n15331), .A(n15330), .B(n15329), .ZN(
        n15367) );
  INV_X1 U16938 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15332) );
  AOI22_X1 U16939 ( .A1(n15364), .A2(n15367), .B1(n15332), .B2(n15362), .ZN(
        P2_U3439) );
  INV_X1 U16940 ( .A(n15333), .ZN(n15338) );
  OAI211_X1 U16941 ( .C1(n15336), .C2(n15342), .A(n15335), .B(n15334), .ZN(
        n15337) );
  AOI21_X1 U16942 ( .B1(n15338), .B2(n15339), .A(n15337), .ZN(n15368) );
  AOI22_X1 U16943 ( .A1(n15364), .A2(n15368), .B1(n7812), .B2(n15362), .ZN(
        P2_U3442) );
  AND2_X1 U16944 ( .A1(n15340), .A2(n15339), .ZN(n15345) );
  OAI21_X1 U16945 ( .B1(n15343), .B2(n15342), .A(n15341), .ZN(n15344) );
  NOR3_X1 U16946 ( .A1(n15346), .A2(n15345), .A3(n15344), .ZN(n15369) );
  AOI22_X1 U16947 ( .A1(n15364), .A2(n15369), .B1(n7862), .B2(n15362), .ZN(
        P2_U3448) );
  NOR2_X1 U16948 ( .A1(n15347), .A2(n15360), .ZN(n15352) );
  AND2_X1 U16949 ( .A1(n15348), .A2(n15356), .ZN(n15349) );
  OR2_X1 U16950 ( .A1(n15350), .A2(n15349), .ZN(n15351) );
  NOR3_X1 U16951 ( .A1(n15353), .A2(n15352), .A3(n15351), .ZN(n15370) );
  AOI22_X1 U16952 ( .A1(n15364), .A2(n15370), .B1(n7885), .B2(n15362), .ZN(
        P2_U3451) );
  AOI21_X1 U16953 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n15357) );
  OAI211_X1 U16954 ( .C1(n15360), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        n15361) );
  INV_X1 U16955 ( .A(n15361), .ZN(n15372) );
  INV_X1 U16956 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15363) );
  AOI22_X1 U16957 ( .A1(n15364), .A2(n15372), .B1(n15363), .B2(n15362), .ZN(
        P2_U3457) );
  AOI22_X1 U16958 ( .A1(n13815), .A2(n15365), .B1(n10356), .B2(n15371), .ZN(
        P2_U3500) );
  AOI22_X1 U16959 ( .A1(n13815), .A2(n15366), .B1(n10357), .B2(n15371), .ZN(
        P2_U3501) );
  AOI22_X1 U16960 ( .A1(n13815), .A2(n15367), .B1(n7780), .B2(n15371), .ZN(
        P2_U3502) );
  AOI22_X1 U16961 ( .A1(n13815), .A2(n15368), .B1(n7811), .B2(n15371), .ZN(
        P2_U3503) );
  AOI22_X1 U16962 ( .A1(n13815), .A2(n15369), .B1(n10359), .B2(n15371), .ZN(
        P2_U3505) );
  AOI22_X1 U16963 ( .A1(n13815), .A2(n15370), .B1(n10451), .B2(n15371), .ZN(
        P2_U3506) );
  AOI22_X1 U16964 ( .A1(n13815), .A2(n15372), .B1(n10668), .B2(n15371), .ZN(
        P2_U3508) );
  NOR2_X1 U16965 ( .A1(P3_U3897), .A2(n15460), .ZN(P3_U3150) );
  AOI21_X1 U16966 ( .B1(n15374), .B2(n6715), .A(n15373), .ZN(n15387) );
  INV_X1 U16967 ( .A(n15395), .ZN(n15378) );
  AOI21_X1 U16968 ( .B1(n15376), .B2(n15391), .A(n15375), .ZN(n15377) );
  AOI21_X1 U16969 ( .B1(n15378), .B2(n15391), .A(n15377), .ZN(n15379) );
  OAI22_X1 U16970 ( .A1(n15379), .A2(n15456), .B1(n7028), .B2(n15454), .ZN(
        n15380) );
  AOI211_X1 U16971 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n15460), .A(n15381), .B(
        n15380), .ZN(n15386) );
  OAI21_X1 U16972 ( .B1(n15383), .B2(P3_REG1_REG_5__SCAN_IN), .A(n15382), .ZN(
        n15384) );
  NAND2_X1 U16973 ( .A1(n15463), .A2(n15384), .ZN(n15385) );
  OAI211_X1 U16974 ( .C1(n15387), .C2(n15467), .A(n15386), .B(n15385), .ZN(
        P3_U3187) );
  AOI21_X1 U16975 ( .B1(n15390), .B2(n15389), .A(n15388), .ZN(n15407) );
  INV_X1 U16976 ( .A(n15391), .ZN(n15392) );
  NOR2_X1 U16977 ( .A1(n15393), .A2(n15392), .ZN(n15396) );
  INV_X1 U16978 ( .A(n15414), .ZN(n15394) );
  AOI21_X1 U16979 ( .B1(n15396), .B2(n15395), .A(n15394), .ZN(n15398) );
  OAI22_X1 U16980 ( .A1(n15398), .A2(n15456), .B1(n15397), .B2(n15454), .ZN(
        n15399) );
  AOI211_X1 U16981 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n15460), .A(n15400), .B(
        n15399), .ZN(n15406) );
  OAI21_X1 U16982 ( .B1(n15403), .B2(n15402), .A(n15401), .ZN(n15404) );
  NAND2_X1 U16983 ( .A1(n15463), .A2(n15404), .ZN(n15405) );
  OAI211_X1 U16984 ( .C1(n15407), .C2(n15467), .A(n15406), .B(n15405), .ZN(
        P3_U3188) );
  AOI21_X1 U16985 ( .B1(n11303), .B2(n15409), .A(n15408), .ZN(n15425) );
  INV_X1 U16986 ( .A(n15410), .ZN(n15411) );
  NOR2_X1 U16987 ( .A1(n15412), .A2(n15411), .ZN(n15415) );
  INV_X1 U16988 ( .A(n15433), .ZN(n15413) );
  AOI21_X1 U16989 ( .B1(n15415), .B2(n15414), .A(n15413), .ZN(n15417) );
  OAI22_X1 U16990 ( .A1(n15417), .A2(n15456), .B1(n15416), .B2(n15454), .ZN(
        n15418) );
  AOI211_X1 U16991 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n15460), .A(n15419), .B(
        n15418), .ZN(n15424) );
  OAI21_X1 U16992 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n15421), .A(n15420), .ZN(
        n15422) );
  NAND2_X1 U16993 ( .A1(n15422), .A2(n15463), .ZN(n15423) );
  OAI211_X1 U16994 ( .C1(n15425), .C2(n15467), .A(n15424), .B(n15423), .ZN(
        P3_U3189) );
  AOI21_X1 U16995 ( .B1(n15428), .B2(n15427), .A(n15426), .ZN(n15445) );
  INV_X1 U16996 ( .A(n15429), .ZN(n15430) );
  NOR2_X1 U16997 ( .A1(n15431), .A2(n15430), .ZN(n15434) );
  INV_X1 U16998 ( .A(n15452), .ZN(n15432) );
  AOI21_X1 U16999 ( .B1(n15434), .B2(n15433), .A(n15432), .ZN(n15436) );
  OAI22_X1 U17000 ( .A1(n15436), .A2(n15456), .B1(n15435), .B2(n15454), .ZN(
        n15437) );
  AOI211_X1 U17001 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n15460), .A(n15438), .B(
        n15437), .ZN(n15444) );
  OAI21_X1 U17002 ( .B1(n15441), .B2(n15440), .A(n15439), .ZN(n15442) );
  NAND2_X1 U17003 ( .A1(n15442), .A2(n15463), .ZN(n15443) );
  OAI211_X1 U17004 ( .C1(n15445), .C2(n15467), .A(n15444), .B(n15443), .ZN(
        P3_U3190) );
  AOI21_X1 U17005 ( .B1(n11851), .B2(n15447), .A(n15446), .ZN(n15468) );
  INV_X1 U17006 ( .A(n15448), .ZN(n15449) );
  NOR2_X1 U17007 ( .A1(n15450), .A2(n15449), .ZN(n15453) );
  AOI21_X1 U17008 ( .B1(n15453), .B2(n15452), .A(n15451), .ZN(n15457) );
  OAI22_X1 U17009 ( .A1(n15457), .A2(n15456), .B1(n15455), .B2(n15454), .ZN(
        n15458) );
  AOI211_X1 U17010 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15460), .A(n15459), .B(
        n15458), .ZN(n15466) );
  OAI21_X1 U17011 ( .B1(n15462), .B2(P3_REG1_REG_9__SCAN_IN), .A(n15461), .ZN(
        n15464) );
  NAND2_X1 U17012 ( .A1(n15464), .A2(n15463), .ZN(n15465) );
  OAI211_X1 U17013 ( .C1(n15468), .C2(n15467), .A(n15466), .B(n15465), .ZN(
        P3_U3191) );
  XNOR2_X1 U17014 ( .A(n15469), .B(n15470), .ZN(n15477) );
  INV_X1 U17015 ( .A(n15477), .ZN(n15552) );
  XNOR2_X1 U17016 ( .A(n15471), .B(n6673), .ZN(n15475) );
  OAI22_X1 U17017 ( .A1(n15473), .A2(n15509), .B1(n15472), .B2(n15507), .ZN(
        n15474) );
  AOI21_X1 U17018 ( .B1(n15475), .B2(n15511), .A(n15474), .ZN(n15476) );
  OAI21_X1 U17019 ( .B1(n15477), .B2(n15514), .A(n15476), .ZN(n15550) );
  AOI21_X1 U17020 ( .B1(n15498), .B2(n15552), .A(n15550), .ZN(n15485) );
  NOR2_X1 U17021 ( .A1(n15478), .A2(n15545), .ZN(n15551) );
  INV_X1 U17022 ( .A(n15551), .ZN(n15481) );
  OAI22_X1 U17023 ( .A1(n15482), .A2(n15481), .B1(n15480), .B2(n15479), .ZN(
        n15483) );
  INV_X1 U17024 ( .A(n15483), .ZN(n15484) );
  OAI221_X1 U17025 ( .B1(n13166), .B2(n15485), .C1(n15501), .C2(n11303), .A(
        n15484), .ZN(P3_U3226) );
  OAI21_X1 U17026 ( .B1(n15487), .B2(n12627), .A(n15486), .ZN(n15527) );
  OAI22_X1 U17027 ( .A1(n6848), .A2(n15509), .B1(n15488), .B2(n15507), .ZN(
        n15494) );
  NAND3_X1 U17028 ( .A1(n15505), .A2(n12627), .A3(n15489), .ZN(n15491) );
  AOI21_X1 U17029 ( .B1(n15492), .B2(n15491), .A(n15490), .ZN(n15493) );
  AOI211_X1 U17030 ( .C1(n15495), .C2(n15527), .A(n15494), .B(n15493), .ZN(
        n15496) );
  INV_X1 U17031 ( .A(n15496), .ZN(n15525) );
  NOR2_X1 U17032 ( .A1(n15497), .A2(n15545), .ZN(n15526) );
  AOI22_X1 U17033 ( .A1(n15527), .A2(n15498), .B1(n15526), .B2(n15515), .ZN(
        n15499) );
  INV_X1 U17034 ( .A(n15499), .ZN(n15500) );
  AOI211_X1 U17035 ( .C1(n15517), .C2(P3_REG3_REG_2__SCAN_IN), .A(n15525), .B(
        n15500), .ZN(n15502) );
  AOI22_X1 U17036 ( .A1(n13166), .A2(n9549), .B1(n15502), .B2(n15501), .ZN(
        P3_U3231) );
  NOR2_X1 U17037 ( .A1(n9568), .A2(n15545), .ZN(n15522) );
  XNOR2_X1 U17038 ( .A(n11008), .B(n15504), .ZN(n15516) );
  OAI21_X1 U17039 ( .B1(n15506), .B2(n11008), .A(n15505), .ZN(n15512) );
  OAI22_X1 U17040 ( .A1(n9978), .A2(n15509), .B1(n15508), .B2(n15507), .ZN(
        n15510) );
  AOI21_X1 U17041 ( .B1(n15512), .B2(n15511), .A(n15510), .ZN(n15513) );
  OAI21_X1 U17042 ( .B1(n15516), .B2(n15514), .A(n15513), .ZN(n15521) );
  AOI21_X1 U17043 ( .B1(n15522), .B2(n15515), .A(n15521), .ZN(n15520) );
  INV_X1 U17044 ( .A(n15516), .ZN(n15523) );
  AOI22_X1 U17045 ( .A1(n15523), .A2(n15518), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15517), .ZN(n15519) );
  OAI221_X1 U17046 ( .B1(n13166), .B2(n15520), .C1(n15501), .C2(n10826), .A(
        n15519), .ZN(P3_U3232) );
  AOI211_X1 U17047 ( .C1(n15566), .C2(n15523), .A(n15522), .B(n15521), .ZN(
        n15571) );
  INV_X1 U17048 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15524) );
  AOI22_X1 U17049 ( .A1(n15570), .A2(n15571), .B1(n15524), .B2(n15568), .ZN(
        P3_U3393) );
  AOI211_X1 U17050 ( .C1(n15566), .C2(n15527), .A(n15526), .B(n15525), .ZN(
        n15573) );
  INV_X1 U17051 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15528) );
  AOI22_X1 U17052 ( .A1(n15570), .A2(n15573), .B1(n15528), .B2(n15568), .ZN(
        P3_U3396) );
  INV_X1 U17053 ( .A(n15529), .ZN(n15530) );
  AOI211_X1 U17054 ( .C1(n15532), .C2(n15566), .A(n15531), .B(n15530), .ZN(
        n15575) );
  INV_X1 U17055 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15533) );
  AOI22_X1 U17056 ( .A1(n15570), .A2(n15575), .B1(n15533), .B2(n15568), .ZN(
        P3_U3399) );
  NOR2_X1 U17057 ( .A1(n15534), .A2(n15545), .ZN(n15536) );
  AOI211_X1 U17058 ( .C1(n15566), .C2(n15537), .A(n15536), .B(n15535), .ZN(
        n15576) );
  INV_X1 U17059 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15538) );
  AOI22_X1 U17060 ( .A1(n15570), .A2(n15576), .B1(n15538), .B2(n15568), .ZN(
        P3_U3402) );
  INV_X1 U17061 ( .A(n15539), .ZN(n15540) );
  AOI211_X1 U17062 ( .C1(n15542), .C2(n15566), .A(n15541), .B(n15540), .ZN(
        n15578) );
  INV_X1 U17063 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15543) );
  AOI22_X1 U17064 ( .A1(n15570), .A2(n15578), .B1(n15543), .B2(n15568), .ZN(
        P3_U3405) );
  INV_X1 U17065 ( .A(n15544), .ZN(n15549) );
  NOR2_X1 U17066 ( .A1(n15546), .A2(n15545), .ZN(n15548) );
  AOI211_X1 U17067 ( .C1(n15549), .C2(n15566), .A(n15548), .B(n15547), .ZN(
        n15579) );
  AOI22_X1 U17068 ( .A1(n15570), .A2(n15579), .B1(n9628), .B2(n15568), .ZN(
        P3_U3408) );
  AOI211_X1 U17069 ( .C1(n15552), .C2(n15566), .A(n15551), .B(n15550), .ZN(
        n15580) );
  INV_X1 U17070 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15553) );
  AOI22_X1 U17071 ( .A1(n15570), .A2(n15580), .B1(n15553), .B2(n15568), .ZN(
        P3_U3411) );
  AOI21_X1 U17072 ( .B1(n15555), .B2(n15566), .A(n15554), .ZN(n15556) );
  INV_X1 U17073 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15558) );
  AOI22_X1 U17074 ( .A1(n15570), .A2(n15581), .B1(n15558), .B2(n15568), .ZN(
        P3_U3414) );
  AOI21_X1 U17075 ( .B1(n15560), .B2(n15566), .A(n15559), .ZN(n15561) );
  AND2_X1 U17076 ( .A1(n15562), .A2(n15561), .ZN(n15582) );
  INV_X1 U17077 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U17078 ( .A1(n15570), .A2(n15582), .B1(n15563), .B2(n15568), .ZN(
        P3_U3417) );
  AOI211_X1 U17079 ( .C1(n15567), .C2(n15566), .A(n15565), .B(n15564), .ZN(
        n15584) );
  INV_X1 U17080 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15569) );
  AOI22_X1 U17081 ( .A1(n15570), .A2(n15584), .B1(n15569), .B2(n15568), .ZN(
        P3_U3420) );
  AOI22_X1 U17082 ( .A1(n15585), .A2(n15571), .B1(n10898), .B2(n15583), .ZN(
        P3_U3460) );
  INV_X1 U17083 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U17084 ( .A1(n15585), .A2(n15573), .B1(n15572), .B2(n15583), .ZN(
        P3_U3461) );
  INV_X1 U17085 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U17086 ( .A1(n15585), .A2(n15575), .B1(n15574), .B2(n15583), .ZN(
        P3_U3462) );
  AOI22_X1 U17087 ( .A1(n15585), .A2(n15576), .B1(n9598), .B2(n15583), .ZN(
        P3_U3463) );
  AOI22_X1 U17088 ( .A1(n15585), .A2(n15578), .B1(n15577), .B2(n15583), .ZN(
        P3_U3464) );
  AOI22_X1 U17089 ( .A1(n15585), .A2(n15579), .B1(n11295), .B2(n15583), .ZN(
        P3_U3465) );
  AOI22_X1 U17090 ( .A1(n15585), .A2(n15580), .B1(n11302), .B2(n15583), .ZN(
        P3_U3466) );
  AOI22_X1 U17091 ( .A1(n15585), .A2(n15581), .B1(n11309), .B2(n15583), .ZN(
        P3_U3467) );
  AOI22_X1 U17092 ( .A1(n15585), .A2(n15582), .B1(n11316), .B2(n15583), .ZN(
        P3_U3468) );
  AOI22_X1 U17093 ( .A1(n15585), .A2(n15584), .B1(n11322), .B2(n15583), .ZN(
        P3_U3469) );
  AOI21_X1 U17094 ( .B1(n15588), .B2(n15587), .A(n15586), .ZN(SUB_1596_U59) );
  OAI21_X1 U17095 ( .B1(n15591), .B2(n15590), .A(n15589), .ZN(SUB_1596_U58) );
  XOR2_X1 U17096 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15592), .Z(SUB_1596_U53) );
  AOI21_X1 U17097 ( .B1(n15595), .B2(n15594), .A(n15593), .ZN(SUB_1596_U56) );
  AOI21_X1 U17098 ( .B1(n15598), .B2(n15597), .A(n15596), .ZN(n15600) );
  XNOR2_X1 U17099 ( .A(n15600), .B(n15599), .ZN(SUB_1596_U60) );
  AOI21_X1 U17100 ( .B1(n15603), .B2(n15602), .A(n15601), .ZN(SUB_1596_U5) );
  AND2_X1 U7487 ( .A1(n8579), .A2(n8527), .ZN(n8620) );
  XNOR2_X1 U9656 ( .A(n7688), .B(n8497), .ZN(n9299) );
  BUF_X2 U7394 ( .A(n7990), .Z(n6690) );
  AND2_X1 U7401 ( .A1(n12626), .A2(n11383), .ZN(n9596) );
  OAI21_X1 U7432 ( .B1(n12518), .B2(n7249), .A(n7246), .ZN(n12482) );
  CLKBUF_X1 U7448 ( .A(n9569), .Z(n6689) );
  XNOR2_X1 U7457 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9554) );
  CLKBUF_X1 U7463 ( .A(n7929), .Z(n8412) );
  CLKBUF_X1 U7474 ( .A(n7810), .Z(n6671) );
  NAND2_X1 U7480 ( .A1(n8384), .A2(n8383), .ZN(n13511) );
  CLKBUF_X1 U7500 ( .A(n7727), .Z(n7752) );
  NAND2_X1 U7508 ( .A1(n14389), .A2(n15026), .ZN(n8848) );
  CLKBUF_X1 U7516 ( .A(n14139), .Z(n6854) );
  NAND2_X1 U7521 ( .A1(n8545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8546) );
  NOR2_X2 U7549 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8579) );
  CLKBUF_X1 U7551 ( .A(n9867), .Z(n6683) );
  OR2_X1 U7552 ( .A1(n7334), .A2(n9720), .ZN(n9456) );
  CLKBUF_X2 U7557 ( .A(n8431), .Z(n6672) );
  CLKBUF_X1 U7576 ( .A(n9162), .Z(n14376) );
  CLKBUF_X1 U7585 ( .A(n7708), .Z(n11719) );
  XNOR2_X1 U7590 ( .A(n9407), .B(n9406), .ZN(n14786) );
  AND3_X1 U7603 ( .A1(n9560), .A2(n9558), .A3(n9561), .ZN(n15607) );
endmodule

