

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225;

  OR2_X1 U4764 ( .A1(n7181), .A2(n4630), .ZN(n7194) );
  CLKBUF_X2 U4765 ( .A(n6975), .Z(n7900) );
  CLKBUF_X2 U4766 ( .A(n5729), .Z(n5915) );
  NAND2_X1 U4767 ( .A1(n4631), .A2(n4630), .ZN(n7200) );
  CLKBUF_X1 U4768 ( .A(n6879), .Z(n7986) );
  INV_X1 U4769 ( .A(n8435), .ZN(n4954) );
  NAND2_X1 U4771 ( .A1(n4441), .A2(n4440), .ZN(n9081) );
  INV_X1 U4772 ( .A(n5247), .ZN(n5729) );
  AND2_X1 U4773 ( .A1(n6281), .A2(n6280), .ZN(n6533) );
  NAND2_X1 U4774 ( .A1(n7678), .A2(n6454), .ZN(n6519) );
  NAND2_X1 U4775 ( .A1(n7678), .A2(n6455), .ZN(n9049) );
  NAND2_X2 U4776 ( .A1(n7607), .A2(n8794), .ZN(n5247) );
  AND4_X1 U4777 ( .A1(n10051), .A2(n5141), .A3(n5150), .A4(n4956), .ZN(n4977)
         );
  CLKBUF_X2 U4778 ( .A(n5218), .Z(n6454) );
  INV_X4 U4779 ( .A(n9589), .ZN(n9566) );
  OR2_X1 U4780 ( .A1(n9065), .A2(n9039), .ZN(n9248) );
  NAND2_X1 U4781 ( .A1(n6960), .A2(n5054), .ZN(n7473) );
  INV_X1 U4782 ( .A(n9974), .ZN(n4630) );
  NAND2_X1 U4783 ( .A1(n5288), .A2(n5287), .ZN(n7193) );
  AND2_X1 U4784 ( .A1(n4494), .A2(n8959), .ZN(n8956) );
  INV_X1 U4785 ( .A(n7875), .ZN(n6975) );
  INV_X1 U4786 ( .A(n9227), .ZN(n9057) );
  AND2_X1 U4787 ( .A1(n4936), .A2(n4937), .ZN(n7977) );
  NAND2_X1 U4788 ( .A1(n4750), .A2(n4748), .ZN(n4843) );
  INV_X1 U4789 ( .A(n8505), .ZN(n8086) );
  INV_X1 U4790 ( .A(n5269), .ZN(n6715) );
  NAND2_X1 U4791 ( .A1(n6053), .A2(n6038), .ZN(n8488) );
  NOR2_X1 U4792 ( .A1(n8976), .A2(n5084), .ZN(n5086) );
  CLKBUF_X3 U4793 ( .A(n6975), .Z(n7892) );
  INV_X1 U4794 ( .A(n9224), .ZN(n9259) );
  OR2_X1 U4795 ( .A1(n9612), .A2(n9390), .ZN(n9249) );
  XNOR2_X1 U4796 ( .A(n5177), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5181) );
  XNOR2_X1 U4797 ( .A(n5147), .B(n5141), .ZN(n7278) );
  OR2_X1 U4798 ( .A1(n9271), .A2(n9270), .ZN(n4666) );
  INV_X2 U4800 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5141) );
  XNOR2_X1 U4802 ( .A(n6307), .B(n6306), .ZN(n6320) );
  XNOR2_X2 U4803 ( .A(n6210), .B(n6209), .ZN(n6213) );
  AOI21_X2 U4804 ( .B1(n5067), .B2(n4718), .A(n4343), .ZN(n4717) );
  XNOR2_X2 U4805 ( .A(n4843), .B(n4960), .ZN(n8126) );
  OAI21_X2 U4806 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10010), .ZN(n10212) );
  OR2_X1 U4807 ( .A1(n8888), .A2(n8982), .ZN(n4384) );
  AOI21_X2 U4808 ( .B1(n8286), .B2(n8285), .A(n8284), .ZN(n8297) );
  OAI21_X2 U4809 ( .B1(n8248), .B2(n8263), .A(n6653), .ZN(n8286) );
  OAI211_X2 U4810 ( .C1(n5217), .C2(n6501), .A(n5174), .B(n5173), .ZN(n9915)
         );
  BUF_X4 U4811 ( .A(n5463), .Z(n4260) );
  INV_X1 U4812 ( .A(n5217), .ZN(n5463) );
  NAND2_X4 U4813 ( .A1(n6356), .A2(n6482), .ZN(n7875) );
  NOR2_X2 U4814 ( .A1(n8488), .A2(n5051), .ZN(n5050) );
  AND2_X1 U4815 ( .A1(n7806), .A2(n7805), .ZN(n8962) );
  NOR2_X1 U4816 ( .A1(n4482), .A2(n7732), .ZN(n4481) );
  NAND2_X1 U4817 ( .A1(n5693), .A2(n5692), .ZN(n8691) );
  INV_X1 U4818 ( .A(n9573), .ZN(n8987) );
  INV_X1 U4819 ( .A(n4450), .ZN(n9190) );
  NAND2_X1 U4820 ( .A1(n5313), .A2(n5312), .ZN(n7378) );
  INV_X2 U4821 ( .A(n7898), .ZN(n4732) );
  INV_X2 U4822 ( .A(n7890), .ZN(n7763) );
  NAND2_X1 U4823 ( .A1(n5986), .A2(n5990), .ZN(n7058) );
  INV_X2 U4824 ( .A(n6715), .ZN(n5322) );
  NAND2_X2 U4825 ( .A1(n6482), .A2(n6463), .ZN(n6524) );
  NAND2_X4 U4826 ( .A1(n6464), .A2(n6463), .ZN(n7890) );
  NAND4_X1 U4827 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n9281)
         );
  INV_X2 U4828 ( .A(n4259), .ZN(n9261) );
  INV_X2 U4829 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5532) );
  AOI211_X1 U4830 ( .C1(n9607), .C2(n9581), .A(n9401), .B(n9400), .ZN(n9402)
         );
  OR2_X1 U4831 ( .A1(n8673), .A2(n8651), .ZN(n4647) );
  AND2_X1 U4832 ( .A1(n8401), .A2(n8400), .ZN(n8673) );
  AOI21_X1 U4833 ( .B1(n9393), .B2(n9577), .A(n9392), .ZN(n9609) );
  AOI21_X1 U4834 ( .B1(n9415), .B2(n9416), .A(n9414), .ZN(n9614) );
  NAND2_X1 U4835 ( .A1(n4494), .A2(n7844), .ZN(n4729) );
  OR2_X1 U4836 ( .A1(n8382), .A2(n5030), .ZN(n8383) );
  AOI21_X1 U4837 ( .B1(n4680), .B2(n9577), .A(n4677), .ZN(n9619) );
  NAND2_X1 U4838 ( .A1(n8458), .A2(n8464), .ZN(n8457) );
  AOI21_X1 U4839 ( .B1(n8671), .B2(n8629), .A(n8402), .ZN(n4646) );
  NAND2_X1 U4840 ( .A1(n4753), .A2(n4755), .ZN(n8157) );
  OAI21_X1 U4841 ( .B1(n8823), .B2(n5068), .A(n4481), .ZN(n7913) );
  OR2_X1 U4842 ( .A1(n8072), .A2(n4758), .ZN(n4753) );
  NAND2_X1 U4843 ( .A1(n7912), .A2(n7911), .ZN(n7916) );
  NAND2_X1 U4844 ( .A1(n5902), .A2(n5901), .ZN(n8666) );
  NAND2_X1 U4845 ( .A1(n9606), .A2(n9413), .ZN(n9062) );
  NAND2_X1 U4846 ( .A1(n8074), .A2(n8073), .ZN(n8072) );
  OAI21_X1 U4847 ( .B1(n8117), .B2(n8116), .A(n5568), .ZN(n8175) );
  XNOR2_X1 U4848 ( .A(n5895), .B(n5894), .ZN(n9736) );
  NAND2_X1 U4849 ( .A1(n5726), .A2(n5725), .ZN(n8688) );
  AND2_X1 U4850 ( .A1(n7874), .A2(n7873), .ZN(n9390) );
  AND2_X1 U4851 ( .A1(n7994), .A2(n7883), .ZN(n9395) );
  NAND2_X1 U4852 ( .A1(n7810), .A2(n7809), .ZN(n9628) );
  OR2_X1 U4853 ( .A1(n7882), .A2(n7881), .ZN(n7994) );
  NAND2_X1 U4854 ( .A1(n4399), .A2(n4971), .ZN(n4968) );
  NAND2_X1 U4855 ( .A1(n7824), .A2(n7823), .ZN(n9631) );
  NAND2_X1 U4856 ( .A1(n5763), .A2(n5762), .ZN(n8206) );
  INV_X1 U4857 ( .A(n5044), .ZN(n5043) );
  NAND2_X1 U4858 ( .A1(n4588), .A2(n4587), .ZN(n5770) );
  AND2_X1 U4859 ( .A1(n4961), .A2(n4775), .ZN(n4774) );
  NAND2_X1 U4860 ( .A1(n5663), .A2(n5662), .ZN(n8703) );
  OAI21_X1 U4861 ( .B1(n4766), .B2(n4398), .A(n4396), .ZN(n7335) );
  NAND2_X1 U4862 ( .A1(n8638), .A2(n4311), .ZN(n8620) );
  NAND2_X1 U4863 ( .A1(n5886), .A2(n5055), .ZN(n8638) );
  NAND2_X1 U4864 ( .A1(n7736), .A2(n7735), .ZN(n9651) );
  AND2_X1 U4865 ( .A1(n4969), .A2(n4967), .ZN(n4966) );
  NAND2_X1 U4866 ( .A1(n7429), .A2(n6014), .ZN(n5886) );
  OR2_X1 U4867 ( .A1(n8608), .A2(n8110), .ZN(n6032) );
  AOI21_X1 U4868 ( .B1(n4971), .B2(n4970), .A(n4308), .ZN(n4969) );
  AND2_X1 U4869 ( .A1(n7668), .A2(n7667), .ZN(n9559) );
  NAND2_X1 U4870 ( .A1(n4444), .A2(n4442), .ZN(n9866) );
  AND2_X1 U4871 ( .A1(n7726), .A2(n7725), .ZN(n8905) );
  XNOR2_X1 U4872 ( .A(n4601), .B(n4600), .ZN(n7213) );
  NAND2_X1 U4873 ( .A1(n5883), .A2(n5884), .ZN(n6960) );
  NAND2_X1 U4874 ( .A1(n5664), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5706) );
  OR2_X1 U4875 ( .A1(n5402), .A2(n5401), .ZN(n4973) );
  NAND2_X1 U4876 ( .A1(n5441), .A2(n5440), .ZN(n8002) );
  AND2_X1 U4877 ( .A1(n6009), .A2(n6004), .ZN(n7499) );
  OR2_X1 U4878 ( .A1(n7455), .A2(n7615), .ZN(n7525) );
  NAND2_X1 U4879 ( .A1(n7628), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U4880 ( .A1(n5393), .A2(n5392), .ZN(n8759) );
  NAND2_X1 U4881 ( .A1(n7284), .A2(n7283), .ZN(n9694) );
  XNOR2_X1 U4882 ( .A(n4388), .B(n5462), .ZN(n7511) );
  NAND2_X1 U4883 ( .A1(n4577), .A2(n5481), .ZN(n5500) );
  NAND2_X1 U4884 ( .A1(n7156), .A2(n7155), .ZN(n9699) );
  XNOR2_X1 U4885 ( .A(n5426), .B(n5424), .ZN(n7285) );
  OR2_X1 U4886 ( .A1(n7378), .A2(n7206), .ZN(n5997) );
  AND2_X1 U4887 ( .A1(n5268), .A2(n5267), .ZN(n9974) );
  AND3_X1 U4888 ( .A1(n5246), .A2(n5245), .A3(n5244), .ZN(n9965) );
  AND2_X1 U4889 ( .A1(n5350), .A2(n4348), .ZN(n5885) );
  OR2_X1 U4890 ( .A1(n9909), .A2(n7054), .ZN(n5986) );
  INV_X1 U4891 ( .A(n8214), .ZN(n4631) );
  INV_X2 U4892 ( .A(n5236), .ZN(n5802) );
  AND3_X1 U4893 ( .A1(n6739), .A2(n6738), .A3(n6737), .ZN(n6985) );
  NAND2_X1 U4894 ( .A1(n5264), .A2(n4548), .ZN(n4547) );
  AND2_X2 U4895 ( .A1(n6200), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND4_X1 U4896 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n8214)
         );
  AND4_X1 U4897 ( .A1(n6883), .A2(n6882), .A3(n6881), .A4(n6880), .ZN(n9080)
         );
  NAND4_X2 U4898 ( .A1(n6332), .A2(n6331), .A3(n6330), .A4(n6329), .ZN(n9285)
         );
  AND4_X1 U4899 ( .A1(n6285), .A2(n6282), .A3(n6283), .A4(n6284), .ZN(n6360)
         );
  NAND2_X1 U4900 ( .A1(n9259), .A2(n7276), .ZN(n6463) );
  NAND4_X1 U4901 ( .A1(n6538), .A2(n6537), .A3(n6536), .A4(n6535), .ZN(n9282)
         );
  AND3_X2 U4903 ( .A1(n6456), .A2(n6458), .A3(n6457), .ZN(n9821) );
  INV_X1 U4904 ( .A(n9915), .ZN(n9948) );
  INV_X1 U4905 ( .A(n9049), .ZN(n7734) );
  CLKBUF_X1 U4906 ( .A(n5909), .Z(n5927) );
  BUF_X4 U4907 ( .A(n6533), .Z(n4264) );
  NAND2_X1 U4908 ( .A1(n4501), .A2(n6152), .ZN(n6482) );
  NAND2_X1 U4909 ( .A1(n6119), .A2(n6118), .ZN(n9224) );
  CLKBUF_X3 U4910 ( .A(n5225), .Z(n5909) );
  CLKBUF_X1 U4911 ( .A(n5140), .Z(n6554) );
  NAND2_X1 U4912 ( .A1(n6455), .A2(n6401), .ZN(n5217) );
  OAI211_X1 U4913 ( .C1(n6104), .C2(n6108), .A(n6103), .B(n6102), .ZN(n7606)
         );
  XNOR2_X1 U4914 ( .A(n5144), .B(n5143), .ZN(n7554) );
  INV_X1 U4915 ( .A(n5180), .ZN(n8794) );
  XNOR2_X1 U4916 ( .A(n5283), .B(SI_5_), .ZN(n5280) );
  NAND2_X1 U4917 ( .A1(n6108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6116) );
  INV_X1 U4918 ( .A(n5181), .ZN(n7607) );
  NAND2_X1 U4919 ( .A1(n4634), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U4920 ( .A1(n5155), .A2(n5175), .ZN(n6619) );
  XNOR2_X1 U4921 ( .A(n5331), .B(SI_7_), .ZN(n5328) );
  NAND2_X2 U4922 ( .A1(n6455), .A2(P2_U3152), .ZN(n8799) );
  INV_X2 U4923 ( .A(n9735), .ZN(n4261) );
  NAND2_X1 U4924 ( .A1(n5072), .A2(n5116), .ZN(n6108) );
  NAND2_X2 U4925 ( .A1(n6455), .A2(P1_U3084), .ZN(n9743) );
  NAND2_X1 U4926 ( .A1(n4840), .A2(n4838), .ZN(n5155) );
  NAND2_X1 U4927 ( .A1(n8790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5177) );
  INV_X1 U4928 ( .A(n5075), .ZN(n5072) );
  AND2_X1 U4929 ( .A1(n5172), .A2(n5226), .ZN(n6557) );
  NOR2_X1 U4930 ( .A1(n4507), .A2(n4504), .ZN(n5145) );
  CLKBUF_X1 U4931 ( .A(n6165), .Z(n6301) );
  BUF_X4 U4932 ( .A(n5218), .Z(n5504) );
  NAND2_X2 U4933 ( .A1(n5002), .A2(n5000), .ZN(n5218) );
  AND2_X1 U4934 ( .A1(n4271), .A2(n10051), .ZN(n4505) );
  AND2_X2 U4935 ( .A1(n4747), .A2(n4746), .ZN(n5117) );
  NAND2_X1 U4936 ( .A1(n5193), .A2(n5192), .ZN(n6417) );
  AND4_X1 U4937 ( .A1(n4977), .A2(n4839), .A3(n5136), .A4(n5266), .ZN(n4976)
         );
  AND4_X1 U4938 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n10084), .ZN(n4265)
         );
  AND2_X1 U4939 ( .A1(n6096), .A2(n6095), .ZN(n4746) );
  AND4_X1 U4940 ( .A1(n6303), .A2(n6299), .A3(n6094), .A4(n10076), .ZN(n4747)
         );
  AND3_X1 U4941 ( .A1(n5090), .A2(n5089), .A3(n6090), .ZN(n6093) );
  AND2_X1 U4942 ( .A1(n6092), .A2(n6091), .ZN(n6133) );
  NAND3_X1 U4943 ( .A1(n5001), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5000) );
  NAND3_X1 U4944 ( .A1(n5005), .A2(n5004), .A3(n5003), .ZN(n5002) );
  NOR2_X1 U4945 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6091) );
  NOR2_X1 U4946 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6092) );
  NOR2_X1 U4947 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6095) );
  NOR2_X1 U4948 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n6094) );
  INV_X4 U4949 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4950 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10084) );
  NOR2_X1 U4951 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5090) );
  INV_X1 U4952 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5004) );
  NOR2_X1 U4953 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5089) );
  INV_X1 U4954 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5003) );
  INV_X1 U4955 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5001) );
  NOR2_X2 U4956 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5167) );
  INV_X1 U4957 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6207) );
  NOR2_X1 U4958 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5135) );
  NOR2_X1 U4959 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5130) );
  NOR2_X4 U4960 ( .A1(n7171), .A2(n9699), .ZN(n7619) );
  AOI21_X2 U4961 ( .B1(n7165), .B2(n4274), .A(n4332), .ZN(n7166) );
  NOR2_X2 U4962 ( .A1(n6593), .A2(n6859), .ZN(n6902) );
  NAND2_X2 U4963 ( .A1(n5672), .A2(n5671), .ZN(n8505) );
  AND2_X4 U4964 ( .A1(n7607), .A2(n5180), .ZN(n5314) );
  INV_X1 U4965 ( .A(n6524), .ZN(n4262) );
  NOR2_X2 U4966 ( .A1(n7194), .A2(n7193), .ZN(n6949) );
  NOR2_X2 U4967 ( .A1(n9518), .A2(n4565), .ZN(n4564) );
  AOI211_X2 U4968 ( .C1(n9834), .C2(n9628), .A(n9627), .B(n9626), .ZN(n9629)
         );
  NOR2_X2 U4969 ( .A1(n9636), .A2(n9484), .ZN(n9464) );
  NAND2_X2 U4970 ( .A1(n9502), .A2(n8879), .ZN(n9484) );
  NAND4_X2 U4971 ( .A1(n6518), .A2(n6517), .A3(n6516), .A4(n6515), .ZN(n9283)
         );
  CLKBUF_X1 U4972 ( .A(n6533), .Z(n4263) );
  AND2_X4 U4973 ( .A1(n6281), .A2(n9732), .ZN(n6743) );
  INV_X1 U4974 ( .A(n6213), .ZN(n6281) );
  OR2_X1 U4975 ( .A1(n9628), .A2(n9448), .ZN(n7970) );
  AND2_X1 U4976 ( .A1(n9929), .A2(n5842), .ZN(n6543) );
  NAND2_X1 U4977 ( .A1(n4572), .A2(n4287), .ZN(n4567) );
  AOI21_X1 U4978 ( .B1(n4855), .B2(n4273), .A(n4341), .ZN(n4854) );
  OR2_X1 U4979 ( .A1(n8666), .A2(n6068), .ZN(n5033) );
  OR2_X1 U4980 ( .A1(n9631), .A2(n7957), .ZN(n9157) );
  INV_X1 U4981 ( .A(n7949), .ZN(n4421) );
  NAND2_X1 U4982 ( .A1(n7107), .A2(n9187), .ZN(n4444) );
  AND2_X1 U4983 ( .A1(n5640), .A2(n5623), .ZN(n5638) );
  INV_X1 U4984 ( .A(n5794), .ZN(n5782) );
  NAND2_X1 U4985 ( .A1(n5033), .A2(n5954), .ZN(n8027) );
  NAND2_X1 U4986 ( .A1(n4708), .A2(n4707), .ZN(n8487) );
  AOI21_X1 U4987 ( .B1(n4269), .B2(n4712), .A(n4323), .ZN(n4707) );
  NAND2_X1 U4988 ( .A1(n4269), .A2(n8532), .ZN(n4708) );
  INV_X1 U4989 ( .A(n6532), .ZN(n7990) );
  AOI21_X1 U4990 ( .B1(n4938), .B2(n4943), .A(n4326), .ZN(n4937) );
  CLKBUF_X1 U4991 ( .A(n9049), .Z(n4635) );
  INV_X1 U4992 ( .A(n9185), .ZN(n4558) );
  NAND2_X1 U4993 ( .A1(n4480), .A2(n4479), .ZN(n4476) );
  NAND2_X1 U4994 ( .A1(n9124), .A2(n4426), .ZN(n4480) );
  OR2_X1 U4995 ( .A1(n8703), .A2(n8086), .ZN(n6053) );
  INV_X1 U4996 ( .A(n8216), .ZN(n6938) );
  NOR2_X1 U4997 ( .A1(n4566), .A2(n5456), .ZN(n4570) );
  NAND2_X1 U4998 ( .A1(n5425), .A2(n5429), .ZN(n4566) );
  NAND2_X1 U4999 ( .A1(n5431), .A2(n5430), .ZN(n5455) );
  INV_X1 U5000 ( .A(SI_12_), .ZN(n5430) );
  INV_X1 U5001 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5360) );
  INV_X1 U5002 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U5003 ( .A1(n5333), .A2(n4286), .ZN(n5406) );
  NAND2_X1 U5004 ( .A1(n5335), .A2(n10085), .ZN(n5403) );
  NAND2_X1 U5005 ( .A1(n5261), .A2(n4574), .ZN(n5264) );
  NAND2_X1 U5006 ( .A1(n4963), .A2(n5497), .ZN(n4961) );
  OR2_X1 U5007 ( .A1(n4776), .A2(n4966), .ZN(n4775) );
  OR2_X1 U5008 ( .A1(n8659), .A2(n8377), .ZN(n6075) );
  OR2_X1 U5009 ( .A1(n8675), .A2(n5893), .ZN(n5958) );
  INV_X1 U5010 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5435) );
  AOI21_X1 U5011 ( .B1(n5050), .B2(n5048), .A(n5047), .ZN(n5046) );
  INV_X1 U5012 ( .A(n6053), .ZN(n5047) );
  INV_X1 U5013 ( .A(n8510), .ZN(n5048) );
  AND2_X1 U5014 ( .A1(n5050), .A2(n4818), .ZN(n4817) );
  OR2_X1 U5015 ( .A1(n8746), .A2(n8639), .ZN(n6028) );
  OR2_X1 U5016 ( .A1(n6544), .A2(n6543), .ZN(n6919) );
  AND2_X1 U5017 ( .A1(n5143), .A2(n5141), .ZN(n5138) );
  AND4_X1 U5018 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5130), .ZN(n5137)
         );
  NOR2_X1 U5019 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5132) );
  NOR2_X1 U5020 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5131) );
  INV_X1 U5021 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5464) );
  AND2_X1 U5022 ( .A1(n5077), .A2(n7791), .ZN(n5076) );
  NOR2_X1 U5023 ( .A1(n7000), .A2(n5083), .ZN(n5082) );
  INV_X1 U5024 ( .A(n6991), .ZN(n5083) );
  INV_X1 U5025 ( .A(n7008), .ZN(n4492) );
  NOR2_X1 U5026 ( .A1(n9376), .A2(n9052), .ZN(n9180) );
  OR2_X1 U5027 ( .A1(n7610), .A2(n9877), .ZN(n6188) );
  NAND2_X1 U5028 ( .A1(n4873), .A2(n4365), .ZN(n4544) );
  OR2_X1 U5029 ( .A1(n7998), .A2(n9391), .ZN(n9171) );
  OR2_X1 U5030 ( .A1(n9648), .A2(n9483), .ZN(n9185) );
  NAND2_X1 U5031 ( .A1(n5921), .A2(n4370), .ZN(n4590) );
  NAND2_X1 U5032 ( .A1(n5117), .A2(n6309), .ZN(n5075) );
  INV_X1 U5033 ( .A(n5503), .ZN(n4866) );
  OR2_X1 U5034 ( .A1(n8181), .A2(n4273), .ZN(n4857) );
  AND2_X1 U5035 ( .A1(n6401), .A2(n5504), .ZN(n5225) );
  NOR2_X1 U5036 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5134) );
  NAND2_X1 U5037 ( .A1(n5137), .A2(n5266), .ZN(n4507) );
  AND2_X1 U5038 ( .A1(n4956), .A2(n5150), .ZN(n4271) );
  NOR2_X1 U5039 ( .A1(n8703), .A2(n4990), .ZN(n4989) );
  INV_X1 U5040 ( .A(n4991), .ZN(n4990) );
  NAND2_X1 U5041 ( .A1(n8504), .A2(n8510), .ZN(n5052) );
  AOI21_X1 U5042 ( .B1(n4714), .B2(n4711), .A(n4299), .ZN(n4710) );
  INV_X1 U5043 ( .A(n8014), .ZN(n4711) );
  NAND2_X1 U5044 ( .A1(n4896), .A2(n4394), .ZN(n8532) );
  AOI21_X1 U5045 ( .B1(n4898), .B2(n8011), .A(n4324), .ZN(n4896) );
  NAND2_X1 U5046 ( .A1(n4898), .A2(n8576), .ZN(n4394) );
  NAND2_X1 U5047 ( .A1(n8620), .A2(n6028), .ZN(n8593) );
  NAND2_X1 U5048 ( .A1(n6550), .A2(n6549), .ZN(n9913) );
  INV_X1 U5049 ( .A(n9985), .ZN(n9956) );
  NAND2_X1 U5050 ( .A1(n4955), .A2(n7278), .ZN(n9986) );
  NAND2_X1 U5051 ( .A1(n5831), .A2(n9932), .ZN(n7145) );
  NAND2_X1 U5052 ( .A1(n4726), .A2(n5061), .ZN(n4725) );
  INV_X1 U5053 ( .A(n7345), .ZN(n4726) );
  AND3_X1 U5054 ( .A1(n4382), .A2(n4358), .A3(n4384), .ZN(n7693) );
  AND2_X1 U5055 ( .A1(n4385), .A2(n4383), .ZN(n4382) );
  NAND2_X1 U5056 ( .A1(n4722), .A2(n4724), .ZN(n4719) );
  AND2_X1 U5057 ( .A1(n9261), .A2(n7276), .ZN(n9267) );
  INV_X1 U5058 ( .A(n9180), .ZN(n9258) );
  AND2_X1 U5059 ( .A1(n4881), .A2(n4878), .ZN(n4877) );
  INV_X1 U5060 ( .A(n6346), .ZN(n4878) );
  XNOR2_X1 U5061 ( .A(n4407), .B(n7739), .ZN(n9370) );
  NAND2_X1 U5062 ( .A1(n9366), .A2(n4368), .ZN(n4407) );
  NAND2_X1 U5063 ( .A1(n7983), .A2(n4573), .ZN(n9415) );
  NOR2_X1 U5064 ( .A1(n9410), .A2(n9038), .ZN(n4573) );
  AOI21_X1 U5065 ( .B1(n4942), .B2(n4941), .A(n4339), .ZN(n4940) );
  NAND2_X1 U5066 ( .A1(n9249), .A2(n9163), .ZN(n9410) );
  NAND2_X1 U5067 ( .A1(n7971), .A2(n7970), .ZN(n9442) );
  NAND2_X1 U5068 ( .A1(n4417), .A2(n4416), .ZN(n7971) );
  AND2_X1 U5069 ( .A1(n4418), .A2(n7969), .ZN(n4416) );
  AOI21_X1 U5070 ( .B1(n5099), .B2(n5101), .A(n5098), .ZN(n5097) );
  NOR2_X1 U5071 ( .A1(n5106), .A2(n9068), .ZN(n5099) );
  AND2_X1 U5072 ( .A1(n7833), .A2(n7832), .ZN(n7957) );
  NAND2_X1 U5073 ( .A1(n9470), .A2(n4420), .ZN(n4417) );
  AOI21_X1 U5074 ( .B1(n9479), .B2(n9184), .A(n9475), .ZN(n9478) );
  NOR2_X1 U5075 ( .A1(n4330), .A2(n4948), .ZN(n4947) );
  INV_X1 U5076 ( .A(n7924), .ZN(n4948) );
  NOR2_X1 U5077 ( .A1(n4555), .A2(n9122), .ZN(n4551) );
  AOI21_X1 U5078 ( .B1(n4782), .B2(n4780), .A(n4327), .ZN(n4779) );
  INV_X1 U5079 ( .A(n4785), .ZN(n4780) );
  AND2_X1 U5080 ( .A1(n4931), .A2(n7330), .ZN(n4930) );
  AOI21_X1 U5081 ( .B1(n7072), .B2(n9195), .A(n7071), .ZN(n7073) );
  AND2_X1 U5082 ( .A1(n6467), .A2(n6466), .ZN(n9496) );
  OR2_X1 U5083 ( .A1(n9226), .A2(n9780), .ZN(n9501) );
  INV_X1 U5084 ( .A(n9574), .ZN(n9499) );
  INV_X1 U5085 ( .A(n9496), .ZN(n9577) );
  NOR2_X1 U5086 ( .A1(n6150), .A2(n7606), .ZN(n4501) );
  XNOR2_X1 U5087 ( .A(n5908), .B(n5907), .ZN(n9044) );
  NAND2_X1 U5088 ( .A1(n5921), .A2(n5920), .ZN(n5908) );
  XNOR2_X1 U5089 ( .A(n6212), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6280) );
  INV_X1 U5090 ( .A(n4580), .ZN(n5639) );
  AOI21_X1 U5091 ( .B1(n4586), .B2(n4584), .A(n4583), .ZN(n4580) );
  NAND2_X1 U5092 ( .A1(n5556), .A2(n5555), .ZN(n5569) );
  NAND2_X1 U5093 ( .A1(n10036), .A2(n6138), .ZN(n6174) );
  NAND2_X1 U5094 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n10036) );
  INV_X1 U5095 ( .A(n8186), .ZN(n8195) );
  XNOR2_X1 U5096 ( .A(n4900), .B(n8027), .ZN(n8669) );
  AOI21_X1 U5097 ( .B1(n8390), .B2(n4825), .A(n8026), .ZN(n4900) );
  NAND2_X1 U5098 ( .A1(n7864), .A2(n7863), .ZN(n9612) );
  OAI21_X1 U5099 ( .B1(n9229), .B2(n9226), .A(n9260), .ZN(n4454) );
  AND2_X1 U5100 ( .A1(n9086), .A2(n4741), .ZN(n4740) );
  INV_X1 U5101 ( .A(n9089), .ZN(n4742) );
  AOI21_X1 U5102 ( .B1(n5989), .B2(n4514), .A(n4807), .ZN(n4806) );
  INV_X1 U5103 ( .A(n5992), .ZN(n4807) );
  NAND2_X1 U5104 ( .A1(n5984), .A2(n4515), .ZN(n4514) );
  OAI211_X1 U5105 ( .C1(n9091), .C2(n9098), .A(n9090), .B(n9095), .ZN(n4739)
         );
  AND2_X1 U5106 ( .A1(n4456), .A2(n9177), .ZN(n4455) );
  OR2_X1 U5107 ( .A1(n4462), .A2(n4738), .ZN(n4456) );
  AND2_X1 U5108 ( .A1(n9101), .A2(n9092), .ZN(n4738) );
  NAND2_X1 U5109 ( .A1(n4460), .A2(n4281), .ZN(n4459) );
  NAND2_X1 U5110 ( .A1(n4462), .A2(n9177), .ZN(n4460) );
  INV_X1 U5111 ( .A(n6020), .ZN(n4794) );
  NAND2_X1 U5112 ( .A1(n9109), .A2(n4735), .ZN(n9108) );
  AND2_X1 U5113 ( .A1(n9104), .A2(n9105), .ZN(n4735) );
  AND2_X1 U5114 ( .A1(n9211), .A2(n9131), .ZN(n4479) );
  MUX2_X1 U5115 ( .A(n9143), .B(n9142), .S(n9177), .Z(n9152) );
  NAND2_X1 U5116 ( .A1(n4512), .A2(n4309), .ZN(n4511) );
  NAND2_X1 U5117 ( .A1(n4509), .A2(n4508), .ZN(n4512) );
  NOR2_X1 U5118 ( .A1(n4513), .A2(n4277), .ZN(n4508) );
  NAND2_X1 U5119 ( .A1(n4801), .A2(n4800), .ZN(n4651) );
  INV_X1 U5120 ( .A(n6066), .ZN(n4800) );
  OR2_X1 U5121 ( .A1(n4802), .A2(n5035), .ZN(n4801) );
  INV_X1 U5122 ( .A(n6073), .ZN(n4612) );
  INV_X1 U5123 ( .A(n6074), .ZN(n4611) );
  NAND2_X1 U5124 ( .A1(n4578), .A2(n4571), .ZN(n4577) );
  NAND2_X1 U5125 ( .A1(n4568), .A2(n4567), .ZN(n4571) );
  AOI21_X1 U5126 ( .B1(n5014), .B2(n5016), .A(n5462), .ZN(n4578) );
  NOR2_X1 U5127 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  NAND2_X1 U5128 ( .A1(n5459), .A2(n5458), .ZN(n5481) );
  INV_X1 U5129 ( .A(SI_13_), .ZN(n5458) );
  NAND2_X1 U5130 ( .A1(n5386), .A2(n5385), .ZN(n5408) );
  NAND2_X1 U5131 ( .A1(n5363), .A2(SI_9_), .ZN(n5407) );
  OAI21_X1 U5132 ( .B1(n5504), .B2(n4629), .A(n4628), .ZN(n5307) );
  NAND2_X1 U5133 ( .A1(n5504), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4628) );
  OAI21_X1 U5134 ( .B1(n5504), .B2(n4676), .A(n4675), .ZN(n5262) );
  XNOR2_X1 U5135 ( .A(n7054), .B(n5802), .ZN(n5235) );
  AND2_X1 U5136 ( .A1(n5269), .A2(n8216), .ZN(n5211) );
  NOR2_X1 U5137 ( .A1(n5755), .A2(n8183), .ZN(n4682) );
  NAND2_X1 U5138 ( .A1(n4338), .A2(n5454), .ZN(n4776) );
  OAI21_X1 U5139 ( .B1(n4810), .B2(n4809), .A(n6055), .ZN(n6057) );
  NOR2_X1 U5140 ( .A1(n6040), .A2(n6079), .ZN(n4809) );
  INV_X1 U5141 ( .A(n8680), .ZN(n4978) );
  INV_X1 U5142 ( .A(n5665), .ZN(n5664) );
  AND2_X1 U5143 ( .A1(n8517), .A2(n4715), .ZN(n4714) );
  NAND2_X1 U5144 ( .A1(n8015), .A2(n8014), .ZN(n4715) );
  NAND2_X1 U5145 ( .A1(n5013), .A2(n8563), .ZN(n6041) );
  OR2_X1 U5146 ( .A1(n8731), .A2(n8111), .ZN(n5963) );
  INV_X1 U5147 ( .A(n6032), .ZN(n5045) );
  OAI21_X1 U5148 ( .B1(n8594), .B2(n5045), .A(n5966), .ZN(n5044) );
  AND2_X1 U5149 ( .A1(n5963), .A2(n5962), .ZN(n8010) );
  NOR2_X1 U5150 ( .A1(n8608), .A2(n4987), .ZN(n4986) );
  INV_X1 U5151 ( .A(n4988), .ZN(n4987) );
  NOR2_X1 U5152 ( .A1(n8652), .A2(n8746), .ZN(n4988) );
  NOR2_X1 U5153 ( .A1(n8002), .A2(n8207), .ZN(n4699) );
  OR2_X1 U5154 ( .A1(n8002), .A2(n8642), .ZN(n6015) );
  NOR2_X1 U5155 ( .A1(n5938), .A2(n4835), .ZN(n4834) );
  INV_X1 U5156 ( .A(n6001), .ZN(n4835) );
  AND2_X1 U5157 ( .A1(n4391), .A2(n4390), .ZN(n7380) );
  OR2_X1 U5158 ( .A1(n8764), .A2(n8210), .ZN(n4390) );
  NAND2_X1 U5159 ( .A1(n4331), .A2(n4392), .ZN(n4391) );
  NAND2_X1 U5160 ( .A1(n7471), .A2(n5885), .ZN(n6001) );
  AND2_X1 U5161 ( .A1(n7467), .A2(n5997), .ZN(n5054) );
  AOI21_X1 U5162 ( .B1(n4704), .B2(n4703), .A(n4321), .ZN(n4702) );
  OR2_X1 U5163 ( .A1(n7179), .A2(n4631), .ZN(n5126) );
  NAND2_X1 U5164 ( .A1(n6942), .A2(n9898), .ZN(n5985) );
  NAND2_X1 U5165 ( .A1(n4884), .A2(n4887), .ZN(n5975) );
  AND2_X1 U5166 ( .A1(n4885), .A2(n5036), .ZN(n4884) );
  AND2_X1 U5167 ( .A1(n8218), .A2(n6931), .ZN(n6934) );
  NAND2_X1 U5168 ( .A1(n9941), .A2(n9911), .ZN(n7024) );
  AND2_X1 U5169 ( .A1(n5168), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4400) );
  NOR2_X1 U5170 ( .A1(n5364), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5438) );
  XNOR2_X1 U5171 ( .A(n4387), .B(n7890), .ZN(n7686) );
  AOI21_X1 U5172 ( .B1(n9682), .B2(n7893), .A(n4322), .ZN(n4387) );
  INV_X1 U5173 ( .A(n9043), .ZN(n4656) );
  INV_X1 U5174 ( .A(n9251), .ZN(n4657) );
  OR2_X1 U5175 ( .A1(n9383), .A2(n9053), .ZN(n9175) );
  AND2_X1 U5176 ( .A1(n9171), .A2(n9064), .ZN(n4625) );
  INV_X1 U5177 ( .A(n6344), .ZN(n4876) );
  NAND2_X1 U5178 ( .A1(n4544), .A2(n9311), .ZN(n9297) );
  OR2_X1 U5179 ( .A1(n9616), .A2(n9412), .ZN(n9165) );
  NOR2_X1 U5180 ( .A1(n5108), .A2(n4555), .ZN(n4553) );
  NOR2_X1 U5181 ( .A1(n4307), .A2(n4783), .ZN(n4782) );
  INV_X1 U5182 ( .A(n4950), .ZN(n4783) );
  NAND2_X1 U5183 ( .A1(n9678), .A2(n7662), .ZN(n9114) );
  NOR2_X1 U5184 ( .A1(n7455), .A2(n9694), .ZN(n4912) );
  INV_X1 U5185 ( .A(n7328), .ZN(n4935) );
  NAND2_X1 U5186 ( .A1(n7166), .A2(n9090), .ZN(n7280) );
  NOR2_X1 U5187 ( .A1(n4916), .A2(n7108), .ZN(n4915) );
  NAND2_X1 U5188 ( .A1(n9845), .A2(n9851), .ZN(n4916) );
  AND2_X1 U5189 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  NAND2_X1 U5190 ( .A1(n4588), .A2(n5691), .ZN(n5742) );
  OAI21_X1 U5191 ( .B1(n5654), .B2(n5653), .A(n5657), .ZN(n5682) );
  NAND2_X1 U5192 ( .A1(n5593), .A2(n5592), .ZN(n4586) );
  AND2_X1 U5193 ( .A1(n5555), .A2(n5529), .ZN(n5553) );
  AOI21_X1 U5194 ( .B1(n4865), .B2(n5499), .A(n4863), .ZN(n4862) );
  INV_X1 U5195 ( .A(n5522), .ZN(n4863) );
  NAND2_X1 U5196 ( .A1(n5502), .A2(SI_14_), .ZN(n5503) );
  NOR2_X1 U5197 ( .A1(n4570), .A2(n5015), .ZN(n5014) );
  NAND2_X1 U5198 ( .A1(n5455), .A2(n5433), .ZN(n5456) );
  XNOR2_X1 U5199 ( .A(n5427), .B(SI_11_), .ZN(n5424) );
  NAND2_X1 U5200 ( .A1(n4567), .A2(n5408), .ZN(n5426) );
  NAND2_X1 U5201 ( .A1(n5362), .A2(n5361), .ZN(n5404) );
  INV_X1 U5202 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U5203 ( .A1(n5403), .A2(n5337), .ZN(n5357) );
  NAND2_X1 U5204 ( .A1(n4380), .A2(n4378), .ZN(n5333) );
  NAND2_X1 U5205 ( .A1(n4381), .A2(n5308), .ZN(n4380) );
  INV_X1 U5206 ( .A(n4379), .ZN(n4378) );
  INV_X1 U5207 ( .A(n4547), .ZN(n4381) );
  INV_X1 U5208 ( .A(n5280), .ZN(n5281) );
  NAND2_X1 U5209 ( .A1(n5264), .A2(n5263), .ZN(n5282) );
  XNOR2_X1 U5210 ( .A(n5262), .B(n4995), .ZN(n5261) );
  INV_X1 U5211 ( .A(SI_4_), .ZN(n4995) );
  NAND2_X1 U5212 ( .A1(n4965), .A2(n5480), .ZN(n4964) );
  INV_X1 U5213 ( .A(n7573), .ZN(n4965) );
  INV_X1 U5214 ( .A(n4765), .ZN(n4764) );
  OAI21_X1 U5215 ( .B1(n4769), .B2(n4767), .A(n6909), .ZN(n4765) );
  NAND2_X1 U5216 ( .A1(n6831), .A2(n4761), .ZN(n4766) );
  AND2_X1 U5217 ( .A1(n6832), .A2(n5327), .ZN(n4761) );
  NAND2_X1 U5218 ( .A1(n4682), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5792) );
  INV_X1 U5219 ( .A(n4854), .ZN(n4851) );
  AOI21_X1 U5220 ( .B1(n4854), .B2(n4856), .A(n5857), .ZN(n4850) );
  INV_X1 U5221 ( .A(n4973), .ZN(n4970) );
  INV_X1 U5222 ( .A(n7335), .ZN(n4399) );
  NAND2_X1 U5223 ( .A1(n8137), .A2(n5260), .ZN(n6794) );
  NAND2_X1 U5224 ( .A1(n6794), .A2(n6795), .ZN(n6793) );
  OAI21_X1 U5225 ( .B1(n8157), .B2(n4337), .A(n4959), .ZN(n8124) );
  NAND2_X1 U5226 ( .A1(n4749), .A2(n5705), .ZN(n4959) );
  AND2_X1 U5227 ( .A1(n5380), .A2(n5355), .ZN(n4957) );
  NAND2_X1 U5228 ( .A1(n6793), .A2(n5279), .ZN(n6831) );
  NAND2_X1 U5229 ( .A1(n5027), .A2(n5029), .ZN(n5022) );
  INV_X1 U5230 ( .A(n7554), .ZN(n5972) );
  INV_X1 U5231 ( .A(n5314), .ZN(n5862) );
  OR2_X1 U5232 ( .A1(n7210), .A2(n4602), .ZN(n4601) );
  NOR2_X1 U5233 ( .A1(n7214), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4602) );
  NOR2_X1 U5234 ( .A1(n8410), .A2(n5035), .ZN(n5034) );
  NAND2_X1 U5235 ( .A1(n4893), .A2(n4267), .ZN(n4892) );
  INV_X1 U5236 ( .A(n8019), .ZN(n4893) );
  NAND2_X1 U5237 ( .A1(n4290), .A2(n4267), .ZN(n4891) );
  NAND2_X1 U5238 ( .A1(n8021), .A2(n8018), .ZN(n8019) );
  NAND2_X1 U5239 ( .A1(n6064), .A2(n6063), .ZN(n8426) );
  NAND2_X1 U5240 ( .A1(n8699), .A2(n8017), .ZN(n8463) );
  AND2_X1 U5241 ( .A1(n8424), .A2(n5959), .ZN(n8464) );
  OAI21_X1 U5242 ( .B1(n5049), .B2(n4815), .A(n5046), .ZN(n4814) );
  XNOR2_X1 U5243 ( .A(n8696), .B(n8165), .ZN(n8482) );
  INV_X1 U5244 ( .A(n4714), .ZN(n4712) );
  NAND2_X1 U5245 ( .A1(n8549), .A2(n4993), .ZN(n8524) );
  AND2_X1 U5246 ( .A1(n6041), .A2(n6044), .ZN(n8554) );
  NAND2_X1 U5247 ( .A1(n4837), .A2(n5963), .ZN(n8546) );
  NAND2_X1 U5248 ( .A1(n8562), .A2(n8010), .ZN(n4837) );
  INV_X1 U5249 ( .A(n8010), .ZN(n8561) );
  NAND2_X1 U5250 ( .A1(n8600), .A2(n8008), .ZN(n8576) );
  OR2_X1 U5251 ( .A1(n8576), .A2(n8575), .ZN(n8578) );
  NAND2_X1 U5252 ( .A1(n8593), .A2(n8594), .ZN(n8592) );
  NAND2_X1 U5253 ( .A1(n4695), .A2(n4694), .ZN(n8600) );
  AOI21_X1 U5254 ( .B1(n4697), .B2(n4700), .A(n8594), .ZN(n4694) );
  NAND2_X1 U5255 ( .A1(n8004), .A2(n4697), .ZN(n4695) );
  INV_X1 U5256 ( .A(n8623), .ZN(n5057) );
  NAND2_X1 U5257 ( .A1(n8638), .A2(n6021), .ZN(n8622) );
  NAND2_X1 U5258 ( .A1(n7373), .A2(n6010), .ZN(n7429) );
  AND2_X1 U5259 ( .A1(n6010), .A2(n7428), .ZN(n7383) );
  AND2_X1 U5260 ( .A1(n7380), .A2(n7389), .ZN(n4906) );
  AND2_X1 U5261 ( .A1(n5992), .A2(n6957), .ZN(n7191) );
  NAND2_X1 U5262 ( .A1(n6946), .A2(n5126), .ZN(n7192) );
  AOI21_X1 U5263 ( .B1(n7058), .B2(n4895), .A(n4333), .ZN(n4894) );
  NAND2_X1 U5264 ( .A1(n6940), .A2(n6939), .ZN(n7052) );
  NAND2_X1 U5265 ( .A1(n6937), .A2(n9923), .ZN(n6940) );
  NAND2_X1 U5266 ( .A1(n5811), .A2(n5810), .ZN(n8670) );
  NAND2_X1 U5267 ( .A1(n9736), .A2(n5216), .ZN(n5811) );
  INV_X1 U5268 ( .A(n8687), .ZN(n4663) );
  NOR2_X1 U5269 ( .A1(n6919), .A2(n6546), .ZN(n7146) );
  AND2_X1 U5270 ( .A1(n5830), .A2(n8806), .ZN(n9929) );
  AND2_X1 U5271 ( .A1(n4839), .A2(n5176), .ZN(n5053) );
  NOR2_X1 U5272 ( .A1(n5816), .A2(n5819), .ZN(n5823) );
  NAND2_X1 U5273 ( .A1(n7006), .A2(n7005), .ZN(n7007) );
  AOI21_X1 U5274 ( .B1(n5086), .B2(n8881), .A(n4342), .ZN(n5085) );
  NAND2_X1 U5275 ( .A1(n4729), .A2(n4292), .ZN(n4728) );
  INV_X2 U5276 ( .A(n6524), .ZN(n7893) );
  NAND2_X1 U5277 ( .A1(n7007), .A2(n7008), .ZN(n7238) );
  OR2_X1 U5278 ( .A1(n6489), .A2(n7763), .ZN(n6490) );
  INV_X1 U5279 ( .A(n7772), .ZN(n5080) );
  NAND2_X1 U5280 ( .A1(n5065), .A2(n7698), .ZN(n4718) );
  INV_X1 U5281 ( .A(n7665), .ZN(n5070) );
  NAND2_X1 U5282 ( .A1(n4672), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7703) );
  XNOR2_X1 U5283 ( .A(n4603), .B(n7890), .ZN(n8914) );
  NAND2_X1 U5284 ( .A1(n4605), .A2(n4604), .ZN(n4603) );
  NAND2_X1 U5285 ( .A1(n9448), .A2(n7892), .ZN(n4604) );
  NAND2_X1 U5286 ( .A1(n9628), .A2(n7893), .ZN(n4605) );
  NOR2_X1 U5287 ( .A1(n6979), .A2(n4488), .ZN(n4487) );
  INV_X1 U5288 ( .A(n6514), .ZN(n4488) );
  INV_X1 U5289 ( .A(n6980), .ZN(n4486) );
  NAND2_X1 U5290 ( .A1(n7654), .A2(n7653), .ZN(n4483) );
  INV_X1 U5291 ( .A(n7344), .ZN(n4724) );
  OAI21_X1 U5292 ( .B1(n7006), .B2(n4492), .A(n4490), .ZN(n5058) );
  NOR2_X1 U5293 ( .A1(n4491), .A2(n5059), .ZN(n4490) );
  NOR2_X1 U5294 ( .A1(n7005), .A2(n4492), .ZN(n4491) );
  INV_X1 U5295 ( .A(n7445), .ZN(n4723) );
  AND2_X1 U5296 ( .A1(n6188), .A2(n6187), .ZN(n6223) );
  XNOR2_X1 U5297 ( .A(n6503), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U5298 ( .A1(n4414), .A2(n4413), .ZN(n6257) );
  NAND2_X1 U5299 ( .A1(n6521), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4413) );
  OR2_X1 U5300 ( .A1(n6521), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4414) );
  NAND2_X1 U5301 ( .A1(n6383), .A2(n4412), .ZN(n6198) );
  OR2_X1 U5302 ( .A1(n6194), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4412) );
  NOR2_X1 U5303 ( .A1(n6198), .A2(n6197), .ZN(n6239) );
  OR2_X1 U5304 ( .A1(n9794), .A2(n9795), .ZN(n4880) );
  NAND2_X1 U5305 ( .A1(n4543), .A2(n4542), .ZN(n9798) );
  INV_X1 U5306 ( .A(n6270), .ZN(n4542) );
  INV_X1 U5307 ( .A(n6269), .ZN(n4543) );
  AOI21_X1 U5308 ( .B1(n6344), .B2(n9795), .A(n4325), .ZN(n4881) );
  OR2_X1 U5309 ( .A1(n7255), .A2(n7253), .ZN(n4874) );
  NAND2_X1 U5310 ( .A1(n4617), .A2(n4363), .ZN(n4873) );
  OR2_X1 U5311 ( .A1(n7134), .A2(n7135), .ZN(n7254) );
  NAND2_X1 U5312 ( .A1(n9310), .A2(n4405), .ZN(n9322) );
  OR2_X1 U5313 ( .A1(n9311), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4405) );
  OR2_X1 U5314 ( .A1(n9327), .A2(n9326), .ZN(n4409) );
  NOR2_X1 U5315 ( .A1(n9334), .A2(n4540), .ZN(n9337) );
  AND2_X1 U5316 ( .A1(n9340), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4540) );
  OR2_X1 U5317 ( .A1(n9337), .A2(n9336), .ZN(n4539) );
  AND2_X1 U5318 ( .A1(n4539), .A2(n4538), .ZN(n9352) );
  NAND2_X1 U5319 ( .A1(n9355), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4538) );
  NOR2_X1 U5320 ( .A1(n9352), .A2(n9351), .ZN(n9364) );
  NAND2_X1 U5321 ( .A1(n7631), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n7882) );
  INV_X1 U5322 ( .A(n7866), .ZN(n7631) );
  INV_X1 U5323 ( .A(n4923), .ZN(n4921) );
  OR2_X1 U5324 ( .A1(n9436), .A2(n4924), .ZN(n9404) );
  INV_X1 U5325 ( .A(n9612), .ZN(n9409) );
  AND2_X1 U5326 ( .A1(n9165), .A2(n9162), .ZN(n9426) );
  NOR2_X1 U5327 ( .A1(n9436), .A2(n9616), .ZN(n9423) );
  INV_X1 U5328 ( .A(n9426), .ZN(n4681) );
  NAND2_X1 U5329 ( .A1(n9422), .A2(n9572), .ZN(n4679) );
  NOR2_X1 U5330 ( .A1(n9628), .A2(n9450), .ZN(n9435) );
  NAND2_X1 U5331 ( .A1(n9183), .A2(n9155), .ZN(n5107) );
  AOI21_X1 U5332 ( .B1(n5106), .B2(n5103), .A(n5102), .ZN(n5101) );
  AOI21_X1 U5333 ( .B1(n4420), .B2(n4419), .A(n4317), .ZN(n4418) );
  INV_X1 U5334 ( .A(n4289), .ZN(n4419) );
  OR2_X1 U5335 ( .A1(n7950), .A2(n7968), .ZN(n9216) );
  INV_X1 U5336 ( .A(n9214), .ZN(n9456) );
  AND2_X1 U5337 ( .A1(n9468), .A2(n9447), .ZN(n9183) );
  NAND2_X1 U5338 ( .A1(n7946), .A2(n7945), .ZN(n9470) );
  NAND2_X1 U5339 ( .A1(n4429), .A2(n4310), .ZN(n7946) );
  AOI21_X1 U5340 ( .B1(n7940), .B2(n4431), .A(n4303), .ZN(n4430) );
  INV_X1 U5341 ( .A(n7938), .ZN(n4431) );
  AND2_X1 U5342 ( .A1(n7742), .A2(n7741), .ZN(n9498) );
  NOR2_X1 U5343 ( .A1(n7954), .A2(n9535), .ZN(n4565) );
  AOI21_X1 U5344 ( .B1(n4564), .B2(n7954), .A(n4563), .ZN(n4562) );
  AND2_X1 U5345 ( .A1(n9185), .A2(n9184), .ZN(n9495) );
  NAND2_X1 U5346 ( .A1(n9534), .A2(n7936), .ZN(n9519) );
  AND2_X1 U5347 ( .A1(n7935), .A2(n7926), .ZN(n4789) );
  NAND2_X1 U5348 ( .A1(n9560), .A2(n9561), .ZN(n7925) );
  OR2_X1 U5349 ( .A1(n9128), .A2(n9127), .ZN(n9546) );
  INV_X1 U5350 ( .A(n5108), .ZN(n4556) );
  NAND2_X1 U5351 ( .A1(n9570), .A2(n9571), .ZN(n9569) );
  INV_X1 U5352 ( .A(n4782), .ZN(n4781) );
  NAND2_X1 U5353 ( .A1(n9021), .A2(n9114), .ZN(n7588) );
  AND3_X1 U5354 ( .A1(n7596), .A2(n7595), .A3(n7594), .ZN(n7952) );
  NOR2_X1 U5355 ( .A1(n7585), .A2(n9678), .ZN(n9578) );
  OR2_X1 U5356 ( .A1(n9682), .A2(n9275), .ZN(n4950) );
  NOR2_X1 U5357 ( .A1(n7580), .A2(n4786), .ZN(n4785) );
  INV_X1 U5358 ( .A(n7515), .ZN(n4786) );
  NAND2_X1 U5359 ( .A1(n7280), .A2(n9092), .ZN(n7614) );
  AND2_X1 U5360 ( .A1(n9101), .A2(n9093), .ZN(n9203) );
  NAND2_X1 U5361 ( .A1(n9866), .A2(n7152), .ZN(n7327) );
  NAND2_X1 U5362 ( .A1(n7010), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7096) );
  INV_X1 U5363 ( .A(n7012), .ZN(n7010) );
  AND4_X1 U5364 ( .A1(n7101), .A2(n7100), .A3(n7099), .A4(n7098), .ZN(n7618)
         );
  NAND2_X1 U5365 ( .A1(n9242), .A2(n9073), .ZN(n9187) );
  AOI21_X1 U5366 ( .B1(n4438), .B2(n6868), .A(n4436), .ZN(n4440) );
  NAND2_X1 U5367 ( .A1(n6867), .A2(n7087), .ZN(n4441) );
  NOR2_X1 U5368 ( .A1(n4438), .A2(n4437), .ZN(n4436) );
  AND2_X1 U5369 ( .A1(n6469), .A2(n9780), .ZN(n9574) );
  NAND2_X1 U5370 ( .A1(n7948), .A2(n7947), .ZN(n9636) );
  INV_X1 U5371 ( .A(n9869), .ZN(n9835) );
  INV_X1 U5372 ( .A(n9868), .ZN(n9834) );
  OR2_X1 U5373 ( .A1(n6519), .A2(n7609), .ZN(n6458) );
  AND3_X1 U5374 ( .A1(n6322), .A2(n6437), .A3(n6321), .ZN(n6606) );
  XNOR2_X1 U5375 ( .A(n4589), .B(n5926), .ZN(n9048) );
  NAND2_X1 U5376 ( .A1(n4590), .A2(n5924), .ZN(n4589) );
  XNOR2_X1 U5377 ( .A(n5905), .B(n5900), .ZN(n8793) );
  XNOR2_X1 U5378 ( .A(n6107), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6152) );
  XNOR2_X1 U5379 ( .A(n4642), .B(n4641), .ZN(n8804) );
  INV_X1 U5380 ( .A(n5767), .ZN(n4641) );
  NAND2_X1 U5381 ( .A1(n5770), .A2(n5768), .ZN(n4642) );
  NOR2_X1 U5382 ( .A1(n5075), .A2(n5073), .ZN(n6105) );
  NAND2_X1 U5383 ( .A1(n5116), .A2(n5074), .ZN(n5073) );
  INV_X1 U5384 ( .A(n6104), .ZN(n5074) );
  AND2_X1 U5385 ( .A1(n5691), .A2(n5686), .ZN(n5689) );
  INV_X1 U5386 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U5387 ( .A1(n6173), .A2(n6139), .ZN(n6176) );
  INV_X1 U5388 ( .A(n6174), .ZN(n6173) );
  NOR2_X1 U5389 ( .A1(n9760), .A2(n9759), .ZN(n9761) );
  NAND2_X1 U5390 ( .A1(n4591), .A2(n9764), .ZN(n9765) );
  OAI21_X1 U5391 ( .B1(n5739), .B2(n4403), .A(n4401), .ZN(n4404) );
  AOI21_X1 U5392 ( .B1(n8181), .B2(n4402), .A(n4273), .ZN(n4401) );
  INV_X1 U5393 ( .A(n8181), .ZN(n4403) );
  INV_X1 U5394 ( .A(n5738), .ZN(n4402) );
  NAND2_X1 U5395 ( .A1(n5643), .A2(n5642), .ZN(n8709) );
  NAND2_X1 U5396 ( .A1(n5625), .A2(n5624), .ZN(n8714) );
  INV_X1 U5397 ( .A(n8192), .ZN(n8167) );
  AND2_X1 U5398 ( .A1(n5872), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8186) );
  INV_X1 U5399 ( .A(n8115), .ZN(n8197) );
  NAND2_X1 U5400 ( .A1(n5801), .A2(n5800), .ZN(n8205) );
  NAND2_X1 U5401 ( .A1(n5734), .A2(n5733), .ZN(n8459) );
  NAND2_X1 U5402 ( .A1(n5911), .A2(n5910), .ZN(n5030) );
  NAND2_X1 U5403 ( .A1(n9044), .A2(n5216), .ZN(n5911) );
  NAND2_X1 U5404 ( .A1(n5136), .A2(n4271), .ZN(n4503) );
  NAND2_X1 U5405 ( .A1(n8447), .A2(n8446), .ZN(n8686) );
  NAND2_X1 U5406 ( .A1(n5052), .A2(n5050), .ZN(n8491) );
  NAND2_X1 U5407 ( .A1(n4713), .A2(n8014), .ZN(n8515) );
  OR2_X1 U5408 ( .A1(n8532), .A2(n8015), .ZN(n4713) );
  OAI211_X1 U5409 ( .C1(n8669), .C2(n8751), .A(n4692), .B(n8668), .ZN(n8771)
         );
  AND2_X1 U5410 ( .A1(n7818), .A2(n7817), .ZN(n8849) );
  AND4_X1 U5411 ( .A1(n7296), .A2(n7295), .A3(n7294), .A4(n7293), .ZN(n7615)
         );
  INV_X1 U5412 ( .A(n4448), .ZN(n4447) );
  OAI22_X1 U5413 ( .A1(n4449), .A2(n6519), .B1(n9049), .B2(n6522), .ZN(n4448)
         );
  AND2_X1 U5414 ( .A1(n7760), .A2(n7759), .ZN(n9483) );
  NAND2_X1 U5415 ( .A1(n9736), .A2(n7087), .ZN(n7880) );
  NAND2_X1 U5416 ( .A1(n7975), .A2(n7973), .ZN(n9622) );
  INV_X1 U5417 ( .A(n9559), .ZN(n9668) );
  NAND2_X1 U5418 ( .A1(n7701), .A2(n7700), .ZN(n9663) );
  OR2_X1 U5419 ( .A1(n8882), .A2(n7868), .ZN(n7853) );
  NAND2_X1 U5420 ( .A1(n8927), .A2(n8926), .ZN(n8925) );
  AND3_X1 U5421 ( .A1(n7707), .A2(n7706), .A3(n7705), .ZN(n8896) );
  OR2_X1 U5422 ( .A1(n6448), .A2(n6441), .ZN(n8993) );
  NAND2_X1 U5423 ( .A1(n9266), .A2(n9265), .ZN(n4623) );
  NAND2_X1 U5424 ( .A1(n4744), .A2(n9170), .ZN(n4743) );
  NAND2_X1 U5425 ( .A1(n9264), .A2(n4371), .ZN(n4452) );
  INV_X1 U5426 ( .A(n9390), .ZN(n9422) );
  INV_X1 U5427 ( .A(n8849), .ZN(n9448) );
  INV_X1 U5428 ( .A(n9483), .ZN(n9511) );
  INV_X1 U5429 ( .A(n9498), .ZN(n9524) );
  INV_X1 U5430 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4869) );
  INV_X1 U5431 ( .A(n6261), .ZN(n4536) );
  INV_X1 U5432 ( .A(n9798), .ZN(n9794) );
  AOI21_X1 U5433 ( .B1(n9808), .B2(n6341), .A(n9809), .ZN(n9806) );
  AOI21_X1 U5434 ( .B1(n6777), .B2(n6776), .A(n4410), .ZN(n7130) );
  NOR2_X1 U5435 ( .A1(n7282), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4410) );
  NAND2_X1 U5436 ( .A1(n9288), .A2(n9289), .ZN(n9310) );
  XNOR2_X1 U5437 ( .A(n9322), .B(n9323), .ZN(n9313) );
  OAI21_X1 U5438 ( .B1(n9309), .B2(n4871), .A(n4870), .ZN(n9334) );
  NAND2_X1 U5439 ( .A1(n4872), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4871) );
  NAND2_X1 U5440 ( .A1(n9319), .A2(n4872), .ZN(n4870) );
  INV_X1 U5441 ( .A(n9321), .ZN(n4872) );
  OR2_X1 U5442 ( .A1(n9373), .A2(n9372), .ZN(n4534) );
  OAI21_X1 U5443 ( .B1(n9370), .B2(n9807), .A(n4530), .ZN(n4529) );
  NAND2_X1 U5444 ( .A1(n4446), .A2(n9388), .ZN(n4445) );
  INV_X1 U5445 ( .A(n7977), .ZN(n4446) );
  AND2_X1 U5446 ( .A1(n9415), .A2(n9249), .ZN(n9389) );
  NAND2_X1 U5447 ( .A1(n4939), .A2(n4940), .ZN(n9403) );
  OR2_X1 U5448 ( .A1(n9442), .A2(n4943), .ZN(n4939) );
  INV_X1 U5449 ( .A(n9490), .ZN(n9586) );
  NAND2_X1 U5450 ( .A1(n6418), .A2(n9530), .ZN(n9589) );
  NAND2_X1 U5451 ( .A1(n4616), .A2(n9865), .ZN(n4615) );
  NAND2_X1 U5452 ( .A1(n9728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6210) );
  XNOR2_X1 U5453 ( .A(n6115), .B(n6114), .ZN(n9227) );
  NOR2_X1 U5454 ( .A1(n10031), .A2(n4377), .ZN(n10030) );
  NOR2_X1 U5455 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  OR2_X1 U5456 ( .A1(n9088), .A2(n9859), .ZN(n4741) );
  INV_X1 U5457 ( .A(n4516), .ZN(n4515) );
  NAND2_X1 U5458 ( .A1(n4812), .A2(n4811), .ZN(n5994) );
  NAND2_X1 U5459 ( .A1(n6956), .A2(n6079), .ZN(n4811) );
  NAND2_X1 U5460 ( .A1(n9094), .A2(n9093), .ZN(n4462) );
  OAI21_X1 U5461 ( .B1(n4806), .B2(n4302), .A(n4805), .ZN(n5999) );
  AND2_X1 U5462 ( .A1(n4907), .A2(n4304), .ZN(n4805) );
  NAND3_X1 U5463 ( .A1(n4458), .A2(n4457), .A3(n4461), .ZN(n9109) );
  NOR2_X1 U5464 ( .A1(n4315), .A2(n4459), .ZN(n4461) );
  AND2_X1 U5465 ( .A1(n6026), .A2(n4520), .ZN(n4519) );
  INV_X1 U5466 ( .A(n6025), .ZN(n4520) );
  NAND2_X1 U5467 ( .A1(n4522), .A2(n8631), .ZN(n4521) );
  NAND2_X1 U5468 ( .A1(n4523), .A2(n6019), .ZN(n4522) );
  NAND2_X1 U5469 ( .A1(n4795), .A2(n4316), .ZN(n4523) );
  NAND2_X1 U5470 ( .A1(n4319), .A2(n4278), .ZN(n4518) );
  NAND2_X1 U5471 ( .A1(n6041), .A2(n5012), .ZN(n5011) );
  AND2_X1 U5472 ( .A1(n5963), .A2(n6070), .ZN(n5012) );
  OR2_X1 U5473 ( .A1(n5964), .A2(n6070), .ZN(n5010) );
  OAI21_X1 U5474 ( .B1(n9125), .B2(n4477), .A(n4475), .ZN(n9139) );
  NAND2_X1 U5475 ( .A1(n9571), .A2(n4479), .ZN(n4477) );
  AND2_X1 U5476 ( .A1(n9132), .A2(n4476), .ZN(n4475) );
  NAND2_X1 U5477 ( .A1(n9139), .A2(n4478), .ZN(n9136) );
  AND2_X1 U5478 ( .A1(n9133), .A2(n9134), .ZN(n4478) );
  NAND2_X1 U5479 ( .A1(n6052), .A2(n6046), .ZN(n4513) );
  OAI21_X1 U5480 ( .B1(n4793), .B2(n4792), .A(n6036), .ZN(n6042) );
  NAND2_X1 U5481 ( .A1(n6035), .A2(n8010), .ZN(n4792) );
  NAND2_X1 U5482 ( .A1(n5011), .A2(n5010), .ZN(n6036) );
  AOI21_X1 U5483 ( .B1(n4521), .B2(n4519), .A(n4518), .ZN(n4793) );
  AOI21_X1 U5484 ( .B1(n6061), .B2(n6059), .A(n4803), .ZN(n4802) );
  MUX2_X1 U5485 ( .A(n5961), .B(n5960), .S(n6070), .Z(n6061) );
  NOR2_X1 U5486 ( .A1(n4467), .A2(n4301), .ZN(n4466) );
  INV_X1 U5487 ( .A(n9146), .ZN(n4467) );
  AOI21_X1 U5488 ( .B1(n9145), .B2(n9144), .A(n4734), .ZN(n4733) );
  NAND2_X1 U5489 ( .A1(n9157), .A2(n9153), .ZN(n4734) );
  NAND2_X1 U5490 ( .A1(n5455), .A2(n5408), .ZN(n4569) );
  AOI21_X1 U5491 ( .B1(n5029), .B2(n5033), .A(n5030), .ZN(n5028) );
  AOI211_X1 U5492 ( .C1(n4999), .C2(n6070), .A(n8482), .B(n4320), .ZN(n4810)
         );
  OAI21_X1 U5493 ( .B1(n8027), .B2(n6074), .A(n9913), .ZN(n4827) );
  INV_X1 U5494 ( .A(n7499), .ZN(n4392) );
  INV_X1 U5495 ( .A(n7203), .ZN(n4703) );
  INV_X1 U5496 ( .A(n6947), .ZN(n4705) );
  INV_X1 U5497 ( .A(n6956), .ZN(n5981) );
  NAND2_X1 U5498 ( .A1(n4464), .A2(n4463), .ZN(n4474) );
  AOI21_X1 U5499 ( .B1(n4466), .B2(n5098), .A(n9177), .ZN(n4463) );
  OR2_X1 U5500 ( .A1(n4733), .A2(n4465), .ZN(n4464) );
  INV_X1 U5501 ( .A(n4466), .ZN(n4465) );
  NOR2_X1 U5502 ( .A1(n4471), .A2(n9068), .ZN(n4470) );
  OAI21_X1 U5503 ( .B1(n9234), .B2(n9235), .A(n4926), .ZN(n9241) );
  OR2_X1 U5504 ( .A1(n9606), .A2(n9413), .ZN(n9064) );
  INV_X1 U5505 ( .A(n5555), .ZN(n5007) );
  INV_X1 U5506 ( .A(n5570), .ZN(n5009) );
  NOR2_X1 U5507 ( .A1(n4861), .A2(n4576), .ZN(n4575) );
  INV_X1 U5508 ( .A(n5481), .ZN(n4576) );
  INV_X1 U5509 ( .A(n4862), .ZN(n4861) );
  INV_X1 U5510 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5334) );
  OAI21_X1 U5511 ( .B1(n4997), .B2(n4545), .A(n5329), .ZN(n4379) );
  OAI21_X1 U5512 ( .B1(n5504), .B2(n4627), .A(n4626), .ZN(n5283) );
  INV_X1 U5513 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5514 ( .A1(n5504), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4626) );
  NAND2_X1 U5515 ( .A1(n4597), .A2(n4618), .ZN(n5240) );
  NAND2_X1 U5516 ( .A1(n5218), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4618) );
  INV_X1 U5517 ( .A(n5208), .ZN(n5199) );
  AND2_X1 U5518 ( .A1(n5207), .A2(n5206), .ZN(n6610) );
  NOR2_X1 U5519 ( .A1(n5443), .A2(n5442), .ZN(n4685) );
  AOI21_X1 U5520 ( .B1(n4774), .B2(n4776), .A(n4298), .ZN(n4772) );
  NOR2_X1 U5521 ( .A1(n5626), .A2(n8150), .ZN(n4684) );
  XNOR2_X1 U5522 ( .A(n8703), .B(n5802), .ZN(n5673) );
  AND2_X1 U5523 ( .A1(n4756), .A2(n8083), .ZN(n4755) );
  NAND2_X1 U5524 ( .A1(n4757), .A2(n5637), .ZN(n4756) );
  INV_X1 U5525 ( .A(n4759), .ZN(n4757) );
  NAND2_X1 U5526 ( .A1(n9911), .A2(n5269), .ZN(n5208) );
  OR3_X1 U5527 ( .A1(n7145), .A2(n6543), .A3(n6917), .ZN(n5869) );
  AND2_X1 U5528 ( .A1(n5935), .A2(n5033), .ZN(n5027) );
  NAND2_X1 U5529 ( .A1(n5026), .A2(n5024), .ZN(n5023) );
  INV_X1 U5530 ( .A(n5028), .ZN(n5024) );
  NAND2_X1 U5531 ( .A1(n4799), .A2(n6067), .ZN(n4798) );
  NAND2_X1 U5532 ( .A1(n4651), .A2(n4650), .ZN(n4799) );
  NOR2_X1 U5533 ( .A1(n4804), .A2(n4335), .ZN(n4527) );
  OAI21_X1 U5534 ( .B1(n8027), .B2(n5952), .A(n6073), .ZN(n4797) );
  AND2_X1 U5535 ( .A1(n4610), .A2(n6072), .ZN(n4599) );
  NAND2_X1 U5536 ( .A1(n4612), .A2(n4611), .ZN(n4610) );
  XNOR2_X1 U5537 ( .A(n5030), .B(n8204), .ZN(n4613) );
  NAND2_X1 U5538 ( .A1(n5757), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4393) );
  OR2_X1 U5539 ( .A1(n8670), .A2(n8413), .ZN(n6074) );
  NAND2_X1 U5540 ( .A1(n4818), .A2(n4821), .ZN(n4815) );
  NAND2_X1 U5541 ( .A1(n4684), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5665) );
  INV_X1 U5542 ( .A(n6046), .ZN(n4821) );
  AOI21_X1 U5543 ( .B1(n6046), .B2(n4820), .A(n4819), .ZN(n4818) );
  INV_X1 U5544 ( .A(n6050), .ZN(n4819) );
  INV_X1 U5545 ( .A(n6043), .ZN(n4820) );
  OR2_X1 U5546 ( .A1(n8714), .A2(n8085), .ZN(n6046) );
  NOR2_X1 U5547 ( .A1(n8714), .A2(n8721), .ZN(n4993) );
  INV_X1 U5548 ( .A(n4899), .ZN(n4898) );
  OAI21_X1 U5549 ( .B1(n4288), .B2(n8011), .A(n8013), .ZN(n4899) );
  NOR2_X1 U5550 ( .A1(n5516), .A2(n5515), .ZN(n4686) );
  NOR2_X1 U5551 ( .A1(n5560), .A2(n10193), .ZN(n4609) );
  INV_X1 U5552 ( .A(n4686), .ZN(n5539) );
  OR2_X1 U5553 ( .A1(n5486), .A2(n6850), .ZN(n5516) );
  OAI21_X1 U5554 ( .B1(n4906), .B2(n4905), .A(n7435), .ZN(n4904) );
  NAND2_X1 U5555 ( .A1(n4607), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5415) );
  INV_X1 U5556 ( .A(n5395), .ZN(n4607) );
  INV_X1 U5557 ( .A(n5882), .ZN(n6955) );
  INV_X1 U5558 ( .A(n6939), .ZN(n4895) );
  OR2_X1 U5559 ( .A1(n9899), .A2(n9898), .ZN(n7181) );
  OR2_X1 U5560 ( .A1(n5342), .A2(n5341), .ZN(n5364) );
  INV_X1 U5561 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5338) );
  INV_X1 U5562 ( .A(n8959), .ZN(n8957) );
  NAND2_X1 U5563 ( .A1(n7692), .A2(n7691), .ZN(n4385) );
  INV_X1 U5564 ( .A(n7237), .ZN(n5060) );
  NOR2_X1 U5565 ( .A1(n7263), .A2(n5062), .ZN(n5063) );
  INV_X1 U5566 ( .A(n5087), .ZN(n5084) );
  NOR2_X1 U5567 ( .A1(n7592), .A2(n7591), .ZN(n4672) );
  NOR2_X1 U5568 ( .A1(n4665), .A2(n5122), .ZN(n4664) );
  INV_X1 U5569 ( .A(n9166), .ZN(n4665) );
  AND2_X1 U5570 ( .A1(n9410), .A2(n4940), .ZN(n4938) );
  NOR2_X1 U5571 ( .A1(n4924), .A2(n9606), .ZN(n4923) );
  NOR2_X1 U5572 ( .A1(n9399), .A2(n5122), .ZN(n5121) );
  NAND2_X1 U5573 ( .A1(n9409), .A2(n4925), .ZN(n4924) );
  NAND2_X1 U5574 ( .A1(n7630), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7848) );
  INV_X1 U5575 ( .A(n7846), .ZN(n7630) );
  NOR2_X1 U5576 ( .A1(n5096), .A2(n9068), .ZN(n5095) );
  INV_X1 U5577 ( .A(n5101), .ZN(n5096) );
  NOR2_X1 U5578 ( .A1(n7825), .A2(n8846), .ZN(n4671) );
  NAND2_X1 U5579 ( .A1(n4430), .A2(n4432), .ZN(n4428) );
  NAND2_X1 U5580 ( .A1(n7939), .A2(n4430), .ZN(n4429) );
  NAND2_X1 U5581 ( .A1(n4920), .A2(n9517), .ZN(n4919) );
  NOR2_X1 U5582 ( .A1(n9656), .A2(n9663), .ZN(n4920) );
  NAND2_X1 U5583 ( .A1(n9106), .A2(n9206), .ZN(n5109) );
  NAND2_X1 U5584 ( .A1(n7527), .A2(n5110), .ZN(n4554) );
  NOR2_X1 U5585 ( .A1(n7588), .A2(n7589), .ZN(n5110) );
  OR2_X1 U5586 ( .A1(n7527), .A2(n9206), .ZN(n5111) );
  NAND2_X1 U5587 ( .A1(n4934), .A2(n7328), .ZN(n4933) );
  INV_X1 U5588 ( .A(n7326), .ZN(n4934) );
  NAND2_X1 U5589 ( .A1(n4283), .A2(n4935), .ZN(n4931) );
  AOI21_X1 U5590 ( .B1(n9203), .B2(n5094), .A(n5093), .ZN(n5092) );
  INV_X1 U5591 ( .A(n9092), .ZN(n5094) );
  NOR2_X1 U5592 ( .A1(n5114), .A2(n5113), .ZN(n5112) );
  NAND2_X1 U5593 ( .A1(n9232), .A2(n4926), .ZN(n7076) );
  NAND2_X1 U5594 ( .A1(n6455), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U5595 ( .A1(n4928), .A2(n4927), .ZN(n4926) );
  INV_X1 U5596 ( .A(n9081), .ZN(n4927) );
  NAND2_X1 U5597 ( .A1(n9007), .A2(n9004), .ZN(n9189) );
  OR2_X1 U5598 ( .A1(n5905), .A2(n5904), .ZN(n5921) );
  AND2_X1 U5599 ( .A1(n5806), .A2(n5777), .ZN(n5804) );
  AND2_X1 U5600 ( .A1(n5771), .A2(n5752), .ZN(n5767) );
  AND2_X1 U5601 ( .A1(n4362), .A2(n5691), .ZN(n4587) );
  INV_X1 U5602 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U5603 ( .B1(n4586), .B2(n4583), .A(n4581), .ZN(n5641) );
  INV_X1 U5604 ( .A(n4582), .ZN(n4581) );
  OAI21_X1 U5605 ( .B1(n4584), .B2(n4583), .A(n5638), .ZN(n4582) );
  NOR2_X1 U5606 ( .A1(n5618), .A2(n4585), .ZN(n4584) );
  INV_X1 U5607 ( .A(n5595), .ZN(n4585) );
  INV_X1 U5608 ( .A(n5617), .ZN(n4583) );
  NOR2_X2 U5609 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6299) );
  NAND2_X1 U5610 ( .A1(n4579), .A2(n4859), .ZN(n5556) );
  AOI21_X1 U5611 ( .B1(n4862), .B2(n4864), .A(n4860), .ZN(n4859) );
  NAND2_X1 U5612 ( .A1(n4577), .A2(n4575), .ZN(n4579) );
  INV_X1 U5613 ( .A(n5553), .ZN(n4860) );
  OR2_X1 U5614 ( .A1(n6351), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6802) );
  OR2_X1 U5615 ( .A1(n6291), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6351) );
  AOI21_X1 U5616 ( .B1(n5280), .B2(n5284), .A(n5306), .ZN(n4997) );
  NOR2_X1 U5617 ( .A1(n4998), .A2(n4549), .ZN(n4548) );
  INV_X1 U5618 ( .A(n5263), .ZN(n4549) );
  OR2_X1 U5619 ( .A1(n6143), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U5620 ( .A1(n5291), .A2(n5290), .ZN(n5316) );
  AND2_X1 U5621 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5290) );
  INV_X1 U5622 ( .A(n5294), .ZN(n5291) );
  NAND2_X1 U5623 ( .A1(n5315), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5347) );
  INV_X1 U5624 ( .A(n5316), .ZN(n5315) );
  NOR2_X1 U5625 ( .A1(n4285), .A2(n4752), .ZN(n4751) );
  INV_X1 U5626 ( .A(n4755), .ZN(n4752) );
  INV_X1 U5627 ( .A(n5637), .ZN(n4758) );
  XNOR2_X1 U5628 ( .A(n5235), .B(n4300), .ZN(n8066) );
  NOR2_X1 U5629 ( .A1(n8148), .A2(n4760), .ZN(n4759) );
  INV_X1 U5630 ( .A(n5616), .ZN(n4760) );
  NAND2_X1 U5631 ( .A1(n4606), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5443) );
  INV_X1 U5632 ( .A(n5415), .ZN(n4606) );
  INV_X1 U5633 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5442) );
  INV_X1 U5634 ( .A(n4685), .ZN(n5470) );
  INV_X1 U5635 ( .A(n7485), .ZN(n4967) );
  NAND2_X1 U5636 ( .A1(n4952), .A2(n4313), .ZN(n8137) );
  NAND2_X1 U5637 ( .A1(n4766), .A2(n4764), .ZN(n4958) );
  OR2_X1 U5638 ( .A1(n5604), .A2(n5603), .ZN(n5626) );
  INV_X1 U5639 ( .A(n4684), .ZN(n5644) );
  AND2_X1 U5640 ( .A1(n5209), .A2(n5208), .ZN(n6720) );
  NAND2_X1 U5641 ( .A1(n4609), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U5642 ( .A1(n6831), .A2(n6832), .ZN(n6830) );
  OAI21_X1 U5643 ( .B1(n4968), .B2(n4776), .A(n4774), .ZN(n8099) );
  AND2_X1 U5644 ( .A1(n6075), .A2(n5930), .ZN(n5032) );
  OAI21_X1 U5645 ( .B1(n4526), .B2(n4525), .A(n4524), .ZN(n6078) );
  AND2_X1 U5646 ( .A1(n4599), .A2(n4613), .ZN(n4524) );
  INV_X1 U5647 ( .A(n4797), .ZN(n4525) );
  AOI21_X1 U5648 ( .B1(n6060), .B2(n4527), .A(n4798), .ZN(n4526) );
  AND2_X1 U5649 ( .A1(n5038), .A2(n5197), .ZN(n5036) );
  OR2_X1 U5650 ( .A1(n5247), .A2(n5039), .ZN(n5038) );
  NAND2_X1 U5651 ( .A1(n5314), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5037) );
  AND3_X1 U5652 ( .A1(n6414), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6423) );
  OR2_X1 U5653 ( .A1(n6686), .A2(n6687), .ZN(n6705) );
  INV_X1 U5654 ( .A(n4601), .ZN(n8322) );
  INV_X1 U5655 ( .A(SI_8_), .ZN(n10085) );
  NOR2_X1 U5656 ( .A1(n4825), .A2(n8027), .ZN(n4826) );
  NAND2_X1 U5657 ( .A1(n8415), .A2(n5958), .ZN(n8397) );
  NAND2_X1 U5658 ( .A1(n8439), .A2(n4279), .ZN(n8404) );
  NAND2_X1 U5659 ( .A1(n8439), .A2(n4266), .ZN(n8432) );
  OR2_X1 U5660 ( .A1(n8688), .A2(n8132), .ZN(n8425) );
  NAND2_X1 U5661 ( .A1(n8439), .A2(n8452), .ZN(n8440) );
  AND2_X1 U5662 ( .A1(n5708), .A2(n5707), .ZN(n8478) );
  NOR2_X1 U5663 ( .A1(n4992), .A2(n8709), .ZN(n4991) );
  INV_X1 U5664 ( .A(n4993), .ZN(n4992) );
  INV_X1 U5665 ( .A(n6049), .ZN(n5051) );
  NAND2_X1 U5666 ( .A1(n5052), .A2(n6049), .ZN(n8489) );
  OAI21_X1 U5667 ( .B1(n8534), .B2(n4821), .A(n4818), .ZN(n8504) );
  NAND2_X1 U5668 ( .A1(n8549), .A2(n8081), .ZN(n8537) );
  NAND2_X1 U5669 ( .A1(n8534), .A2(n6043), .ZN(n8516) );
  INV_X1 U5670 ( .A(n6041), .ZN(n4836) );
  NAND2_X1 U5671 ( .A1(n4686), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5560) );
  INV_X1 U5672 ( .A(n4609), .ZN(n5579) );
  AOI21_X1 U5673 ( .B1(n5043), .B2(n5045), .A(n5042), .ZN(n5041) );
  NAND2_X1 U5674 ( .A1(n8593), .A2(n5043), .ZN(n5040) );
  NAND2_X1 U5675 ( .A1(n8034), .A2(n4276), .ZN(n8584) );
  NAND2_X1 U5676 ( .A1(n8034), .A2(n4986), .ZN(n8603) );
  AND2_X1 U5677 ( .A1(n4698), .A2(n8007), .ZN(n4697) );
  NAND2_X1 U5678 ( .A1(n4270), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U5679 ( .A1(n4270), .A2(n7430), .ZN(n4700) );
  NAND2_X1 U5680 ( .A1(n8034), .A2(n8753), .ZN(n8648) );
  OAI21_X1 U5681 ( .B1(n8004), .B2(n8003), .A(n4696), .ZN(n8632) );
  INV_X1 U5682 ( .A(n4699), .ZN(n4696) );
  INV_X1 U5683 ( .A(n8595), .ZN(n8639) );
  NAND2_X1 U5684 ( .A1(n5886), .A2(n6015), .ZN(n8636) );
  NOR2_X1 U5685 ( .A1(n8635), .A2(n5056), .ZN(n5055) );
  INV_X1 U5686 ( .A(n6015), .ZN(n5056) );
  INV_X1 U5687 ( .A(n7383), .ZN(n7435) );
  NAND2_X1 U5688 ( .A1(n6008), .A2(n6009), .ZN(n4829) );
  INV_X1 U5689 ( .A(n4832), .ZN(n4831) );
  OAI21_X1 U5690 ( .B1(n4834), .B2(n4833), .A(n6005), .ZN(n4832) );
  AND2_X1 U5691 ( .A1(n6949), .A2(n4979), .ZN(n7397) );
  NOR2_X1 U5692 ( .A1(n4981), .A2(n8759), .ZN(n4979) );
  NAND2_X1 U5693 ( .A1(n4830), .A2(n6009), .ZN(n7392) );
  NAND2_X1 U5694 ( .A1(n7473), .A2(n4834), .ZN(n4830) );
  NAND2_X1 U5695 ( .A1(n7381), .A2(n7380), .ZN(n7390) );
  NAND2_X1 U5696 ( .A1(n4608), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5368) );
  INV_X1 U5697 ( .A(n5347), .ZN(n4608) );
  INV_X1 U5698 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5367) );
  OR2_X1 U5699 ( .A1(n5368), .A2(n5367), .ZN(n5395) );
  NAND2_X1 U5700 ( .A1(n7473), .A2(n6001), .ZN(n7498) );
  NAND2_X1 U5701 ( .A1(n6961), .A2(n5997), .ZN(n7475) );
  NAND2_X1 U5702 ( .A1(n6949), .A2(n4272), .ZN(n7506) );
  CLKBUF_X1 U5703 ( .A(n6960), .Z(n6961) );
  INV_X1 U5704 ( .A(n9919), .ZN(n8649) );
  NAND2_X1 U5705 ( .A1(n6944), .A2(n6943), .ZN(n7179) );
  NAND2_X1 U5706 ( .A1(n9902), .A2(n9893), .ZN(n6944) );
  NAND2_X1 U5707 ( .A1(n4689), .A2(n5985), .ZN(n9893) );
  NAND2_X1 U5708 ( .A1(n9907), .A2(n5977), .ZN(n7059) );
  AND2_X1 U5709 ( .A1(n7024), .A2(n7029), .ZN(n9908) );
  NAND2_X1 U5710 ( .A1(n9922), .A2(n9908), .ZN(n9907) );
  NAND2_X1 U5711 ( .A1(n7036), .A2(n6936), .ZN(n9923) );
  NOR2_X1 U5712 ( .A1(n9916), .A2(n9915), .ZN(n9917) );
  NAND2_X1 U5713 ( .A1(n6397), .A2(n9938), .ZN(n6394) );
  NAND2_X1 U5714 ( .A1(n4886), .A2(n5975), .ZN(n7037) );
  NAND2_X1 U5715 ( .A1(n4883), .A2(n9941), .ZN(n4886) );
  NAND2_X1 U5716 ( .A1(n4887), .A2(n5036), .ZN(n4883) );
  OR2_X1 U5717 ( .A1(n6920), .A2(n6919), .ZN(n6930) );
  NAND2_X1 U5718 ( .A1(n8793), .A2(n4260), .ZN(n5902) );
  NAND2_X1 U5719 ( .A1(n5485), .A2(n5484), .ZN(n8746) );
  CLKBUF_X1 U5720 ( .A(n5867), .Z(n6410) );
  NAND2_X1 U5721 ( .A1(n4839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4838) );
  AOI21_X1 U5722 ( .B1(n4282), .B2(n4296), .A(n4400), .ZN(n4840) );
  INV_X1 U5723 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U5724 ( .A1(n4505), .A2(n5136), .ZN(n4504) );
  OR2_X1 U5725 ( .A1(n4507), .A2(n4506), .ZN(n5574) );
  NAND2_X1 U5726 ( .A1(n5136), .A2(n4956), .ZN(n4506) );
  OR2_X1 U5727 ( .A1(n5438), .A2(n5168), .ZN(n5390) );
  OAI21_X1 U5728 ( .B1(n4949), .B2(n6165), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4791) );
  OR2_X1 U5729 ( .A1(n8827), .A2(n8826), .ZN(n8889) );
  INV_X1 U5730 ( .A(n7771), .ZN(n5078) );
  NAND2_X1 U5731 ( .A1(n7965), .A2(n7087), .ZN(n7975) );
  NAND2_X1 U5732 ( .A1(n7263), .A2(n5062), .ZN(n5061) );
  NAND2_X1 U5733 ( .A1(n4670), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7158) );
  INV_X1 U5734 ( .A(n7096), .ZN(n4670) );
  AND2_X1 U5735 ( .A1(n6359), .A2(n6358), .ZN(n6365) );
  NAND2_X1 U5736 ( .A1(n6364), .A2(n6363), .ZN(n6489) );
  OR2_X1 U5737 ( .A1(n6360), .A2(n7875), .ZN(n6364) );
  AND2_X1 U5738 ( .A1(n7686), .A2(n7687), .ZN(n8946) );
  OR2_X1 U5739 ( .A1(n8823), .A2(n8944), .ZN(n8947) );
  OR2_X1 U5740 ( .A1(n7314), .A2(n7313), .ZN(n7519) );
  NAND2_X1 U5741 ( .A1(n7298), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7314) );
  INV_X1 U5742 ( .A(n7300), .ZN(n7298) );
  OR2_X1 U5743 ( .A1(n7794), .A2(n8967), .ZN(n7825) );
  NAND2_X1 U5744 ( .A1(n7289), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7300) );
  INV_X1 U5745 ( .A(n7291), .ZN(n7289) );
  OR2_X1 U5746 ( .A1(n7898), .A2(n4731), .ZN(n6508) );
  NAND2_X1 U5747 ( .A1(n4717), .A2(n5068), .ZN(n4386) );
  INV_X1 U5748 ( .A(n4717), .ZN(n4482) );
  NAND2_X1 U5749 ( .A1(n8925), .A2(n6991), .ZN(n7116) );
  NAND3_X1 U5750 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6746) );
  OR2_X1 U5751 ( .A1(n7858), .A2(n7857), .ZN(n5087) );
  OR2_X1 U5752 ( .A1(n8880), .A2(n8881), .ZN(n5088) );
  NAND2_X1 U5753 ( .A1(n7517), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7592) );
  INV_X1 U5754 ( .A(n7519), .ZN(n7517) );
  INV_X1 U5755 ( .A(n4672), .ZN(n7670) );
  AND2_X1 U5756 ( .A1(n9258), .A2(n9259), .ZN(n4620) );
  AOI21_X1 U5757 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n6230), .A(n6226), .ZN(
        n6374) );
  NOR2_X1 U5758 ( .A1(n6374), .A2(n6373), .ZN(n6372) );
  NOR2_X1 U5759 ( .A1(n6239), .A2(n4294), .ZN(n6241) );
  NAND2_X1 U5760 ( .A1(n6340), .A2(n4411), .ZN(n9808) );
  OR2_X1 U5761 ( .A1(n6969), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4411) );
  AOI21_X1 U5762 ( .B1(n9798), .B2(n4877), .A(n4541), .ZN(n6577) );
  INV_X1 U5763 ( .A(n4875), .ZN(n4541) );
  AOI21_X1 U5764 ( .B1(n4877), .B2(n4876), .A(n4291), .ZN(n4875) );
  AOI21_X1 U5765 ( .B1(n7282), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6778), .ZN(
        n6782) );
  INV_X1 U5766 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U5767 ( .A1(n9295), .A2(n9294), .ZN(n9296) );
  INV_X1 U5768 ( .A(n4544), .ZN(n9295) );
  NOR2_X1 U5769 ( .A1(n9298), .A2(n9299), .ZN(n9306) );
  NOR2_X1 U5770 ( .A1(n9306), .A2(n9307), .ZN(n9317) );
  INV_X1 U5771 ( .A(n9297), .ZN(n9307) );
  NOR2_X1 U5772 ( .A1(n9317), .A2(n9323), .ZN(n9319) );
  AND2_X1 U5773 ( .A1(n4409), .A2(n4408), .ZN(n9342) );
  NAND2_X1 U5774 ( .A1(n9340), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n4408) );
  NOR2_X1 U5775 ( .A1(n9342), .A2(n9341), .ZN(n9354) );
  AOI21_X1 U5776 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9367), .A(n9364), .ZN(
        n9365) );
  NAND2_X1 U5777 ( .A1(n9051), .A2(n9050), .ZN(n9376) );
  OR2_X1 U5778 ( .A1(n9436), .A2(n4922), .ZN(n9382) );
  NAND2_X1 U5779 ( .A1(n9603), .A2(n4923), .ZN(n4922) );
  NAND2_X1 U5780 ( .A1(n9047), .A2(n9046), .ZN(n9383) );
  NAND2_X1 U5781 ( .A1(n9171), .A2(n9253), .ZN(n9061) );
  AOI21_X1 U5782 ( .B1(n5121), .B2(n9410), .A(n5120), .ZN(n5119) );
  INV_X1 U5783 ( .A(n9062), .ZN(n5120) );
  OR2_X1 U5784 ( .A1(n8817), .A2(n7868), .ZN(n7874) );
  NAND2_X1 U5785 ( .A1(n9415), .A2(n5121), .ZN(n9387) );
  NAND2_X1 U5786 ( .A1(n4671), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7846) );
  INV_X1 U5787 ( .A(n4671), .ZN(n7827) );
  NAND2_X1 U5788 ( .A1(n4673), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7794) );
  INV_X1 U5789 ( .A(n4673), .ZN(n7776) );
  INV_X1 U5790 ( .A(n7940), .ZN(n4432) );
  INV_X1 U5791 ( .A(n7720), .ZN(n7628) );
  NOR2_X1 U5792 ( .A1(n5125), .A2(n4918), .ZN(n9526) );
  INV_X1 U5793 ( .A(n4920), .ZN(n4918) );
  NOR2_X1 U5794 ( .A1(n5125), .A2(n9663), .ZN(n9542) );
  AND2_X1 U5795 ( .A1(n5111), .A2(n5110), .ZN(n7951) );
  NAND2_X1 U5796 ( .A1(n7619), .A2(n4280), .ZN(n7585) );
  AND4_X1 U5797 ( .A1(n7524), .A2(n7523), .A3(n7522), .A4(n7521), .ZN(n7662)
         );
  NAND2_X1 U5798 ( .A1(n7516), .A2(n7515), .ZN(n7581) );
  NAND2_X1 U5799 ( .A1(n7619), .A2(n4268), .ZN(n7533) );
  NAND2_X1 U5800 ( .A1(n7619), .A2(n4912), .ZN(n7361) );
  AND2_X1 U5801 ( .A1(n7619), .A2(n7624), .ZN(n7620) );
  AOI21_X1 U5802 ( .B1(n7327), .B2(n7326), .A(n4935), .ZN(n4932) );
  AND4_X1 U5803 ( .A1(n7163), .A2(n7162), .A3(n7161), .A4(n7160), .ZN(n7364)
         );
  NAND2_X1 U5804 ( .A1(n6875), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7012) );
  INV_X1 U5805 ( .A(n6877), .ZN(n6875) );
  NAND2_X1 U5806 ( .A1(n4914), .A2(n4275), .ZN(n7171) );
  INV_X1 U5807 ( .A(n9015), .ZN(n9091) );
  NAND2_X1 U5808 ( .A1(n4914), .A2(n4915), .ZN(n7105) );
  NOR2_X1 U5809 ( .A1(n6818), .A2(n4916), .ZN(n7080) );
  NOR2_X1 U5810 ( .A1(n6818), .A2(n7048), .ZN(n6887) );
  NAND2_X1 U5811 ( .A1(n9821), .A2(n6477), .ZN(n6593) );
  NOR2_X1 U5812 ( .A1(n9199), .A2(n4443), .ZN(n4442) );
  INV_X1 U5813 ( .A(n7109), .ZN(n4443) );
  INV_X1 U5814 ( .A(n6985), .ZN(n9833) );
  OR2_X1 U5815 ( .A1(n6440), .A2(n9263), .ZN(n9869) );
  XNOR2_X1 U5816 ( .A(n5805), .B(n5804), .ZN(n8801) );
  XNOR2_X1 U5817 ( .A(n5724), .B(n5743), .ZN(n7965) );
  OAI21_X1 U5818 ( .B1(n5742), .B2(n5741), .A(n5744), .ZN(n5724) );
  NAND2_X1 U5819 ( .A1(n4586), .A2(n5595), .ZN(n5619) );
  NAND2_X1 U5820 ( .A1(n4858), .A2(n4862), .ZN(n5554) );
  NAND2_X1 U5821 ( .A1(n5500), .A2(n4865), .ZN(n4858) );
  NAND2_X1 U5822 ( .A1(n4868), .A2(n5498), .ZN(n4867) );
  INV_X1 U5823 ( .A(n5500), .ZN(n4868) );
  XNOR2_X1 U5824 ( .A(n5500), .B(n5498), .ZN(n7582) );
  AOI21_X1 U5825 ( .B1(n5426), .B2(n5017), .A(n4389), .ZN(n4388) );
  INV_X1 U5826 ( .A(n5014), .ZN(n4389) );
  OAI21_X1 U5827 ( .B1(n5426), .B2(n5425), .A(n5429), .ZN(n5457) );
  XNOR2_X1 U5828 ( .A(n5389), .B(n5124), .ZN(n7281) );
  XNOR2_X1 U5829 ( .A(n5356), .B(n5357), .ZN(n7088) );
  NAND2_X1 U5830 ( .A1(n4434), .A2(n4433), .ZN(n6867) );
  INV_X1 U5831 ( .A(n5261), .ZN(n4994) );
  NOR2_X1 U5832 ( .A1(n10208), .A2(n9762), .ZN(n9763) );
  NAND2_X1 U5833 ( .A1(n4592), .A2(n9766), .ZN(n9767) );
  NAND2_X1 U5834 ( .A1(n6830), .A2(n5305), .ZN(n6824) );
  AND2_X1 U5835 ( .A1(n4964), .A2(n4293), .ZN(n8050) );
  NAND2_X1 U5836 ( .A1(n4964), .A2(n4962), .ZN(n8049) );
  NAND2_X1 U5837 ( .A1(n5688), .A2(n5687), .ZN(n8696) );
  INV_X1 U5838 ( .A(n4397), .ZN(n4396) );
  OAI21_X1 U5839 ( .B1(n4764), .B2(n4398), .A(n5381), .ZN(n4397) );
  INV_X1 U5840 ( .A(n4957), .ZN(n4398) );
  AND2_X1 U5841 ( .A1(n5858), .A2(n5793), .ZN(n8392) );
  AND2_X1 U5842 ( .A1(n4849), .A2(n4848), .ZN(n4847) );
  AOI21_X1 U5843 ( .B1(n4850), .B2(n4851), .A(n4297), .ZN(n4848) );
  NAND2_X1 U5844 ( .A1(n4852), .A2(n4856), .ZN(n4849) );
  OAI21_X1 U5845 ( .B1(n6831), .B2(n4763), .A(n4762), .ZN(n6910) );
  AOI21_X1 U5846 ( .B1(n4768), .B2(n4769), .A(n4767), .ZN(n4762) );
  INV_X1 U5847 ( .A(n4769), .ZN(n4763) );
  INV_X1 U5848 ( .A(n6832), .ZN(n4768) );
  NAND2_X1 U5849 ( .A1(n4754), .A2(n5637), .ZN(n8082) );
  NAND2_X1 U5850 ( .A1(n8072), .A2(n4759), .ZN(n4754) );
  NAND2_X1 U5851 ( .A1(n4966), .A2(n4968), .ZN(n7488) );
  NAND2_X1 U5852 ( .A1(n4969), .A2(n4968), .ZN(n7486) );
  NAND2_X1 U5853 ( .A1(n5702), .A2(n5703), .ZN(n4841) );
  NAND2_X1 U5854 ( .A1(n8126), .A2(n5716), .ZN(n4842) );
  AND2_X1 U5855 ( .A1(n5755), .A2(n5728), .ZN(n8450) );
  AND2_X1 U5856 ( .A1(n5866), .A2(n5870), .ZN(n8143) );
  NAND2_X1 U5857 ( .A1(n4958), .A2(n5355), .ZN(n7226) );
  AND2_X1 U5858 ( .A1(n8143), .A2(n9910), .ZN(n8192) );
  NAND2_X1 U5859 ( .A1(n8072), .A2(n5616), .ZN(n8149) );
  NAND2_X1 U5860 ( .A1(n7488), .A2(n5454), .ZN(n7573) );
  AND2_X1 U5861 ( .A1(n8143), .A2(n8596), .ZN(n8191) );
  NAND2_X1 U5862 ( .A1(n5739), .A2(n5738), .ZN(n8180) );
  AND2_X1 U5863 ( .A1(n5780), .A2(n5756), .ZN(n8433) );
  NAND2_X1 U5864 ( .A1(n5701), .A2(n5700), .ZN(n8474) );
  OR2_X1 U5865 ( .A1(n8465), .A2(n5782), .ZN(n5701) );
  OR2_X1 U5866 ( .A1(n8497), .A2(n5782), .ZN(n5672) );
  INV_X1 U5867 ( .A(n5885), .ZN(n8211) );
  NAND2_X1 U5868 ( .A1(n5729), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5183) );
  NAND4_X2 U5869 ( .A1(n5205), .A2(n5204), .A3(n5203), .A4(n5202), .ZN(n8218)
         );
  NAND2_X1 U5870 ( .A1(n5729), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5204) );
  AOI21_X1 U5871 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n6427), .A(n6423), .ZN(
        n6425) );
  INV_X1 U5872 ( .A(n4639), .ZN(n8310) );
  NAND2_X1 U5873 ( .A1(n8313), .A2(n5414), .ZN(n4638) );
  INV_X1 U5874 ( .A(n8330), .ZN(n4600) );
  XNOR2_X1 U5875 ( .A(n8350), .B(n8360), .ZN(n8344) );
  INV_X1 U5876 ( .A(n10194), .ZN(n8359) );
  NAND2_X1 U5877 ( .A1(n5929), .A2(n5928), .ZN(n8659) );
  OAI21_X1 U5878 ( .B1(n8385), .B2(n8384), .A(n8383), .ZN(n8664) );
  NAND2_X1 U5879 ( .A1(n5892), .A2(n6063), .ZN(n8411) );
  NAND2_X1 U5880 ( .A1(n4888), .A2(n4891), .ZN(n8403) );
  OR2_X1 U5881 ( .A1(n8463), .A2(n4892), .ZN(n4888) );
  OAI21_X1 U5882 ( .B1(n8463), .B2(n8019), .A(n8420), .ZN(n8422) );
  NAND2_X1 U5883 ( .A1(n5754), .A2(n5753), .ZN(n8680) );
  AND2_X1 U5884 ( .A1(n8461), .A2(n8460), .ZN(n8694) );
  NAND2_X1 U5885 ( .A1(n8483), .A2(n8482), .ZN(n8699) );
  NAND2_X1 U5886 ( .A1(n4709), .A2(n4710), .ZN(n8511) );
  OR2_X1 U5887 ( .A1(n8532), .A2(n4712), .ZN(n4709) );
  NAND2_X1 U5888 ( .A1(n4897), .A2(n8012), .ZN(n8555) );
  NAND2_X1 U5889 ( .A1(n8576), .A2(n4288), .ZN(n4897) );
  NAND2_X1 U5890 ( .A1(n5559), .A2(n5558), .ZN(n8731) );
  NAND2_X1 U5891 ( .A1(n8592), .A2(n6032), .ZN(n8574) );
  NAND2_X1 U5892 ( .A1(n4902), .A2(n7382), .ZN(n7436) );
  NAND2_X1 U5893 ( .A1(n7381), .A2(n4906), .ZN(n4902) );
  NAND2_X1 U5894 ( .A1(n4706), .A2(n6947), .ZN(n7376) );
  NAND2_X1 U5895 ( .A1(n7192), .A2(n7203), .ZN(n4706) );
  NAND2_X1 U5896 ( .A1(n6930), .A2(n9919), .ZN(n8606) );
  INV_X1 U5897 ( .A(n8629), .ZN(n9921) );
  OR2_X1 U5898 ( .A1(n6394), .A2(n6545), .ZN(n9919) );
  NAND2_X1 U5899 ( .A1(n8606), .A2(n6929), .ZN(n9925) );
  INV_X1 U5900 ( .A(n9925), .ZN(n8653) );
  NOR2_X1 U5901 ( .A1(n8686), .A2(n4661), .ZN(n8689) );
  NAND2_X1 U5902 ( .A1(n4663), .A2(n4662), .ZN(n4661) );
  NAND2_X1 U5903 ( .A1(n8688), .A2(n9956), .ZN(n4662) );
  OR2_X1 U5904 ( .A1(n8708), .A2(n8707), .ZN(n8778) );
  OR2_X1 U5905 ( .A1(n8719), .A2(n8718), .ZN(n8780) );
  INV_X1 U5906 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4909) );
  AND2_X1 U5907 ( .A1(n5829), .A2(n5828), .ZN(n8806) );
  XNOR2_X1 U5908 ( .A(n5814), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7603) );
  INV_X1 U5909 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6337) );
  INV_X1 U5910 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6295) );
  INV_X1 U5911 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10129) );
  INV_X1 U5912 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6221) );
  INV_X1 U5913 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10127) );
  MUX2_X1 U5914 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5191), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5193) );
  AND4_X1 U5915 ( .A1(n7017), .A2(n7016), .A3(n7015), .A4(n7014), .ZN(n7239)
         );
  AND4_X1 U5916 ( .A1(n7319), .A2(n7318), .A3(n7317), .A4(n7316), .ZN(n8834)
         );
  INV_X1 U5917 ( .A(n4720), .ZN(n7446) );
  AOI21_X1 U5918 ( .B1(n5058), .B2(n4721), .A(n4724), .ZN(n4720) );
  INV_X1 U5919 ( .A(n4725), .ZN(n4721) );
  NAND2_X1 U5920 ( .A1(n6628), .A2(n6514), .ZN(n6981) );
  NAND2_X1 U5921 ( .A1(n7913), .A2(n7916), .ZN(n8865) );
  AND2_X1 U5922 ( .A1(n7897), .A2(n8964), .ZN(n4645) );
  NAND2_X1 U5923 ( .A1(n5064), .A2(n7241), .ZN(n7264) );
  NAND2_X1 U5924 ( .A1(n7238), .A2(n7237), .ZN(n5064) );
  AND2_X1 U5925 ( .A1(n7647), .A2(n7646), .ZN(n9412) );
  AOI21_X1 U5926 ( .B1(n4493), .B2(n8959), .A(n7843), .ZN(n8880) );
  INV_X1 U5927 ( .A(n4729), .ZN(n4493) );
  OAI21_X1 U5928 ( .B1(n8823), .B2(n5071), .A(n5069), .ZN(n8903) );
  INV_X1 U5929 ( .A(n4718), .ZN(n5069) );
  NAND2_X1 U5930 ( .A1(n4486), .A2(n4489), .ZN(n4484) );
  NAND2_X1 U5931 ( .A1(n6628), .A2(n4487), .ZN(n4485) );
  INV_X1 U5932 ( .A(n6979), .ZN(n4489) );
  NAND2_X1 U5933 ( .A1(n5058), .A2(n5061), .ZN(n7346) );
  NAND2_X1 U5934 ( .A1(n7751), .A2(n7750), .ZN(n9648) );
  NAND2_X1 U5935 ( .A1(n5058), .A2(n4722), .ZN(n4648) );
  NAND2_X1 U5936 ( .A1(n5081), .A2(n7450), .ZN(n7456) );
  OAI21_X1 U5937 ( .B1(n5058), .B2(n4724), .A(n4722), .ZN(n5081) );
  INV_X1 U5938 ( .A(n8968), .ZN(n8984) );
  OR2_X1 U5939 ( .A1(n6531), .A2(n9056), .ZN(n8968) );
  NAND2_X1 U5940 ( .A1(n8804), .A2(n7087), .ZN(n7639) );
  NAND2_X1 U5941 ( .A1(n4499), .A2(n8976), .ZN(n4498) );
  NAND2_X1 U5942 ( .A1(n5088), .A2(n5087), .ZN(n4499) );
  AOI21_X1 U5943 ( .B1(n5088), .B2(n5086), .A(n8993), .ZN(n4500) );
  NAND2_X1 U5944 ( .A1(n6488), .A2(n6487), .ZN(n8991) );
  INV_X1 U5945 ( .A(n9412), .ZN(n9433) );
  INV_X1 U5946 ( .A(n7662), .ZN(n9575) );
  NAND2_X1 U5947 ( .A1(n4263), .A2(n6903), .ZN(n6517) );
  NOR2_X1 U5948 ( .A1(n6227), .A2(n6366), .ZN(n6226) );
  INV_X1 U5949 ( .A(n4537), .ZN(n6262) );
  NOR2_X1 U5950 ( .A1(n6260), .A2(n4328), .ZN(n6382) );
  NAND2_X1 U5951 ( .A1(n6382), .A2(n6381), .ZN(n6380) );
  OAI21_X1 U5952 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n6194), .A(n6380), .ZN(
        n6247) );
  AND2_X1 U5953 ( .A1(n6241), .A2(n6240), .ZN(n6274) );
  OAI21_X1 U5954 ( .B1(n6274), .B2(n6272), .A(n6273), .ZN(n6340) );
  NAND2_X1 U5955 ( .A1(n4880), .A2(n6344), .ZN(n9801) );
  NAND2_X1 U5956 ( .A1(n4879), .A2(n4881), .ZN(n6345) );
  NAND2_X1 U5957 ( .A1(n9794), .A2(n6344), .ZN(n4879) );
  OAI22_X1 U5958 ( .A1(n9806), .A2(n6574), .B1(n7154), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n6777) );
  AND2_X1 U5959 ( .A1(n7254), .A2(n7253), .ZN(n7256) );
  NAND2_X1 U5960 ( .A1(n4873), .A2(n4874), .ZN(n9292) );
  AOI22_X1 U5961 ( .A1(n7252), .A2(n7251), .B1(n7250), .B2(n7249), .ZN(n9287)
         );
  OAI21_X1 U5962 ( .B1(n9287), .B2(n9286), .A(n4406), .ZN(n9288) );
  OR2_X1 U5963 ( .A1(n9293), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4406) );
  XNOR2_X1 U5964 ( .A(n9317), .B(n9323), .ZN(n9309) );
  NOR2_X1 U5965 ( .A1(n9309), .A2(n9308), .ZN(n9318) );
  NOR2_X1 U5966 ( .A1(n9324), .A2(n9325), .ZN(n9327) );
  INV_X1 U5967 ( .A(n4409), .ZN(n9339) );
  INV_X1 U5968 ( .A(n4539), .ZN(n9349) );
  NAND2_X1 U5969 ( .A1(n7980), .A2(n7979), .ZN(n7998) );
  NAND2_X1 U5970 ( .A1(n4944), .A2(n7976), .ZN(n9427) );
  NAND2_X1 U5971 ( .A1(n9442), .A2(n9431), .ZN(n4944) );
  NAND2_X1 U5972 ( .A1(n4679), .A2(n4678), .ZN(n4677) );
  XNOR2_X1 U5973 ( .A(n9421), .B(n4681), .ZN(n4680) );
  NAND2_X1 U5974 ( .A1(n7972), .A2(n9574), .ZN(n4678) );
  OAI21_X1 U5975 ( .B1(n9461), .B2(n5104), .A(n5101), .ZN(n7982) );
  NAND2_X1 U5976 ( .A1(n4417), .A2(n4418), .ZN(n7967) );
  NAND2_X1 U5977 ( .A1(n4422), .A2(n7949), .ZN(n9457) );
  NAND2_X1 U5978 ( .A1(n4423), .A2(n4289), .ZN(n4422) );
  INV_X1 U5979 ( .A(n9470), .ZN(n4423) );
  NAND2_X1 U5980 ( .A1(n5105), .A2(n9155), .ZN(n9446) );
  OR2_X1 U5981 ( .A1(n9461), .A2(n9183), .ZN(n5105) );
  AND2_X1 U5982 ( .A1(n7948), .A2(n7947), .ZN(n9468) );
  NAND2_X1 U5983 ( .A1(n7944), .A2(n7941), .ZN(n9643) );
  NAND2_X1 U5984 ( .A1(n4561), .A2(n4562), .ZN(n9494) );
  NAND2_X1 U5985 ( .A1(n7939), .A2(n7938), .ZN(n9493) );
  AOI21_X1 U5986 ( .B1(n9523), .B2(n9535), .A(n7954), .ZN(n9510) );
  INV_X1 U5987 ( .A(n4947), .ZN(n4427) );
  AND2_X1 U5988 ( .A1(n4789), .A2(n4425), .ZN(n4424) );
  NAND2_X1 U5989 ( .A1(n4947), .A2(n4426), .ZN(n4425) );
  NAND2_X1 U5990 ( .A1(n4790), .A2(n7926), .ZN(n9536) );
  NAND2_X1 U5991 ( .A1(n7925), .A2(n4947), .ZN(n4790) );
  NAND2_X1 U5992 ( .A1(n7925), .A2(n7924), .ZN(n9547) );
  NAND2_X1 U5993 ( .A1(n9569), .A2(n9122), .ZN(n9551) );
  OAI21_X1 U5994 ( .B1(n7516), .B2(n4781), .A(n4779), .ZN(n9568) );
  NAND2_X1 U5995 ( .A1(n4784), .A2(n4950), .ZN(n7922) );
  NAND2_X1 U5996 ( .A1(n7516), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U5997 ( .A1(n7614), .A2(n9203), .ZN(n7613) );
  NAND2_X1 U5998 ( .A1(n6812), .A2(n9011), .ZN(n7075) );
  OR2_X1 U5999 ( .A1(n7324), .A2(n9869), .ZN(n7995) );
  INV_X1 U6000 ( .A(n9821), .ZN(n6642) );
  AND2_X1 U6001 ( .A1(n9589), .A2(n6447), .ZN(n9490) );
  INV_X1 U6002 ( .A(n7995), .ZN(n9581) );
  AND2_X2 U6003 ( .A1(n6606), .A2(n6605), .ZN(n9891) );
  OAI211_X1 U6004 ( .C1(n9697), .C2(n9610), .A(n9608), .B(n9609), .ZN(n9708)
         );
  AND2_X1 U6005 ( .A1(n6482), .A2(n6149), .ZN(n9816) );
  INV_X1 U6006 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6208) );
  OR2_X1 U6007 ( .A1(n6105), .A2(n9727), .ZN(n6098) );
  INV_X1 U6008 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6805) );
  INV_X1 U6009 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6352) );
  INV_X1 U6010 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10071) );
  INV_X1 U6011 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6293) );
  INV_X1 U6012 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6238) );
  INV_X1 U6013 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6219) );
  AND2_X1 U6014 ( .A1(n6166), .A2(n6301), .ZN(n9805) );
  NAND2_X1 U6015 ( .A1(n6176), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U6016 ( .A1(n6176), .A2(n6175), .ZN(n6503) );
  XNOR2_X1 U6017 ( .A(n10036), .B(n4535), .ZN(n7610) );
  OAI21_X1 U6018 ( .B1(n10005), .B2(n9754), .A(n10007), .ZN(n10218) );
  AND2_X1 U6019 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9761), .ZN(n10207) );
  NOR2_X1 U6020 ( .A1(n9771), .A2(n10215), .ZN(n10033) );
  NOR2_X1 U6021 ( .A1(n10028), .A2(n4376), .ZN(n10027) );
  NAND2_X1 U6022 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  OAI21_X1 U6023 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10025), .ZN(n10023) );
  NAND2_X1 U6024 ( .A1(n10023), .A2(n10024), .ZN(n10022) );
  NAND2_X1 U6025 ( .A1(n10022), .A2(n4593), .ZN(n10020) );
  NAND2_X1 U6026 ( .A1(n4594), .A2(n10162), .ZN(n4593) );
  INV_X1 U6027 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n4594) );
  OAI21_X1 U6028 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10019), .ZN(n10017) );
  NAND2_X1 U6029 ( .A1(n10017), .A2(n10018), .ZN(n10016) );
  NAND2_X1 U6030 ( .A1(n10016), .A2(n4595), .ZN(n10014) );
  NAND2_X1 U6031 ( .A1(n7220), .A2(n10098), .ZN(n4595) );
  XNOR2_X1 U6032 ( .A(n4404), .B(n8043), .ZN(n8048) );
  OR2_X1 U6033 ( .A1(n6087), .A2(n4660), .ZN(n4659) );
  AND2_X1 U6034 ( .A1(n6089), .A2(n6086), .ZN(n4502) );
  NAND2_X1 U6035 ( .A1(n4637), .A2(n4636), .ZN(P2_U3264) );
  AOI21_X1 U6036 ( .B1(n8372), .B2(n4954), .A(n8376), .ZN(n4636) );
  NAND2_X1 U6037 ( .A1(n8373), .A2(n8435), .ZN(n4637) );
  NAND2_X1 U6038 ( .A1(n10002), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U6039 ( .A1(n8771), .A2(n10004), .ZN(n4975) );
  NAND2_X1 U6040 ( .A1(n9992), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U6041 ( .A1(n8771), .A2(n9994), .ZN(n4691) );
  NAND2_X1 U6042 ( .A1(n4497), .A2(n4495), .ZN(P1_U3238) );
  NOR2_X1 U6043 ( .A1(n8977), .A2(n4496), .ZN(n4495) );
  NAND2_X1 U6044 ( .A1(n4500), .A2(n4498), .ZN(n4497) );
  AND2_X1 U6045 ( .A1(n9616), .A2(n8978), .ZN(n4496) );
  AOI21_X1 U6046 ( .B1(n4453), .B2(n4451), .A(n4666), .ZN(P1_U3240) );
  AOI21_X1 U6047 ( .B1(n9229), .B2(n9228), .A(n4452), .ZN(n4451) );
  NAND2_X1 U6048 ( .A1(n4454), .A2(n4259), .ZN(n4453) );
  AOI21_X1 U6049 ( .B1(n9375), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9374), .ZN(
        n4882) );
  INV_X1 U6050 ( .A(n4652), .ZN(n9418) );
  OAI21_X1 U6051 ( .B1(n9614), .B2(n9566), .A(n4653), .ZN(n4652) );
  AOI21_X1 U6052 ( .B1(n9611), .B2(n9564), .A(n9417), .ZN(n4653) );
  INV_X1 U6053 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4632) );
  OAI21_X1 U6054 ( .B1(n8001), .B2(n4261), .A(n4945), .ZN(P1_U3323) );
  INV_X1 U6055 ( .A(n4946), .ZN(n4945) );
  OAI21_X1 U6056 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9775), .A(n10211), .ZN(
        n9777) );
  INV_X1 U6057 ( .A(n7241), .ZN(n5062) );
  AND2_X1 U6058 ( .A1(n8452), .A2(n4978), .ZN(n4266) );
  OR2_X1 U6059 ( .A1(n8023), .A2(n8426), .ZN(n4267) );
  XNOR2_X1 U6060 ( .A(n5501), .B(SI_14_), .ZN(n5498) );
  AND2_X1 U6061 ( .A1(n4912), .A2(n4911), .ZN(n4268) );
  INV_X1 U6062 ( .A(n5705), .ZN(n4960) );
  AND2_X1 U6063 ( .A1(n4710), .A2(n4329), .ZN(n4269) );
  AND2_X1 U6064 ( .A1(n8623), .A2(n8614), .ZN(n4270) );
  INV_X1 U6065 ( .A(n9155), .ZN(n5103) );
  INV_X1 U6066 ( .A(n4943), .ZN(n4942) );
  NAND2_X1 U6067 ( .A1(n4340), .A2(n7976), .ZN(n4943) );
  AND2_X1 U6068 ( .A1(n6948), .A2(n4983), .ZN(n4272) );
  INV_X1 U6069 ( .A(n9431), .ZN(n4941) );
  NAND2_X1 U6070 ( .A1(n5577), .A2(n5576), .ZN(n8725) );
  INV_X1 U6071 ( .A(n8725), .ZN(n5013) );
  AND2_X1 U6072 ( .A1(n5766), .A2(n5765), .ZN(n4273) );
  XNOR2_X1 U6073 ( .A(n7981), .B(n9061), .ZN(n9602) );
  NOR2_X1 U6074 ( .A1(n9187), .A2(n9091), .ZN(n4274) );
  AND2_X1 U6075 ( .A1(n4915), .A2(n4913), .ZN(n4275) );
  AND2_X1 U6076 ( .A1(n4986), .A2(n4985), .ZN(n4276) );
  NOR2_X1 U6077 ( .A1(n6037), .A2(n6047), .ZN(n4277) );
  AND2_X1 U6078 ( .A1(n6034), .A2(n8575), .ZN(n4278) );
  AND2_X1 U6079 ( .A1(n8409), .A2(n4266), .ZN(n4279) );
  AND2_X1 U6080 ( .A1(n4268), .A2(n4910), .ZN(n4280) );
  NAND2_X1 U6081 ( .A1(n4890), .A2(n6065), .ZN(n4804) );
  INV_X1 U6082 ( .A(n4804), .ZN(n4650) );
  NAND2_X1 U6083 ( .A1(n5093), .A2(n9170), .ZN(n4281) );
  INV_X1 U6084 ( .A(n7377), .ZN(n4907) );
  AND2_X2 U6085 ( .A1(n5137), .A2(n4347), .ZN(n4282) );
  AND2_X1 U6086 ( .A1(n9227), .A2(n4259), .ZN(n9170) );
  NAND2_X1 U6087 ( .A1(n4674), .A2(n7089), .ZN(n9867) );
  NAND2_X1 U6088 ( .A1(n4483), .A2(n7658), .ZN(n8823) );
  NAND2_X1 U6089 ( .A1(n7880), .A2(n7879), .ZN(n9606) );
  INV_X1 U6090 ( .A(n4264), .ZN(n7868) );
  AND2_X1 U6091 ( .A1(n7329), .A2(n4933), .ZN(n4283) );
  NAND2_X1 U6092 ( .A1(n7584), .A2(n7583), .ZN(n9678) );
  INV_X1 U6093 ( .A(n4737), .ZN(n9827) );
  NAND2_X1 U6094 ( .A1(n6523), .A2(n4447), .ZN(n4737) );
  NAND2_X1 U6095 ( .A1(n7681), .A2(n7680), .ZN(n9672) );
  XNOR2_X1 U6096 ( .A(n4415), .B(n6140), .ZN(n6521) );
  AND2_X1 U6097 ( .A1(n4639), .A2(n4638), .ZN(n4284) );
  AND2_X1 U6098 ( .A1(n5673), .A2(n8161), .ZN(n4285) );
  AND2_X1 U6099 ( .A1(n5358), .A2(n5332), .ZN(n4286) );
  AND2_X1 U6100 ( .A1(n5124), .A2(n5407), .ZN(n4287) );
  AND2_X1 U6101 ( .A1(n8561), .A2(n8559), .ZN(n4288) );
  INV_X1 U6102 ( .A(n5504), .ZN(n6455) );
  CLKBUF_X3 U6103 ( .A(n5504), .Z(n5808) );
  NAND2_X1 U6104 ( .A1(n9636), .A2(n9447), .ZN(n4289) );
  INV_X1 U6105 ( .A(n9130), .ZN(n4555) );
  INV_X1 U6106 ( .A(n5679), .ZN(n4749) );
  AND2_X1 U6107 ( .A1(n4972), .A2(n7404), .ZN(n4971) );
  NAND2_X1 U6108 ( .A1(n8420), .A2(n8022), .ZN(n4290) );
  NAND2_X1 U6109 ( .A1(n5779), .A2(n5778), .ZN(n8675) );
  AND2_X1 U6110 ( .A1(n7154), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4291) );
  INV_X1 U6111 ( .A(n9561), .ZN(n4426) );
  AND2_X1 U6112 ( .A1(n5086), .A2(n4730), .ZN(n4292) );
  NAND2_X1 U6113 ( .A1(n5479), .A2(n5478), .ZN(n4293) );
  AND2_X1 U6114 ( .A1(n6731), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4294) );
  NAND2_X1 U6115 ( .A1(n5467), .A2(n5466), .ZN(n8652) );
  INV_X1 U6116 ( .A(n9159), .ZN(n5098) );
  AND2_X1 U6117 ( .A1(n6733), .A2(n6732), .ZN(n9845) );
  INV_X1 U6118 ( .A(n9156), .ZN(n5102) );
  NAND2_X1 U6119 ( .A1(n5235), .A2(n4300), .ZN(n4295) );
  AND4_X1 U6120 ( .A1(n5266), .A2(n5136), .A3(n4977), .A4(
        P2_IR_REG_27__SCAN_IN), .ZN(n4296) );
  AND2_X1 U6121 ( .A1(n5853), .A2(n8202), .ZN(n4297) );
  INV_X1 U6122 ( .A(n9135), .ZN(n4563) );
  INV_X1 U6123 ( .A(n6165), .ZN(n5115) );
  INV_X1 U6124 ( .A(n9011), .ZN(n5113) );
  AND2_X1 U6125 ( .A1(n8100), .A2(n5544), .ZN(n4298) );
  AND2_X1 U6126 ( .A1(n8714), .A2(n8535), .ZN(n4299) );
  NAND2_X1 U6127 ( .A1(n5283), .A2(SI_5_), .ZN(n5284) );
  INV_X1 U6128 ( .A(n5284), .ZN(n4998) );
  INV_X1 U6129 ( .A(n9249), .ZN(n5122) );
  AND2_X1 U6130 ( .A1(n5269), .A2(n9909), .ZN(n4300) );
  AND2_X1 U6131 ( .A1(n9159), .A2(n5102), .ZN(n4301) );
  AND4_X1 U6132 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n9079)
         );
  INV_X1 U6133 ( .A(n9079), .ZN(n4928) );
  AND2_X1 U6134 ( .A1(n5995), .A2(n6079), .ZN(n4302) );
  AND2_X1 U6135 ( .A1(n9648), .A2(n9511), .ZN(n4303) );
  OR2_X1 U6136 ( .A1(n6957), .A2(n6070), .ZN(n4304) );
  AOI21_X1 U6137 ( .B1(n4725), .B2(n7344), .A(n4723), .ZN(n4722) );
  NOR2_X1 U6138 ( .A1(n9318), .A2(n9319), .ZN(n4305) );
  NAND2_X1 U6139 ( .A1(n7639), .A2(n7638), .ZN(n9616) );
  INV_X1 U6140 ( .A(n9616), .ZN(n4925) );
  NOR2_X1 U6141 ( .A1(n9631), .A2(n9462), .ZN(n4306) );
  NOR2_X1 U6142 ( .A1(n9678), .A2(n9575), .ZN(n4307) );
  INV_X1 U6143 ( .A(n7430), .ZN(n8003) );
  AND2_X1 U6144 ( .A1(n5423), .A2(n5422), .ZN(n4308) );
  NAND2_X1 U6145 ( .A1(n8666), .A2(n6068), .ZN(n5954) );
  INV_X1 U6146 ( .A(n5954), .ZN(n5029) );
  NAND2_X1 U6147 ( .A1(n5602), .A2(n5601), .ZN(n8721) );
  NAND2_X1 U6148 ( .A1(n5514), .A2(n5513), .ZN(n8608) );
  AND2_X1 U6149 ( .A1(n6038), .A2(n6049), .ZN(n4309) );
  INV_X1 U6150 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4956) );
  INV_X1 U6151 ( .A(n5017), .ZN(n5016) );
  NOR2_X1 U6152 ( .A1(n5456), .A2(n5018), .ZN(n5017) );
  INV_X1 U6153 ( .A(n4865), .ZN(n4864) );
  NOR2_X1 U6154 ( .A1(n5523), .A2(n4866), .ZN(n4865) );
  AND2_X1 U6155 ( .A1(n4428), .A2(n9475), .ZN(n4310) );
  AND2_X1 U6156 ( .A1(n5057), .A2(n6021), .ZN(n4311) );
  INV_X1 U6157 ( .A(n7455), .ZN(n7466) );
  NAND2_X1 U6158 ( .A1(n7288), .A2(n7287), .ZN(n7455) );
  AND2_X1 U6159 ( .A1(n5936), .A2(n5935), .ZN(n4312) );
  NOR2_X1 U6160 ( .A1(n4306), .A2(n4421), .ZN(n4420) );
  AND2_X1 U6161 ( .A1(n8138), .A2(n4295), .ZN(n4313) );
  INV_X1 U6162 ( .A(n6009), .ZN(n4833) );
  OR2_X1 U6163 ( .A1(n8764), .A2(n6912), .ZN(n6009) );
  AND2_X1 U6164 ( .A1(n7458), .A2(n7450), .ZN(n4314) );
  NAND2_X1 U6165 ( .A1(n9110), .A2(n9102), .ZN(n4315) );
  AND2_X1 U6166 ( .A1(n4794), .A2(n8003), .ZN(n4316) );
  AND2_X1 U6167 ( .A1(n9631), .A2(n9462), .ZN(n4317) );
  NAND2_X1 U6168 ( .A1(n8027), .A2(n6074), .ZN(n4318) );
  NAND2_X1 U6169 ( .A1(n8594), .A2(n6031), .ZN(n4319) );
  AND2_X1 U6170 ( .A1(n6039), .A2(n6079), .ZN(n4320) );
  OR2_X1 U6171 ( .A1(n5063), .A2(n5060), .ZN(n5059) );
  INV_X1 U6172 ( .A(n5429), .ZN(n5018) );
  NAND2_X1 U6173 ( .A1(n5428), .A2(SI_11_), .ZN(n5429) );
  INV_X1 U6174 ( .A(n7843), .ZN(n4730) );
  INV_X1 U6175 ( .A(n4856), .ZN(n4855) );
  NAND2_X1 U6176 ( .A1(n4857), .A2(n8043), .ZN(n4856) );
  OR2_X1 U6177 ( .A1(n8680), .A2(n8412), .ZN(n6064) );
  INV_X1 U6178 ( .A(n6064), .ZN(n4803) );
  AND2_X1 U6179 ( .A1(n9015), .A2(n9095), .ZN(n9199) );
  NOR2_X1 U6180 ( .A1(n7378), .A2(n8212), .ZN(n4321) );
  NOR2_X1 U6181 ( .A1(n8834), .A2(n7875), .ZN(n4322) );
  NOR2_X1 U6182 ( .A1(n8709), .A2(n8520), .ZN(n4323) );
  NOR2_X1 U6183 ( .A1(n8725), .A2(n8563), .ZN(n4324) );
  NOR2_X1 U6184 ( .A1(n9805), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4325) );
  NOR2_X1 U6185 ( .A1(n9612), .A2(n9422), .ZN(n4326) );
  INV_X1 U6186 ( .A(n5106), .ZN(n5104) );
  AND2_X1 U6187 ( .A1(n9157), .A2(n5107), .ZN(n5106) );
  AND2_X1 U6188 ( .A1(n9678), .A2(n9575), .ZN(n4327) );
  AND2_X1 U6189 ( .A1(n9628), .A2(n8849), .ZN(n9068) );
  AND2_X1 U6190 ( .A1(n6193), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4328) );
  INV_X1 U6191 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5394) );
  INV_X1 U6192 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5346) );
  INV_X1 U6193 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7095) );
  NAND2_X1 U6194 ( .A1(n8709), .A2(n8520), .ZN(n4329) );
  INV_X1 U6195 ( .A(n4981), .ZN(n4980) );
  NAND2_X1 U6196 ( .A1(n4272), .A2(n4982), .ZN(n4981) );
  AND2_X1 U6197 ( .A1(n9663), .A2(n9553), .ZN(n4330) );
  NOR2_X1 U6198 ( .A1(n7474), .A2(n7495), .ZN(n4331) );
  NOR2_X1 U6199 ( .A1(n9091), .A2(n8998), .ZN(n4332) );
  INV_X1 U6200 ( .A(n5939), .ZN(n4689) );
  AND2_X1 U6201 ( .A1(n6941), .A2(n7054), .ZN(n4333) );
  AND2_X1 U6202 ( .A1(n6032), .A2(n6033), .ZN(n8594) );
  NAND2_X1 U6203 ( .A1(n5958), .A2(n5955), .ZN(n8410) );
  INV_X1 U6204 ( .A(n8410), .ZN(n4890) );
  OR2_X1 U6205 ( .A1(n9559), .A2(n9573), .ZN(n7953) );
  INV_X1 U6206 ( .A(n5455), .ZN(n5015) );
  OR2_X1 U6207 ( .A1(n4507), .A2(n4503), .ZN(n4334) );
  NAND2_X1 U6208 ( .A1(n6063), .A2(n6059), .ZN(n4335) );
  NAND2_X1 U6209 ( .A1(n5079), .A2(n5077), .ZN(n4336) );
  OR2_X1 U6210 ( .A1(n4285), .A2(n4960), .ZN(n4337) );
  AND2_X1 U6211 ( .A1(n5480), .A2(n5497), .ZN(n4338) );
  AND2_X1 U6212 ( .A1(n9123), .A2(n9122), .ZN(n9571) );
  AND2_X1 U6213 ( .A1(n9616), .A2(n9433), .ZN(n4339) );
  OR2_X1 U6214 ( .A1(n9616), .A2(n9433), .ZN(n4340) );
  AND2_X1 U6215 ( .A1(n5790), .A2(n5789), .ZN(n4341) );
  AND2_X1 U6216 ( .A1(n7860), .A2(n7861), .ZN(n4342) );
  AND2_X1 U6217 ( .A1(n7714), .A2(n7713), .ZN(n4343) );
  OAI21_X1 U6218 ( .B1(n7939), .B2(n4432), .A(n4430), .ZN(n9474) );
  INV_X1 U6219 ( .A(n4963), .ZN(n4962) );
  NAND2_X1 U6220 ( .A1(n8051), .A2(n4293), .ZN(n4963) );
  INV_X1 U6221 ( .A(n5424), .ZN(n5425) );
  AND4_X1 U6222 ( .A1(n7305), .A2(n7304), .A3(n7303), .A4(n7302), .ZN(n8951)
         );
  NAND2_X1 U6223 ( .A1(n7437), .A2(n8208), .ZN(n4344) );
  AND2_X1 U6224 ( .A1(n5306), .A2(n4998), .ZN(n4345) );
  INV_X1 U6225 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5168) );
  OR2_X1 U6226 ( .A1(n8735), .A2(n8119), .ZN(n5965) );
  INV_X1 U6227 ( .A(n5965), .ZN(n5042) );
  AND3_X1 U6228 ( .A1(n6124), .A2(n6207), .A3(n6208), .ZN(n4346) );
  AND3_X1 U6229 ( .A1(n5153), .A2(n5152), .A3(n5151), .ZN(n4347) );
  AND2_X1 U6230 ( .A1(n7853), .A2(n7852), .ZN(n8921) );
  AND3_X1 U6231 ( .A1(n5351), .A2(n5349), .A3(n4393), .ZN(n4348) );
  AND2_X1 U6232 ( .A1(n7783), .A2(n7782), .ZN(n9500) );
  XNOR2_X1 U6233 ( .A(n5307), .B(SI_6_), .ZN(n5306) );
  AND2_X1 U6234 ( .A1(n8549), .A2(n4991), .ZN(n4349) );
  AND2_X1 U6235 ( .A1(n6074), .A2(n5956), .ZN(n8396) );
  INV_X1 U6236 ( .A(n8396), .ZN(n4825) );
  NOR2_X1 U6237 ( .A1(n9672), .A2(n9552), .ZN(n4350) );
  AND2_X1 U6238 ( .A1(n5974), .A2(n5977), .ZN(n4351) );
  AND2_X1 U6239 ( .A1(n9219), .A2(n9253), .ZN(n4352) );
  AND2_X1 U6240 ( .A1(n6124), .A2(n6207), .ZN(n4353) );
  AND2_X1 U6241 ( .A1(n9426), .A2(n9161), .ZN(n4354) );
  NOR2_X1 U6242 ( .A1(n4907), .A2(n4705), .ZN(n4704) );
  INV_X1 U6243 ( .A(n5327), .ZN(n4767) );
  AND2_X1 U6244 ( .A1(n6377), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4355) );
  AND2_X1 U6245 ( .A1(n4647), .A2(n4646), .ZN(n4356) );
  INV_X1 U6246 ( .A(n9399), .ZN(n9388) );
  NAND2_X1 U6247 ( .A1(n9064), .A2(n9062), .ZN(n9399) );
  INV_X1 U6248 ( .A(n5936), .ZN(n6077) );
  OR2_X1 U6249 ( .A1(n9678), .A2(n7662), .ZN(n9021) );
  AND2_X1 U6250 ( .A1(n4719), .A2(n4314), .ZN(n4357) );
  NAND2_X1 U6251 ( .A1(n8893), .A2(n8892), .ZN(n4358) );
  INV_X1 U6252 ( .A(n6063), .ZN(n5035) );
  INV_X1 U6253 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n10051) );
  INV_X1 U6254 ( .A(n4494), .ZN(n8958) );
  OR2_X1 U6255 ( .A1(n7806), .A2(n7805), .ZN(n4494) );
  AND2_X1 U6256 ( .A1(n5053), .A2(n4909), .ZN(n4359) );
  INV_X1 U6257 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4839) );
  INV_X1 U6258 ( .A(n7382), .ZN(n4905) );
  INV_X1 U6259 ( .A(n4853), .ZN(n4852) );
  NAND2_X1 U6260 ( .A1(n4854), .A2(n5856), .ZN(n4853) );
  INV_X2 U6261 ( .A(n8606), .ZN(n8651) );
  INV_X1 U6262 ( .A(n5217), .ZN(n5216) );
  NOR2_X1 U6263 ( .A1(n6823), .A2(n4770), .ZN(n4769) );
  NAND2_X1 U6264 ( .A1(n5881), .A2(n5986), .ZN(n6954) );
  INV_X1 U6265 ( .A(n10004), .ZN(n10002) );
  OAI21_X1 U6266 ( .B1(n9560), .B2(n4427), .A(n4424), .ZN(n9534) );
  AND2_X1 U6267 ( .A1(n6949), .A2(n6948), .ZN(n4360) );
  AND2_X1 U6268 ( .A1(n8034), .A2(n4988), .ZN(n4361) );
  NAND2_X1 U6269 ( .A1(n7962), .A2(n7554), .ZN(n6088) );
  INV_X1 U6270 ( .A(n6088), .ZN(n4955) );
  NAND2_X1 U6271 ( .A1(n4669), .A2(n7923), .ZN(n9560) );
  NAND2_X1 U6272 ( .A1(n4693), .A2(n4282), .ZN(n5828) );
  OR2_X1 U6273 ( .A1(n9694), .A2(n7364), .ZN(n9101) );
  INV_X1 U6274 ( .A(n9101), .ZN(n5093) );
  NOR2_X1 U6275 ( .A1(n5741), .A2(n5747), .ZN(n4362) );
  NOR2_X1 U6276 ( .A1(n7255), .A2(n7135), .ZN(n4363) );
  XNOR2_X1 U6277 ( .A(n6098), .B(n10084), .ZN(n6150) );
  NAND2_X1 U6278 ( .A1(n6949), .A2(n4980), .ZN(n4984) );
  NAND2_X1 U6279 ( .A1(n9293), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4364) );
  AND2_X1 U6280 ( .A1(n4874), .A2(n4364), .ZN(n4365) );
  AND2_X1 U6281 ( .A1(n4958), .A2(n4957), .ZN(n4366) );
  INV_X1 U6282 ( .A(n4917), .ZN(n9513) );
  NOR2_X1 U6283 ( .A1(n5125), .A2(n4919), .ZN(n4917) );
  NAND2_X1 U6284 ( .A1(n5145), .A2(n5138), .ZN(n5816) );
  INV_X1 U6285 ( .A(n4932), .ZN(n7357) );
  OR2_X1 U6286 ( .A1(n5064), .A2(n7241), .ZN(n4367) );
  AND2_X2 U6287 ( .A1(n7146), .A2(n7145), .ZN(n9994) );
  INV_X1 U6288 ( .A(n7471), .ZN(n4983) );
  INV_X1 U6289 ( .A(n9799), .ZN(n4531) );
  AND3_X1 U6290 ( .A1(n6592), .A2(n6591), .A3(n6590), .ZN(n6586) );
  NAND2_X1 U6291 ( .A1(n7513), .A2(n7512), .ZN(n9682) );
  INV_X1 U6292 ( .A(n9682), .ZN(n4910) );
  NAND2_X1 U6293 ( .A1(n5537), .A2(n5536), .ZN(n8735) );
  INV_X1 U6294 ( .A(n8735), .ZN(n4985) );
  NAND2_X1 U6295 ( .A1(n5366), .A2(n5365), .ZN(n8764) );
  INV_X1 U6296 ( .A(n8764), .ZN(n4982) );
  AND2_X1 U6297 ( .A1(n9601), .A2(n9839), .ZN(n9697) );
  OR2_X1 U6298 ( .A1(n9367), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4368) );
  INV_X1 U6299 ( .A(n9283), .ZN(n4736) );
  NAND2_X1 U6300 ( .A1(n7322), .A2(n7321), .ZN(n9688) );
  INV_X1 U6301 ( .A(n9688), .ZN(n4911) );
  OR2_X1 U6302 ( .A1(n9876), .A2(n4632), .ZN(n4369) );
  INV_X1 U6303 ( .A(n9867), .ZN(n4913) );
  OR2_X1 U6304 ( .A1(n6901), .A2(n9833), .ZN(n6818) );
  INV_X1 U6305 ( .A(n6818), .ZN(n4914) );
  NAND2_X1 U6306 ( .A1(n4444), .A2(n7109), .ZN(n7110) );
  AND2_X1 U6307 ( .A1(n5920), .A2(n5919), .ZN(n4370) );
  AND2_X1 U6308 ( .A1(n9266), .A2(n9263), .ZN(n4371) );
  AND2_X1 U6309 ( .A1(n4879), .A2(n4877), .ZN(n4372) );
  OR2_X1 U6310 ( .A1(n6895), .A2(n6894), .ZN(n4373) );
  OR2_X1 U6311 ( .A1(n9891), .A2(n7634), .ZN(n4374) );
  NAND2_X1 U6312 ( .A1(n8377), .A2(n5972), .ZN(n4375) );
  INV_X1 U6313 ( .A(n6520), .ZN(n4449) );
  XNOR2_X1 U6314 ( .A(n5139), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8435) );
  NAND4_X1 U6315 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n9284)
         );
  INV_X1 U6316 ( .A(n9284), .ZN(n4731) );
  AND2_X1 U6317 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4376) );
  AND2_X1 U6318 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n4377) );
  INV_X1 U6319 ( .A(n7278), .ZN(n6553) );
  INV_X1 U6320 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4619) );
  INV_X1 U6321 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4676) );
  INV_X1 U6322 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4629) );
  INV_X1 U6323 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5005) );
  INV_X1 U6324 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U6325 ( .A1(n5982), .A2(n6070), .ZN(n4812) );
  NAND2_X1 U6326 ( .A1(n4351), .A2(n6070), .ZN(n4517) );
  OAI211_X1 U6327 ( .C1(n5980), .C2(n6070), .A(n5983), .B(n4517), .ZN(n4516)
         );
  INV_X1 U6328 ( .A(n6070), .ZN(n6079) );
  OR3_X2 U6329 ( .A1(n6554), .A2(n7554), .A3(n4954), .ZN(n6070) );
  OAI21_X2 U6330 ( .B1(n5066), .B2(n7693), .A(n8902), .ZN(n5068) );
  NAND2_X1 U6331 ( .A1(n7690), .A2(n7689), .ZN(n4383) );
  NAND3_X1 U6332 ( .A1(n4716), .A2(n4386), .A3(n7732), .ZN(n7912) );
  OR2_X2 U6333 ( .A1(n8962), .A2(n8960), .ZN(n8959) );
  NAND3_X1 U6334 ( .A1(n4901), .A2(n4344), .A3(n4395), .ZN(n8004) );
  OR2_X1 U6335 ( .A1(n4904), .A2(n7382), .ZN(n4395) );
  INV_X1 U6336 ( .A(n4904), .ZN(n4903) );
  NAND3_X1 U6337 ( .A1(n4693), .A2(n4282), .A3(n4359), .ZN(n8790) );
  AND3_X2 U6338 ( .A1(n5266), .A2(n5136), .A3(n4977), .ZN(n4693) );
  AOI21_X1 U6339 ( .B1(n4996), .B2(n4439), .A(n4345), .ZN(n4433) );
  NAND2_X1 U6340 ( .A1(n4435), .A2(n5306), .ZN(n4434) );
  INV_X1 U6341 ( .A(n4996), .ZN(n4435) );
  INV_X2 U6342 ( .A(n7678), .ZN(n4438) );
  NOR2_X1 U6343 ( .A1(n5306), .A2(n4998), .ZN(n4439) );
  NAND2_X1 U6344 ( .A1(n7074), .A2(n7073), .ZN(n7107) );
  NAND2_X1 U6345 ( .A1(n4445), .A2(n9398), .ZN(n9610) );
  INV_X2 U6346 ( .A(n6519), .ZN(n7087) );
  NAND2_X1 U6347 ( .A1(n9009), .A2(n9230), .ZN(n4450) );
  NAND2_X1 U6348 ( .A1(n6894), .A2(n4450), .ZN(n6765) );
  AND2_X1 U6349 ( .A1(n4450), .A2(n9189), .ZN(n5123) );
  XNOR2_X1 U6350 ( .A(n4373), .B(n9190), .ZN(n6900) );
  NAND2_X1 U6351 ( .A1(n4739), .A2(n4455), .ZN(n4458) );
  NAND3_X1 U6352 ( .A1(n9100), .A2(n9170), .A3(n9099), .ZN(n4457) );
  NAND2_X1 U6353 ( .A1(n4468), .A2(n4354), .ZN(n9167) );
  NAND2_X1 U6354 ( .A1(n4474), .A2(n4469), .ZN(n4468) );
  AOI22_X1 U6355 ( .A1(n4473), .A2(n4470), .B1(n9147), .B2(n9177), .ZN(n4469)
         );
  NAND3_X1 U6356 ( .A1(n9456), .A2(n9159), .A3(n4472), .ZN(n4471) );
  NAND2_X1 U6357 ( .A1(n9155), .A2(n9170), .ZN(n4472) );
  NAND3_X1 U6358 ( .A1(n9154), .A2(n9153), .A3(n9177), .ZN(n4473) );
  NAND2_X1 U6359 ( .A1(n6641), .A2(n6509), .ZN(n6628) );
  NAND2_X1 U6360 ( .A1(n4485), .A2(n4484), .ZN(n8927) );
  NAND3_X1 U6361 ( .A1(n4659), .A2(n4649), .A3(n4502), .ZN(P2_U3244) );
  NAND3_X1 U6362 ( .A1(n6042), .A2(n4510), .A3(n6044), .ZN(n4509) );
  INV_X1 U6363 ( .A(n6037), .ZN(n4510) );
  NAND2_X1 U6364 ( .A1(n4511), .A2(n6053), .ZN(n4999) );
  NAND3_X1 U6365 ( .A1(n4532), .A2(n4882), .A3(n4528), .ZN(P1_U3260) );
  NAND2_X1 U6366 ( .A1(n4529), .A2(n9261), .ZN(n4528) );
  NAND2_X1 U6367 ( .A1(n9373), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U6368 ( .A1(n4533), .A2(n4259), .ZN(n4532) );
  NAND2_X1 U6369 ( .A1(n9371), .A2(n4534), .ZN(n4533) );
  XNOR2_X1 U6370 ( .A(n7610), .B(n4869), .ZN(n6227) );
  INV_X1 U6371 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4535) );
  AND2_X1 U6372 ( .A1(n4537), .A2(n4536), .ZN(n6260) );
  OR2_X1 U6373 ( .A1(n6372), .A2(n4355), .ZN(n4537) );
  INV_X1 U6374 ( .A(n5308), .ZN(n4545) );
  NAND2_X1 U6375 ( .A1(n4546), .A2(n5308), .ZN(n5330) );
  NAND2_X1 U6376 ( .A1(n4547), .A2(n4997), .ZN(n4546) );
  AND2_X2 U6377 ( .A1(n4552), .A2(n4550), .ZN(n9540) );
  NOR2_X1 U6378 ( .A1(n4551), .A2(n9129), .ZN(n4550) );
  NAND3_X1 U6379 ( .A1(n9571), .A2(n4553), .A3(n4554), .ZN(n4552) );
  AND2_X1 U6380 ( .A1(n4556), .A2(n4554), .ZN(n9570) );
  OAI21_X2 U6381 ( .B1(n9523), .B2(n4560), .A(n4557), .ZN(n9479) );
  AOI21_X1 U6382 ( .B1(n4562), .B2(n4559), .A(n4558), .ZN(n4557) );
  INV_X1 U6383 ( .A(n4564), .ZN(n4559) );
  INV_X1 U6384 ( .A(n4562), .ZN(n4560) );
  NAND2_X1 U6385 ( .A1(n9523), .A2(n4564), .ZN(n4561) );
  NAND2_X1 U6386 ( .A1(n5406), .A2(n5405), .ZN(n4572) );
  NAND2_X1 U6387 ( .A1(n7983), .A2(n9162), .ZN(n9411) );
  XNOR2_X1 U6388 ( .A(n4994), .B(n4574), .ZN(n6734) );
  NAND2_X1 U6389 ( .A1(n5242), .A2(n5241), .ZN(n4574) );
  NAND2_X1 U6390 ( .A1(n5770), .A2(n5769), .ZN(n5772) );
  NAND2_X1 U6391 ( .A1(n5690), .A2(n5689), .ZN(n4588) );
  NAND2_X1 U6392 ( .A1(n5772), .A2(n5771), .ZN(n5805) );
  NAND2_X1 U6393 ( .A1(n5899), .A2(n5898), .ZN(n5905) );
  OAI21_X1 U6394 ( .B1(n5682), .B2(n5681), .A(n5680), .ZN(n5690) );
  NAND2_X1 U6395 ( .A1(n5504), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4675) );
  NAND2_X1 U6396 ( .A1(n10210), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n4591) );
  NAND2_X1 U6397 ( .A1(n10221), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n4592) );
  NOR2_X1 U6398 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10207), .ZN(n9762) );
  NAND2_X1 U6399 ( .A1(n5239), .A2(n5238), .ZN(n5242) );
  NAND2_X1 U6400 ( .A1(n7977), .A2(n9399), .ZN(n9398) );
  INV_X1 U6401 ( .A(n9602), .ZN(n4616) );
  NAND2_X1 U6402 ( .A1(n4788), .A2(n4615), .ZN(n9707) );
  NAND2_X1 U6403 ( .A1(n7514), .A2(n9186), .ZN(n7516) );
  NAND2_X1 U6404 ( .A1(n4823), .A2(n4318), .ZN(n4822) );
  NAND2_X1 U6405 ( .A1(n4736), .A2(n4737), .ZN(n9230) );
  NAND2_X1 U6406 ( .A1(n4930), .A2(n4929), .ZN(n7514) );
  AOI21_X1 U6407 ( .B1(n6807), .B2(n6810), .A(n6766), .ZN(n6767) );
  NAND2_X1 U6408 ( .A1(n4598), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4597) );
  NAND2_X1 U6409 ( .A1(n8106), .A2(n5552), .ZN(n8117) );
  NAND2_X1 U6410 ( .A1(n8124), .A2(n5704), .ZN(n4844) );
  INV_X1 U6411 ( .A(n5050), .ZN(n5049) );
  NAND2_X1 U6412 ( .A1(n4596), .A2(n5224), .ZN(n5238) );
  NAND2_X1 U6413 ( .A1(n5222), .A2(n5221), .ZN(n4596) );
  NAND2_X1 U6414 ( .A1(n5807), .A2(n5806), .ZN(n5895) );
  NAND2_X1 U6415 ( .A1(n5641), .A2(n5640), .ZN(n5654) );
  NOR2_X1 U6416 ( .A1(n5009), .A2(n5007), .ZN(n5006) );
  AOI21_X1 U6417 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6193), .A(n6254), .ZN(
        n6385) );
  OAI22_X1 U6418 ( .A1(n7130), .A2(n7129), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n7286), .ZN(n7252) );
  AOI21_X1 U6419 ( .B1(n9355), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9354), .ZN(
        n9356) );
  XNOR2_X1 U6420 ( .A(n5240), .B(SI_3_), .ZN(n5237) );
  INV_X1 U6421 ( .A(n5218), .ZN(n4598) );
  NAND2_X1 U6422 ( .A1(n6812), .A2(n5112), .ZN(n9075) );
  NAND2_X1 U6423 ( .A1(n9238), .A2(n9190), .ZN(n6896) );
  NOR2_X2 U6424 ( .A1(n9478), .A2(n7955), .ZN(n9461) );
  AOI21_X1 U6425 ( .B1(n5028), .B2(n5031), .A(n4375), .ZN(n5026) );
  OAI21_X1 U6426 ( .B1(n9248), .B2(n9040), .A(n4625), .ZN(n9254) );
  NOR2_X1 U6427 ( .A1(n5026), .A2(n5027), .ZN(n5025) );
  INV_X1 U6428 ( .A(n4827), .ZN(n4823) );
  NAND2_X1 U6429 ( .A1(n4624), .A2(n4623), .ZN(n9270) );
  INV_X1 U6430 ( .A(n9256), .ZN(n4744) );
  NAND2_X1 U6431 ( .A1(n9048), .A2(n5216), .ZN(n5929) );
  NAND2_X1 U6432 ( .A1(n9432), .A2(n9160), .ZN(n9420) );
  NAND2_X1 U6433 ( .A1(n5100), .A2(n5097), .ZN(n9432) );
  NOR2_X1 U6434 ( .A1(n6425), .A2(n6424), .ZN(n8224) );
  NAND2_X1 U6435 ( .A1(n8309), .A2(n8308), .ZN(n4639) );
  AOI21_X1 U6436 ( .B1(n8222), .B2(n6570), .A(n6569), .ZN(n6650) );
  NOR2_X1 U6437 ( .A1(n8323), .A2(n8324), .ZN(n8327) );
  NOR2_X1 U6438 ( .A1(n6839), .A2(n6838), .ZN(n6842) );
  NAND2_X2 U6439 ( .A1(n6186), .A2(n9055), .ZN(n7678) );
  NAND2_X1 U6440 ( .A1(n5008), .A2(n5573), .ZN(n5593) );
  NOR2_X1 U6441 ( .A1(n9600), .A2(n9605), .ZN(n4788) );
  NAND2_X1 U6442 ( .A1(n5694), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U6443 ( .A1(n4685), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5486) );
  INV_X1 U6444 ( .A(n4682), .ZN(n5780) );
  OAI21_X2 U6445 ( .B1(n8406), .B2(n5782), .A(n5787), .ZN(n8398) );
  NOR2_X4 U6446 ( .A1(n8691), .A2(n8477), .ZN(n8439) );
  NOR2_X4 U6447 ( .A1(n7438), .A2(n8002), .ZN(n8034) );
  INV_X1 U6448 ( .A(n8665), .ZN(n4692) );
  NAND2_X1 U6449 ( .A1(n4614), .A2(n4822), .ZN(n4622) );
  NAND2_X1 U6450 ( .A1(n4824), .A2(n8397), .ZN(n4614) );
  INV_X1 U6451 ( .A(n7134), .ZN(n4617) );
  AOI21_X1 U6452 ( .B1(n4779), .B2(n4781), .A(n4350), .ZN(n4778) );
  XNOR2_X1 U6453 ( .A(n9365), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U6454 ( .A1(n9398), .A2(n7978), .ZN(n7981) );
  NAND2_X1 U6455 ( .A1(n4648), .A2(n4357), .ZN(n7559) );
  INV_X1 U6456 ( .A(n6630), .ZN(n6641) );
  AOI21_X1 U6457 ( .B1(n4751), .B2(n4758), .A(n4749), .ZN(n4748) );
  NOR2_X1 U6458 ( .A1(n5025), .A2(n8028), .ZN(n5020) );
  NAND2_X1 U6459 ( .A1(n4657), .A2(n4656), .ZN(n4655) );
  NAND2_X1 U6460 ( .A1(n4621), .A2(n4620), .ZN(n9262) );
  NAND2_X1 U6461 ( .A1(n9257), .A2(n9256), .ZN(n4621) );
  AOI21_X1 U6462 ( .B1(n6078), .B2(n5032), .A(n6077), .ZN(n6080) );
  NAND2_X1 U6463 ( .A1(n4622), .A2(n4828), .ZN(n8033) );
  NOR2_X1 U6464 ( .A1(n4827), .A2(n4825), .ZN(n4824) );
  OAI21_X1 U6465 ( .B1(n5020), .B2(n5021), .A(n5936), .ZN(n5019) );
  NAND3_X1 U6466 ( .A1(n9268), .A2(n9266), .A3(n9267), .ZN(n4624) );
  AOI21_X1 U6467 ( .B1(n4891), .B2(n4892), .A(n4890), .ZN(n4889) );
  NAND2_X1 U6468 ( .A1(n7334), .A2(n4973), .ZN(n4972) );
  INV_X1 U6469 ( .A(n4774), .ZN(n4773) );
  NAND2_X1 U6470 ( .A1(n5876), .A2(n7191), .ZN(n5882) );
  OAI21_X2 U6471 ( .B1(n8473), .B2(n8482), .A(n6040), .ZN(n8423) );
  NAND2_X1 U6472 ( .A1(n4633), .A2(n4369), .ZN(P1_U3520) );
  NAND2_X1 U6473 ( .A1(n9707), .A2(n9876), .ZN(n4633) );
  NAND3_X1 U6474 ( .A1(n5117), .A2(n4265), .A3(n5115), .ZN(n4634) );
  NAND2_X1 U6475 ( .A1(n6813), .A2(n9231), .ZN(n6812) );
  OAI21_X2 U6476 ( .B1(n9540), .B2(n9128), .A(n9126), .ZN(n9523) );
  NAND3_X1 U6477 ( .A1(n5117), .A2(n4265), .A3(n6124), .ZN(n4949) );
  NAND2_X1 U6478 ( .A1(n9461), .A2(n5095), .ZN(n5100) );
  NOR2_X1 U6479 ( .A1(n7213), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8323) );
  NOR2_X1 U6480 ( .A1(n5167), .A2(n5168), .ZN(n5169) );
  NOR2_X1 U6481 ( .A1(n6701), .A2(n6702), .ZN(n6838) );
  NOR2_X1 U6482 ( .A1(n6841), .A2(n6842), .ZN(n7210) );
  NAND3_X1 U6483 ( .A1(n6082), .A2(n6087), .A3(n7540), .ZN(n4649) );
  NAND2_X1 U6484 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  NAND2_X1 U6485 ( .A1(n8344), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8363) );
  XNOR2_X1 U6486 ( .A(n4640), .B(n4954), .ZN(n5951) );
  NAND3_X1 U6487 ( .A1(n5032), .A2(n4312), .A3(n4683), .ZN(n4640) );
  OAI21_X1 U6488 ( .B1(n4644), .B2(n7901), .A(n4643), .ZN(n7906) );
  NAND2_X1 U6489 ( .A1(n7901), .A2(n7907), .ZN(n4643) );
  AND2_X1 U6490 ( .A1(n7908), .A2(n4645), .ZN(n4644) );
  NAND2_X1 U6491 ( .A1(n5892), .A2(n5034), .ZN(n8415) );
  NAND2_X1 U6492 ( .A1(n8395), .A2(n6074), .ZN(n8028) );
  INV_X1 U6493 ( .A(n4814), .ZN(n4813) );
  NAND2_X1 U6494 ( .A1(n8659), .A2(n8377), .ZN(n5936) );
  NAND2_X1 U6495 ( .A1(n6081), .A2(n6070), .ZN(n4658) );
  NAND3_X1 U6496 ( .A1(n7166), .A2(n9090), .A3(n9203), .ZN(n5091) );
  NAND2_X1 U6497 ( .A1(n5091), .A2(n5092), .ZN(n7362) );
  NAND3_X1 U6498 ( .A1(n9182), .A2(n4745), .A3(n4743), .ZN(n9229) );
  NAND2_X1 U6499 ( .A1(n4654), .A2(n4352), .ZN(n9054) );
  NAND2_X1 U6500 ( .A1(n9042), .A2(n4655), .ZN(n4654) );
  NAND3_X1 U6501 ( .A1(n4658), .A2(n4808), .A3(n7278), .ZN(n6087) );
  NAND3_X1 U6502 ( .A1(n7540), .A2(n6088), .A3(n6550), .ZN(n4660) );
  XNOR2_X1 U6503 ( .A(n5682), .B(n5681), .ZN(n7792) );
  INV_X1 U6504 ( .A(n8423), .ZN(n8458) );
  NAND2_X1 U6505 ( .A1(n4816), .A2(n4813), .ZN(n8473) );
  NAND3_X1 U6506 ( .A1(n9167), .A2(n9388), .A3(n4664), .ZN(n9168) );
  NAND2_X1 U6507 ( .A1(n9707), .A2(n9891), .ZN(n4787) );
  NAND2_X1 U6508 ( .A1(n4867), .A2(n5503), .ZN(n5524) );
  INV_X1 U6509 ( .A(n5066), .ZN(n7698) );
  NAND2_X1 U6510 ( .A1(n4668), .A2(n4667), .ZN(n5066) );
  NAND2_X1 U6511 ( .A1(n7695), .A2(n8888), .ZN(n4667) );
  NAND2_X1 U6512 ( .A1(n7696), .A2(n7697), .ZN(n4668) );
  INV_X1 U6513 ( .A(n5068), .ZN(n5067) );
  XNOR2_X1 U6514 ( .A(n4791), .B(n6207), .ZN(n6186) );
  NAND2_X1 U6515 ( .A1(n4777), .A2(n4778), .ZN(n4669) );
  NAND2_X1 U6516 ( .A1(n6744), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6877) );
  INV_X1 U6517 ( .A(n7878), .ZN(n8816) );
  AOI21_X2 U6518 ( .B1(n7526), .B2(n9017), .A(n9016), .ZN(n7527) );
  NOR2_X2 U6519 ( .A1(n7753), .A2(n7629), .ZN(n4673) );
  NAND2_X1 U6520 ( .A1(n4691), .A2(n4690), .ZN(P2_U3517) );
  NAND2_X1 U6521 ( .A1(n4975), .A2(n4974), .ZN(P2_U3549) );
  NAND2_X1 U6522 ( .A1(n6497), .A2(n6498), .ZN(n6640) );
  NAND2_X1 U6523 ( .A1(n7088), .A2(n7087), .ZN(n4674) );
  NAND2_X1 U6524 ( .A1(n5333), .A2(n5332), .ZN(n5356) );
  OAI21_X2 U6525 ( .B1(n9075), .B2(n7077), .A(n9236), .ZN(n7164) );
  OAI21_X1 U6526 ( .B1(n6752), .B2(n9285), .A(n9821), .ZN(n6754) );
  OAI21_X2 U6527 ( .B1(n8297), .B2(n8292), .A(n6655), .ZN(n8295) );
  XNOR2_X2 U6528 ( .A(n5227), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U6529 ( .A1(n6490), .A2(n6491), .ZN(n6497) );
  NAND2_X1 U6530 ( .A1(n5079), .A2(n5076), .ZN(n7806) );
  NAND4_X1 U6531 ( .A1(n5117), .A2(n5115), .A3(n4346), .A4(n4265), .ZN(n9728)
         );
  NAND2_X1 U6532 ( .A1(n4787), .A2(n4374), .ZN(P1_U3552) );
  NAND2_X1 U6533 ( .A1(n6080), .A2(n6079), .ZN(n4808) );
  NOR2_X2 U6534 ( .A1(n5706), .A2(n8059), .ZN(n5694) );
  NOR2_X1 U6535 ( .A1(n5950), .A2(n8027), .ZN(n4683) );
  NAND2_X1 U6536 ( .A1(n8463), .A2(n4891), .ZN(n4687) );
  NAND2_X1 U6537 ( .A1(n4687), .A2(n4889), .ZN(n8025) );
  INV_X1 U6538 ( .A(n9922), .ZN(n6937) );
  NAND2_X1 U6539 ( .A1(n4894), .A2(n4688), .ZN(n9902) );
  NAND3_X1 U6540 ( .A1(n6937), .A2(n9923), .A3(n7058), .ZN(n4688) );
  INV_X1 U6541 ( .A(n9893), .ZN(n9903) );
  NAND3_X1 U6542 ( .A1(n4282), .A2(n4693), .A3(n5053), .ZN(n4908) );
  OAI21_X1 U6543 ( .B1(n8004), .B2(n4700), .A(n4697), .ZN(n8602) );
  NAND3_X1 U6544 ( .A1(n6946), .A2(n5126), .A3(n4704), .ZN(n4701) );
  NAND2_X1 U6545 ( .A1(n4701), .A2(n4702), .ZN(n7468) );
  NAND2_X1 U6546 ( .A1(n8823), .A2(n4717), .ZN(n4716) );
  NAND3_X1 U6547 ( .A1(n4728), .A2(n5085), .A3(n4727), .ZN(n7878) );
  NAND2_X1 U6548 ( .A1(n8957), .A2(n4292), .ZN(n4727) );
  NAND2_X2 U6549 ( .A1(n4262), .A2(n6355), .ZN(n7898) );
  NAND3_X1 U6550 ( .A1(n7893), .A2(n6355), .A3(n6643), .ZN(n6359) );
  NAND2_X1 U6551 ( .A1(n4732), .A2(n9285), .ZN(n6496) );
  NAND2_X1 U6552 ( .A1(n4732), .A2(n9283), .ZN(n6529) );
  NAND2_X1 U6553 ( .A1(n4732), .A2(n9282), .ZN(n6987) );
  NAND2_X1 U6554 ( .A1(n4732), .A2(n9281), .ZN(n6998) );
  AOI22_X1 U6555 ( .A1(n9280), .A2(n4732), .B1(n7900), .B2(n7108), .ZN(n7235)
         );
  NAND2_X1 U6556 ( .A1(n7932), .A2(n4732), .ZN(n7730) );
  NAND2_X1 U6557 ( .A1(n9511), .A2(n4732), .ZN(n7765) );
  NAND2_X1 U6558 ( .A1(n9447), .A2(n4732), .ZN(n7802) );
  NAND2_X1 U6559 ( .A1(n9462), .A2(n4732), .ZN(n7834) );
  NAND2_X1 U6560 ( .A1(n9448), .A2(n4732), .ZN(n7819) );
  NAND3_X1 U6561 ( .A1(n9087), .A2(n4742), .A3(n4740), .ZN(n9098) );
  NAND4_X1 U6562 ( .A1(n9174), .A2(n9256), .A3(n9252), .A4(n9173), .ZN(n4745)
         );
  NAND4_X1 U6563 ( .A1(n5115), .A2(n4265), .A3(n4353), .A4(n5117), .ZN(n6211)
         );
  NAND2_X1 U6564 ( .A1(n8072), .A2(n4751), .ZN(n4750) );
  INV_X1 U6565 ( .A(n5305), .ZN(n4770) );
  INV_X1 U6566 ( .A(n4968), .ZN(n4771) );
  OAI21_X1 U6567 ( .B1(n4771), .B2(n4773), .A(n4772), .ZN(n5548) );
  NAND2_X2 U6568 ( .A1(n6619), .A2(n5867), .ZN(n6401) );
  NOR2_X2 U6569 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6303) );
  NAND2_X1 U6570 ( .A1(n7516), .A2(n4779), .ZN(n4777) );
  NAND4_X1 U6571 ( .A1(n4796), .A2(n6007), .A3(n6008), .A4(n6009), .ZN(n4795)
         );
  NAND3_X1 U6572 ( .A1(n6003), .A2(n6002), .A3(n6004), .ZN(n4796) );
  NAND2_X1 U6573 ( .A1(n5985), .A2(n7200), .ZN(n6956) );
  NAND2_X1 U6574 ( .A1(n8534), .A2(n4817), .ZN(n4816) );
  OAI21_X2 U6575 ( .B1(n8423), .B2(n5891), .A(n5890), .ZN(n5892) );
  NAND2_X1 U6576 ( .A1(n8397), .A2(n4826), .ZN(n4828) );
  NAND2_X1 U6577 ( .A1(n8397), .A2(n8396), .ZN(n8395) );
  OAI22_X2 U6578 ( .A1(n7473), .A2(n4829), .B1(n4831), .B2(n5943), .ZN(n7373)
         );
  AOI21_X2 U6579 ( .B1(n8546), .B2(n8554), .A(n4836), .ZN(n5129) );
  INV_X2 U6580 ( .A(n4885), .ZN(n9941) );
  NAND3_X1 U6581 ( .A1(n5194), .A2(n5196), .A3(n5195), .ZN(n4885) );
  NAND3_X1 U6582 ( .A1(n4844), .A2(n4842), .A3(n4841), .ZN(n8092) );
  OR2_X1 U6583 ( .A1(n8180), .A2(n4853), .ZN(n4846) );
  NAND3_X1 U6584 ( .A1(n4846), .A2(n4845), .A3(n4847), .ZN(n5875) );
  NAND2_X1 U6585 ( .A1(n8180), .A2(n4850), .ZN(n4845) );
  AND2_X1 U6586 ( .A1(n5198), .A2(n5037), .ZN(n4887) );
  NAND2_X1 U6587 ( .A1(n4887), .A2(n5036), .ZN(n9911) );
  NAND2_X1 U6588 ( .A1(n7381), .A2(n4903), .ZN(n4901) );
  NAND2_X1 U6589 ( .A1(n4908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5178) );
  AOI21_X1 U6590 ( .B1(n8487), .B2(n8488), .A(n8016), .ZN(n8483) );
  OAI21_X1 U6591 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7286), .A(n7132), .ZN(
        n7134) );
  NAND2_X1 U6592 ( .A1(n9297), .A2(n9296), .ZN(n9298) );
  INV_X1 U6593 ( .A(n6945), .ZN(n6946) );
  NOR3_X4 U6594 ( .A1(n5125), .A2(n9648), .A3(n4919), .ZN(n9502) );
  NOR2_X1 U6595 ( .A1(n9436), .A2(n4921), .ZN(n9394) );
  NAND2_X1 U6596 ( .A1(n9239), .A2(n4926), .ZN(n9195) );
  NAND4_X1 U6597 ( .A1(n9077), .A2(n9242), .A3(n9170), .A4(n4926), .ZN(n9087)
         );
  NAND2_X1 U6598 ( .A1(n7327), .A2(n4283), .ZN(n4929) );
  NAND2_X1 U6599 ( .A1(n9442), .A2(n4938), .ZN(n4936) );
  AND2_X2 U6600 ( .A1(n6213), .A2(n6280), .ZN(n6532) );
  AND2_X2 U6601 ( .A1(n6213), .A2(n9732), .ZN(n6879) );
  OAI22_X1 U6602 ( .A1(n6213), .A2(P1_U3084), .B1(n9743), .B2(n9045), .ZN(
        n4946) );
  NAND2_X1 U6603 ( .A1(n4951), .A2(n4953), .ZN(n4952) );
  INV_X1 U6604 ( .A(n8067), .ZN(n4951) );
  AND2_X1 U6605 ( .A1(n4952), .A2(n4295), .ZN(n8139) );
  INV_X1 U6606 ( .A(n8066), .ZN(n4953) );
  NAND3_X1 U6607 ( .A1(n4955), .A2(n7278), .A3(n4954), .ZN(n5269) );
  NAND3_X1 U6608 ( .A1(n5137), .A2(n5266), .A3(n5136), .ZN(n5149) );
  AOI21_X2 U6609 ( .B1(n8175), .B2(n8174), .A(n5590), .ZN(n8074) );
  OAI21_X1 U6610 ( .B1(n7335), .B2(n7334), .A(n4973), .ZN(n7405) );
  NAND2_X1 U6611 ( .A1(n4282), .A2(n4976), .ZN(n5175) );
  INV_X1 U6612 ( .A(n4984), .ZN(n7505) );
  NAND2_X1 U6613 ( .A1(n8549), .A2(n4989), .ZN(n8496) );
  INV_X1 U6614 ( .A(n7930), .ZN(n7910) );
  NAND2_X1 U6615 ( .A1(n7930), .A2(n4260), .ZN(n5577) );
  NAND2_X1 U6616 ( .A1(n5282), .A2(n5281), .ZN(n4996) );
  NAND2_X1 U6617 ( .A1(n5556), .A2(n5006), .ZN(n5008) );
  XNOR2_X1 U6618 ( .A(n5019), .B(n8435), .ZN(n5934) );
  NAND3_X1 U6619 ( .A1(n5023), .A2(n5032), .A3(n5022), .ZN(n5021) );
  INV_X1 U6620 ( .A(n5033), .ZN(n5031) );
  NAND2_X1 U6621 ( .A1(n5129), .A2(n5887), .ZN(n8534) );
  NAND2_X1 U6622 ( .A1(n5040), .A2(n5041), .ZN(n8562) );
  NAND2_X1 U6623 ( .A1(n7693), .A2(n5070), .ZN(n5065) );
  INV_X1 U6624 ( .A(n7693), .ZN(n5071) );
  NAND2_X1 U6625 ( .A1(n5116), .A2(n5117), .ZN(n6308) );
  NAND2_X1 U6626 ( .A1(n8872), .A2(n5078), .ZN(n5077) );
  NAND4_X1 U6627 ( .A1(n7916), .A2(n7913), .A3(n8872), .A4(n5080), .ZN(n5079)
         );
  NAND2_X1 U6628 ( .A1(n8925), .A2(n5082), .ZN(n7006) );
  NAND2_X1 U6629 ( .A1(n6360), .A2(n6476), .ZN(n6752) );
  OAI21_X1 U6630 ( .B1(n5109), .B2(n7588), .A(n9021), .ZN(n5108) );
  INV_X1 U6631 ( .A(n5111), .ZN(n7590) );
  INV_X1 U6632 ( .A(n9012), .ZN(n5114) );
  INV_X1 U6633 ( .A(n6165), .ZN(n5116) );
  NAND2_X1 U6634 ( .A1(n9411), .A2(n5121), .ZN(n5118) );
  NAND2_X1 U6635 ( .A1(n5118), .A2(n5119), .ZN(n7984) );
  AND2_X1 U6636 ( .A1(n7928), .A2(n7931), .ZN(n9528) );
  INV_X1 U6637 ( .A(n9622), .ZN(n9441) );
  CLKBUF_X1 U6638 ( .A(n6186), .Z(n9056) );
  NAND2_X1 U6639 ( .A1(n9435), .A2(n9441), .ZN(n9436) );
  INV_X1 U6640 ( .A(n8099), .ZN(n8101) );
  OR2_X1 U6641 ( .A1(n6088), .A2(n5870), .ZN(n9985) );
  OR2_X1 U6642 ( .A1(n9986), .A2(n4954), .ZN(n6545) );
  NAND2_X1 U6643 ( .A1(n5805), .A2(n5804), .ZN(n5807) );
  NAND2_X1 U6644 ( .A1(n5895), .A2(n5894), .ZN(n5899) );
  CLKBUF_X1 U6645 ( .A(n7473), .Z(n7477) );
  XNOR2_X1 U6646 ( .A(n5742), .B(n5717), .ZN(n7807) );
  NAND2_X1 U6647 ( .A1(n6365), .A2(n6489), .ZN(n6491) );
  XNOR2_X1 U6648 ( .A(n8659), .B(n8383), .ZN(n8661) );
  AND2_X1 U6649 ( .A1(n5408), .A2(n5388), .ZN(n5124) );
  OR2_X2 U6650 ( .A1(n9579), .A2(n9668), .ZN(n5125) );
  INV_X1 U6651 ( .A(n8596), .ZN(n8640) );
  AND2_X1 U6652 ( .A1(n5874), .A2(n5873), .ZN(n5127) );
  INV_X1 U6653 ( .A(n8533), .ZN(n5887) );
  AND2_X1 U6654 ( .A1(n9816), .A2(n6447), .ZN(n5128) );
  INV_X1 U6655 ( .A(n8021), .ZN(n8444) );
  NAND2_X1 U6656 ( .A1(n8425), .A2(n6062), .ZN(n8021) );
  NAND3_X1 U6657 ( .A1(n6550), .A2(n6088), .A3(n7554), .ZN(n5148) );
  INV_X1 U6658 ( .A(n8464), .ZN(n8018) );
  AND2_X1 U6659 ( .A1(n9165), .A2(n9419), .ZN(n9040) );
  AND2_X1 U6660 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NAND2_X2 U6661 ( .A1(n5148), .A2(n6923), .ZN(n5236) );
  INV_X1 U6662 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10076) );
  AND2_X1 U6663 ( .A1(n9195), .A2(n7069), .ZN(n7067) );
  INV_X1 U6664 ( .A(n5498), .ZN(n5499) );
  INV_X1 U6665 ( .A(SI_10_), .ZN(n5385) );
  INV_X1 U6666 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U6667 ( .A1(n7025), .A2(n5975), .ZN(n7029) );
  INV_X1 U6668 ( .A(n8573), .ZN(n8575) );
  INV_X1 U6669 ( .A(n7191), .ZN(n7203) );
  INV_X1 U6670 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5176) );
  INV_X1 U6671 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7157) );
  INV_X1 U6672 ( .A(n6746), .ZN(n6744) );
  NAND2_X1 U6673 ( .A1(n7297), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7253) );
  OR2_X1 U6674 ( .A1(n9628), .A2(n8849), .ZN(n9159) );
  INV_X1 U6675 ( .A(n9535), .ZN(n7935) );
  INV_X1 U6676 ( .A(n7998), .ZN(n9603) );
  OR2_X1 U6677 ( .A1(n5747), .A2(n5746), .ZN(n5768) );
  NAND2_X1 U6678 ( .A1(n5507), .A2(n5506), .ZN(n5522) );
  INV_X1 U6679 ( .A(n8206), .ZN(n8412) );
  INV_X1 U6680 ( .A(n8474), .ZN(n8061) );
  INV_X1 U6681 ( .A(n8459), .ZN(n8132) );
  INV_X1 U6682 ( .A(n8492), .ZN(n8165) );
  OR2_X1 U6683 ( .A1(n6715), .A2(n6548), .ZN(n5932) );
  INV_X1 U6684 ( .A(n8594), .ZN(n8601) );
  INV_X1 U6685 ( .A(n8209), .ZN(n7375) );
  INV_X1 U6686 ( .A(n9913), .ZN(n9892) );
  NAND2_X1 U6687 ( .A1(n5145), .A2(n5141), .ZN(n5142) );
  NAND2_X1 U6688 ( .A1(n6640), .A2(n6638), .ZN(n6635) );
  INV_X1 U6689 ( .A(n7254), .ZN(n7133) );
  AND2_X1 U6690 ( .A1(n9628), .A2(n9448), .ZN(n7968) );
  INV_X1 U6691 ( .A(n9081), .ZN(n9851) );
  NAND2_X1 U6692 ( .A1(n5522), .A2(n5509), .ZN(n5523) );
  INV_X1 U6693 ( .A(n8202), .ZN(n8162) );
  NOR2_X1 U6694 ( .A1(n5869), .A2(n6394), .ZN(n5866) );
  INV_X1 U6695 ( .A(n5289), .ZN(n5797) );
  INV_X1 U6696 ( .A(n10204), .ZN(n8335) );
  INV_X1 U6697 ( .A(n8370), .ZN(n10190) );
  AND2_X1 U6698 ( .A1(n8634), .A2(n8633), .ZN(n8752) );
  INV_X1 U6699 ( .A(n9924), .ZN(n8611) );
  AND2_X1 U6700 ( .A1(n8581), .A2(n9984), .ZN(n8751) );
  INV_X1 U6701 ( .A(n8751), .ZN(n9981) );
  INV_X1 U6702 ( .A(n8993), .ZN(n8964) );
  NAND2_X1 U6703 ( .A1(n6446), .A2(n9530), .ZN(n8978) );
  INV_X1 U6704 ( .A(n9056), .ZN(n9780) );
  AND2_X1 U6705 ( .A1(n9368), .A2(n9056), .ZN(n9369) );
  INV_X1 U6706 ( .A(n9813), .ZN(n9375) );
  INV_X1 U6707 ( .A(n9501), .ZN(n9572) );
  INV_X1 U6708 ( .A(n9845), .ZN(n7048) );
  INV_X1 U6709 ( .A(n9530), .ZN(n9582) );
  OR2_X1 U6710 ( .A1(n6440), .A2(n9267), .ZN(n9868) );
  AND2_X1 U6711 ( .A1(n9170), .A2(n7276), .ZN(n9856) );
  AND2_X1 U6712 ( .A1(n6292), .A2(n6351), .ZN(n7297) );
  INV_X1 U6713 ( .A(n8375), .ZN(n10200) );
  AND2_X1 U6714 ( .A1(n5850), .A2(n9919), .ZN(n8115) );
  INV_X1 U6715 ( .A(n8191), .ZN(n8166) );
  NAND2_X1 U6716 ( .A1(n5866), .A2(n5852), .ZN(n8202) );
  NAND2_X1 U6717 ( .A1(n8606), .A2(n6924), .ZN(n9924) );
  AND2_X2 U6718 ( .A1(n7146), .A2(n6547), .ZN(n10004) );
  INV_X1 U6719 ( .A(n9994), .ZN(n9992) );
  INV_X1 U6720 ( .A(n9931), .ZN(n9935) );
  INV_X1 U6721 ( .A(n9930), .ZN(n9938) );
  INV_X1 U6722 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6354) );
  INV_X1 U6723 ( .A(n7108), .ZN(n9859) );
  INV_X1 U6724 ( .A(n8978), .ZN(n8988) );
  AOI21_X1 U6725 ( .B1(n7636), .B2(n4264), .A(n7635), .ZN(n9391) );
  INV_X1 U6726 ( .A(n7957), .ZN(n9462) );
  INV_X1 U6727 ( .A(P1_U4006), .ZN(n9274) );
  INV_X1 U6728 ( .A(n9376), .ZN(n9595) );
  INV_X1 U6729 ( .A(n9891), .ZN(n9888) );
  INV_X1 U6730 ( .A(n9876), .ZN(n9874) );
  INV_X1 U6731 ( .A(n9817), .ZN(n9818) );
  INV_X1 U6732 ( .A(n6152), .ZN(n9746) );
  INV_X1 U6733 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7677) );
  NOR2_X1 U6734 ( .A1(n10217), .A2(n10216), .ZN(n10215) );
  NOR2_X1 U6735 ( .A1(n10033), .A2(n10032), .ZN(n10031) );
  NOR2_X1 U6736 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5133) );
  AND2_X2 U6737 ( .A1(n5167), .A2(n5134), .ZN(n5266) );
  NAND2_X1 U6738 ( .A1(n5816), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5812) );
  XNOR2_X1 U6739 ( .A(n5812), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6740 ( .A1(n4334), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6741 ( .A1(n5140), .A2(n8435), .ZN(n6550) );
  INV_X1 U6742 ( .A(n5140), .ZN(n7962) );
  NAND2_X1 U6743 ( .A1(n5142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5144) );
  INV_X1 U6744 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U6745 ( .A1(n5146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5147) );
  INV_X1 U6746 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5150) );
  NOR2_X1 U6747 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5153) );
  NOR2_X1 U6748 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5152) );
  NOR2_X1 U6749 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5151) );
  NAND2_X1 U6750 ( .A1(n5175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5154) );
  XNOR2_X1 U6751 ( .A(n5154), .B(n5176), .ZN(n5867) );
  NOR2_X1 U6752 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5158) );
  AND2_X1 U6753 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5186) );
  INV_X1 U6754 ( .A(n5186), .ZN(n5157) );
  NAND2_X1 U6755 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5156) );
  OAI21_X1 U6756 ( .B1(n5158), .B2(n5157), .A(n5156), .ZN(n5159) );
  NAND2_X1 U6757 ( .A1(n6454), .A2(n5159), .ZN(n5164) );
  NOR2_X1 U6758 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6759 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6760 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5160) );
  OAI21_X1 U6761 ( .B1(n5161), .B2(n5187), .A(n5160), .ZN(n5162) );
  NAND2_X1 U6762 ( .A1(n4598), .A2(n5162), .ZN(n5163) );
  NAND2_X1 U6763 ( .A1(n5164), .A2(n5163), .ZN(n5221) );
  INV_X1 U6764 ( .A(SI_2_), .ZN(n5219) );
  XNOR2_X1 U6765 ( .A(n5221), .B(n5219), .ZN(n5166) );
  MUX2_X1 U6766 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5504), .Z(n5165) );
  XNOR2_X1 U6767 ( .A(n5166), .B(n5165), .ZN(n6501) );
  NAND2_X1 U6768 ( .A1(n5225), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5174) );
  INV_X4 U6769 ( .A(n6401), .ZN(n5600) );
  NAND2_X1 U6770 ( .A1(n5169), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5172) );
  INV_X1 U6771 ( .A(n5169), .ZN(n5171) );
  INV_X1 U6772 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6773 ( .A1(n5171), .A2(n5170), .ZN(n5226) );
  NAND2_X1 U6774 ( .A1(n5600), .A2(n6557), .ZN(n5173) );
  XNOR2_X1 U6775 ( .A(n5236), .B(n9915), .ZN(n5210) );
  MUX2_X1 U6776 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5178), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5179) );
  AND2_X2 U6777 ( .A1(n5179), .A2(n8790), .ZN(n5180) );
  NAND2_X1 U6778 ( .A1(n5314), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5185) );
  AND2_X2 U6779 ( .A1(n5181), .A2(n8794), .ZN(n5289) );
  NAND2_X1 U6780 ( .A1(n5289), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5184) );
  AND2_X4 U6781 ( .A1(n5181), .A2(n5180), .ZN(n5794) );
  NAND2_X1 U6782 ( .A1(n5794), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5182) );
  NAND4_X2 U6783 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n8216)
         );
  NAND2_X1 U6784 ( .A1(n5210), .A2(n5211), .ZN(n6723) );
  NAND2_X1 U6785 ( .A1(n5504), .A2(n5186), .ZN(n6326) );
  OAI21_X1 U6786 ( .B1(n5504), .B2(n5187), .A(n6326), .ZN(n5188) );
  XNOR2_X1 U6787 ( .A(n5188), .B(SI_1_), .ZN(n5190) );
  MUX2_X1 U6788 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5504), .Z(n5189) );
  XNOR2_X1 U6789 ( .A(n5190), .B(n5189), .ZN(n6127) );
  NAND2_X1 U6790 ( .A1(n5216), .A2(n6127), .ZN(n5196) );
  NAND2_X1 U6791 ( .A1(n5225), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6792 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5191) );
  INV_X1 U6793 ( .A(n5167), .ZN(n5192) );
  INV_X1 U6794 ( .A(n6417), .ZN(n6427) );
  NAND2_X1 U6795 ( .A1(n5600), .A2(n6427), .ZN(n5194) );
  XNOR2_X1 U6796 ( .A(n5236), .B(n9941), .ZN(n5209) );
  INV_X1 U6797 ( .A(n5209), .ZN(n5200) );
  NAND2_X1 U6798 ( .A1(n5794), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6799 ( .A1(n5289), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6800 ( .A1(n5200), .A2(n5199), .ZN(n6611) );
  NAND2_X1 U6801 ( .A1(n6455), .A2(SI_0_), .ZN(n5201) );
  XNOR2_X1 U6802 ( .A(n5201), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8812) );
  MUX2_X1 U6803 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8812), .S(n6401), .Z(n6931) );
  OR2_X1 U6804 ( .A1(n5236), .A2(n6931), .ZN(n5207) );
  NAND2_X1 U6805 ( .A1(n5314), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6806 ( .A1(n5289), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6807 ( .A1(n5794), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U6808 ( .A1(n6934), .A2(n5269), .ZN(n5206) );
  NAND3_X1 U6809 ( .A1(n6723), .A2(n6611), .A3(n6610), .ZN(n5215) );
  NAND2_X1 U6810 ( .A1(n6720), .A2(n6723), .ZN(n5214) );
  INV_X1 U6811 ( .A(n5210), .ZN(n5213) );
  INV_X1 U6812 ( .A(n5211), .ZN(n5212) );
  NAND2_X1 U6813 ( .A1(n5213), .A2(n5212), .ZN(n6722) );
  NAND3_X1 U6814 ( .A1(n5215), .A2(n5214), .A3(n6722), .ZN(n8067) );
  INV_X1 U6815 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U6816 ( .A1(n6454), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5220) );
  OAI211_X1 U6817 ( .C1(n6454), .C2(n6147), .A(n5220), .B(n5219), .ZN(n5222)
         );
  INV_X1 U6818 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U6819 ( .A1(n6454), .A2(n6502), .ZN(n5223) );
  OAI211_X1 U6820 ( .C1(n6454), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5223), .B(
        SI_2_), .ZN(n5224) );
  XNOR2_X1 U6821 ( .A(n5237), .B(n5238), .ZN(n6520) );
  NAND2_X1 U6822 ( .A1(n4260), .A2(n6520), .ZN(n5230) );
  NAND2_X1 U6823 ( .A1(n5909), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6824 ( .A1(n5226), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6825 ( .A1(n5600), .A2(n8225), .ZN(n5228) );
  AND3_X2 U6826 ( .A1(n5230), .A2(n5229), .A3(n5228), .ZN(n7054) );
  INV_X1 U6827 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6828 ( .A1(n5794), .A2(n5249), .ZN(n5234) );
  NAND2_X1 U6829 ( .A1(n5314), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6831 ( .A1(n5289), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6832 ( .A1(n5729), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5231) );
  INV_X1 U6833 ( .A(n5237), .ZN(n5239) );
  NAND2_X1 U6834 ( .A1(n5240), .A2(SI_3_), .ZN(n5241) );
  NAND2_X1 U6835 ( .A1(n6734), .A2(n4260), .ZN(n5246) );
  OR2_X1 U6836 ( .A1(n5266), .A2(n5168), .ZN(n5243) );
  XNOR2_X1 U6837 ( .A(n5243), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U6838 ( .A1(n5600), .A2(n6663), .ZN(n5245) );
  NAND2_X1 U6839 ( .A1(n5909), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5244) );
  XNOR2_X1 U6840 ( .A(n5236), .B(n9965), .ZN(n5255) );
  NAND2_X1 U6841 ( .A1(n5729), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6842 ( .A1(n5314), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5253) );
  INV_X1 U6843 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6844 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  AND2_X1 U6846 ( .A1(n5250), .A2(n5294), .ZN(n9900) );
  NAND2_X1 U6847 ( .A1(n5794), .A2(n9900), .ZN(n5252) );
  BUF_X1 U6848 ( .A(n5289), .Z(n5757) );
  NAND2_X1 U6849 ( .A1(n5757), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5251) );
  NAND4_X1 U6850 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n8215)
         );
  NAND2_X1 U6851 ( .A1(n5269), .A2(n8215), .ZN(n5256) );
  NAND2_X1 U6852 ( .A1(n5255), .A2(n5256), .ZN(n5260) );
  INV_X1 U6853 ( .A(n5255), .ZN(n5258) );
  INV_X1 U6854 ( .A(n5256), .ZN(n5257) );
  NAND2_X1 U6855 ( .A1(n5258), .A2(n5257), .ZN(n5259) );
  AND2_X1 U6856 ( .A1(n5260), .A2(n5259), .ZN(n8138) );
  NAND2_X1 U6857 ( .A1(n5262), .A2(SI_4_), .ZN(n5263) );
  XNOR2_X1 U6858 ( .A(n5282), .B(n5280), .ZN(n6730) );
  NAND2_X1 U6859 ( .A1(n6730), .A2(n4260), .ZN(n5268) );
  INV_X1 U6860 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6861 ( .A1(n5266), .A2(n5265), .ZN(n5342) );
  NAND2_X1 U6862 ( .A1(n5342), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5285) );
  XNOR2_X1 U6863 ( .A(n5285), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8239) );
  AOI22_X1 U6864 ( .A1(n5909), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5600), .B2(
        n8239), .ZN(n5267) );
  XNOR2_X1 U6865 ( .A(n5236), .B(n9974), .ZN(n5274) );
  NAND2_X1 U6866 ( .A1(n5314), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6867 ( .A1(n5757), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5272) );
  XNOR2_X1 U6868 ( .A(n5294), .B(P2_REG3_REG_5__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U6869 ( .A1(n5794), .A2(n6791), .ZN(n5271) );
  NAND2_X1 U6870 ( .A1(n5729), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6871 ( .A1(n5322), .A2(n8214), .ZN(n5275) );
  NAND2_X1 U6872 ( .A1(n5274), .A2(n5275), .ZN(n5279) );
  INV_X1 U6873 ( .A(n5274), .ZN(n5277) );
  INV_X1 U6874 ( .A(n5275), .ZN(n5276) );
  NAND2_X1 U6875 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  AND2_X1 U6876 ( .A1(n5279), .A2(n5278), .ZN(n6795) );
  NAND2_X1 U6877 ( .A1(n6867), .A2(n4260), .ZN(n5288) );
  NAND2_X1 U6878 ( .A1(n5285), .A2(n5338), .ZN(n5286) );
  NAND2_X1 U6879 ( .A1(n5286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5309) );
  XNOR2_X1 U6880 ( .A(n5309), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8253) );
  AOI22_X1 U6881 ( .A1(n5909), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5600), .B2(
        n8253), .ZN(n5287) );
  XNOR2_X1 U6882 ( .A(n7193), .B(n5802), .ZN(n5300) );
  NAND2_X1 U6883 ( .A1(n5314), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6884 ( .A1(n5289), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5298) );
  INV_X1 U6885 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5293) );
  INV_X1 U6886 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5292) );
  OAI21_X1 U6887 ( .B1(n5294), .B2(n5293), .A(n5292), .ZN(n5295) );
  AND2_X1 U6888 ( .A1(n5316), .A2(n5295), .ZN(n7197) );
  NAND2_X1 U6889 ( .A1(n5794), .A2(n7197), .ZN(n5297) );
  NAND2_X1 U6890 ( .A1(n5729), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5296) );
  NAND4_X1 U6891 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n8213)
         );
  NAND2_X1 U6892 ( .A1(n5322), .A2(n8213), .ZN(n5301) );
  NAND2_X1 U6893 ( .A1(n5300), .A2(n5301), .ZN(n5305) );
  INV_X1 U6894 ( .A(n5300), .ZN(n5303) );
  INV_X1 U6895 ( .A(n5301), .ZN(n5302) );
  NAND2_X1 U6896 ( .A1(n5303), .A2(n5302), .ZN(n5304) );
  AND2_X1 U6897 ( .A1(n5305), .A2(n5304), .ZN(n6832) );
  NAND2_X1 U6898 ( .A1(n5307), .A2(SI_6_), .ZN(n5308) );
  MUX2_X1 U6899 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5504), .Z(n5331) );
  XNOR2_X1 U6900 ( .A(n5330), .B(n5328), .ZN(n6968) );
  NAND2_X1 U6901 ( .A1(n6968), .A2(n4260), .ZN(n5313) );
  INV_X1 U6902 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6903 ( .A1(n5309), .A2(n5339), .ZN(n5310) );
  NAND2_X1 U6904 ( .A1(n5310), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5311) );
  XNOR2_X1 U6905 ( .A(n5311), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8268) );
  AOI22_X1 U6906 ( .A1(n5909), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5600), .B2(
        n8268), .ZN(n5312) );
  XNOR2_X1 U6907 ( .A(n7378), .B(n5802), .ZN(n5323) );
  NAND2_X1 U6908 ( .A1(n5729), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6909 ( .A1(n5314), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5320) );
  INV_X1 U6910 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U6911 ( .A1(n5316), .A2(n10171), .ZN(n5317) );
  AND2_X1 U6912 ( .A1(n5347), .A2(n5317), .ZN(n6950) );
  NAND2_X1 U6913 ( .A1(n5794), .A2(n6950), .ZN(n5319) );
  NAND2_X1 U6914 ( .A1(n5289), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5318) );
  NAND4_X1 U6915 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), .ZN(n8212)
         );
  NAND2_X1 U6916 ( .A1(n5322), .A2(n8212), .ZN(n5324) );
  XNOR2_X1 U6917 ( .A(n5323), .B(n5324), .ZN(n6823) );
  INV_X1 U6918 ( .A(n5323), .ZN(n5326) );
  INV_X1 U6919 ( .A(n5324), .ZN(n5325) );
  NAND2_X1 U6920 ( .A1(n5326), .A2(n5325), .ZN(n5327) );
  NAND2_X1 U6921 ( .A1(n5331), .A2(SI_7_), .ZN(n5332) );
  MUX2_X1 U6922 ( .A(n10127), .B(n5334), .S(n5504), .Z(n5335) );
  INV_X1 U6923 ( .A(n5335), .ZN(n5336) );
  NAND2_X1 U6924 ( .A1(n5336), .A2(SI_8_), .ZN(n5337) );
  NAND2_X1 U6925 ( .A1(n7088), .A2(n4260), .ZN(n5345) );
  INV_X1 U6926 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5340) );
  NAND3_X1 U6927 ( .A1(n5340), .A2(n5339), .A3(n5338), .ZN(n5341) );
  NAND2_X1 U6928 ( .A1(n5364), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5343) );
  XNOR2_X1 U6929 ( .A(n5343), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6672) );
  AOI22_X1 U6930 ( .A1(n5909), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5600), .B2(
        n6672), .ZN(n5344) );
  NAND2_X1 U6931 ( .A1(n5345), .A2(n5344), .ZN(n7471) );
  XNOR2_X1 U6932 ( .A(n7471), .B(n5236), .ZN(n5354) );
  NAND2_X1 U6933 ( .A1(n5729), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U6934 ( .A1(n5314), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6935 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  AND2_X1 U6936 ( .A1(n5368), .A2(n5348), .ZN(n7470) );
  NAND2_X1 U6937 ( .A1(n5794), .A2(n7470), .ZN(n5349) );
  NAND2_X1 U6938 ( .A1(n5322), .A2(n8211), .ZN(n5352) );
  XNOR2_X1 U6939 ( .A(n5354), .B(n5352), .ZN(n6909) );
  INV_X1 U6940 ( .A(n5352), .ZN(n5353) );
  NAND2_X1 U6941 ( .A1(n5354), .A2(n5353), .ZN(n5355) );
  INV_X1 U6942 ( .A(n5357), .ZN(n5358) );
  NAND2_X1 U6943 ( .A1(n5406), .A2(n5403), .ZN(n5383) );
  MUX2_X1 U6944 ( .A(n5360), .B(n5359), .S(n5504), .Z(n5362) );
  INV_X1 U6945 ( .A(SI_9_), .ZN(n5361) );
  INV_X1 U6946 ( .A(n5362), .ZN(n5363) );
  AND2_X1 U6947 ( .A1(n5404), .A2(n5407), .ZN(n5382) );
  XNOR2_X1 U6948 ( .A(n5383), .B(n5382), .ZN(n7153) );
  NAND2_X1 U6949 ( .A1(n7153), .A2(n4260), .ZN(n5366) );
  XNOR2_X1 U6950 ( .A(n5390), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8303) );
  AOI22_X1 U6951 ( .A1(n5909), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5600), .B2(
        n8303), .ZN(n5365) );
  XNOR2_X1 U6952 ( .A(n8764), .B(n5802), .ZN(n5375) );
  NAND2_X1 U6953 ( .A1(n5729), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6954 ( .A1(n5314), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6955 ( .A1(n5368), .A2(n5367), .ZN(n5369) );
  NAND2_X1 U6956 ( .A1(n5395), .A2(n5369), .ZN(n7507) );
  INV_X1 U6957 ( .A(n7507), .ZN(n5370) );
  NAND2_X1 U6958 ( .A1(n5794), .A2(n5370), .ZN(n5372) );
  NAND2_X1 U6959 ( .A1(n5289), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5371) );
  NAND4_X1 U6960 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n8210)
         );
  NAND2_X1 U6961 ( .A1(n5322), .A2(n8210), .ZN(n5376) );
  NAND2_X1 U6962 ( .A1(n5375), .A2(n5376), .ZN(n5381) );
  INV_X1 U6963 ( .A(n5375), .ZN(n5378) );
  INV_X1 U6964 ( .A(n5376), .ZN(n5377) );
  NAND2_X1 U6965 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  NAND2_X1 U6966 ( .A1(n5381), .A2(n5379), .ZN(n7225) );
  INV_X1 U6967 ( .A(n7225), .ZN(n5380) );
  NAND2_X1 U6968 ( .A1(n5383), .A2(n5382), .ZN(n5384) );
  NAND2_X1 U6969 ( .A1(n5384), .A2(n5404), .ZN(n5389) );
  MUX2_X1 U6970 ( .A(n6221), .B(n6219), .S(n5808), .Z(n5386) );
  INV_X1 U6971 ( .A(n5386), .ZN(n5387) );
  NAND2_X1 U6972 ( .A1(n5387), .A2(SI_10_), .ZN(n5388) );
  NAND2_X1 U6973 ( .A1(n7281), .A2(n4260), .ZN(n5393) );
  NAND2_X1 U6974 ( .A1(n5390), .A2(n5435), .ZN(n5391) );
  NAND2_X1 U6975 ( .A1(n5391), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5409) );
  XNOR2_X1 U6976 ( .A(n5409), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6689) );
  AOI22_X1 U6977 ( .A1(n5909), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5600), .B2(
        n6689), .ZN(n5392) );
  XNOR2_X1 U6978 ( .A(n8759), .B(n5802), .ZN(n5402) );
  NAND2_X1 U6979 ( .A1(n5314), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6980 ( .A1(n5289), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6981 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  AND2_X1 U6982 ( .A1(n5415), .A2(n5396), .ZN(n7398) );
  NAND2_X1 U6983 ( .A1(n5794), .A2(n7398), .ZN(n5398) );
  NAND2_X1 U6984 ( .A1(n5915), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5397) );
  NAND4_X1 U6985 ( .A1(n5400), .A2(n5399), .A3(n5398), .A4(n5397), .ZN(n8209)
         );
  NAND2_X1 U6986 ( .A1(n5322), .A2(n8209), .ZN(n5401) );
  XNOR2_X1 U6987 ( .A(n5402), .B(n5401), .ZN(n7334) );
  MUX2_X1 U6988 ( .A(n10129), .B(n6238), .S(n5504), .Z(n5427) );
  NAND2_X1 U6989 ( .A1(n7285), .A2(n4260), .ZN(n5413) );
  INV_X1 U6990 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6991 ( .A1(n5409), .A2(n5436), .ZN(n5410) );
  NAND2_X1 U6992 ( .A1(n5410), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5411) );
  XNOR2_X1 U6993 ( .A(n5411), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6690) );
  AOI22_X1 U6994 ( .A1(n6690), .A2(n5600), .B1(n5909), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6995 ( .A1(n5413), .A2(n5412), .ZN(n7437) );
  XNOR2_X1 U6996 ( .A(n7437), .B(n5236), .ZN(n5423) );
  NAND2_X1 U6997 ( .A1(n5314), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5420) );
  INV_X1 U6998 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5414) );
  OR2_X1 U6999 ( .A1(n5797), .A2(n5414), .ZN(n5419) );
  INV_X1 U7000 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U7001 ( .A1(n5415), .A2(n8312), .ZN(n5416) );
  AND2_X1 U7002 ( .A1(n5443), .A2(n5416), .ZN(n7406) );
  NAND2_X1 U7003 ( .A1(n5794), .A2(n7406), .ZN(n5418) );
  NAND2_X1 U7004 ( .A1(n5915), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5417) );
  NAND4_X1 U7005 ( .A1(n5420), .A2(n5419), .A3(n5418), .A4(n5417), .ZN(n8208)
         );
  NAND2_X1 U7006 ( .A1(n5322), .A2(n8208), .ZN(n5421) );
  XNOR2_X1 U7007 ( .A(n5423), .B(n5421), .ZN(n7404) );
  INV_X1 U7008 ( .A(n5421), .ZN(n5422) );
  INV_X1 U7009 ( .A(n5427), .ZN(n5428) );
  MUX2_X1 U7010 ( .A(n6295), .B(n6293), .S(n5808), .Z(n5431) );
  INV_X1 U7011 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U7012 ( .A1(n5432), .A2(SI_12_), .ZN(n5433) );
  XNOR2_X1 U7013 ( .A(n5457), .B(n5456), .ZN(n7308) );
  NAND2_X1 U7014 ( .A1(n7308), .A2(n4260), .ZN(n5441) );
  INV_X1 U7015 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5434) );
  AND3_X1 U7016 ( .A1(n5436), .A2(n5435), .A3(n5434), .ZN(n5437) );
  AND2_X1 U7017 ( .A1(n5438), .A2(n5437), .ZN(n5465) );
  OR2_X1 U7018 ( .A1(n5465), .A2(n5168), .ZN(n5439) );
  XNOR2_X1 U7019 ( .A(n5439), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6703) );
  AOI22_X1 U7020 ( .A1(n5909), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5600), .B2(
        n6703), .ZN(n5440) );
  XNOR2_X1 U7021 ( .A(n8002), .B(n5802), .ZN(n5449) );
  NAND2_X1 U7022 ( .A1(n5915), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U7023 ( .A1(n5314), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U7024 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  AND2_X1 U7025 ( .A1(n5470), .A2(n5444), .ZN(n7490) );
  NAND2_X1 U7026 ( .A1(n5794), .A2(n7490), .ZN(n5446) );
  NAND2_X1 U7027 ( .A1(n5757), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5445) );
  NAND4_X1 U7028 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(n8207)
         );
  NAND2_X1 U7029 ( .A1(n5322), .A2(n8207), .ZN(n5450) );
  NAND2_X1 U7030 ( .A1(n5449), .A2(n5450), .ZN(n5454) );
  INV_X1 U7031 ( .A(n5449), .ZN(n5452) );
  INV_X1 U7032 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U7033 ( .A1(n5452), .A2(n5451), .ZN(n5453) );
  NAND2_X1 U7034 ( .A1(n5454), .A2(n5453), .ZN(n7485) );
  MUX2_X1 U7035 ( .A(n6337), .B(n10071), .S(n5504), .Z(n5459) );
  INV_X1 U7036 ( .A(n5459), .ZN(n5460) );
  NAND2_X1 U7037 ( .A1(n5460), .A2(SI_13_), .ZN(n5461) );
  NAND2_X1 U7038 ( .A1(n5481), .A2(n5461), .ZN(n5462) );
  NAND2_X1 U7039 ( .A1(n7511), .A2(n4260), .ZN(n5467) );
  NAND2_X1 U7040 ( .A1(n5465), .A2(n5464), .ZN(n5534) );
  NAND2_X1 U7041 ( .A1(n5534), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5482) );
  XNOR2_X1 U7042 ( .A(n5482), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6845) );
  AOI22_X1 U7043 ( .A1(n5909), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6845), .B2(
        n5600), .ZN(n5466) );
  XNOR2_X1 U7044 ( .A(n8652), .B(n5802), .ZN(n5476) );
  NAND2_X1 U7045 ( .A1(n5915), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7046 ( .A1(n5314), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5474) );
  INV_X1 U7047 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5468) );
  OR2_X1 U7048 ( .A1(n5797), .A2(n5468), .ZN(n5473) );
  INV_X1 U7049 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7050 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  AND2_X1 U7051 ( .A1(n5486), .A2(n5471), .ZN(n8650) );
  NAND2_X1 U7052 ( .A1(n5794), .A2(n8650), .ZN(n5472) );
  NAND4_X1 U7053 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n8619)
         );
  NAND2_X1 U7054 ( .A1(n5322), .A2(n8619), .ZN(n5477) );
  XNOR2_X1 U7055 ( .A(n5476), .B(n5477), .ZN(n7572) );
  INV_X1 U7056 ( .A(n7572), .ZN(n5480) );
  INV_X1 U7057 ( .A(n5476), .ZN(n5479) );
  INV_X1 U7058 ( .A(n5477), .ZN(n5478) );
  MUX2_X1 U7059 ( .A(n6354), .B(n6352), .S(n5504), .Z(n5501) );
  NAND2_X1 U7060 ( .A1(n7582), .A2(n4260), .ZN(n5485) );
  INV_X1 U7061 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7062 ( .A1(n5482), .A2(n5531), .ZN(n5483) );
  NAND2_X1 U7063 ( .A1(n5483), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5510) );
  XNOR2_X1 U7064 ( .A(n5510), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7214) );
  AOI22_X1 U7065 ( .A1(n7214), .A2(n5600), .B1(n5909), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5484) );
  XNOR2_X1 U7066 ( .A(n8746), .B(n5802), .ZN(n5492) );
  INV_X1 U7067 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U7068 ( .A1(n5486), .A2(n6850), .ZN(n5487) );
  AND2_X1 U7069 ( .A1(n5516), .A2(n5487), .ZN(n8616) );
  NAND2_X1 U7070 ( .A1(n8616), .A2(n5794), .ZN(n5491) );
  NAND2_X1 U7071 ( .A1(n5314), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5490) );
  INV_X1 U7072 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7211) );
  OR2_X1 U7073 ( .A1(n5797), .A2(n7211), .ZN(n5489) );
  NAND2_X1 U7074 ( .A1(n5915), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5488) );
  NAND4_X1 U7075 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n8595)
         );
  NAND2_X1 U7076 ( .A1(n5269), .A2(n8595), .ZN(n5493) );
  NAND2_X1 U7077 ( .A1(n5492), .A2(n5493), .ZN(n5497) );
  INV_X1 U7078 ( .A(n5492), .ZN(n5495) );
  INV_X1 U7079 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U7080 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  AND2_X1 U7081 ( .A1(n5497), .A2(n5496), .ZN(n8051) );
  INV_X1 U7082 ( .A(n5501), .ZN(n5502) );
  INV_X1 U7083 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5505) );
  MUX2_X1 U7084 ( .A(n5505), .B(n7677), .S(n5808), .Z(n5507) );
  INV_X1 U7085 ( .A(SI_15_), .ZN(n5506) );
  INV_X1 U7086 ( .A(n5507), .ZN(n5508) );
  NAND2_X1 U7087 ( .A1(n5508), .A2(SI_15_), .ZN(n5509) );
  XNOR2_X1 U7088 ( .A(n5524), .B(n5523), .ZN(n7676) );
  NAND2_X1 U7089 ( .A1(n7676), .A2(n4260), .ZN(n5514) );
  INV_X1 U7090 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7091 ( .A1(n5510), .A2(n5530), .ZN(n5511) );
  NAND2_X1 U7092 ( .A1(n5511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5512) );
  XNOR2_X1 U7093 ( .A(n5512), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8330) );
  AOI22_X1 U7094 ( .A1(n8330), .A2(n5600), .B1(n5909), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5513) );
  XNOR2_X1 U7095 ( .A(n8608), .B(n5802), .ZN(n8100) );
  INV_X1 U7096 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U7097 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  NAND2_X1 U7098 ( .A1(n5539), .A2(n5517), .ZN(n8604) );
  NAND2_X1 U7099 ( .A1(n5314), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7100 ( .A1(n5289), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5518) );
  AND2_X1 U7101 ( .A1(n5519), .A2(n5518), .ZN(n5521) );
  NAND2_X1 U7102 ( .A1(n5915), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5520) );
  OAI211_X1 U7103 ( .C1(n8604), .C2(n5782), .A(n5521), .B(n5520), .ZN(n8626)
         );
  NAND2_X1 U7104 ( .A1(n5269), .A2(n8626), .ZN(n5544) );
  INV_X1 U7105 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5525) );
  MUX2_X1 U7106 ( .A(n5525), .B(n6805), .S(n5808), .Z(n5527) );
  INV_X1 U7107 ( .A(SI_16_), .ZN(n5526) );
  NAND2_X1 U7108 ( .A1(n5527), .A2(n5526), .ZN(n5555) );
  INV_X1 U7109 ( .A(n5527), .ZN(n5528) );
  NAND2_X1 U7110 ( .A1(n5528), .A2(SI_16_), .ZN(n5529) );
  XNOR2_X1 U7111 ( .A(n5554), .B(n5553), .ZN(n7666) );
  NAND2_X1 U7112 ( .A1(n7666), .A2(n4260), .ZN(n5537) );
  NAND3_X1 U7113 ( .A1(n5532), .A2(n5531), .A3(n5530), .ZN(n5533) );
  OAI21_X1 U7114 ( .B1(n5534), .B2(n5533), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5535) );
  XNOR2_X1 U7115 ( .A(n5535), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8346) );
  AOI22_X1 U7116 ( .A1(n8346), .A2(n5600), .B1(n5909), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n5536) );
  XNOR2_X1 U7117 ( .A(n8735), .B(n5236), .ZN(n5549) );
  INV_X1 U7118 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5543) );
  INV_X1 U7119 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7120 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  NAND2_X1 U7121 ( .A1(n5560), .A2(n5540), .ZN(n8109) );
  OR2_X1 U7122 ( .A1(n8109), .A2(n5782), .ZN(n5542) );
  AOI22_X1 U7123 ( .A1(n5314), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n5915), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n5541) );
  OAI211_X1 U7124 ( .C1(n5797), .C2(n5543), .A(n5542), .B(n5541), .ZN(n8597)
         );
  NAND2_X1 U7125 ( .A1(n8597), .A2(n5322), .ZN(n5550) );
  XNOR2_X1 U7126 ( .A(n5549), .B(n5550), .ZN(n8104) );
  INV_X1 U7127 ( .A(n8100), .ZN(n5545) );
  INV_X1 U7128 ( .A(n5544), .ZN(n8102) );
  NAND2_X1 U7129 ( .A1(n5545), .A2(n8102), .ZN(n5546) );
  AND2_X1 U7130 ( .A1(n8104), .A2(n5546), .ZN(n5547) );
  NAND2_X1 U7131 ( .A1(n5548), .A2(n5547), .ZN(n8106) );
  INV_X1 U7132 ( .A(n5549), .ZN(n5551) );
  NAND2_X1 U7133 ( .A1(n5551), .A2(n5550), .ZN(n5552) );
  INV_X1 U7134 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6857) );
  INV_X1 U7135 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10037) );
  MUX2_X1 U7136 ( .A(n6857), .B(n10037), .S(n5808), .Z(n5571) );
  XNOR2_X1 U7137 ( .A(n5571), .B(SI_17_), .ZN(n5570) );
  XNOR2_X1 U7138 ( .A(n5569), .B(n5570), .ZN(n7699) );
  NAND2_X1 U7139 ( .A1(n7699), .A2(n4260), .ZN(n5559) );
  NAND2_X1 U7140 ( .A1(n5149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5557) );
  XNOR2_X1 U7141 ( .A(n5557), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8347) );
  AOI22_X1 U7142 ( .A1(n5909), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5600), .B2(
        n8347), .ZN(n5558) );
  XNOR2_X1 U7143 ( .A(n8731), .B(n5802), .ZN(n5564) );
  INV_X1 U7144 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10193) );
  NAND2_X1 U7145 ( .A1(n5560), .A2(n10193), .ZN(n5561) );
  NAND2_X1 U7146 ( .A1(n5579), .A2(n5561), .ZN(n8569) );
  AOI22_X1 U7147 ( .A1(n5314), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n5757), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7148 ( .A1(n5915), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5562) );
  OAI211_X1 U7149 ( .C1(n8569), .C2(n5782), .A(n5563), .B(n5562), .ZN(n8579)
         );
  NAND2_X1 U7150 ( .A1(n8579), .A2(n5322), .ZN(n5565) );
  XNOR2_X1 U7151 ( .A(n5564), .B(n5565), .ZN(n8116) );
  INV_X1 U7152 ( .A(n5564), .ZN(n5567) );
  INV_X1 U7153 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7154 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  INV_X1 U7155 ( .A(n5571), .ZN(n5572) );
  NAND2_X1 U7156 ( .A1(n5572), .A2(SI_17_), .ZN(n5573) );
  MUX2_X1 U7157 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5808), .Z(n5594) );
  XNOR2_X1 U7158 ( .A(n5594), .B(SI_18_), .ZN(n5591) );
  XNOR2_X1 U7159 ( .A(n5593), .B(n5591), .ZN(n7930) );
  NAND2_X1 U7160 ( .A1(n5574), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5575) );
  XNOR2_X1 U7161 ( .A(n5575), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8361) );
  AOI22_X1 U7162 ( .A1(n5909), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5600), .B2(
        n8361), .ZN(n5576) );
  XNOR2_X1 U7163 ( .A(n8725), .B(n5236), .ZN(n5589) );
  INV_X1 U7164 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7165 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  NAND2_X1 U7166 ( .A1(n5604), .A2(n5580), .ZN(n8551) );
  OR2_X1 U7167 ( .A1(n8551), .A2(n5782), .ZN(n5586) );
  INV_X1 U7168 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7169 ( .A1(n5915), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7170 ( .A1(n5314), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5581) );
  OAI211_X1 U7171 ( .C1(n5583), .C2(n5797), .A(n5582), .B(n5581), .ZN(n5584)
         );
  INV_X1 U7172 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7173 ( .A1(n5586), .A2(n5585), .ZN(n8563) );
  NAND2_X1 U7174 ( .A1(n8563), .A2(n5322), .ZN(n5587) );
  XNOR2_X1 U7175 ( .A(n5589), .B(n5587), .ZN(n8174) );
  INV_X1 U7176 ( .A(n5587), .ZN(n5588) );
  AND2_X1 U7177 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  INV_X1 U7178 ( .A(n5591), .ZN(n5592) );
  NAND2_X1 U7179 ( .A1(n5594), .A2(SI_18_), .ZN(n5595) );
  INV_X1 U7180 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7151) );
  INV_X1 U7181 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7178) );
  MUX2_X1 U7182 ( .A(n7151), .B(n7178), .S(n5808), .Z(n5597) );
  INV_X1 U7183 ( .A(SI_19_), .ZN(n5596) );
  NAND2_X1 U7184 ( .A1(n5597), .A2(n5596), .ZN(n5617) );
  INV_X1 U7185 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7186 ( .A1(n5598), .A2(SI_19_), .ZN(n5599) );
  NAND2_X1 U7187 ( .A1(n5617), .A2(n5599), .ZN(n5618) );
  XNOR2_X1 U7188 ( .A(n5619), .B(n5618), .ZN(n7733) );
  NAND2_X1 U7189 ( .A1(n7733), .A2(n4260), .ZN(n5602) );
  AOI22_X1 U7190 ( .A1(n5909), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5600), .B2(
        n8435), .ZN(n5601) );
  XNOR2_X1 U7191 ( .A(n8721), .B(n5802), .ZN(n5611) );
  INV_X1 U7192 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7193 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U7194 ( .A1(n5626), .A2(n5605), .ZN(n8076) );
  OR2_X1 U7195 ( .A1(n8076), .A2(n5782), .ZN(n5610) );
  INV_X1 U7196 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U7197 ( .A1(n5757), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7198 ( .A1(n5915), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5606) );
  OAI211_X1 U7199 ( .C1(n5862), .C2(n10056), .A(n5607), .B(n5606), .ZN(n5608)
         );
  INV_X1 U7200 ( .A(n5608), .ZN(n5609) );
  NAND2_X1 U7201 ( .A1(n5610), .A2(n5609), .ZN(n8547) );
  NAND2_X1 U7202 ( .A1(n8547), .A2(n5269), .ZN(n5612) );
  NAND2_X1 U7203 ( .A1(n5611), .A2(n5612), .ZN(n5616) );
  INV_X1 U7204 ( .A(n5611), .ZN(n5614) );
  INV_X1 U7205 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7206 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  AND2_X1 U7207 ( .A1(n5616), .A2(n5615), .ZN(n8073) );
  INV_X1 U7208 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7279) );
  INV_X1 U7209 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7749) );
  MUX2_X1 U7210 ( .A(n7279), .B(n7749), .S(n5808), .Z(n5621) );
  INV_X1 U7211 ( .A(SI_20_), .ZN(n5620) );
  NAND2_X1 U7212 ( .A1(n5621), .A2(n5620), .ZN(n5640) );
  INV_X1 U7213 ( .A(n5621), .ZN(n5622) );
  NAND2_X1 U7214 ( .A1(n5622), .A2(SI_20_), .ZN(n5623) );
  XNOR2_X1 U7215 ( .A(n5639), .B(n5638), .ZN(n7748) );
  NAND2_X1 U7216 ( .A1(n7748), .A2(n4260), .ZN(n5625) );
  NAND2_X1 U7217 ( .A1(n5927), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5624) );
  XNOR2_X1 U7218 ( .A(n8714), .B(n5802), .ZN(n5633) );
  INV_X1 U7219 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U7220 ( .A1(n5626), .A2(n8150), .ZN(n5627) );
  NAND2_X1 U7221 ( .A1(n5644), .A2(n5627), .ZN(n8525) );
  INV_X1 U7222 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7223 ( .A1(n5915), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7224 ( .A1(n5757), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5628) );
  OAI211_X1 U7225 ( .C1(n5862), .C2(n5630), .A(n5629), .B(n5628), .ZN(n5631)
         );
  INV_X1 U7226 ( .A(n5631), .ZN(n5632) );
  OAI21_X1 U7227 ( .B1(n8525), .B2(n5782), .A(n5632), .ZN(n8535) );
  NAND2_X1 U7228 ( .A1(n8535), .A2(n5322), .ZN(n5634) );
  XNOR2_X1 U7229 ( .A(n5633), .B(n5634), .ZN(n8148) );
  INV_X1 U7230 ( .A(n5633), .ZN(n5636) );
  INV_X1 U7231 ( .A(n5634), .ZN(n5635) );
  NAND2_X1 U7232 ( .A1(n5636), .A2(n5635), .ZN(n5637) );
  INV_X1 U7233 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7555) );
  INV_X1 U7234 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7774) );
  MUX2_X1 U7235 ( .A(n7555), .B(n7774), .S(n5808), .Z(n5655) );
  XNOR2_X1 U7236 ( .A(n5655), .B(SI_21_), .ZN(n5652) );
  XNOR2_X1 U7237 ( .A(n5654), .B(n5652), .ZN(n7773) );
  NAND2_X1 U7238 ( .A1(n7773), .A2(n4260), .ZN(n5643) );
  NAND2_X1 U7239 ( .A1(n5927), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5642) );
  XNOR2_X1 U7240 ( .A(n8709), .B(n5236), .ZN(n5676) );
  INV_X1 U7241 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U7242 ( .A1(n5644), .A2(n10083), .ZN(n5645) );
  AND2_X1 U7243 ( .A1(n5665), .A2(n5645), .ZN(n8507) );
  NAND2_X1 U7244 ( .A1(n8507), .A2(n5794), .ZN(n5651) );
  INV_X1 U7245 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7246 ( .A1(n5915), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7247 ( .A1(n5289), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5646) );
  OAI211_X1 U7248 ( .C1(n5862), .C2(n5648), .A(n5647), .B(n5646), .ZN(n5649)
         );
  INV_X1 U7249 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7250 ( .A1(n5651), .A2(n5650), .ZN(n8520) );
  NAND2_X1 U7251 ( .A1(n8520), .A2(n5269), .ZN(n5675) );
  XNOR2_X1 U7252 ( .A(n5676), .B(n5675), .ZN(n8083) );
  INV_X1 U7253 ( .A(n5652), .ZN(n5653) );
  INV_X1 U7254 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U7255 ( .A1(n5656), .A2(SI_21_), .ZN(n5657) );
  INV_X1 U7256 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7964) );
  INV_X1 U7257 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7793) );
  MUX2_X1 U7258 ( .A(n7964), .B(n7793), .S(n5808), .Z(n5659) );
  INV_X1 U7259 ( .A(SI_22_), .ZN(n5658) );
  NAND2_X1 U7260 ( .A1(n5659), .A2(n5658), .ZN(n5680) );
  INV_X1 U7261 ( .A(n5659), .ZN(n5660) );
  NAND2_X1 U7262 ( .A1(n5660), .A2(SI_22_), .ZN(n5661) );
  NAND2_X1 U7263 ( .A1(n5680), .A2(n5661), .ZN(n5681) );
  NAND2_X1 U7264 ( .A1(n7792), .A2(n4260), .ZN(n5663) );
  NAND2_X1 U7265 ( .A1(n5927), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5662) );
  INV_X1 U7266 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U7267 ( .A1(n5665), .A2(n8164), .ZN(n5666) );
  NAND2_X1 U7268 ( .A1(n5706), .A2(n5666), .ZN(n8497) );
  INV_X1 U7269 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7270 ( .A1(n5289), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7271 ( .A1(n5915), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5667) );
  OAI211_X1 U7272 ( .C1(n5862), .C2(n5669), .A(n5668), .B(n5667), .ZN(n5670)
         );
  INV_X1 U7273 ( .A(n5670), .ZN(n5671) );
  NAND2_X1 U7274 ( .A1(n8505), .A2(n5269), .ZN(n8161) );
  INV_X1 U7275 ( .A(n5673), .ZN(n8158) );
  INV_X1 U7276 ( .A(n5675), .ZN(n5674) );
  NAND2_X1 U7277 ( .A1(n5676), .A2(n5674), .ZN(n8156) );
  NAND2_X1 U7278 ( .A1(n8156), .A2(n8161), .ZN(n5678) );
  NOR2_X1 U7279 ( .A1(n8086), .A2(n5675), .ZN(n5677) );
  AOI22_X1 U7280 ( .A1(n8158), .A2(n5678), .B1(n5677), .B2(n5676), .ZN(n5679)
         );
  INV_X1 U7281 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5683) );
  INV_X1 U7282 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7822) );
  MUX2_X1 U7283 ( .A(n5683), .B(n7822), .S(n5808), .Z(n5684) );
  INV_X1 U7284 ( .A(SI_23_), .ZN(n10142) );
  NAND2_X1 U7285 ( .A1(n5684), .A2(n10142), .ZN(n5691) );
  INV_X1 U7286 ( .A(n5684), .ZN(n5685) );
  NAND2_X1 U7287 ( .A1(n5685), .A2(SI_23_), .ZN(n5686) );
  XNOR2_X1 U7288 ( .A(n5690), .B(n5689), .ZN(n7821) );
  NAND2_X1 U7289 ( .A1(n7821), .A2(n5216), .ZN(n5688) );
  NAND2_X1 U7290 ( .A1(n5927), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5687) );
  XNOR2_X1 U7291 ( .A(n8696), .B(n5236), .ZN(n5705) );
  INV_X1 U7292 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10169) );
  INV_X1 U7293 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7808) );
  MUX2_X1 U7294 ( .A(n10169), .B(n7808), .S(n5808), .Z(n5718) );
  XNOR2_X1 U7295 ( .A(n5718), .B(SI_24_), .ZN(n5717) );
  NAND2_X1 U7296 ( .A1(n7807), .A2(n4260), .ZN(n5693) );
  NAND2_X1 U7297 ( .A1(n5927), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5692) );
  XNOR2_X1 U7298 ( .A(n8691), .B(n5802), .ZN(n8128) );
  INV_X1 U7299 ( .A(n5694), .ZN(n5708) );
  INV_X1 U7300 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8131) );
  NAND2_X1 U7301 ( .A1(n5708), .A2(n8131), .ZN(n5695) );
  NAND2_X1 U7302 ( .A1(n5727), .A2(n5695), .ZN(n8465) );
  INV_X1 U7303 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7304 ( .A1(n5757), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7305 ( .A1(n5915), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5696) );
  OAI211_X1 U7306 ( .C1(n5862), .C2(n5698), .A(n5697), .B(n5696), .ZN(n5699)
         );
  INV_X1 U7307 ( .A(n5699), .ZN(n5700) );
  NAND2_X1 U7308 ( .A1(n8474), .A2(n5269), .ZN(n8127) );
  NAND2_X1 U7309 ( .A1(n8128), .A2(n8127), .ZN(n5704) );
  INV_X1 U7310 ( .A(n8127), .ZN(n5703) );
  INV_X1 U7311 ( .A(n8128), .ZN(n5702) );
  INV_X1 U7312 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U7313 ( .A1(n5706), .A2(n8059), .ZN(n5707) );
  NAND2_X1 U7314 ( .A1(n8478), .A2(n5794), .ZN(n5715) );
  INV_X1 U7315 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7316 ( .A1(n5915), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7317 ( .A1(n5289), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5710) );
  OAI211_X1 U7318 ( .C1(n5862), .C2(n5712), .A(n5711), .B(n5710), .ZN(n5713)
         );
  INV_X1 U7319 ( .A(n5713), .ZN(n5714) );
  NAND2_X1 U7320 ( .A1(n5715), .A2(n5714), .ZN(n8492) );
  NAND2_X1 U7321 ( .A1(n8492), .A2(n5269), .ZN(n8058) );
  AOI21_X1 U7322 ( .B1(n8128), .B2(n8061), .A(n8058), .ZN(n5716) );
  INV_X1 U7323 ( .A(n5717), .ZN(n5741) );
  INV_X1 U7324 ( .A(n5718), .ZN(n5719) );
  NAND2_X1 U7325 ( .A1(n5719), .A2(SI_24_), .ZN(n5744) );
  INV_X1 U7326 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8810) );
  INV_X1 U7327 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7966) );
  MUX2_X1 U7328 ( .A(n8810), .B(n7966), .S(n5808), .Z(n5721) );
  INV_X1 U7329 ( .A(SI_25_), .ZN(n5720) );
  NAND2_X1 U7330 ( .A1(n5721), .A2(n5720), .ZN(n5740) );
  INV_X1 U7331 ( .A(n5721), .ZN(n5722) );
  NAND2_X1 U7332 ( .A1(n5722), .A2(SI_25_), .ZN(n5723) );
  NAND2_X1 U7333 ( .A1(n5740), .A2(n5723), .ZN(n5743) );
  NAND2_X1 U7334 ( .A1(n7965), .A2(n4260), .ZN(n5726) );
  NAND2_X1 U7335 ( .A1(n5927), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5725) );
  XNOR2_X1 U7336 ( .A(n8688), .B(n5236), .ZN(n5737) );
  INV_X1 U7337 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8094) );
  OR2_X2 U7338 ( .A1(n5727), .A2(n8094), .ZN(n5755) );
  NAND2_X1 U7339 ( .A1(n5727), .A2(n8094), .ZN(n5728) );
  NAND2_X1 U7340 ( .A1(n8450), .A2(n5794), .ZN(n5734) );
  INV_X1 U7341 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10163) );
  NAND2_X1 U7342 ( .A1(n5757), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U7343 ( .A1(n5314), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5730) );
  OAI211_X1 U7344 ( .C1(n5247), .C2(n10163), .A(n5731), .B(n5730), .ZN(n5732)
         );
  INV_X1 U7345 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U7346 ( .A1(n8459), .A2(n5322), .ZN(n5735) );
  XNOR2_X1 U7347 ( .A(n5737), .B(n5735), .ZN(n8091) );
  NAND2_X1 U7348 ( .A1(n8092), .A2(n8091), .ZN(n5739) );
  INV_X1 U7349 ( .A(n5735), .ZN(n5736) );
  NAND2_X1 U7350 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  INV_X1 U7351 ( .A(n5740), .ZN(n5747) );
  INV_X1 U7352 ( .A(n5743), .ZN(n5745) );
  AND2_X1 U7353 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  INV_X1 U7354 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5748) );
  INV_X1 U7355 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9744) );
  MUX2_X1 U7356 ( .A(n5748), .B(n9744), .S(n5808), .Z(n5750) );
  INV_X1 U7357 ( .A(SI_26_), .ZN(n5749) );
  NAND2_X1 U7358 ( .A1(n5750), .A2(n5749), .ZN(n5771) );
  INV_X1 U7359 ( .A(n5750), .ZN(n5751) );
  NAND2_X1 U7360 ( .A1(n5751), .A2(SI_26_), .ZN(n5752) );
  NAND2_X1 U7361 ( .A1(n8804), .A2(n4260), .ZN(n5754) );
  NAND2_X1 U7362 ( .A1(n5927), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5753) );
  XNOR2_X1 U7363 ( .A(n8680), .B(n5236), .ZN(n5766) );
  INV_X1 U7364 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U7365 ( .A1(n5755), .A2(n8183), .ZN(n5756) );
  NAND2_X1 U7366 ( .A1(n8433), .A2(n5794), .ZN(n5763) );
  INV_X1 U7367 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U7368 ( .A1(n5757), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U7369 ( .A1(n5915), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5758) );
  OAI211_X1 U7370 ( .C1(n5862), .C2(n5760), .A(n5759), .B(n5758), .ZN(n5761)
         );
  INV_X1 U7371 ( .A(n5761), .ZN(n5762) );
  NAND2_X1 U7372 ( .A1(n8206), .A2(n5269), .ZN(n5764) );
  XNOR2_X1 U7373 ( .A(n5766), .B(n5764), .ZN(n8181) );
  INV_X1 U7374 ( .A(n5764), .ZN(n5765) );
  INV_X1 U7375 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5773) );
  INV_X1 U7376 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7862) );
  MUX2_X1 U7377 ( .A(n5773), .B(n7862), .S(n5808), .Z(n5775) );
  INV_X1 U7378 ( .A(SI_27_), .ZN(n5774) );
  NAND2_X1 U7379 ( .A1(n5775), .A2(n5774), .ZN(n5806) );
  INV_X1 U7380 ( .A(n5775), .ZN(n5776) );
  NAND2_X1 U7381 ( .A1(n5776), .A2(SI_27_), .ZN(n5777) );
  NAND2_X1 U7382 ( .A1(n8801), .A2(n5216), .ZN(n5779) );
  NAND2_X1 U7383 ( .A1(n5927), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5778) );
  XNOR2_X1 U7384 ( .A(n8675), .B(n5236), .ZN(n5790) );
  INV_X1 U7385 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8044) );
  NAND2_X1 U7386 ( .A1(n5780), .A2(n8044), .ZN(n5781) );
  NAND2_X1 U7387 ( .A1(n5792), .A2(n5781), .ZN(n8406) );
  INV_X1 U7388 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7389 ( .A1(n5915), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7390 ( .A1(n5314), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5783) );
  OAI211_X1 U7391 ( .C1(n5785), .C2(n5797), .A(n5784), .B(n5783), .ZN(n5786)
         );
  INV_X1 U7392 ( .A(n5786), .ZN(n5787) );
  NAND2_X1 U7393 ( .A1(n8398), .A2(n5269), .ZN(n5788) );
  XNOR2_X1 U7394 ( .A(n5790), .B(n5788), .ZN(n8043) );
  INV_X1 U7395 ( .A(n5788), .ZN(n5789) );
  INV_X1 U7396 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5791) );
  OR2_X2 U7397 ( .A1(n5792), .A2(n5791), .ZN(n5858) );
  NAND2_X1 U7398 ( .A1(n5792), .A2(n5791), .ZN(n5793) );
  NAND2_X1 U7399 ( .A1(n8392), .A2(n5794), .ZN(n5801) );
  INV_X1 U7400 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7401 ( .A1(n5915), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7402 ( .A1(n5314), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5795) );
  OAI211_X1 U7403 ( .C1(n5798), .C2(n5797), .A(n5796), .B(n5795), .ZN(n5799)
         );
  INV_X1 U7404 ( .A(n5799), .ZN(n5800) );
  NAND2_X1 U7405 ( .A1(n8205), .A2(n5322), .ZN(n5803) );
  XNOR2_X1 U7406 ( .A(n5803), .B(n5802), .ZN(n5855) );
  INV_X1 U7407 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5809) );
  INV_X1 U7408 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10133) );
  MUX2_X1 U7409 ( .A(n5809), .B(n10133), .S(n5808), .Z(n5897) );
  XNOR2_X1 U7410 ( .A(n5897), .B(SI_28_), .ZN(n5894) );
  NAND2_X1 U7411 ( .A1(n5927), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5810) );
  INV_X1 U7412 ( .A(n8670), .ZN(n8394) );
  INV_X1 U7413 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7414 ( .A1(n5812), .A2(n5818), .ZN(n5813) );
  NAND2_X1 U7415 ( .A1(n5813), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5847) );
  INV_X1 U7416 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U7417 ( .A1(n5847), .A2(n5846), .ZN(n5849) );
  NAND2_X1 U7418 ( .A1(n5849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5814) );
  INV_X1 U7419 ( .A(P2_B_REG_SCAN_IN), .ZN(n5815) );
  XNOR2_X1 U7420 ( .A(n7603), .B(n5815), .ZN(n5825) );
  INV_X1 U7421 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5817) );
  NAND3_X1 U7422 ( .A1(n5818), .A2(n5846), .A3(n5817), .ZN(n5819) );
  INV_X1 U7423 ( .A(n5823), .ZN(n5820) );
  NAND2_X1 U7424 ( .A1(n5820), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5821) );
  MUX2_X1 U7425 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5821), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5824) );
  INV_X1 U7426 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7427 ( .A1(n5823), .A2(n5822), .ZN(n5826) );
  NAND2_X1 U7428 ( .A1(n5824), .A2(n5826), .ZN(n8808) );
  NAND2_X1 U7429 ( .A1(n5825), .A2(n8808), .ZN(n5830) );
  NAND2_X1 U7430 ( .A1(n5826), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5827) );
  MUX2_X1 U7431 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5827), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5829) );
  INV_X1 U7432 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U7433 ( .A1(n9929), .A2(n9933), .ZN(n5831) );
  OR2_X1 U7434 ( .A1(n8806), .A2(n7603), .ZN(n9932) );
  NOR4_X1 U7435 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5835) );
  NOR4_X1 U7436 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5834) );
  NOR4_X1 U7437 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5833) );
  NOR4_X1 U7438 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5832) );
  AND4_X1 U7439 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n5841)
         );
  NOR2_X1 U7440 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5839) );
  NOR4_X1 U7441 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5838) );
  NOR4_X1 U7442 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5837) );
  NOR4_X1 U7443 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5836) );
  AND4_X1 U7444 ( .A1(n5839), .A2(n5838), .A3(n5837), .A4(n5836), .ZN(n5840)
         );
  NAND2_X1 U7445 ( .A1(n5841), .A2(n5840), .ZN(n5842) );
  INV_X1 U7446 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U7447 ( .A1(n9929), .A2(n9936), .ZN(n5844) );
  INV_X1 U7448 ( .A(n8808), .ZN(n5845) );
  NOR2_X1 U7449 ( .A1(n8806), .A2(n5845), .ZN(n9937) );
  INV_X1 U7450 ( .A(n9937), .ZN(n5843) );
  NAND2_X1 U7451 ( .A1(n5844), .A2(n5843), .ZN(n6917) );
  NAND3_X1 U7452 ( .A1(n8806), .A2(n7603), .A3(n5845), .ZN(n6397) );
  OR2_X1 U7453 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  NAND2_X1 U7454 ( .A1(n5849), .A2(n5848), .ZN(n5931) );
  NAND2_X1 U7455 ( .A1(n5931), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9930) );
  AND2_X1 U7456 ( .A1(n4955), .A2(n6553), .ZN(n6929) );
  NAND2_X1 U7457 ( .A1(n5866), .A2(n6929), .ZN(n5850) );
  NOR3_X1 U7458 ( .A1(n8394), .A2(n5855), .A3(n8197), .ZN(n5851) );
  AOI21_X1 U7459 ( .B1(n5855), .B2(n8394), .A(n5851), .ZN(n5857) );
  NAND2_X1 U7460 ( .A1(n8670), .A2(n8197), .ZN(n5853) );
  AND2_X1 U7461 ( .A1(n7278), .A2(n4954), .ZN(n5870) );
  NAND2_X1 U7462 ( .A1(n6554), .A2(n5972), .ZN(n6204) );
  AND2_X1 U7463 ( .A1(n9985), .A2(n6204), .ZN(n5852) );
  NAND3_X1 U7464 ( .A1(n8670), .A2(n5855), .A3(n8115), .ZN(n5854) );
  OAI21_X1 U7465 ( .B1(n8670), .B2(n5855), .A(n5854), .ZN(n5856) );
  INV_X1 U7466 ( .A(n5858), .ZN(n8037) );
  NAND2_X1 U7467 ( .A1(n8037), .A2(n5794), .ZN(n5865) );
  INV_X1 U7468 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7469 ( .A1(n5915), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7470 ( .A1(n5289), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5859) );
  OAI211_X1 U7471 ( .C1(n5862), .C2(n5861), .A(n5860), .B(n5859), .ZN(n5863)
         );
  INV_X1 U7472 ( .A(n5863), .ZN(n5864) );
  NAND2_X1 U7473 ( .A1(n5865), .A2(n5864), .ZN(n8399) );
  INV_X1 U7474 ( .A(n6204), .ZN(n6393) );
  AND2_X2 U7475 ( .A1(n6393), .A2(n6410), .ZN(n8596) );
  INV_X1 U7476 ( .A(n6410), .ZN(n5868) );
  AND2_X2 U7477 ( .A1(n6393), .A2(n5868), .ZN(n9910) );
  AOI22_X1 U7478 ( .A1(n8399), .A2(n8191), .B1(n8398), .B2(n8192), .ZN(n5874)
         );
  NAND2_X1 U7479 ( .A1(n5869), .A2(n6545), .ZN(n6609) );
  OR2_X1 U7480 ( .A1(n6204), .A2(n5870), .ZN(n6083) );
  AND3_X1 U7481 ( .A1(n6397), .A2(n5931), .A3(n6083), .ZN(n5871) );
  NAND2_X1 U7482 ( .A1(n6609), .A2(n5871), .ZN(n5872) );
  INV_X2 U7483 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AOI22_X1 U7484 ( .A1(n8392), .A2(n8186), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5873) );
  NAND2_X1 U7485 ( .A1(n5875), .A2(n5127), .ZN(P2_U3222) );
  INV_X1 U7486 ( .A(n8215), .ZN(n6942) );
  INV_X1 U7487 ( .A(n9965), .ZN(n9898) );
  AND2_X1 U7488 ( .A1(n8215), .A2(n9965), .ZN(n5939) );
  AND2_X1 U7489 ( .A1(n9974), .A2(n8214), .ZN(n7201) );
  AOI21_X1 U7490 ( .B1(n5939), .B2(n7200), .A(n7201), .ZN(n5876) );
  INV_X1 U7491 ( .A(n8213), .ZN(n6825) );
  OR2_X1 U7492 ( .A1(n6825), .A2(n7193), .ZN(n5992) );
  NAND2_X1 U7493 ( .A1(n7193), .A2(n6825), .ZN(n6957) );
  INV_X1 U7494 ( .A(n8212), .ZN(n7206) );
  NAND2_X1 U7495 ( .A1(n7378), .A2(n7206), .ZN(n5996) );
  INV_X1 U7497 ( .A(n6957), .ZN(n5877) );
  NOR2_X1 U7498 ( .A1(n7377), .A2(n5877), .ZN(n5878) );
  OAI21_X1 U7499 ( .B1(n5981), .B2(n5882), .A(n5878), .ZN(n5879) );
  INV_X1 U7500 ( .A(n5879), .ZN(n5884) );
  INV_X1 U7501 ( .A(n8218), .ZN(n5880) );
  NAND2_X1 U7502 ( .A1(n5880), .A2(n6931), .ZN(n7025) );
  NAND2_X1 U7503 ( .A1(n6938), .A2(n9915), .ZN(n5977) );
  NAND2_X1 U7504 ( .A1(n8216), .A2(n9948), .ZN(n5978) );
  AND2_X2 U7505 ( .A1(n5977), .A2(n5978), .ZN(n9922) );
  NAND2_X1 U7506 ( .A1(n9909), .A2(n7054), .ZN(n5990) );
  INV_X1 U7507 ( .A(n7058), .ZN(n5983) );
  NAND2_X1 U7508 ( .A1(n7059), .A2(n5983), .ZN(n5881) );
  NAND2_X1 U7509 ( .A1(n6954), .A2(n6955), .ZN(n5883) );
  OR2_X1 U7510 ( .A1(n7471), .A2(n5885), .ZN(n6000) );
  NAND2_X1 U7511 ( .A1(n6000), .A2(n6001), .ZN(n7474) );
  INV_X1 U7512 ( .A(n8210), .ZN(n6912) );
  AND2_X1 U7513 ( .A1(n8764), .A2(n6912), .ZN(n5938) );
  NAND2_X1 U7514 ( .A1(n8759), .A2(n7375), .ZN(n6005) );
  NOR2_X1 U7515 ( .A1(n8759), .A2(n7375), .ZN(n5943) );
  INV_X1 U7516 ( .A(n8208), .ZN(n7434) );
  OR2_X1 U7517 ( .A1(n7437), .A2(n7434), .ZN(n6010) );
  INV_X1 U7518 ( .A(n8207), .ZN(n8642) );
  NAND2_X1 U7519 ( .A1(n8002), .A2(n8642), .ZN(n6012) );
  NAND2_X1 U7520 ( .A1(n7437), .A2(n7434), .ZN(n7428) );
  AND2_X1 U7521 ( .A1(n6012), .A2(n7428), .ZN(n6014) );
  INV_X1 U7522 ( .A(n8619), .ZN(n7433) );
  OR2_X1 U7523 ( .A1(n8652), .A2(n7433), .ZN(n6022) );
  NAND2_X1 U7524 ( .A1(n8652), .A2(n7433), .ZN(n6021) );
  NAND2_X1 U7525 ( .A1(n6022), .A2(n6021), .ZN(n8635) );
  NAND2_X1 U7526 ( .A1(n8746), .A2(n8639), .ZN(n6027) );
  NAND2_X1 U7527 ( .A1(n6028), .A2(n6027), .ZN(n8623) );
  INV_X1 U7528 ( .A(n8626), .ZN(n8110) );
  NAND2_X1 U7529 ( .A1(n8608), .A2(n8110), .ZN(n6033) );
  INV_X1 U7530 ( .A(n8597), .ZN(n8119) );
  NAND2_X1 U7531 ( .A1(n8735), .A2(n8119), .ZN(n5966) );
  INV_X1 U7532 ( .A(n8579), .ZN(n8111) );
  NAND2_X1 U7533 ( .A1(n8731), .A2(n8111), .ZN(n5962) );
  INV_X1 U7534 ( .A(n8563), .ZN(n8118) );
  NAND2_X1 U7535 ( .A1(n8725), .A2(n8118), .ZN(n6044) );
  INV_X1 U7536 ( .A(n8547), .ZN(n8151) );
  OR2_X1 U7537 ( .A1(n8721), .A2(n8151), .ZN(n6047) );
  NAND2_X1 U7538 ( .A1(n8721), .A2(n8151), .ZN(n6043) );
  NAND2_X1 U7539 ( .A1(n6047), .A2(n6043), .ZN(n8533) );
  INV_X1 U7540 ( .A(n8535), .ZN(n8085) );
  NAND2_X1 U7541 ( .A1(n8714), .A2(n8085), .ZN(n6050) );
  XNOR2_X1 U7542 ( .A(n8709), .B(n8520), .ZN(n8510) );
  INV_X1 U7543 ( .A(n8520), .ZN(n8168) );
  NAND2_X1 U7544 ( .A1(n8709), .A2(n8168), .ZN(n6049) );
  NAND2_X1 U7545 ( .A1(n8703), .A2(n8086), .ZN(n6038) );
  NAND2_X1 U7546 ( .A1(n8696), .A2(n8165), .ZN(n6040) );
  NAND2_X1 U7547 ( .A1(n8688), .A2(n8132), .ZN(n6062) );
  NAND2_X1 U7548 ( .A1(n8691), .A2(n8061), .ZN(n5959) );
  NAND2_X1 U7549 ( .A1(n6062), .A2(n5959), .ZN(n5891) );
  NAND2_X1 U7550 ( .A1(n8680), .A2(n8412), .ZN(n6063) );
  NOR2_X1 U7551 ( .A1(n8691), .A2(n8061), .ZN(n5937) );
  NAND2_X1 U7552 ( .A1(n6062), .A2(n5937), .ZN(n5888) );
  NAND2_X1 U7553 ( .A1(n5888), .A2(n8425), .ZN(n5889) );
  NOR2_X1 U7554 ( .A1(n8426), .A2(n5889), .ZN(n5890) );
  INV_X1 U7555 ( .A(n8398), .ZN(n5893) );
  NAND2_X1 U7556 ( .A1(n8675), .A2(n5893), .ZN(n5955) );
  INV_X2 U7557 ( .A(n8205), .ZN(n8413) );
  NAND2_X1 U7558 ( .A1(n8670), .A2(n8413), .ZN(n5956) );
  INV_X1 U7559 ( .A(SI_28_), .ZN(n5896) );
  NAND2_X1 U7560 ( .A1(n5897), .A2(n5896), .ZN(n5898) );
  INV_X1 U7561 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9734) );
  INV_X1 U7562 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8796) );
  MUX2_X1 U7563 ( .A(n9734), .B(n8796), .S(n6455), .Z(n5903) );
  XNOR2_X1 U7564 ( .A(n5903), .B(SI_29_), .ZN(n5900) );
  NAND2_X1 U7565 ( .A1(n5927), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5901) );
  INV_X1 U7566 ( .A(n8399), .ZN(n6068) );
  INV_X1 U7567 ( .A(n5903), .ZN(n5906) );
  NOR2_X1 U7568 ( .A1(n5906), .A2(SI_29_), .ZN(n5904) );
  NAND2_X1 U7569 ( .A1(n5906), .A2(SI_29_), .ZN(n5920) );
  MUX2_X1 U7570 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6455), .Z(n5922) );
  XNOR2_X1 U7571 ( .A(n5922), .B(SI_30_), .ZN(n5907) );
  NAND2_X1 U7572 ( .A1(n5909), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7573 ( .A1(n5314), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5914) );
  NAND2_X1 U7574 ( .A1(n5289), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7575 ( .A1(n5915), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5912) );
  AND3_X1 U7576 ( .A1(n5914), .A2(n5913), .A3(n5912), .ZN(n8377) );
  NAND2_X1 U7577 ( .A1(n5314), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7578 ( .A1(n5757), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7579 ( .A1(n5915), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5916) );
  AND3_X1 U7580 ( .A1(n5918), .A2(n5917), .A3(n5916), .ZN(n8030) );
  OR2_X1 U7581 ( .A1(n5030), .A2(n8030), .ZN(n5935) );
  NAND2_X1 U7582 ( .A1(n5922), .A2(SI_30_), .ZN(n5919) );
  INV_X1 U7583 ( .A(n5922), .ZN(n5923) );
  INV_X1 U7584 ( .A(SI_30_), .ZN(n10055) );
  NAND2_X1 U7585 ( .A1(n5923), .A2(n10055), .ZN(n5924) );
  MUX2_X1 U7586 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6455), .Z(n5925) );
  INV_X1 U7587 ( .A(SI_31_), .ZN(n10070) );
  XNOR2_X1 U7588 ( .A(n5925), .B(n10070), .ZN(n5926) );
  NAND2_X1 U7589 ( .A1(n5927), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7590 ( .A1(n5030), .A2(n8030), .ZN(n5930) );
  NOR2_X1 U7591 ( .A1(n7554), .A2(n7278), .ZN(n6548) );
  NOR2_X1 U7592 ( .A1(n5931), .A2(P2_U3152), .ZN(n7540) );
  AND2_X1 U7593 ( .A1(n5932), .A2(n7540), .ZN(n5933) );
  NAND2_X1 U7594 ( .A1(n5934), .A2(n5933), .ZN(n6089) );
  INV_X1 U7595 ( .A(n5937), .ZN(n8424) );
  INV_X1 U7596 ( .A(n8488), .ZN(n8486) );
  NAND2_X1 U7597 ( .A1(n6046), .A2(n6050), .ZN(n8517) );
  INV_X1 U7598 ( .A(n8554), .ZN(n8545) );
  NAND2_X1 U7599 ( .A1(n5965), .A2(n5966), .ZN(n8573) );
  NOR2_X1 U7600 ( .A1(n8601), .A2(n8623), .ZN(n6026) );
  NAND2_X1 U7601 ( .A1(n6015), .A2(n6012), .ZN(n7430) );
  INV_X1 U7602 ( .A(n7474), .ZN(n7467) );
  INV_X1 U7603 ( .A(n5938), .ZN(n6004) );
  INV_X1 U7604 ( .A(n6931), .ZN(n7032) );
  NAND2_X1 U7605 ( .A1(n8218), .A2(n7032), .ZN(n6716) );
  NAND2_X1 U7606 ( .A1(n7025), .A2(n6716), .ZN(n6925) );
  NOR4_X1 U7607 ( .A1(n6937), .A2(n6925), .A3(n7037), .A4(n7278), .ZN(n5940)
         );
  NAND3_X1 U7608 ( .A1(n5940), .A2(n5983), .A3(n9903), .ZN(n5941) );
  INV_X1 U7609 ( .A(n7201), .ZN(n5991) );
  NAND2_X1 U7610 ( .A1(n7200), .A2(n5991), .ZN(n7184) );
  NOR4_X1 U7611 ( .A1(n5941), .A2(n7377), .A3(n7203), .A4(n7184), .ZN(n5942)
         );
  NAND4_X1 U7612 ( .A1(n7383), .A2(n7467), .A3(n7499), .A4(n5942), .ZN(n5944)
         );
  INV_X1 U7613 ( .A(n5943), .ZN(n6008) );
  NAND2_X1 U7614 ( .A1(n6008), .A2(n6005), .ZN(n7389) );
  NOR4_X1 U7615 ( .A1(n8635), .A2(n7430), .A3(n5944), .A4(n7389), .ZN(n5945)
         );
  NAND4_X1 U7616 ( .A1(n8010), .A2(n8575), .A3(n6026), .A4(n5945), .ZN(n5946)
         );
  NOR4_X1 U7617 ( .A1(n8517), .A2(n8533), .A3(n8545), .A4(n5946), .ZN(n5947)
         );
  NAND4_X1 U7618 ( .A1(n8464), .A2(n8486), .A3(n5947), .A4(n8510), .ZN(n5948)
         );
  NOR4_X1 U7619 ( .A1(n8426), .A2(n8021), .A3(n5948), .A4(n8482), .ZN(n5949)
         );
  NAND3_X1 U7620 ( .A1(n8396), .A2(n4890), .A3(n5949), .ZN(n5950) );
  OAI22_X1 U7621 ( .A1(n5951), .A2(n5972), .B1(n6553), .B2(n6550), .ZN(n6082)
         );
  NAND2_X1 U7622 ( .A1(n6074), .A2(n6070), .ZN(n5952) );
  AND2_X1 U7623 ( .A1(n5956), .A2(n6079), .ZN(n5953) );
  NAND2_X1 U7624 ( .A1(n5954), .A2(n5953), .ZN(n6073) );
  AND2_X1 U7625 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  MUX2_X1 U7626 ( .A(n5958), .B(n5957), .S(n6070), .Z(n6067) );
  NAND2_X1 U7627 ( .A1(n8425), .A2(n8424), .ZN(n5961) );
  INV_X1 U7628 ( .A(n5959), .ZN(n5960) );
  INV_X1 U7629 ( .A(n6038), .ZN(n6039) );
  INV_X1 U7630 ( .A(n5962), .ZN(n5964) );
  INV_X1 U7631 ( .A(n5966), .ZN(n5967) );
  MUX2_X1 U7632 ( .A(n5042), .B(n5967), .S(n6070), .Z(n5968) );
  INV_X1 U7633 ( .A(n5968), .ZN(n6035) );
  INV_X1 U7634 ( .A(n8635), .ZN(n8631) );
  NAND2_X1 U7635 ( .A1(n7428), .A2(n6005), .ZN(n5971) );
  NAND2_X1 U7636 ( .A1(n6005), .A2(n4833), .ZN(n5969) );
  NAND3_X1 U7637 ( .A1(n5969), .A2(n6008), .A3(n6010), .ZN(n5970) );
  MUX2_X1 U7638 ( .A(n5971), .B(n5970), .S(n6070), .Z(n6020) );
  AND2_X1 U7639 ( .A1(n6716), .A2(n5972), .ZN(n5973) );
  OAI211_X1 U7640 ( .C1(n7029), .C2(n5973), .A(n7024), .B(n5978), .ZN(n5974)
         );
  NAND2_X1 U7641 ( .A1(n6716), .A2(n7024), .ZN(n5976) );
  NAND3_X1 U7642 ( .A1(n5977), .A2(n5976), .A3(n5975), .ZN(n5979) );
  NAND2_X1 U7643 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  NAND2_X1 U7644 ( .A1(n5991), .A2(n4689), .ZN(n5982) );
  INV_X1 U7645 ( .A(n5994), .ZN(n5984) );
  AND2_X1 U7646 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  OAI211_X1 U7647 ( .C1(n5994), .C2(n5987), .A(n7200), .B(n6957), .ZN(n5988)
         );
  NAND2_X1 U7648 ( .A1(n5988), .A2(n6070), .ZN(n5989) );
  AND2_X1 U7649 ( .A1(n4689), .A2(n5990), .ZN(n5993) );
  OAI211_X1 U7650 ( .C1(n5994), .C2(n5993), .A(n5992), .B(n5991), .ZN(n5995)
         );
  MUX2_X1 U7651 ( .A(n5997), .B(n5996), .S(n6070), .Z(n5998) );
  NAND3_X1 U7652 ( .A1(n5999), .A2(n7467), .A3(n5998), .ZN(n6003) );
  MUX2_X1 U7653 ( .A(n6001), .B(n6000), .S(n6070), .Z(n6002) );
  NAND2_X1 U7654 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  NAND2_X1 U7655 ( .A1(n6006), .A2(n6070), .ZN(n6007) );
  INV_X1 U7656 ( .A(n6010), .ZN(n6011) );
  NAND2_X1 U7657 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  AND2_X1 U7658 ( .A1(n6013), .A2(n6015), .ZN(n6018) );
  INV_X1 U7659 ( .A(n6014), .ZN(n6016) );
  NAND2_X1 U7660 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  MUX2_X1 U7661 ( .A(n6018), .B(n6017), .S(n6070), .Z(n6019) );
  INV_X1 U7662 ( .A(n6021), .ZN(n6024) );
  INV_X1 U7663 ( .A(n6022), .ZN(n6023) );
  MUX2_X1 U7664 ( .A(n6024), .B(n6023), .S(n6079), .Z(n6025) );
  INV_X1 U7665 ( .A(n6027), .ZN(n6030) );
  INV_X1 U7666 ( .A(n6028), .ZN(n6029) );
  MUX2_X1 U7667 ( .A(n6030), .B(n6029), .S(n6070), .Z(n6031) );
  MUX2_X1 U7668 ( .A(n6033), .B(n6032), .S(n6070), .Z(n6034) );
  NAND2_X1 U7669 ( .A1(n6050), .A2(n6043), .ZN(n6037) );
  OR2_X1 U7670 ( .A1(n8709), .A2(n8168), .ZN(n6052) );
  NAND2_X1 U7671 ( .A1(n6042), .A2(n6041), .ZN(n6045) );
  NAND3_X1 U7672 ( .A1(n6045), .A2(n6044), .A3(n6043), .ZN(n6048) );
  NAND3_X1 U7673 ( .A1(n6048), .A2(n6047), .A3(n6046), .ZN(n6051) );
  NAND3_X1 U7674 ( .A1(n6051), .A2(n6050), .A3(n6049), .ZN(n6054) );
  NAND4_X1 U7675 ( .A1(n6054), .A2(n6053), .A3(n6079), .A4(n6052), .ZN(n6055)
         );
  OR3_X1 U7676 ( .A1(n8696), .A2(n8165), .A3(n6070), .ZN(n6056) );
  AOI21_X1 U7677 ( .B1(n6057), .B2(n6056), .A(n8018), .ZN(n6060) );
  OAI21_X1 U7678 ( .B1(n8425), .B2(n6079), .A(n6062), .ZN(n6058) );
  INV_X1 U7679 ( .A(n6058), .ZN(n6059) );
  AOI21_X1 U7680 ( .B1(n6063), .B2(n6062), .A(n6079), .ZN(n6066) );
  NAND2_X1 U7681 ( .A1(n4803), .A2(n6070), .ZN(n6065) );
  INV_X1 U7682 ( .A(n8030), .ZN(n8204) );
  NAND3_X1 U7683 ( .A1(n8666), .A2(n6068), .A3(n6070), .ZN(n6069) );
  OAI21_X1 U7684 ( .B1(n5033), .B2(n6070), .A(n6069), .ZN(n6071) );
  INV_X1 U7685 ( .A(n6071), .ZN(n6072) );
  INV_X1 U7686 ( .A(n6075), .ZN(n6076) );
  AOI21_X1 U7687 ( .B1(n6078), .B2(n4312), .A(n6076), .ZN(n6081) );
  INV_X1 U7688 ( .A(n7540), .ZN(n6395) );
  INV_X1 U7689 ( .A(n6083), .ZN(n6084) );
  NOR2_X1 U7690 ( .A1(n6394), .A2(n6084), .ZN(n6608) );
  NOR2_X1 U7691 ( .A1(n6619), .A2(P2_U3152), .ZN(n8802) );
  NAND3_X1 U7692 ( .A1(n6608), .A2(n9910), .A3(n8802), .ZN(n6085) );
  OAI211_X1 U7693 ( .C1(n6554), .C2(n6395), .A(n6085), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6086) );
  NAND2_X1 U7694 ( .A1(n6093), .A2(n6133), .ZN(n6165) );
  NOR2_X1 U7695 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6096) );
  NOR2_X1 U7696 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6123) );
  INV_X1 U7697 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6097) );
  NAND3_X1 U7698 ( .A1(n6123), .A2(n6113), .A3(n6097), .ZN(n6104) );
  NAND3_X1 U7699 ( .A1(n6108), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_24__SCAN_IN), .ZN(n6103) );
  INV_X1 U7700 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7701 ( .A1(n6113), .A2(n6114), .ZN(n6109) );
  INV_X1 U7702 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7703 ( .A1(n6099), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n6101) );
  XNOR2_X1 U7704 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_24__SCAN_IN), .ZN(
        n6100) );
  OAI21_X1 U7705 ( .B1(n6109), .B2(n6101), .A(n6100), .ZN(n6102) );
  NAND2_X1 U7706 ( .A1(n6105), .A2(n10084), .ZN(n6106) );
  NAND2_X1 U7707 ( .A1(n6106), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7708 ( .A1(n6109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7709 ( .A1(n6116), .A2(n6110), .ZN(n6111) );
  XNOR2_X1 U7710 ( .A(n6111), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7551) );
  INV_X1 U7711 ( .A(n7551), .ZN(n6112) );
  NOR2_X1 U7712 ( .A1(n6482), .A2(n6112), .ZN(n6200) );
  NOR2_X2 U7713 ( .A1(n6397), .A2(n9930), .ZN(P2_U3966) );
  NAND2_X1 U7714 ( .A1(n6116), .A2(n6113), .ZN(n6118) );
  NAND2_X1 U7715 ( .A1(n6118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6115) );
  INV_X1 U7716 ( .A(n6116), .ZN(n6117) );
  NAND2_X1 U7717 ( .A1(n6117), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7718 ( .A1(n9057), .A2(n9259), .ZN(n9226) );
  NAND2_X1 U7719 ( .A1(n6482), .A2(n9226), .ZN(n6120) );
  NAND2_X1 U7720 ( .A1(n6120), .A2(n7551), .ZN(n6196) );
  NOR2_X1 U7721 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n6122) );
  NOR2_X1 U7722 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6121) );
  INV_X1 U7723 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6124) );
  XNOR2_X2 U7724 ( .A(n6125), .B(n6124), .ZN(n9055) );
  NAND2_X1 U7725 ( .A1(n6196), .A2(n7678), .ZN(n6126) );
  NAND2_X1 U7726 ( .A1(n6126), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7727 ( .A(n6127), .ZN(n7609) );
  INV_X1 U7728 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6128) );
  NOR2_X1 U7729 ( .A1(n6455), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8805) );
  INV_X1 U7730 ( .A(n8805), .ZN(n8811) );
  OAI222_X1 U7731 ( .A1(n6417), .A2(P2_U3152), .B1(n8799), .B2(n7609), .C1(
        n6128), .C2(n8811), .ZN(P2_U3357) );
  INV_X1 U7732 ( .A(n8225), .ZN(n6129) );
  OAI222_X1 U7733 ( .A1(n8811), .A2(n4619), .B1(n8799), .B2(n4449), .C1(
        P2_U3152), .C2(n6129), .ZN(P2_U3355) );
  INV_X1 U7734 ( .A(n6734), .ZN(n6135) );
  INV_X1 U7735 ( .A(n6663), .ZN(n6648) );
  OAI222_X1 U7736 ( .A1(n8811), .A2(n4676), .B1(n8799), .B2(n6135), .C1(
        P2_U3152), .C2(n6648), .ZN(P2_U3354) );
  INV_X1 U7737 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6736) );
  AND2_X1 U7738 ( .A1(n5808), .A2(P1_U3084), .ZN(n9735) );
  INV_X1 U7739 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9727) );
  NOR2_X1 U7740 ( .A1(n6133), .A2(n9727), .ZN(n6130) );
  MUX2_X1 U7741 ( .A(n9727), .B(n6130), .S(P1_IR_REG_4__SCAN_IN), .Z(n6131) );
  INV_X1 U7742 ( .A(n6131), .ZN(n6134) );
  INV_X1 U7743 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7744 ( .A1(n6133), .A2(n6132), .ZN(n6143) );
  NAND2_X1 U7745 ( .A1(n6134), .A2(n6143), .ZN(n6735) );
  OAI222_X1 U7746 ( .A1(n9743), .A2(n6736), .B1(n4261), .B2(n6135), .C1(
        P1_U3084), .C2(n6735), .ZN(P1_U3349) );
  INV_X1 U7747 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6137) );
  INV_X1 U7748 ( .A(n6730), .ZN(n6142) );
  NAND2_X1 U7749 ( .A1(n6143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6136) );
  XNOR2_X1 U7750 ( .A(n6136), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6731) );
  INV_X1 U7751 ( .A(n6731), .ZN(n6244) );
  OAI222_X1 U7752 ( .A1(n9743), .A2(n6137), .B1(n4261), .B2(n6142), .C1(
        P1_U3084), .C2(n6244), .ZN(P1_U3348) );
  INV_X1 U7753 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U7754 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6138) );
  INV_X1 U7755 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6139) );
  INV_X1 U7756 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6140) );
  OAI222_X1 U7757 ( .A1(n9743), .A2(n6522), .B1(n4261), .B2(n4449), .C1(
        P1_U3084), .C2(n6521), .ZN(P1_U3350) );
  AOI22_X1 U7758 ( .A1(n8239), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8805), .ZN(n6141) );
  OAI21_X1 U7759 ( .B1(n6142), .B2(n8799), .A(n6141), .ZN(P2_U3353) );
  INV_X1 U7760 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6145) );
  INV_X1 U7761 ( .A(n6867), .ZN(n6146) );
  NAND2_X1 U7762 ( .A1(n6161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6144) );
  XNOR2_X1 U7763 ( .A(n6144), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6868) );
  INV_X1 U7764 ( .A(n6868), .ZN(n6267) );
  OAI222_X1 U7765 ( .A1(n9743), .A2(n6145), .B1(n4261), .B2(n6146), .C1(
        P1_U3084), .C2(n6267), .ZN(P1_U3347) );
  INV_X1 U7766 ( .A(n8253), .ZN(n6652) );
  OAI222_X1 U7767 ( .A1(n8811), .A2(n4629), .B1(n8799), .B2(n6146), .C1(
        P2_U3152), .C2(n6652), .ZN(P2_U3352) );
  INV_X1 U7768 ( .A(n6557), .ZN(n6567) );
  OAI222_X1 U7769 ( .A1(n6567), .A2(P2_U3152), .B1(n8799), .B2(n6501), .C1(
        n6147), .C2(n8811), .ZN(P2_U3356) );
  INV_X1 U7770 ( .A(n6968), .ZN(n6171) );
  AOI22_X1 U7771 ( .A1(n8268), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8805), .ZN(n6148) );
  OAI21_X1 U7772 ( .B1(n6171), .B2(n8799), .A(n6148), .ZN(P2_U3351) );
  AND2_X1 U7773 ( .A1(n7551), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6149) );
  INV_X1 U7774 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6156) );
  NAND3_X1 U7775 ( .A1(n6150), .A2(P1_B_REG_SCAN_IN), .A3(n7606), .ZN(n6151)
         );
  OAI211_X1 U7776 ( .C1(P1_B_REG_SCAN_IN), .C2(n7606), .A(n6152), .B(n6151), 
        .ZN(n9815) );
  OR2_X1 U7777 ( .A1(n9815), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7778 ( .A1(n9746), .A2(n7606), .ZN(n6153) );
  NAND2_X1 U7779 ( .A1(n6154), .A2(n6153), .ZN(n6603) );
  INV_X1 U7780 ( .A(n6603), .ZN(n6438) );
  NAND2_X1 U7781 ( .A1(n6438), .A2(n9816), .ZN(n6155) );
  OAI21_X1 U7782 ( .B1(n9816), .B2(n6156), .A(n6155), .ZN(P1_U3440) );
  INV_X1 U7783 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6160) );
  OR2_X1 U7784 ( .A1(n9815), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7785 ( .A1(n9746), .A2(n6150), .ZN(n6157) );
  NAND2_X1 U7786 ( .A1(n6158), .A2(n6157), .ZN(n6322) );
  INV_X1 U7787 ( .A(n6322), .ZN(n6439) );
  NAND2_X1 U7788 ( .A1(n6439), .A2(n9816), .ZN(n6159) );
  OAI21_X1 U7789 ( .B1(n9816), .B2(n6160), .A(n6159), .ZN(P1_U3441) );
  INV_X1 U7790 ( .A(n7088), .ZN(n6168) );
  INV_X1 U7791 ( .A(n6161), .ZN(n6163) );
  NAND2_X1 U7792 ( .A1(n6163), .A2(n6162), .ZN(n6169) );
  OAI21_X1 U7793 ( .B1(n6169), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6164) );
  MUX2_X1 U7794 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6164), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n6166) );
  INV_X1 U7795 ( .A(n9743), .ZN(n9740) );
  AOI22_X1 U7796 ( .A1(n9805), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9740), .ZN(n6167) );
  OAI21_X1 U7797 ( .B1(n6168), .B2(n4261), .A(n6167), .ZN(P1_U3345) );
  INV_X1 U7798 ( .A(n6672), .ZN(n8278) );
  OAI222_X1 U7799 ( .A1(n8811), .A2(n10127), .B1(n8799), .B2(n6168), .C1(
        P2_U3152), .C2(n8278), .ZN(P2_U3350) );
  INV_X1 U7800 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7801 ( .A1(n6169), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6170) );
  XNOR2_X1 U7802 ( .A(n6170), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6969) );
  INV_X1 U7803 ( .A(n6969), .ZN(n6271) );
  OAI222_X1 U7804 ( .A1(n9743), .A2(n6172), .B1(n4261), .B2(n6171), .C1(
        P1_U3084), .C2(n6271), .ZN(P1_U3346) );
  NAND2_X1 U7805 ( .A1(n6174), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n6175) );
  OAI222_X1 U7806 ( .A1(n6503), .A2(P1_U3084), .B1(n4261), .B2(n6501), .C1(
        n6502), .C2(n9743), .ZN(P1_U3351) );
  INV_X1 U7807 ( .A(n7153), .ZN(n6180) );
  NAND2_X1 U7808 ( .A1(n6301), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6177) );
  XNOR2_X1 U7809 ( .A(n6177), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7154) );
  AOI22_X1 U7810 ( .A1(n7154), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9740), .ZN(n6178) );
  OAI21_X1 U7811 ( .B1(n6180), .B2(n4261), .A(n6178), .ZN(P1_U3344) );
  AOI22_X1 U7812 ( .A1(n8303), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8805), .ZN(n6179) );
  OAI21_X1 U7813 ( .B1(n6180), .B2(n8799), .A(n6179), .ZN(P2_U3349) );
  INV_X1 U7814 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6183) );
  INV_X1 U7815 ( .A(n8377), .ZN(n6181) );
  NAND2_X1 U7816 ( .A1(n6181), .A2(P2_U3966), .ZN(n6182) );
  OAI21_X1 U7817 ( .B1(P2_U3966), .B2(n6183), .A(n6182), .ZN(P2_U3583) );
  INV_X1 U7818 ( .A(n6735), .ZN(n6194) );
  INV_X1 U7819 ( .A(n6521), .ZN(n6193) );
  INV_X1 U7820 ( .A(n6503), .ZN(n6377) );
  INV_X1 U7821 ( .A(n7610), .ZN(n6230) );
  NAND2_X1 U7822 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6366) );
  XOR2_X1 U7823 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6503), .Z(n6373) );
  XOR2_X1 U7824 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6521), .Z(n6261) );
  INV_X1 U7825 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6184) );
  MUX2_X1 U7826 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6184), .S(n6735), .Z(n6185)
         );
  INV_X1 U7827 ( .A(n6185), .ZN(n6381) );
  XOR2_X1 U7828 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6731), .Z(n6246) );
  XOR2_X1 U7829 ( .A(n6247), .B(n6246), .Z(n6203) );
  NOR2_X1 U7830 ( .A1(n9055), .A2(P1_U3084), .ZN(n9739) );
  AND2_X1 U7831 ( .A1(n6196), .A2(n9739), .ZN(n9368) );
  NAND2_X1 U7832 ( .A1(n9368), .A2(n9780), .ZN(n9799) );
  AND2_X1 U7833 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7045) );
  INV_X1 U7834 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U7835 ( .A1(n7610), .A2(n9877), .ZN(n6187) );
  AND2_X1 U7836 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6224) );
  NAND2_X1 U7837 ( .A1(n6223), .A2(n6224), .ZN(n6222) );
  NAND2_X1 U7838 ( .A1(n6222), .A2(n6188), .ZN(n6369) );
  NAND2_X1 U7839 ( .A1(n6369), .A2(n6368), .ZN(n6191) );
  INV_X1 U7840 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6189) );
  OR2_X1 U7841 ( .A1(n6503), .A2(n6189), .ZN(n6190) );
  NAND2_X1 U7842 ( .A1(n6191), .A2(n6190), .ZN(n6256) );
  INV_X1 U7843 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6192) );
  AND2_X1 U7844 ( .A1(n6256), .A2(n6257), .ZN(n6254) );
  INV_X1 U7845 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9880) );
  MUX2_X1 U7846 ( .A(n9880), .B(P1_REG1_REG_4__SCAN_IN), .S(n6735), .Z(n6384)
         );
  NAND2_X1 U7847 ( .A1(n6385), .A2(n6384), .ZN(n6383) );
  INV_X1 U7848 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9882) );
  MUX2_X1 U7849 ( .A(n9882), .B(P1_REG1_REG_5__SCAN_IN), .S(n6731), .Z(n6197)
         );
  OR2_X1 U7850 ( .A1(n9056), .A2(P1_U3084), .ZN(n9737) );
  INV_X1 U7851 ( .A(n9055), .ZN(n9778) );
  NOR2_X1 U7852 ( .A1(n9737), .A2(n9778), .ZN(n6195) );
  NAND2_X1 U7853 ( .A1(n6196), .A2(n6195), .ZN(n9807) );
  AOI211_X1 U7854 ( .C1(n6198), .C2(n6197), .A(n9807), .B(n6239), .ZN(n6199)
         );
  AOI211_X1 U7855 ( .C1(n9369), .C2(n6731), .A(n7045), .B(n6199), .ZN(n6202)
         );
  OR2_X1 U7856 ( .A1(P1_U3083), .A2(n6200), .ZN(n9813) );
  NAND2_X1 U7857 ( .A1(n9375), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6201) );
  OAI211_X1 U7858 ( .C1(n6203), .C2(n9799), .A(n6202), .B(n6201), .ZN(P1_U3246) );
  OAI21_X1 U7859 ( .B1(n6394), .B2(n6204), .A(n6401), .ZN(n6206) );
  NAND2_X1 U7860 ( .A1(n6394), .A2(n6395), .ZN(n6205) );
  NAND2_X1 U7861 ( .A1(n6206), .A2(n6205), .ZN(n8375) );
  NOR2_X1 U7862 ( .A1(n10200), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7863 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6218) );
  INV_X1 U7864 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7865 ( .A1(n6211), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7866 ( .A1(n6532), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6216) );
  INV_X1 U7867 ( .A(n6280), .ZN(n9732) );
  NAND2_X1 U7868 ( .A1(n6743), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7869 ( .A1(n7986), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6214) );
  AND3_X1 U7870 ( .A1(n6216), .A2(n6215), .A3(n6214), .ZN(n9052) );
  INV_X1 U7871 ( .A(n9052), .ZN(n9378) );
  NAND2_X1 U7872 ( .A1(n9378), .A2(P1_U4006), .ZN(n6217) );
  OAI21_X1 U7873 ( .B1(P1_U4006), .B2(n6218), .A(n6217), .ZN(P1_U3586) );
  INV_X1 U7874 ( .A(n7281), .ZN(n6220) );
  NOR2_X1 U7875 ( .A1(n6301), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6289) );
  OR2_X1 U7876 ( .A1(n6289), .A2(n9727), .ZN(n6234) );
  XNOR2_X1 U7877 ( .A(n6234), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7282) );
  INV_X1 U7878 ( .A(n7282), .ZN(n6775) );
  OAI222_X1 U7879 ( .A1(n9743), .A2(n6219), .B1(n4261), .B2(n6220), .C1(n6775), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U7880 ( .A(n6689), .ZN(n6660) );
  OAI222_X1 U7881 ( .A1(n8811), .A2(n6221), .B1(n8799), .B2(n6220), .C1(n6660), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7882 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6232) );
  INV_X1 U7883 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6478) );
  INV_X1 U7884 ( .A(n9807), .ZN(n9790) );
  OAI211_X1 U7885 ( .C1(n6224), .C2(n6223), .A(n9790), .B(n6222), .ZN(n6225)
         );
  OAI21_X1 U7886 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6478), .A(n6225), .ZN(n6229) );
  AOI211_X1 U7887 ( .C1(n6366), .C2(n6227), .A(n6226), .B(n9799), .ZN(n6228)
         );
  AOI211_X1 U7888 ( .C1(n9369), .C2(n6230), .A(n6229), .B(n6228), .ZN(n6231)
         );
  OAI21_X1 U7889 ( .B1(n9813), .B2(n6232), .A(n6231), .ZN(P1_U3242) );
  INV_X1 U7890 ( .A(n7285), .ZN(n6237) );
  INV_X1 U7891 ( .A(n6690), .ZN(n8313) );
  OAI222_X1 U7892 ( .A1(n8811), .A2(n10129), .B1(n8799), .B2(n6237), .C1(n8313), .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7893 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7894 ( .A1(n6234), .A2(n6233), .ZN(n6235) );
  NAND2_X1 U7895 ( .A1(n6235), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6236) );
  XNOR2_X1 U7896 ( .A(n6236), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7286) );
  INV_X1 U7897 ( .A(n7286), .ZN(n6784) );
  OAI222_X1 U7898 ( .A1(n9743), .A2(n6238), .B1(n4261), .B2(n6237), .C1(n6784), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U7899 ( .A(n6241), .ZN(n6243) );
  INV_X1 U7900 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9884) );
  MUX2_X1 U7901 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9884), .S(n6868), .Z(n6240)
         );
  INV_X1 U7902 ( .A(n6240), .ZN(n6242) );
  AOI21_X1 U7903 ( .B1(n6243), .B2(n6242), .A(n6274), .ZN(n6253) );
  INV_X1 U7904 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6245) );
  AOI22_X1 U7905 ( .A1(n6247), .A2(n6246), .B1(n6245), .B2(n6244), .ZN(n6249)
         );
  XOR2_X1 U7906 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6868), .Z(n6248) );
  NAND2_X1 U7907 ( .A1(n6249), .A2(n6248), .ZN(n6266) );
  OAI211_X1 U7908 ( .C1(n6249), .C2(n6248), .A(n6266), .B(n4531), .ZN(n6252)
         );
  INV_X1 U7909 ( .A(n9369), .ZN(n9791) );
  NAND2_X1 U7910 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7122) );
  OAI21_X1 U7911 ( .B1(n9791), .B2(n6267), .A(n7122), .ZN(n6250) );
  AOI21_X1 U7912 ( .B1(n9375), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6250), .ZN(
        n6251) );
  OAI211_X1 U7913 ( .C1(n6253), .C2(n9807), .A(n6252), .B(n6251), .ZN(P1_U3247) );
  INV_X1 U7914 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6903) );
  NOR2_X1 U7915 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6903), .ZN(n6540) );
  INV_X1 U7916 ( .A(n6540), .ZN(n6259) );
  INV_X1 U7917 ( .A(n6254), .ZN(n6255) );
  OAI211_X1 U7918 ( .C1(n6257), .C2(n6256), .A(n9790), .B(n6255), .ZN(n6258)
         );
  OAI211_X1 U7919 ( .C1(n9791), .C2(n6521), .A(n6259), .B(n6258), .ZN(n6264)
         );
  AOI211_X1 U7920 ( .C1(n6262), .C2(n6261), .A(n9799), .B(n6260), .ZN(n6263)
         );
  AOI211_X1 U7921 ( .C1(P1_ADDR_REG_3__SCAN_IN), .C2(n9375), .A(n6264), .B(
        n6263), .ZN(n6265) );
  INV_X1 U7922 ( .A(n6265), .ZN(P1_U3244) );
  XNOR2_X1 U7923 ( .A(n6969), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6270) );
  INV_X1 U7924 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6268) );
  OAI21_X1 U7925 ( .B1(n6268), .B2(n6267), .A(n6266), .ZN(n6269) );
  AOI21_X1 U7926 ( .B1(n6270), .B2(n6269), .A(n9794), .ZN(n6279) );
  NAND2_X1 U7927 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7018) );
  OAI21_X1 U7928 ( .B1(n9791), .B2(n6271), .A(n7018), .ZN(n6277) );
  NOR2_X1 U7929 ( .A1(n6868), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6272) );
  INV_X1 U7930 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9886) );
  MUX2_X1 U7931 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9886), .S(n6969), .Z(n6273)
         );
  OR3_X1 U7932 ( .A1(n6274), .A2(n6273), .A3(n6272), .ZN(n6275) );
  AOI21_X1 U7933 ( .B1(n6340), .B2(n6275), .A(n9807), .ZN(n6276) );
  AOI211_X1 U7934 ( .C1(n9375), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n6277), .B(
        n6276), .ZN(n6278) );
  OAI21_X1 U7935 ( .B1(n6279), .B2(n9799), .A(n6278), .ZN(P1_U3248) );
  INV_X1 U7936 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7937 ( .A1(n6532), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7938 ( .A1(n6743), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7939 ( .A1(n4264), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7940 ( .A1(n6879), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6282) );
  INV_X1 U7941 ( .A(n6360), .ZN(n6643) );
  NAND2_X1 U7942 ( .A1(n6643), .A2(P1_U4006), .ZN(n6286) );
  OAI21_X1 U7943 ( .B1(P1_U4006), .B2(n6287), .A(n6286), .ZN(P1_U3555) );
  INV_X1 U7944 ( .A(n7308), .ZN(n6294) );
  NOR2_X1 U7945 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6288) );
  NAND2_X1 U7946 ( .A1(n6289), .A2(n6288), .ZN(n6291) );
  NAND2_X1 U7947 ( .A1(n6291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6290) );
  MUX2_X1 U7948 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6290), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6292) );
  INV_X1 U7949 ( .A(n7297), .ZN(n7250) );
  OAI222_X1 U7950 ( .A1(n9743), .A2(n6293), .B1(n4261), .B2(n6294), .C1(
        P1_U3084), .C2(n7250), .ZN(P1_U3341) );
  INV_X1 U7951 ( .A(n6703), .ZN(n6693) );
  OAI222_X1 U7952 ( .A1(n8811), .A2(n6295), .B1(n8799), .B2(n6294), .C1(
        P2_U3152), .C2(n6693), .ZN(P2_U3346) );
  NOR2_X1 U7953 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6298) );
  NOR2_X1 U7954 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6297) );
  NOR2_X1 U7955 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6296) );
  NAND4_X1 U7956 ( .A1(n6299), .A2(n6298), .A3(n6297), .A4(n6296), .ZN(n6300)
         );
  OR2_X1 U7957 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  NAND2_X1 U7958 ( .A1(n6302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7716) );
  INV_X1 U7959 ( .A(n6303), .ZN(n6304) );
  NAND2_X1 U7960 ( .A1(n6304), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7961 ( .A1(n7716), .A2(n6305), .ZN(n6307) );
  INV_X1 U7962 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7963 ( .A1(n6308), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6310) );
  INV_X1 U7964 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6309) );
  XNOR2_X1 U7965 ( .A(n6310), .B(n6309), .ZN(n7276) );
  OR2_X1 U7966 ( .A1(n9226), .A2(n9267), .ZN(n6483) );
  NAND2_X1 U7967 ( .A1(n9816), .A2(n6483), .ZN(n6604) );
  NOR2_X1 U7968 ( .A1(n6438), .A2(n6604), .ZN(n6323) );
  NOR4_X1 U7969 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6318) );
  NOR4_X1 U7970 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6317) );
  INV_X1 U7971 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10109) );
  INV_X1 U7972 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10147) );
  INV_X1 U7973 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10172) );
  INV_X1 U7974 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10155) );
  NAND4_X1 U7975 ( .A1(n10109), .A2(n10147), .A3(n10172), .A4(n10155), .ZN(
        n10038) );
  NOR4_X1 U7976 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6314) );
  NOR4_X1 U7977 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6313) );
  NOR4_X1 U7978 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6312) );
  NOR4_X1 U7979 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6311) );
  NAND4_X1 U7980 ( .A1(n6314), .A2(n6313), .A3(n6312), .A4(n6311), .ZN(n6315)
         );
  NOR4_X1 U7981 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n10038), .A4(n6315), .ZN(n6316) );
  AND3_X1 U7982 ( .A1(n6318), .A2(n6317), .A3(n6316), .ZN(n6319) );
  OR2_X1 U7983 ( .A1(n9815), .A2(n6319), .ZN(n6437) );
  NAND2_X1 U7984 ( .A1(n9856), .A2(n9224), .ZN(n6321) );
  AND2_X2 U7985 ( .A1(n6323), .A2(n6606), .ZN(n9876) );
  INV_X1 U7986 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6336) );
  INV_X1 U7987 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9786) );
  INV_X1 U7988 ( .A(SI_0_), .ZN(n6325) );
  INV_X1 U7989 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6324) );
  OAI21_X1 U7990 ( .B1(n6455), .B2(n6325), .A(n6324), .ZN(n6327) );
  NAND2_X1 U7991 ( .A1(n6327), .A2(n6326), .ZN(n9747) );
  MUX2_X1 U7992 ( .A(n9786), .B(n9747), .S(n7678), .Z(n6477) );
  NAND2_X1 U7993 ( .A1(n9227), .A2(n9224), .ZN(n6440) );
  AND2_X1 U7994 ( .A1(n6643), .A2(n6477), .ZN(n9003) );
  INV_X1 U7995 ( .A(n9003), .ZN(n6328) );
  NAND2_X1 U7996 ( .A1(n6752), .A2(n6328), .ZN(n9188) );
  NAND2_X1 U7997 ( .A1(n9057), .A2(n9261), .ZN(n6464) );
  OR2_X1 U7998 ( .A1(n6464), .A2(n6463), .ZN(n6770) );
  AND2_X1 U7999 ( .A1(n6770), .A2(n6440), .ZN(n6334) );
  NAND2_X1 U8000 ( .A1(n6879), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U8001 ( .A1(n4264), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U8002 ( .A1(n6743), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U8003 ( .A1(n6532), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6329) );
  AND2_X1 U8004 ( .A1(n9285), .A2(n9572), .ZN(n6333) );
  AOI21_X1 U8005 ( .B1(n9188), .B2(n6334), .A(n6333), .ZN(n6422) );
  OAI21_X1 U8006 ( .B1(n6477), .B2(n6440), .A(n6422), .ZN(n9704) );
  NAND2_X1 U8007 ( .A1(n9704), .A2(n9876), .ZN(n6335) );
  OAI21_X1 U8008 ( .B1(n9876), .B2(n6336), .A(n6335), .ZN(P1_U3454) );
  INV_X1 U8009 ( .A(n7511), .ZN(n6339) );
  INV_X1 U8010 ( .A(n6845), .ZN(n6708) );
  OAI222_X1 U8011 ( .A1(n8811), .A2(n6337), .B1(n8799), .B2(n6339), .C1(n6708), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  NAND2_X1 U8012 ( .A1(n6351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6338) );
  XNOR2_X1 U8013 ( .A(n6338), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9293) );
  INV_X1 U8014 ( .A(n9293), .ZN(n7258) );
  OAI222_X1 U8015 ( .A1(n9743), .A2(n10071), .B1(n4261), .B2(n6339), .C1(n7258), .C2(P1_U3084), .ZN(P1_U3340) );
  NAND2_X1 U8016 ( .A1(n9805), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6341) );
  NOR2_X1 U8017 ( .A1(n9805), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9809) );
  XNOR2_X1 U8018 ( .A(n7154), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n6574) );
  XNOR2_X1 U8019 ( .A(n9806), .B(n6574), .ZN(n6349) );
  INV_X1 U8020 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U8021 ( .A1(n9369), .A2(n7154), .ZN(n6342) );
  NAND2_X1 U8022 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7269) );
  OAI211_X1 U8023 ( .C1(n9813), .C2(n10217), .A(n6342), .B(n7269), .ZN(n6348)
         );
  XNOR2_X1 U8024 ( .A(n7154), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6346) );
  NOR2_X1 U8025 ( .A1(n6969), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9795) );
  INV_X1 U8026 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6343) );
  MUX2_X1 U8027 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6343), .S(n9805), .Z(n6344)
         );
  AOI211_X1 U8028 ( .C1(n6346), .C2(n6345), .A(n9799), .B(n4372), .ZN(n6347)
         );
  AOI211_X1 U8029 ( .C1(n9790), .C2(n6349), .A(n6348), .B(n6347), .ZN(n6350)
         );
  INV_X1 U8030 ( .A(n6350), .ZN(P1_U3250) );
  INV_X1 U8031 ( .A(n7582), .ZN(n6353) );
  NAND2_X1 U8032 ( .A1(n6802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6582) );
  XNOR2_X1 U8033 ( .A(n6582), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9311) );
  INV_X1 U8034 ( .A(n9311), .ZN(n9294) );
  OAI222_X1 U8035 ( .A1(n9743), .A2(n6352), .B1(n4261), .B2(n6353), .C1(n9294), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8036 ( .A(n7214), .ZN(n7212) );
  OAI222_X1 U8037 ( .A1(n8811), .A2(n6354), .B1(n8799), .B2(n6353), .C1(n7212), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8038 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U8039 ( .A1(n9227), .A2(n9267), .ZN(n6355) );
  INV_X1 U8040 ( .A(n6463), .ZN(n6356) );
  OAI22_X1 U8041 ( .A1(n6477), .A2(n7875), .B1(n9786), .B2(n6482), .ZN(n6357)
         );
  INV_X1 U8042 ( .A(n6357), .ZN(n6358) );
  INV_X1 U8043 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6361) );
  OAI22_X1 U8044 ( .A1(n6477), .A2(n6524), .B1(n6361), .B2(n6482), .ZN(n6362)
         );
  INV_X1 U8045 ( .A(n6362), .ZN(n6363) );
  OAI21_X1 U8046 ( .B1(n6365), .B2(n6489), .A(n6491), .ZN(n6436) );
  MUX2_X1 U8047 ( .A(n6366), .B(n6436), .S(n9055), .Z(n6367) );
  INV_X1 U8048 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6419) );
  AND2_X1 U8049 ( .A1(n9778), .A2(n6419), .ZN(n9779) );
  OAI21_X1 U8050 ( .B1(n9779), .B2(n9056), .A(n9786), .ZN(n9782) );
  OAI211_X1 U8051 ( .C1(n6367), .C2(n9056), .A(P1_U4006), .B(n9782), .ZN(n6391) );
  XNOR2_X1 U8052 ( .A(n6369), .B(n6368), .ZN(n6371) );
  INV_X1 U8053 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6370) );
  OAI22_X1 U8054 ( .A1(n9807), .A2(n6371), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6370), .ZN(n6376) );
  AOI211_X1 U8055 ( .C1(n6374), .C2(n6373), .A(n6372), .B(n9799), .ZN(n6375)
         );
  AOI211_X1 U8056 ( .C1(n9369), .C2(n6377), .A(n6376), .B(n6375), .ZN(n6378)
         );
  OAI211_X1 U8057 ( .C1(n9813), .C2(n6379), .A(n6391), .B(n6378), .ZN(P1_U3243) );
  INV_X1 U8058 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U8059 ( .B1(n6382), .B2(n6381), .A(n6380), .ZN(n6389) );
  OAI21_X1 U8060 ( .B1(n6385), .B2(n6384), .A(n6383), .ZN(n6386) );
  AND2_X1 U8061 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n8928) );
  AOI21_X1 U8062 ( .B1(n9790), .B2(n6386), .A(n8928), .ZN(n6387) );
  OAI21_X1 U8063 ( .B1(n9791), .B2(n6735), .A(n6387), .ZN(n6388) );
  AOI21_X1 U8064 ( .B1(n6389), .B2(n4531), .A(n6388), .ZN(n6390) );
  OAI211_X1 U8065 ( .C1(n6392), .C2(n9813), .A(n6391), .B(n6390), .ZN(P1_U3245) );
  OR2_X1 U8066 ( .A1(n6410), .A2(P2_U3152), .ZN(n8798) );
  OR2_X1 U8067 ( .A1(n6394), .A2(n6393), .ZN(n6396) );
  OAI211_X1 U8068 ( .C1(n6397), .C2(n8798), .A(n6396), .B(n6395), .ZN(n6403)
         );
  NAND2_X1 U8069 ( .A1(n6403), .A2(n6401), .ZN(n6398) );
  INV_X2 U8070 ( .A(P2_U3966), .ZN(n8217) );
  NAND2_X1 U8071 ( .A1(n6398), .A2(n8217), .ZN(n8365) );
  NAND2_X1 U8072 ( .A1(n8365), .A2(n6410), .ZN(n10204) );
  INV_X1 U8073 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7033) );
  NOR2_X1 U8074 ( .A1(n7033), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8075 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6406) );
  XNOR2_X1 U8076 ( .A(n6417), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6400) );
  INV_X1 U8077 ( .A(n6400), .ZN(n6405) );
  AND2_X1 U8078 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6399) );
  NAND2_X1 U8079 ( .A1(n6400), .A2(n6399), .ZN(n6429) );
  INV_X1 U8080 ( .A(n6429), .ZN(n6404) );
  AND2_X1 U8081 ( .A1(n6401), .A2(n6619), .ZN(n6402) );
  NAND2_X1 U8082 ( .A1(n6403), .A2(n6402), .ZN(n10194) );
  AOI211_X1 U8083 ( .C1(n6406), .C2(n6405), .A(n6404), .B(n10194), .ZN(n6407)
         );
  AOI211_X1 U8084 ( .C1(n10200), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6408), .B(
        n6407), .ZN(n6416) );
  XNOR2_X1 U8085 ( .A(n6417), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n6414) );
  INV_X1 U8086 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6409) );
  INV_X1 U8087 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6620) );
  NOR2_X1 U8088 ( .A1(n6409), .A2(n6620), .ZN(n6413) );
  NOR2_X1 U8089 ( .A1(n6410), .A2(n6619), .ZN(n6411) );
  NAND2_X1 U8090 ( .A1(n8365), .A2(n6411), .ZN(n8370) );
  INV_X1 U8091 ( .A(n6423), .ZN(n6412) );
  OAI211_X1 U8092 ( .C1(n6414), .C2(n6413), .A(n10190), .B(n6412), .ZN(n6415)
         );
  OAI211_X1 U8093 ( .C1(n10204), .C2(n6417), .A(n6416), .B(n6415), .ZN(
        P2_U3246) );
  INV_X1 U8094 ( .A(n6604), .ZN(n6449) );
  NAND4_X1 U8095 ( .A1(n6449), .A2(n6439), .A3(n6603), .A4(n6437), .ZN(n6418)
         );
  NAND3_X1 U8096 ( .A1(n9816), .A2(n9856), .A3(n9224), .ZN(n9530) );
  OR2_X1 U8097 ( .A1(n6418), .A2(n4259), .ZN(n7324) );
  INV_X1 U8098 ( .A(n7276), .ZN(n9263) );
  NOR2_X1 U8099 ( .A1(n6440), .A2(n7276), .ZN(n6447) );
  INV_X1 U8100 ( .A(n6477), .ZN(n6476) );
  OAI21_X1 U8101 ( .B1(n9581), .B2(n9490), .A(n6476), .ZN(n6421) );
  AOI22_X1 U8102 ( .A1(n9566), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9582), .ZN(n6420) );
  OAI211_X1 U8103 ( .C1(n9566), .C2(n6422), .A(n6421), .B(n6420), .ZN(P1_U3291) );
  INV_X1 U8104 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9914) );
  MUX2_X1 U8105 ( .A(n9914), .B(P2_REG2_REG_2__SCAN_IN), .S(n6557), .Z(n6424)
         );
  AOI211_X1 U8106 ( .C1(n6425), .C2(n6424), .A(n8224), .B(n8370), .ZN(n6435)
         );
  AOI22_X1 U8107 ( .A1(n10200), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n6433) );
  INV_X1 U8108 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6426) );
  XNOR2_X1 U8109 ( .A(n6557), .B(n6426), .ZN(n6431) );
  NAND2_X1 U8110 ( .A1(n6427), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8111 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  NAND2_X1 U8112 ( .A1(n6431), .A2(n6430), .ZN(n6559) );
  OAI211_X1 U8113 ( .C1(n6431), .C2(n6430), .A(n8359), .B(n6559), .ZN(n6432)
         );
  OAI211_X1 U8114 ( .C1(n10204), .C2(n6567), .A(n6433), .B(n6432), .ZN(n6434)
         );
  OR2_X1 U8115 ( .A1(n6435), .A2(n6434), .ZN(P2_U3247) );
  INV_X1 U8116 ( .A(n6436), .ZN(n6452) );
  NAND3_X1 U8117 ( .A1(n6439), .A2(n6438), .A3(n6437), .ZN(n6448) );
  NAND3_X1 U8118 ( .A1(n9816), .A2(n9226), .A3(n9868), .ZN(n6441) );
  INV_X1 U8119 ( .A(n6770), .ZN(n6442) );
  AND2_X1 U8120 ( .A1(n9816), .A2(n6442), .ZN(n9060) );
  INV_X1 U8121 ( .A(n9060), .ZN(n6443) );
  OR2_X1 U8122 ( .A1(n6448), .A2(n6443), .ZN(n6531) );
  INV_X1 U8123 ( .A(n6531), .ZN(n6444) );
  NAND2_X1 U8124 ( .A1(n6444), .A2(n9056), .ZN(n8986) );
  INV_X1 U8125 ( .A(n8986), .ZN(n8971) );
  NAND2_X1 U8126 ( .A1(n9816), .A2(n6447), .ZN(n6445) );
  OR2_X1 U8127 ( .A1(n6448), .A2(n6445), .ZN(n6446) );
  AOI22_X1 U8128 ( .A1(n8971), .A2(n9285), .B1(n6476), .B2(n8978), .ZN(n6451)
         );
  NAND2_X1 U8129 ( .A1(n6448), .A2(n5128), .ZN(n6487) );
  NAND2_X1 U8130 ( .A1(n6448), .A2(n9868), .ZN(n6484) );
  NAND3_X1 U8131 ( .A1(n6487), .A2(n6484), .A3(n6449), .ZN(n6644) );
  NAND2_X1 U8132 ( .A1(n6644), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6450) );
  OAI211_X1 U8133 ( .C1(n6452), .C2(n8993), .A(n6451), .B(n6450), .ZN(P1_U3230) );
  INV_X1 U8134 ( .A(n7676), .ZN(n6585) );
  AOI22_X1 U8135 ( .A1(n8330), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8805), .ZN(n6453) );
  OAI21_X1 U8136 ( .B1(n6585), .B2(n8799), .A(n6453), .ZN(P2_U3343) );
  INV_X1 U8137 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7608) );
  OR2_X1 U8138 ( .A1(n9049), .A2(n7608), .ZN(n6457) );
  OR2_X1 U8139 ( .A1(n7678), .A2(n7610), .ZN(n6456) );
  XNOR2_X1 U8140 ( .A(n9285), .B(n9821), .ZN(n6459) );
  AND2_X1 U8141 ( .A1(n6643), .A2(n6476), .ZN(n6460) );
  NAND2_X1 U8142 ( .A1(n6459), .A2(n6460), .ZN(n6588) );
  OR2_X1 U8143 ( .A1(n6459), .A2(n6460), .ZN(n6461) );
  NAND2_X1 U8144 ( .A1(n6588), .A2(n6461), .ZN(n9819) );
  NOR2_X1 U8145 ( .A1(n6463), .A2(n9261), .ZN(n6462) );
  NAND2_X1 U8146 ( .A1(n9589), .A2(n6462), .ZN(n7536) );
  NAND3_X1 U8147 ( .A1(n6770), .A2(n7890), .A3(n9261), .ZN(n9601) );
  INV_X1 U8148 ( .A(n6752), .ZN(n6465) );
  INV_X1 U8149 ( .A(n6459), .ZN(n9192) );
  NAND2_X1 U8150 ( .A1(n9192), .A2(n6465), .ZN(n6596) );
  OAI21_X1 U8151 ( .B1(n6465), .B2(n9192), .A(n6596), .ZN(n6468) );
  NAND2_X1 U8152 ( .A1(n9057), .A2(n4259), .ZN(n6467) );
  NAND2_X1 U8153 ( .A1(n9259), .A2(n9263), .ZN(n6466) );
  NAND2_X1 U8154 ( .A1(n6468), .A2(n9577), .ZN(n6475) );
  INV_X1 U8155 ( .A(n9226), .ZN(n6469) );
  NAND2_X1 U8156 ( .A1(n6879), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U8157 ( .A1(n6743), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U8158 ( .A1(n4264), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8159 ( .A1(n6532), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6470) );
  AOI22_X1 U8160 ( .A1(n9574), .A2(n6643), .B1(n9284), .B2(n9572), .ZN(n6474)
         );
  OAI211_X1 U8161 ( .C1(n9819), .C2(n9601), .A(n6475), .B(n6474), .ZN(n9822)
         );
  OAI211_X1 U8162 ( .C1(n9821), .C2(n6477), .A(n9835), .B(n6593), .ZN(n9820)
         );
  OAI22_X1 U8163 ( .A1(n9820), .A2(n4259), .B1(n6478), .B2(n9530), .ZN(n6479)
         );
  OAI21_X1 U8164 ( .B1(n9822), .B2(n6479), .A(n9589), .ZN(n6481) );
  AOI22_X1 U8165 ( .A1(n9490), .A2(n6642), .B1(n9566), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6480) );
  OAI211_X1 U8166 ( .C1(n9819), .C2(n7536), .A(n6481), .B(n6480), .ZN(P1_U3290) );
  AND3_X1 U8167 ( .A1(n6483), .A2(n7551), .A3(n6482), .ZN(n6485) );
  NAND2_X1 U8168 ( .A1(n6485), .A2(n6484), .ZN(n6486) );
  NAND2_X1 U8169 ( .A1(n6486), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6488) );
  INV_X1 U8170 ( .A(n8991), .ZN(n8966) );
  NAND2_X1 U8171 ( .A1(n9285), .A2(n6975), .ZN(n6493) );
  OR2_X1 U8172 ( .A1(n9821), .A2(n6524), .ZN(n6492) );
  NAND2_X1 U8173 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  XNOR2_X1 U8174 ( .A(n6494), .B(n7763), .ZN(n6498) );
  OR2_X1 U8175 ( .A1(n9821), .A2(n7875), .ZN(n6495) );
  NAND2_X1 U8176 ( .A1(n6496), .A2(n6495), .ZN(n6638) );
  INV_X1 U8177 ( .A(n6497), .ZN(n6500) );
  INV_X1 U8178 ( .A(n6498), .ZN(n6499) );
  NAND2_X1 U8179 ( .A1(n6500), .A2(n6499), .ZN(n6636) );
  NAND2_X1 U8180 ( .A1(n6635), .A2(n6636), .ZN(n6630) );
  NAND2_X1 U8181 ( .A1(n9284), .A2(n6975), .ZN(n6505) );
  OR2_X1 U8182 ( .A1(n6519), .A2(n6501), .ZN(n6592) );
  OR2_X1 U8183 ( .A1(n9049), .A2(n6502), .ZN(n6591) );
  OR2_X1 U8184 ( .A1(n7678), .A2(n6503), .ZN(n6590) );
  OR2_X1 U8185 ( .A1(n6586), .A2(n6524), .ZN(n6504) );
  NAND2_X1 U8186 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  XNOR2_X1 U8187 ( .A(n6506), .B(n7890), .ZN(n6510) );
  OR2_X1 U8188 ( .A1(n6586), .A2(n7875), .ZN(n6507) );
  NAND2_X1 U8189 ( .A1(n6508), .A2(n6507), .ZN(n6511) );
  XNOR2_X1 U8190 ( .A(n6510), .B(n6511), .ZN(n6631) );
  INV_X1 U8191 ( .A(n6631), .ZN(n6509) );
  INV_X1 U8192 ( .A(n6510), .ZN(n6513) );
  INV_X1 U8193 ( .A(n6511), .ZN(n6512) );
  NAND2_X1 U8194 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  NAND2_X1 U8195 ( .A1(n6743), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U8196 ( .A1(n6879), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U8197 ( .A1(n6532), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6515) );
  NAND2_X1 U8198 ( .A1(n9283), .A2(n7892), .ZN(n6526) );
  OR2_X1 U8199 ( .A1(n7678), .A2(n6521), .ZN(n6523) );
  OR2_X1 U8200 ( .A1(n9827), .A2(n6524), .ZN(n6525) );
  NAND2_X1 U8201 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  XNOR2_X1 U8202 ( .A(n6527), .B(n7763), .ZN(n6978) );
  OR2_X1 U8203 ( .A1(n9827), .A2(n7875), .ZN(n6528) );
  NAND2_X1 U8204 ( .A1(n6529), .A2(n6528), .ZN(n6976) );
  XNOR2_X1 U8205 ( .A(n6978), .B(n6976), .ZN(n6980) );
  XNOR2_X1 U8206 ( .A(n6981), .B(n6980), .ZN(n6530) );
  NAND2_X1 U8207 ( .A1(n6530), .A2(n8964), .ZN(n6542) );
  NAND2_X1 U8208 ( .A1(n6532), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U8209 ( .A1(n6743), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6537) );
  INV_X1 U8210 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6534) );
  XNOR2_X1 U8211 ( .A(n6534), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U8212 ( .A1(n4264), .A2(n8929), .ZN(n6536) );
  NAND2_X1 U8213 ( .A1(n6879), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6535) );
  INV_X1 U8214 ( .A(n9282), .ZN(n6762) );
  OAI22_X1 U8215 ( .A1(n8968), .A2(n4731), .B1(n6762), .B2(n8986), .ZN(n6539)
         );
  AOI211_X1 U8216 ( .C1(n4737), .C2(n8978), .A(n6540), .B(n6539), .ZN(n6541)
         );
  OAI211_X1 U8217 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8966), .A(n6542), .B(
        n6541), .ZN(P1_U3216) );
  INV_X1 U8218 ( .A(n6608), .ZN(n6544) );
  NAND2_X1 U8219 ( .A1(n6917), .A2(n6545), .ZN(n6546) );
  INV_X1 U8220 ( .A(n7145), .ZN(n6547) );
  INV_X1 U8221 ( .A(n6548), .ZN(n6549) );
  AND2_X1 U8222 ( .A1(n8596), .A2(n9911), .ZN(n6551) );
  AOI21_X1 U8223 ( .B1(n6925), .B2(n9913), .A(n6551), .ZN(n6922) );
  XNOR2_X1 U8224 ( .A(n6554), .B(n6923), .ZN(n6552) );
  NAND2_X1 U8225 ( .A1(n6552), .A2(n4954), .ZN(n8581) );
  OR3_X1 U8226 ( .A1(n6554), .A2(n6553), .A3(n4954), .ZN(n9984) );
  AOI22_X1 U8227 ( .A1(n9981), .A2(n6925), .B1(n6931), .B2(n4955), .ZN(n6555)
         );
  AND2_X1 U8228 ( .A1(n6922), .A2(n6555), .ZN(n9940) );
  NAND2_X1 U8229 ( .A1(n10002), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6556) );
  OAI21_X1 U8230 ( .B1(n10002), .B2(n9940), .A(n6556), .ZN(P2_U3520) );
  INV_X1 U8231 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6565) );
  INV_X1 U8232 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10130) );
  MUX2_X1 U8233 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10130), .S(n6663), .Z(n6563)
         );
  NAND2_X1 U8234 ( .A1(n6557), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U8235 ( .A1(n6559), .A2(n6558), .ZN(n8227) );
  INV_X1 U8236 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6560) );
  XNOR2_X1 U8237 ( .A(n8225), .B(n6560), .ZN(n8228) );
  NAND2_X1 U8238 ( .A1(n8227), .A2(n8228), .ZN(n8226) );
  NAND2_X1 U8239 ( .A1(n8225), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8240 ( .A1(n8226), .A2(n6561), .ZN(n6562) );
  NAND2_X1 U8241 ( .A1(n6562), .A2(n6563), .ZN(n6665) );
  OAI211_X1 U8242 ( .C1(n6563), .C2(n6562), .A(n8359), .B(n6665), .ZN(n6564)
         );
  NAND2_X1 U8243 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8146) );
  OAI211_X1 U8244 ( .C1(n8375), .C2(n6565), .A(n6564), .B(n8146), .ZN(n6566)
         );
  AOI21_X1 U8245 ( .B1(n6663), .B2(n8335), .A(n6566), .ZN(n6573) );
  NOR2_X1 U8246 ( .A1(n6567), .A2(n9914), .ZN(n8219) );
  INV_X1 U8247 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7064) );
  MUX2_X1 U8248 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7064), .S(n8225), .Z(n6568)
         );
  OAI21_X1 U8249 ( .B1(n8224), .B2(n8219), .A(n6568), .ZN(n8222) );
  NAND2_X1 U8250 ( .A1(n8225), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6570) );
  INV_X1 U8251 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9897) );
  MUX2_X1 U8252 ( .A(n9897), .B(P2_REG2_REG_4__SCAN_IN), .S(n6663), .Z(n6569)
         );
  INV_X1 U8253 ( .A(n6650), .ZN(n8237) );
  NAND3_X1 U8254 ( .A1(n8222), .A2(n6570), .A3(n6569), .ZN(n6571) );
  NAND3_X1 U8255 ( .A1(n10190), .A2(n8237), .A3(n6571), .ZN(n6572) );
  NAND2_X1 U8256 ( .A1(n6573), .A2(n6572), .ZN(P2_U3249) );
  XOR2_X1 U8257 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7282), .Z(n6776) );
  XNOR2_X1 U8258 ( .A(n6777), .B(n6776), .ZN(n6580) );
  NAND2_X1 U8259 ( .A1(n9375), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n6575) );
  NAND2_X1 U8260 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7351) );
  OAI211_X1 U8261 ( .C1(n9791), .C2(n6775), .A(n6575), .B(n7351), .ZN(n6579)
         );
  XNOR2_X1 U8262 ( .A(n7282), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6576) );
  NOR2_X1 U8263 ( .A1(n6577), .A2(n6576), .ZN(n6778) );
  AOI211_X1 U8264 ( .C1(n6577), .C2(n6576), .A(n9799), .B(n6778), .ZN(n6578)
         );
  AOI211_X1 U8265 ( .C1(n9790), .C2(n6580), .A(n6579), .B(n6578), .ZN(n6581)
         );
  INV_X1 U8266 ( .A(n6581), .ZN(P1_U3251) );
  INV_X1 U8267 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8268 ( .A1(n6582), .A2(n6799), .ZN(n6583) );
  NAND2_X1 U8269 ( .A1(n6583), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6584) );
  INV_X1 U8270 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6800) );
  XNOR2_X1 U8271 ( .A(n6584), .B(n6800), .ZN(n9323) );
  OAI222_X1 U8272 ( .A1(n9743), .A2(n7677), .B1(n4261), .B2(n6585), .C1(
        P1_U3084), .C2(n9323), .ZN(P1_U3338) );
  OR2_X1 U8273 ( .A1(n9284), .A2(n6586), .ZN(n9007) );
  NAND2_X1 U8274 ( .A1(n9284), .A2(n6586), .ZN(n9004) );
  INV_X1 U8275 ( .A(n9189), .ZN(n6597) );
  NAND2_X1 U8276 ( .A1(n9285), .A2(n6642), .ZN(n6587) );
  AND2_X1 U8277 ( .A1(n6588), .A2(n6587), .ZN(n6806) );
  INV_X1 U8278 ( .A(n6806), .ZN(n6589) );
  NOR2_X1 U8279 ( .A1(n6589), .A2(n6597), .ZN(n6895) );
  AOI21_X1 U8280 ( .B1(n6597), .B2(n6589), .A(n6895), .ZN(n6601) );
  INV_X1 U8281 ( .A(n6601), .ZN(n6864) );
  NAND3_X1 U8282 ( .A1(n6592), .A2(n6591), .A3(n6590), .ZN(n6859) );
  INV_X1 U8283 ( .A(n6593), .ZN(n6595) );
  INV_X1 U8284 ( .A(n6902), .ZN(n6594) );
  OAI21_X1 U8285 ( .B1(n6586), .B2(n6595), .A(n6594), .ZN(n6862) );
  OAI22_X1 U8286 ( .A1(n6862), .A2(n9869), .B1(n6586), .B2(n9868), .ZN(n6602)
         );
  AOI22_X1 U8287 ( .A1(n9574), .A2(n9285), .B1(n9283), .B2(n9572), .ZN(n6600)
         );
  OAI21_X1 U8288 ( .B1(n9821), .B2(n9285), .A(n6596), .ZN(n9006) );
  XNOR2_X1 U8289 ( .A(n9006), .B(n6597), .ZN(n6598) );
  NAND2_X1 U8290 ( .A1(n6598), .A2(n9577), .ZN(n6599) );
  OAI211_X1 U8291 ( .C1(n6601), .C2(n9601), .A(n6600), .B(n6599), .ZN(n6858)
         );
  AOI211_X1 U8292 ( .C1(n9856), .C2(n6864), .A(n6602), .B(n6858), .ZN(n9826)
         );
  NOR2_X1 U8293 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  NAND2_X1 U8294 ( .A1(n9888), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6607) );
  OAI21_X1 U8295 ( .B1(n9826), .B2(n9888), .A(n6607), .ZN(P1_U3525) );
  AOI22_X1 U8296 ( .A1(n8192), .A2(n8218), .B1(n8191), .B2(n8216), .ZN(n6618)
         );
  NAND2_X1 U8297 ( .A1(n6609), .A2(n6608), .ZN(n6726) );
  INV_X1 U8298 ( .A(n6610), .ZN(n6614) );
  INV_X1 U8299 ( .A(n6720), .ZN(n6612) );
  NAND2_X1 U8300 ( .A1(n6612), .A2(n6611), .ZN(n6613) );
  NOR2_X1 U8301 ( .A1(n6613), .A2(n6614), .ZN(n6721) );
  AOI21_X1 U8302 ( .B1(n6614), .B2(n6613), .A(n6721), .ZN(n6615) );
  NOR2_X1 U8303 ( .A1(n8202), .A2(n6615), .ZN(n6616) );
  AOI21_X1 U8304 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6726), .A(n6616), .ZN(
        n6617) );
  OAI211_X1 U8305 ( .C1(n9941), .C2(n8115), .A(n6618), .B(n6617), .ZN(P2_U3224) );
  INV_X1 U8306 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U8307 ( .A1(n10190), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n8359), .ZN(n6624) );
  INV_X1 U8308 ( .A(n6619), .ZN(n8366) );
  NAND3_X1 U8309 ( .A1(n8365), .A2(n8366), .A3(n6620), .ZN(n6621) );
  OAI211_X1 U8310 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10194), .A(n10204), .B(
        n6621), .ZN(n6622) );
  INV_X1 U8311 ( .A(n6622), .ZN(n6623) );
  MUX2_X1 U8312 ( .A(n6624), .B(n6623), .S(P2_IR_REG_0__SCAN_IN), .Z(n6626) );
  NAND2_X1 U8313 ( .A1(P2_U3152), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6625) );
  OAI211_X1 U8314 ( .C1(n8375), .C2(n6627), .A(n6626), .B(n6625), .ZN(P2_U3245) );
  INV_X1 U8315 ( .A(n6628), .ZN(n6629) );
  AOI21_X1 U8316 ( .B1(n6631), .B2(n6630), .A(n6629), .ZN(n6634) );
  AOI22_X1 U8317 ( .A1(n8984), .A2(n9285), .B1(n6859), .B2(n8978), .ZN(n6633)
         );
  AOI22_X1 U8318 ( .A1(n8971), .A2(n9283), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6644), .ZN(n6632) );
  OAI211_X1 U8319 ( .C1(n6634), .C2(n8993), .A(n6633), .B(n6632), .ZN(P1_U3235) );
  INV_X1 U8320 ( .A(n6635), .ZN(n6637) );
  NAND2_X1 U8321 ( .A1(n6637), .A2(n6636), .ZN(n6639) );
  AOI22_X1 U8322 ( .A1(n6641), .A2(n6640), .B1(n6639), .B2(n6638), .ZN(n6647)
         );
  AOI22_X1 U8323 ( .A1(n8984), .A2(n6643), .B1(n6642), .B2(n8978), .ZN(n6646)
         );
  AOI22_X1 U8324 ( .A1(n8971), .A2(n9284), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6644), .ZN(n6645) );
  OAI211_X1 U8325 ( .C1(n6647), .C2(n8993), .A(n6646), .B(n6645), .ZN(P1_U3220) );
  NOR2_X1 U8326 ( .A1(n6648), .A2(n9897), .ZN(n8233) );
  INV_X1 U8327 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n8234) );
  MUX2_X1 U8328 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n8234), .S(n8239), .Z(n6649)
         );
  OAI21_X1 U8329 ( .B1(n6650), .B2(n8233), .A(n6649), .ZN(n8251) );
  NAND2_X1 U8330 ( .A1(n8239), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8250) );
  INV_X1 U8331 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6651) );
  MUX2_X1 U8332 ( .A(n6651), .B(P2_REG2_REG_6__SCAN_IN), .S(n8253), .Z(n8249)
         );
  AOI21_X1 U8333 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8248) );
  NOR2_X1 U8334 ( .A1(n6652), .A2(n6651), .ZN(n8263) );
  INV_X1 U8335 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6965) );
  MUX2_X1 U8336 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6965), .S(n8268), .Z(n6653)
         );
  NAND2_X1 U8337 ( .A1(n8268), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8285) );
  INV_X1 U8338 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6654) );
  MUX2_X1 U8339 ( .A(n6654), .B(P2_REG2_REG_8__SCAN_IN), .S(n6672), .Z(n8284)
         );
  NOR2_X1 U8340 ( .A1(n8278), .A2(n6654), .ZN(n8292) );
  INV_X1 U8341 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7504) );
  MUX2_X1 U8342 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7504), .S(n8303), .Z(n6655)
         );
  NAND2_X1 U8343 ( .A1(n8303), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6658) );
  INV_X1 U8344 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6656) );
  MUX2_X1 U8345 ( .A(n6656), .B(P2_REG2_REG_10__SCAN_IN), .S(n6689), .Z(n6657)
         );
  AOI21_X1 U8346 ( .B1(n8295), .B2(n6658), .A(n6657), .ZN(n6688) );
  NAND3_X1 U8347 ( .A1(n8295), .A2(n6658), .A3(n6657), .ZN(n6659) );
  NAND2_X1 U8348 ( .A1(n6659), .A2(n10190), .ZN(n6680) );
  AND2_X1 U8349 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7336) );
  NOR2_X1 U8350 ( .A1(n10204), .A2(n6660), .ZN(n6661) );
  AOI211_X1 U8351 ( .C1(n10200), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7336), .B(
        n6661), .ZN(n6679) );
  INV_X1 U8352 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6662) );
  XNOR2_X1 U8353 ( .A(n6689), .B(n6662), .ZN(n6677) );
  NAND2_X1 U8354 ( .A1(n6663), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U8355 ( .A1(n6665), .A2(n6664), .ZN(n8242) );
  INV_X1 U8356 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6666) );
  XNOR2_X1 U8357 ( .A(n8239), .B(n6666), .ZN(n8243) );
  NAND2_X1 U8358 ( .A1(n8242), .A2(n8243), .ZN(n8241) );
  NAND2_X1 U8359 ( .A1(n8239), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U8360 ( .A1(n8241), .A2(n6667), .ZN(n8257) );
  INV_X1 U8361 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6668) );
  XNOR2_X1 U8362 ( .A(n8253), .B(n6668), .ZN(n8258) );
  NAND2_X1 U8363 ( .A1(n8257), .A2(n8258), .ZN(n8256) );
  NAND2_X1 U8364 ( .A1(n8253), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8365 ( .A1(n8256), .A2(n6669), .ZN(n8271) );
  INV_X1 U8366 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6670) );
  XNOR2_X1 U8367 ( .A(n8268), .B(n6670), .ZN(n8272) );
  NAND2_X1 U8368 ( .A1(n8271), .A2(n8272), .ZN(n8270) );
  NAND2_X1 U8369 ( .A1(n8268), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8370 ( .A1(n8270), .A2(n6671), .ZN(n8282) );
  INV_X1 U8371 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10141) );
  MUX2_X1 U8372 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10141), .S(n6672), .Z(n8283)
         );
  NAND2_X1 U8373 ( .A1(n8282), .A2(n8283), .ZN(n8281) );
  NAND2_X1 U8374 ( .A1(n6672), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8375 ( .A1(n8281), .A2(n6673), .ZN(n8301) );
  INV_X1 U8376 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6674) );
  XNOR2_X1 U8377 ( .A(n8303), .B(n6674), .ZN(n8302) );
  NAND2_X1 U8378 ( .A1(n8301), .A2(n8302), .ZN(n8300) );
  NAND2_X1 U8379 ( .A1(n8303), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8380 ( .A1(n8300), .A2(n6675), .ZN(n6676) );
  NAND2_X1 U8381 ( .A1(n6676), .A2(n6677), .ZN(n6682) );
  OAI211_X1 U8382 ( .C1(n6677), .C2(n6676), .A(n8359), .B(n6682), .ZN(n6678)
         );
  OAI211_X1 U8383 ( .C1(n6688), .C2(n6680), .A(n6679), .B(n6678), .ZN(P2_U3255) );
  XNOR2_X1 U8384 ( .A(n6703), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n6687) );
  NAND2_X1 U8385 ( .A1(n6689), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6681) );
  NAND2_X1 U8386 ( .A1(n6682), .A2(n6681), .ZN(n8318) );
  INV_X1 U8387 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6683) );
  XNOR2_X1 U8388 ( .A(n6690), .B(n6683), .ZN(n8317) );
  NAND2_X1 U8389 ( .A1(n8318), .A2(n8317), .ZN(n8316) );
  NAND2_X1 U8390 ( .A1(n6690), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U8391 ( .A1(n8316), .A2(n6684), .ZN(n6686) );
  INV_X1 U8392 ( .A(n6705), .ZN(n6685) );
  AOI21_X1 U8393 ( .B1(n6687), .B2(n6686), .A(n6685), .ZN(n6697) );
  AOI21_X1 U8394 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6689), .A(n6688), .ZN(
        n8309) );
  MUX2_X1 U8395 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n5414), .S(n6690), .Z(n8308)
         );
  INV_X1 U8396 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6691) );
  MUX2_X1 U8397 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6691), .S(n6703), .Z(n6692)
         );
  NAND2_X1 U8398 ( .A1(n6703), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6700) );
  OAI211_X1 U8399 ( .C1(n6703), .C2(P2_REG2_REG_12__SCAN_IN), .A(n4284), .B(
        n6700), .ZN(n6699) );
  OAI211_X1 U8400 ( .C1(n4284), .C2(n6692), .A(n6699), .B(n10190), .ZN(n6696)
         );
  AND2_X1 U8401 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7489) );
  NOR2_X1 U8402 ( .A1(n10204), .A2(n6693), .ZN(n6694) );
  AOI211_X1 U8403 ( .C1(n10200), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7489), .B(
        n6694), .ZN(n6695) );
  OAI211_X1 U8404 ( .C1(n6697), .C2(n10194), .A(n6696), .B(n6695), .ZN(
        P2_U3257) );
  NOR2_X1 U8405 ( .A1(n6845), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6839) );
  INV_X1 U8406 ( .A(n6839), .ZN(n6698) );
  OAI21_X1 U8407 ( .B1(n5468), .B2(n6708), .A(n6698), .ZN(n6702) );
  NAND2_X1 U8408 ( .A1(n6700), .A2(n6699), .ZN(n6701) );
  AOI21_X1 U8409 ( .B1(n6702), .B2(n6701), .A(n6838), .ZN(n6712) );
  OR2_X1 U8410 ( .A1(n6703), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6704) );
  NAND2_X1 U8411 ( .A1(n6705), .A2(n6704), .ZN(n6844) );
  INV_X1 U8412 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6706) );
  XNOR2_X1 U8413 ( .A(n6845), .B(n6706), .ZN(n6843) );
  XNOR2_X1 U8414 ( .A(n6844), .B(n6843), .ZN(n6707) );
  NAND2_X1 U8415 ( .A1(n6707), .A2(n8359), .ZN(n6711) );
  AND2_X1 U8416 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7574) );
  NOR2_X1 U8417 ( .A1(n10204), .A2(n6708), .ZN(n6709) );
  AOI211_X1 U8418 ( .C1(n10200), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n7574), .B(
        n6709), .ZN(n6710) );
  OAI211_X1 U8419 ( .C1(n6712), .C2(n8370), .A(n6711), .B(n6710), .ZN(P2_U3258) );
  INV_X1 U8420 ( .A(n7666), .ZN(n6804) );
  AOI22_X1 U8421 ( .A1(n8346), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8805), .ZN(n6713) );
  OAI21_X1 U8422 ( .B1(n6804), .B2(n8799), .A(n6713), .ZN(P2_U3342) );
  INV_X1 U8423 ( .A(n9911), .ZN(n6935) );
  AOI21_X1 U8424 ( .B1(n8218), .B2(n5269), .A(n8202), .ZN(n6714) );
  OAI21_X1 U8425 ( .B1(n6714), .B2(n8197), .A(n6931), .ZN(n6719) );
  NOR2_X1 U8426 ( .A1(n8202), .A2(n6715), .ZN(n8198) );
  INV_X1 U8427 ( .A(n6716), .ZN(n6717) );
  AOI22_X1 U8428 ( .A1(n8198), .A2(n6717), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n6726), .ZN(n6718) );
  OAI211_X1 U8429 ( .C1(n6935), .C2(n8166), .A(n6719), .B(n6718), .ZN(P2_U3234) );
  AOI22_X1 U8430 ( .A1(n9915), .A2(n8197), .B1(n8191), .B2(n9909), .ZN(n6729)
         );
  NOR2_X1 U8431 ( .A1(n6721), .A2(n6720), .ZN(n6725) );
  NAND2_X1 U8432 ( .A1(n6723), .A2(n6722), .ZN(n6724) );
  XNOR2_X1 U8433 ( .A(n6725), .B(n6724), .ZN(n6727) );
  AOI22_X1 U8434 ( .A1(n8162), .A2(n6727), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n6726), .ZN(n6728) );
  OAI211_X1 U8435 ( .C1(n6935), .C2(n8167), .A(n6729), .B(n6728), .ZN(P2_U3239) );
  NAND2_X1 U8436 ( .A1(n6730), .A2(n7087), .ZN(n6733) );
  AOI22_X1 U8437 ( .A1(n7734), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n4438), .B2(
        n6731), .ZN(n6732) );
  NAND2_X1 U8438 ( .A1(n6902), .A2(n9827), .ZN(n6901) );
  NAND2_X1 U8439 ( .A1(n7087), .A2(n6734), .ZN(n6739) );
  OR2_X1 U8440 ( .A1(n7678), .A2(n6735), .ZN(n6738) );
  OR2_X1 U8441 ( .A1(n9049), .A2(n6736), .ZN(n6737) );
  AOI211_X1 U8442 ( .C1(n7048), .C2(n6818), .A(n9869), .B(n6887), .ZN(n9847)
         );
  INV_X1 U8443 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6741) );
  NAND2_X1 U8444 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6740) );
  NAND2_X1 U8445 ( .A1(n6741), .A2(n6740), .ZN(n6742) );
  AND2_X1 U8446 ( .A1(n6746), .A2(n6742), .ZN(n6756) );
  INV_X1 U8447 ( .A(n6756), .ZN(n7051) );
  NOR2_X1 U8448 ( .A1(n9530), .A2(n7051), .ZN(n6763) );
  NAND2_X1 U8449 ( .A1(n6532), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6751) );
  NAND2_X1 U8450 ( .A1(n6743), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6750) );
  INV_X1 U8451 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U8452 ( .A1(n6746), .A2(n6745), .ZN(n6747) );
  AND2_X1 U8453 ( .A1(n6877), .A2(n6747), .ZN(n7126) );
  NAND2_X1 U8454 ( .A1(n4264), .A2(n7126), .ZN(n6749) );
  NAND2_X1 U8455 ( .A1(n6879), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6748) );
  NAND2_X1 U8456 ( .A1(n9283), .A2(n9827), .ZN(n9009) );
  NAND2_X1 U8457 ( .A1(n6752), .A2(n9285), .ZN(n6753) );
  NAND3_X1 U8458 ( .A1(n6754), .A2(n9004), .A3(n6753), .ZN(n6755) );
  NAND2_X1 U8459 ( .A1(n6755), .A2(n9007), .ZN(n9238) );
  NAND2_X1 U8460 ( .A1(n6896), .A2(n9230), .ZN(n6813) );
  NAND2_X1 U8461 ( .A1(n9282), .A2(n6985), .ZN(n9231) );
  OR2_X1 U8462 ( .A1(n9282), .A2(n6985), .ZN(n9011) );
  NAND2_X1 U8463 ( .A1(n6743), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U8464 ( .A1(n6532), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U8465 ( .A1(n4264), .A2(n6756), .ZN(n6758) );
  NAND2_X1 U8466 ( .A1(n6879), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6757) );
  OR2_X1 U8467 ( .A1(n9281), .A2(n9845), .ZN(n9012) );
  NAND2_X1 U8468 ( .A1(n9281), .A2(n9845), .ZN(n9232) );
  NAND2_X1 U8469 ( .A1(n9012), .A2(n9232), .ZN(n9194) );
  INV_X1 U8470 ( .A(n9194), .ZN(n6769) );
  XNOR2_X1 U8471 ( .A(n7075), .B(n9194), .ZN(n6761) );
  OAI222_X1 U8472 ( .A1(n9499), .A2(n6762), .B1(n9501), .B2(n9079), .C1(n6761), 
        .C2(n9496), .ZN(n9849) );
  AOI211_X1 U8473 ( .C1(n9261), .C2(n9847), .A(n6763), .B(n9849), .ZN(n6774)
         );
  AOI22_X1 U8474 ( .A1(n9490), .A2(n7048), .B1(n9566), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U8475 ( .A1(n9011), .A2(n9231), .ZN(n6810) );
  NAND3_X1 U8476 ( .A1(n5123), .A2(n6806), .A3(n6810), .ZN(n6768) );
  NOR2_X1 U8477 ( .A1(n9284), .A2(n6859), .ZN(n6894) );
  OR2_X1 U8478 ( .A1(n9283), .A2(n4737), .ZN(n6764) );
  NAND2_X1 U8479 ( .A1(n6765), .A2(n6764), .ZN(n6807) );
  NOR2_X1 U8480 ( .A1(n9282), .A2(n9833), .ZN(n6766) );
  NAND2_X1 U8481 ( .A1(n6768), .A2(n6767), .ZN(n7068) );
  OR2_X1 U8482 ( .A1(n7068), .A2(n6769), .ZN(n9844) );
  NAND2_X1 U8483 ( .A1(n7068), .A2(n6769), .ZN(n9843) );
  AND2_X1 U8484 ( .A1(n6770), .A2(n7890), .ZN(n6771) );
  NAND2_X1 U8485 ( .A1(n9589), .A2(n6771), .ZN(n9592) );
  INV_X1 U8486 ( .A(n9592), .ZN(n9537) );
  NAND3_X1 U8487 ( .A1(n9844), .A2(n9843), .A3(n9537), .ZN(n6772) );
  OAI211_X1 U8488 ( .C1(n6774), .C2(n9566), .A(n6773), .B(n6772), .ZN(P1_U3286) );
  XNOR2_X1 U8489 ( .A(n7286), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7129) );
  XOR2_X1 U8490 ( .A(n7129), .B(n7130), .Z(n6788) );
  INV_X1 U8491 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6779) );
  MUX2_X1 U8492 ( .A(n6779), .B(P1_REG2_REG_11__SCAN_IN), .S(n7286), .Z(n6780)
         );
  INV_X1 U8493 ( .A(n6780), .ZN(n6781) );
  NAND2_X1 U8494 ( .A1(n6782), .A2(n6781), .ZN(n7132) );
  OAI21_X1 U8495 ( .B1(n6782), .B2(n6781), .A(n7132), .ZN(n6783) );
  NAND2_X1 U8496 ( .A1(n6783), .A2(n4531), .ZN(n6787) );
  NAND2_X1 U8497 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7460) );
  OAI21_X1 U8498 ( .B1(n9791), .B2(n6784), .A(n7460), .ZN(n6785) );
  AOI21_X1 U8499 ( .B1(n9375), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6785), .ZN(
        n6786) );
  OAI211_X1 U8500 ( .C1(n9807), .C2(n6788), .A(n6787), .B(n6786), .ZN(P1_U3252) );
  NAND2_X1 U8501 ( .A1(n8596), .A2(n8213), .ZN(n6790) );
  NAND2_X1 U8502 ( .A1(n9910), .A2(n8215), .ZN(n6789) );
  NAND2_X1 U8503 ( .A1(n6790), .A2(n6789), .ZN(n7185) );
  AND2_X1 U8504 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8240) );
  INV_X1 U8505 ( .A(n6791), .ZN(n7180) );
  OAI22_X1 U8506 ( .A1(n9974), .A2(n8115), .B1(n8195), .B2(n7180), .ZN(n6792)
         );
  AOI211_X1 U8507 ( .C1(n8143), .C2(n7185), .A(n8240), .B(n6792), .ZN(n6798)
         );
  OAI21_X1 U8508 ( .B1(n6795), .B2(n6794), .A(n6793), .ZN(n6796) );
  NAND2_X1 U8509 ( .A1(n6796), .A2(n8162), .ZN(n6797) );
  NAND2_X1 U8510 ( .A1(n6798), .A2(n6797), .ZN(P2_U3229) );
  NAND2_X1 U8511 ( .A1(n6800), .A2(n6799), .ZN(n6801) );
  OAI21_X1 U8512 ( .B1(n6802), .B2(n6801), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6803) );
  XNOR2_X1 U8513 ( .A(n6803), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9340) );
  INV_X1 U8514 ( .A(n9340), .ZN(n9330) );
  OAI222_X1 U8515 ( .A1(n9743), .A2(n6805), .B1(n4261), .B2(n6804), .C1(n9330), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  NAND2_X1 U8516 ( .A1(n6806), .A2(n5123), .ZN(n6809) );
  INV_X1 U8517 ( .A(n6807), .ZN(n6808) );
  NAND2_X1 U8518 ( .A1(n6809), .A2(n6808), .ZN(n6811) );
  INV_X1 U8519 ( .A(n6810), .ZN(n9191) );
  XNOR2_X1 U8520 ( .A(n6811), .B(n9191), .ZN(n9840) );
  OAI22_X1 U8521 ( .A1(n6812), .A2(n5113), .B1(n9191), .B2(n6813), .ZN(n6817)
         );
  INV_X1 U8522 ( .A(n9281), .ZN(n6814) );
  OAI22_X1 U8523 ( .A1(n4736), .A2(n9499), .B1(n6814), .B2(n9501), .ZN(n6816)
         );
  NOR2_X1 U8524 ( .A1(n9840), .A2(n9601), .ZN(n6815) );
  AOI211_X1 U8525 ( .C1(n9577), .C2(n6817), .A(n6816), .B(n6815), .ZN(n9838)
         );
  MUX2_X1 U8526 ( .A(n6184), .B(n9838), .S(n9589), .Z(n6822) );
  AOI21_X1 U8527 ( .B1(n9833), .B2(n6901), .A(n4914), .ZN(n9836) );
  INV_X1 U8528 ( .A(n8929), .ZN(n6819) );
  OAI22_X1 U8529 ( .A1(n9586), .A2(n6985), .B1(n6819), .B2(n9530), .ZN(n6820)
         );
  AOI21_X1 U8530 ( .B1(n9836), .B2(n9581), .A(n6820), .ZN(n6821) );
  OAI211_X1 U8531 ( .C1(n9840), .C2(n7536), .A(n6822), .B(n6821), .ZN(P1_U3287) );
  XNOR2_X1 U8532 ( .A(n6824), .B(n6823), .ZN(n6829) );
  NOR2_X1 U8533 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10171), .ZN(n8269) );
  NOR2_X1 U8534 ( .A1(n8167), .A2(n6825), .ZN(n6826) );
  AOI211_X1 U8535 ( .C1(n8186), .C2(n6950), .A(n8269), .B(n6826), .ZN(n6828)
         );
  AOI22_X1 U8536 ( .A1(n7378), .A2(n8197), .B1(n8191), .B2(n8211), .ZN(n6827)
         );
  OAI211_X1 U8537 ( .C1(n6829), .C2(n8202), .A(n6828), .B(n6827), .ZN(P2_U3215) );
  OAI21_X1 U8538 ( .B1(n6832), .B2(n6831), .A(n6830), .ZN(n6836) );
  INV_X1 U8539 ( .A(n7193), .ZN(n9977) );
  OAI22_X1 U8540 ( .A1(n8166), .A2(n7206), .B1(n9977), .B2(n8115), .ZN(n6835)
         );
  NAND2_X1 U8541 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8254) );
  NAND2_X1 U8542 ( .A1(n8186), .A2(n7197), .ZN(n6833) );
  OAI211_X1 U8543 ( .C1(n8167), .C2(n4631), .A(n8254), .B(n6833), .ZN(n6834)
         );
  AOI211_X1 U8544 ( .C1(n8162), .C2(n6836), .A(n6835), .B(n6834), .ZN(n6837)
         );
  INV_X1 U8545 ( .A(n6837), .ZN(P2_U3241) );
  MUX2_X1 U8546 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n7211), .S(n7214), .Z(n6840)
         );
  INV_X1 U8547 ( .A(n6840), .ZN(n6841) );
  AOI21_X1 U8548 ( .B1(n6842), .B2(n6841), .A(n7210), .ZN(n6854) );
  NAND2_X1 U8549 ( .A1(n6844), .A2(n6843), .ZN(n6847) );
  OR2_X1 U8550 ( .A1(n6845), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U8551 ( .A1(n6847), .A2(n6846), .ZN(n7217) );
  INV_X1 U8552 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6848) );
  XNOR2_X1 U8553 ( .A(n7214), .B(n6848), .ZN(n7216) );
  XNOR2_X1 U8554 ( .A(n7217), .B(n7216), .ZN(n6849) );
  NAND2_X1 U8555 ( .A1(n6849), .A2(n8359), .ZN(n6853) );
  NOR2_X1 U8556 ( .A1(n6850), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8052) );
  NOR2_X1 U8557 ( .A1(n10204), .A2(n7212), .ZN(n6851) );
  AOI211_X1 U8558 ( .C1(n10200), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8052), .B(
        n6851), .ZN(n6852) );
  OAI211_X1 U8559 ( .C1(n6854), .C2(n8370), .A(n6853), .B(n6852), .ZN(P2_U3259) );
  INV_X1 U8560 ( .A(n7699), .ZN(n6856) );
  XNOR2_X1 U8561 ( .A(n7716), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9355) );
  AOI22_X1 U8562 ( .A1(n9355), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9740), .ZN(n6855) );
  OAI21_X1 U8563 ( .B1(n6856), .B2(n4261), .A(n6855), .ZN(P1_U3336) );
  INV_X1 U8564 ( .A(n8347), .ZN(n10203) );
  OAI222_X1 U8565 ( .A1(n8811), .A2(n6857), .B1(n8799), .B2(n6856), .C1(n10203), .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8566 ( .A(n6858), .ZN(n6866) );
  INV_X1 U8567 ( .A(n7536), .ZN(n7426) );
  AOI22_X1 U8568 ( .A1(n9566), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9582), .ZN(n6861) );
  NAND2_X1 U8569 ( .A1(n9490), .A2(n6859), .ZN(n6860) );
  OAI211_X1 U8570 ( .C1(n7995), .C2(n6862), .A(n6861), .B(n6860), .ZN(n6863)
         );
  AOI21_X1 U8571 ( .B1(n6864), .B2(n7426), .A(n6863), .ZN(n6865) );
  OAI21_X1 U8572 ( .B1(n6866), .B2(n9566), .A(n6865), .ZN(P1_U3289) );
  NAND2_X1 U8573 ( .A1(n9281), .A2(n7048), .ZN(n7069) );
  NAND2_X1 U8574 ( .A1(n9844), .A2(n7069), .ZN(n6869) );
  NAND2_X1 U8575 ( .A1(n9081), .A2(n9079), .ZN(n9239) );
  XNOR2_X1 U8576 ( .A(n6869), .B(n9195), .ZN(n6886) );
  INV_X1 U8577 ( .A(n9232), .ZN(n6872) );
  NAND2_X1 U8578 ( .A1(n5113), .A2(n9232), .ZN(n6870) );
  NAND2_X1 U8579 ( .A1(n6870), .A2(n9012), .ZN(n9235) );
  INV_X1 U8580 ( .A(n9235), .ZN(n6871) );
  OAI21_X1 U8581 ( .B1(n6812), .B2(n6872), .A(n6871), .ZN(n9077) );
  INV_X1 U8582 ( .A(n9077), .ZN(n6873) );
  XNOR2_X1 U8583 ( .A(n6873), .B(n9195), .ZN(n6874) );
  NAND2_X1 U8584 ( .A1(n6874), .A2(n9577), .ZN(n6885) );
  NAND2_X1 U8585 ( .A1(n6532), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U8586 ( .A1(n6743), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6882) );
  INV_X1 U8587 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U8588 ( .A1(n6877), .A2(n6876), .ZN(n6878) );
  AND2_X1 U8589 ( .A1(n7012), .A2(n6878), .ZN(n7081) );
  NAND2_X1 U8590 ( .A1(n4264), .A2(n7081), .ZN(n6881) );
  NAND2_X1 U8591 ( .A1(n7986), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6880) );
  INV_X1 U8592 ( .A(n9080), .ZN(n9280) );
  AOI22_X1 U8593 ( .A1(n9280), .A2(n9572), .B1(n9574), .B2(n9281), .ZN(n6884)
         );
  OAI211_X1 U8594 ( .C1(n6886), .C2(n9601), .A(n6885), .B(n6884), .ZN(n9853)
         );
  INV_X1 U8595 ( .A(n9853), .ZN(n6893) );
  INV_X1 U8596 ( .A(n6886), .ZN(n9855) );
  NOR2_X1 U8597 ( .A1(n6887), .A2(n9851), .ZN(n6888) );
  OR2_X1 U8598 ( .A1(n7080), .A2(n6888), .ZN(n9852) );
  AOI22_X1 U8599 ( .A1(n9566), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7126), .B2(
        n9582), .ZN(n6890) );
  NAND2_X1 U8600 ( .A1(n9490), .A2(n9081), .ZN(n6889) );
  OAI211_X1 U8601 ( .C1(n9852), .C2(n7995), .A(n6890), .B(n6889), .ZN(n6891)
         );
  AOI21_X1 U8602 ( .B1(n9855), .B2(n7426), .A(n6891), .ZN(n6892) );
  OAI21_X1 U8603 ( .B1(n6893), .B2(n9566), .A(n6892), .ZN(P1_U3285) );
  AOI22_X1 U8604 ( .A1(n9574), .A2(n9284), .B1(n9282), .B2(n9572), .ZN(n6899)
         );
  OAI21_X1 U8605 ( .B1(n9190), .B2(n9238), .A(n6896), .ZN(n6897) );
  NAND2_X1 U8606 ( .A1(n6897), .A2(n9577), .ZN(n6898) );
  OAI211_X1 U8607 ( .C1(n6900), .C2(n9601), .A(n6899), .B(n6898), .ZN(n9829)
         );
  INV_X1 U8608 ( .A(n9829), .ZN(n6908) );
  INV_X1 U8609 ( .A(n6900), .ZN(n9831) );
  OAI21_X1 U8610 ( .B1(n6902), .B2(n9827), .A(n6901), .ZN(n9828) );
  AOI22_X1 U8611 ( .A1(n9566), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9582), .B2(
        n6903), .ZN(n6905) );
  NAND2_X1 U8612 ( .A1(n9490), .A2(n4737), .ZN(n6904) );
  OAI211_X1 U8613 ( .C1(n7995), .C2(n9828), .A(n6905), .B(n6904), .ZN(n6906)
         );
  AOI21_X1 U8614 ( .B1(n9831), .B2(n7426), .A(n6906), .ZN(n6907) );
  OAI21_X1 U8615 ( .B1(n6908), .B2(n9566), .A(n6907), .ZN(P1_U3288) );
  XNOR2_X1 U8616 ( .A(n6910), .B(n6909), .ZN(n6916) );
  INV_X1 U8617 ( .A(n7470), .ZN(n6911) );
  NAND2_X1 U8618 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8277) );
  OAI21_X1 U8619 ( .B1(n8195), .B2(n6911), .A(n8277), .ZN(n6914) );
  OAI22_X1 U8620 ( .A1(n8166), .A2(n6912), .B1(n4983), .B2(n8115), .ZN(n6913)
         );
  AOI211_X1 U8621 ( .C1(n8192), .C2(n8212), .A(n6914), .B(n6913), .ZN(n6915)
         );
  OAI21_X1 U8622 ( .B1(n8202), .B2(n6916), .A(n6915), .ZN(P2_U3223) );
  INV_X1 U8623 ( .A(n6917), .ZN(n6918) );
  NAND2_X1 U8624 ( .A1(n6918), .A2(n7145), .ZN(n6920) );
  INV_X1 U8625 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6921) );
  OAI22_X1 U8626 ( .A1(n8651), .A2(n6922), .B1(n6921), .B2(n9919), .ZN(n6928)
         );
  OR2_X1 U8627 ( .A1(n6923), .A2(n4954), .ZN(n7053) );
  NAND2_X1 U8628 ( .A1(n8581), .A2(n7053), .ZN(n6924) );
  INV_X1 U8629 ( .A(n6925), .ZN(n6926) );
  NOR2_X1 U8630 ( .A1(n9924), .A2(n6926), .ZN(n6927) );
  AOI211_X1 U8631 ( .C1(n8651), .C2(P2_REG2_REG_0__SCAN_IN), .A(n6928), .B(
        n6927), .ZN(n6933) );
  NOR2_X2 U8632 ( .A1(n6930), .A2(n5322), .ZN(n8629) );
  OAI21_X1 U8633 ( .B1(n8653), .B2(n8629), .A(n6931), .ZN(n6932) );
  NAND2_X1 U8634 ( .A1(n6933), .A2(n6932), .ZN(P2_U3296) );
  INV_X1 U8635 ( .A(n6934), .ZN(n7038) );
  NAND2_X1 U8636 ( .A1(n7038), .A2(n7037), .ZN(n7036) );
  NAND2_X1 U8637 ( .A1(n6935), .A2(n9941), .ZN(n6936) );
  NAND2_X1 U8638 ( .A1(n6938), .A2(n9948), .ZN(n6939) );
  INV_X1 U8639 ( .A(n9909), .ZN(n6941) );
  NAND2_X1 U8640 ( .A1(n6942), .A2(n9965), .ZN(n6943) );
  AOI21_X1 U8641 ( .B1(n7179), .B2(n4631), .A(n9974), .ZN(n6945) );
  NAND2_X1 U8642 ( .A1(n7193), .A2(n8213), .ZN(n6947) );
  XNOR2_X1 U8643 ( .A(n7376), .B(n7377), .ZN(n7143) );
  NAND2_X1 U8644 ( .A1(n9941), .A2(n7032), .ZN(n9916) );
  NAND2_X1 U8645 ( .A1(n9917), .A2(n7054), .ZN(n9899) );
  INV_X1 U8646 ( .A(n6949), .ZN(n7196) );
  INV_X1 U8647 ( .A(n7378), .ZN(n6948) );
  AOI21_X1 U8648 ( .B1(n7378), .B2(n7196), .A(n4360), .ZN(n7140) );
  INV_X1 U8649 ( .A(n7140), .ZN(n6952) );
  INV_X1 U8650 ( .A(n6950), .ZN(n6951) );
  OAI22_X1 U8651 ( .A1(n6952), .A2(n9921), .B1(n6951), .B2(n9919), .ZN(n6953)
         );
  AOI21_X1 U8652 ( .B1(n8653), .B2(n7378), .A(n6953), .ZN(n6967) );
  OAI21_X1 U8653 ( .B1(n6954), .B2(n6956), .A(n6955), .ZN(n6958) );
  NAND2_X1 U8654 ( .A1(n6958), .A2(n6957), .ZN(n6959) );
  NAND2_X1 U8655 ( .A1(n6959), .A2(n7377), .ZN(n6962) );
  NAND3_X1 U8656 ( .A1(n6962), .A2(n6961), .A3(n9913), .ZN(n6964) );
  AOI22_X1 U8657 ( .A1(n8596), .A2(n8211), .B1(n9910), .B2(n8213), .ZN(n6963)
         );
  AND2_X1 U8658 ( .A1(n6964), .A2(n6963), .ZN(n7142) );
  MUX2_X1 U8659 ( .A(n7142), .B(n6965), .S(n8651), .Z(n6966) );
  OAI211_X1 U8660 ( .C1(n7143), .C2(n9924), .A(n6967), .B(n6966), .ZN(P2_U3289) );
  NAND2_X1 U8661 ( .A1(n6968), .A2(n7087), .ZN(n6971) );
  AOI22_X1 U8662 ( .A1(n7734), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4438), .B2(
        n6969), .ZN(n6970) );
  NAND2_X1 U8663 ( .A1(n6971), .A2(n6970), .ZN(n7108) );
  NAND2_X1 U8664 ( .A1(n7108), .A2(n7893), .ZN(n6973) );
  OR2_X1 U8665 ( .A1(n9080), .A2(n7875), .ZN(n6972) );
  NAND2_X1 U8666 ( .A1(n6973), .A2(n6972), .ZN(n6974) );
  XNOR2_X1 U8667 ( .A(n6974), .B(n7890), .ZN(n7234) );
  XNOR2_X1 U8668 ( .A(n7234), .B(n7235), .ZN(n7008) );
  INV_X1 U8669 ( .A(n6976), .ZN(n6977) );
  AND2_X1 U8670 ( .A1(n6978), .A2(n6977), .ZN(n6979) );
  NAND2_X1 U8671 ( .A1(n9282), .A2(n7900), .ZN(n6983) );
  OR2_X1 U8672 ( .A1(n6985), .A2(n6524), .ZN(n6982) );
  NAND2_X1 U8673 ( .A1(n6983), .A2(n6982), .ZN(n6984) );
  XNOR2_X1 U8674 ( .A(n6984), .B(n7763), .ZN(n6988) );
  OR2_X1 U8675 ( .A1(n6985), .A2(n7875), .ZN(n6986) );
  NAND2_X1 U8676 ( .A1(n6987), .A2(n6986), .ZN(n6989) );
  XNOR2_X1 U8677 ( .A(n6988), .B(n6989), .ZN(n8926) );
  INV_X1 U8678 ( .A(n6988), .ZN(n6990) );
  NAND2_X1 U8679 ( .A1(n6990), .A2(n6989), .ZN(n6991) );
  NAND2_X1 U8680 ( .A1(n9081), .A2(n7893), .ZN(n6992) );
  OAI21_X1 U8681 ( .B1(n9079), .B2(n7875), .A(n6992), .ZN(n6993) );
  XNOR2_X1 U8682 ( .A(n6993), .B(n7763), .ZN(n7119) );
  OR2_X1 U8683 ( .A1(n9079), .A2(n7898), .ZN(n6995) );
  NAND2_X1 U8684 ( .A1(n9081), .A2(n7900), .ZN(n6994) );
  AND2_X1 U8685 ( .A1(n6995), .A2(n6994), .ZN(n7118) );
  NAND2_X1 U8686 ( .A1(n9281), .A2(n7900), .ZN(n6996) );
  OAI21_X1 U8687 ( .B1(n9845), .B2(n6524), .A(n6996), .ZN(n6997) );
  XNOR2_X1 U8688 ( .A(n6997), .B(n7763), .ZN(n7041) );
  OR2_X1 U8689 ( .A1(n9845), .A2(n7875), .ZN(n6999) );
  AND2_X1 U8690 ( .A1(n6999), .A2(n6998), .ZN(n7043) );
  OAI22_X1 U8691 ( .A1(n7119), .A2(n7118), .B1(n7041), .B2(n7043), .ZN(n7000)
         );
  INV_X1 U8692 ( .A(n7041), .ZN(n7117) );
  INV_X1 U8693 ( .A(n7043), .ZN(n7001) );
  INV_X1 U8694 ( .A(n7118), .ZN(n7002) );
  OAI21_X1 U8695 ( .B1(n7117), .B2(n7001), .A(n7002), .ZN(n7004) );
  NOR2_X1 U8696 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  AOI22_X1 U8697 ( .A1(n7004), .A2(n7119), .B1(n7041), .B2(n7003), .ZN(n7005)
         );
  OAI21_X1 U8698 ( .B1(n7008), .B2(n7007), .A(n7238), .ZN(n7009) );
  NAND2_X1 U8699 ( .A1(n7009), .A2(n8964), .ZN(n7023) );
  NAND2_X1 U8700 ( .A1(n6532), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7017) );
  NAND2_X1 U8701 ( .A1(n6743), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7016) );
  INV_X1 U8702 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7011) );
  NAND2_X1 U8703 ( .A1(n7012), .A2(n7011), .ZN(n7013) );
  AND2_X1 U8704 ( .A1(n7096), .A2(n7013), .ZN(n7245) );
  NAND2_X1 U8705 ( .A1(n4264), .A2(n7245), .ZN(n7015) );
  NAND2_X1 U8706 ( .A1(n7986), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7014) );
  INV_X1 U8707 ( .A(n7018), .ZN(n7019) );
  AOI21_X1 U8708 ( .B1(n8984), .B2(n4928), .A(n7019), .ZN(n7020) );
  OAI21_X1 U8709 ( .B1(n7239), .B2(n8986), .A(n7020), .ZN(n7021) );
  AOI21_X1 U8710 ( .B1(n7081), .B2(n8991), .A(n7021), .ZN(n7022) );
  OAI211_X1 U8711 ( .C1(n9859), .C2(n8988), .A(n7023), .B(n7022), .ZN(P1_U3211) );
  INV_X1 U8712 ( .A(n7024), .ZN(n7028) );
  INV_X1 U8713 ( .A(n7025), .ZN(n7026) );
  NAND2_X1 U8714 ( .A1(n7026), .A2(n7037), .ZN(n7027) );
  OAI211_X1 U8715 ( .C1(n7029), .C2(n7028), .A(n9913), .B(n7027), .ZN(n7031)
         );
  AOI22_X1 U8716 ( .A1(n9910), .A2(n8218), .B1(n8596), .B2(n8216), .ZN(n7030)
         );
  AND2_X1 U8717 ( .A1(n7031), .A2(n7030), .ZN(n9943) );
  NOR2_X1 U8718 ( .A1(n8651), .A2(n9943), .ZN(n7035) );
  OAI21_X1 U8719 ( .B1(n9941), .B2(n7032), .A(n9916), .ZN(n9942) );
  OAI22_X1 U8720 ( .A1(n9921), .A2(n9942), .B1(n7033), .B2(n9919), .ZN(n7034)
         );
  AOI211_X1 U8721 ( .C1(n8651), .C2(P2_REG2_REG_1__SCAN_IN), .A(n7035), .B(
        n7034), .ZN(n7040) );
  OAI21_X1 U8722 ( .B1(n7038), .B2(n7037), .A(n7036), .ZN(n9946) );
  NAND2_X1 U8723 ( .A1(n8611), .A2(n9946), .ZN(n7039) );
  OAI211_X1 U8724 ( .C1(n9941), .C2(n9925), .A(n7040), .B(n7039), .ZN(P2_U3295) );
  XNOR2_X1 U8725 ( .A(n7116), .B(n7041), .ZN(n7042) );
  NAND2_X1 U8726 ( .A1(n7042), .A2(n7043), .ZN(n7115) );
  OAI21_X1 U8727 ( .B1(n7043), .B2(n7042), .A(n7115), .ZN(n7044) );
  NAND2_X1 U8728 ( .A1(n7044), .A2(n8964), .ZN(n7050) );
  AOI21_X1 U8729 ( .B1(n8984), .B2(n9282), .A(n7045), .ZN(n7046) );
  OAI21_X1 U8730 ( .B1(n9079), .B2(n8986), .A(n7046), .ZN(n7047) );
  AOI21_X1 U8731 ( .B1(n7048), .B2(n8978), .A(n7047), .ZN(n7049) );
  OAI211_X1 U8732 ( .C1(n8966), .C2(n7051), .A(n7050), .B(n7049), .ZN(P1_U3225) );
  XNOR2_X1 U8733 ( .A(n7052), .B(n7058), .ZN(n7063) );
  INV_X1 U8734 ( .A(n7063), .ZN(n9961) );
  OR2_X1 U8735 ( .A1(n8651), .A2(n7053), .ZN(n8588) );
  INV_X1 U8736 ( .A(n7054), .ZN(n9955) );
  OR2_X1 U8737 ( .A1(n9917), .A2(n7054), .ZN(n7055) );
  AND2_X1 U8738 ( .A1(n9899), .A2(n7055), .ZN(n9958) );
  NAND2_X1 U8739 ( .A1(n8629), .A2(n9958), .ZN(n7056) );
  OAI21_X1 U8740 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n9919), .A(n7056), .ZN(
        n7057) );
  AOI21_X1 U8741 ( .B1(n8653), .B2(n9955), .A(n7057), .ZN(n7066) );
  INV_X1 U8742 ( .A(n8581), .ZN(n8645) );
  XNOR2_X1 U8743 ( .A(n7059), .B(n7058), .ZN(n7061) );
  AOI22_X1 U8744 ( .A1(n9910), .A2(n8216), .B1(n8596), .B2(n8215), .ZN(n7060)
         );
  OAI21_X1 U8745 ( .B1(n7061), .B2(n9892), .A(n7060), .ZN(n7062) );
  AOI21_X1 U8746 ( .B1(n8645), .B2(n7063), .A(n7062), .ZN(n9960) );
  MUX2_X1 U8747 ( .A(n9960), .B(n7064), .S(n8651), .Z(n7065) );
  OAI211_X1 U8748 ( .C1(n9961), .C2(n8588), .A(n7066), .B(n7065), .ZN(P2_U3293) );
  NAND2_X1 U8749 ( .A1(n7068), .A2(n7067), .ZN(n7074) );
  INV_X1 U8750 ( .A(n7069), .ZN(n7070) );
  NOR2_X1 U8751 ( .A1(n9194), .A2(n7070), .ZN(n7072) );
  NOR2_X1 U8752 ( .A1(n9081), .A2(n4928), .ZN(n7071) );
  OR2_X1 U8753 ( .A1(n7108), .A2(n9080), .ZN(n9242) );
  NAND2_X1 U8754 ( .A1(n7108), .A2(n9080), .ZN(n9073) );
  XNOR2_X1 U8755 ( .A(n7107), .B(n9187), .ZN(n9862) );
  INV_X1 U8756 ( .A(n9862), .ZN(n7086) );
  AND2_X1 U8757 ( .A1(n9081), .A2(n9079), .ZN(n7077) );
  NAND2_X1 U8758 ( .A1(n7076), .A2(n9239), .ZN(n9236) );
  OR2_X1 U8759 ( .A1(n7164), .A2(n9187), .ZN(n7090) );
  INV_X1 U8760 ( .A(n7090), .ZN(n7078) );
  AOI21_X1 U8761 ( .B1(n9187), .B2(n7164), .A(n7078), .ZN(n7079) );
  OAI222_X1 U8762 ( .A1(n9501), .A2(n7239), .B1(n9499), .B2(n9079), .C1(n9496), 
        .C2(n7079), .ZN(n9860) );
  OAI211_X1 U8763 ( .C1(n7080), .C2(n9859), .A(n9835), .B(n7105), .ZN(n9858)
         );
  AOI22_X1 U8764 ( .A1(n9566), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7081), .B2(
        n9582), .ZN(n7083) );
  NAND2_X1 U8765 ( .A1(n9490), .A2(n7108), .ZN(n7082) );
  OAI211_X1 U8766 ( .C1(n9858), .C2(n7324), .A(n7083), .B(n7082), .ZN(n7084)
         );
  AOI21_X1 U8767 ( .B1(n9860), .B2(n9589), .A(n7084), .ZN(n7085) );
  OAI21_X1 U8768 ( .B1(n7086), .B2(n9592), .A(n7085), .ZN(P1_U3284) );
  AOI22_X1 U8769 ( .A1(n7734), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4438), .B2(
        n9805), .ZN(n7089) );
  NAND2_X1 U8770 ( .A1(n9867), .A2(n7239), .ZN(n9095) );
  AND2_X1 U8771 ( .A1(n9095), .A2(n9073), .ZN(n8998) );
  NAND2_X1 U8772 ( .A1(n7090), .A2(n8998), .ZN(n7094) );
  OR2_X1 U8773 ( .A1(n9867), .A2(n7239), .ZN(n9015) );
  NAND2_X1 U8774 ( .A1(n7090), .A2(n9073), .ZN(n7092) );
  INV_X1 U8775 ( .A(n9199), .ZN(n7091) );
  NAND2_X1 U8776 ( .A1(n7092), .A2(n7091), .ZN(n7093) );
  OAI211_X1 U8777 ( .C1(n7094), .C2(n9091), .A(n7093), .B(n9577), .ZN(n7104)
         );
  NAND2_X1 U8778 ( .A1(n6743), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7101) );
  NAND2_X1 U8779 ( .A1(n6879), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7100) );
  NAND2_X1 U8780 ( .A1(n7096), .A2(n7095), .ZN(n7097) );
  AND2_X1 U8781 ( .A1(n7158), .A2(n7097), .ZN(n7272) );
  NAND2_X1 U8782 ( .A1(n4264), .A2(n7272), .ZN(n7099) );
  NAND2_X1 U8783 ( .A1(n6532), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7098) );
  OAI22_X1 U8784 ( .A1(n9080), .A2(n9499), .B1(n7618), .B2(n9501), .ZN(n7102)
         );
  INV_X1 U8785 ( .A(n7102), .ZN(n7103) );
  NAND2_X1 U8786 ( .A1(n7104), .A2(n7103), .ZN(n9873) );
  MUX2_X1 U8787 ( .A(n9873), .B(P1_REG2_REG_8__SCAN_IN), .S(n9566), .Z(n7114)
         );
  NAND2_X1 U8788 ( .A1(n7105), .A2(n9867), .ZN(n7106) );
  NAND2_X1 U8789 ( .A1(n7171), .A2(n7106), .ZN(n9870) );
  OR2_X1 U8790 ( .A1(n7108), .A2(n9280), .ZN(n7109) );
  NAND2_X1 U8791 ( .A1(n7110), .A2(n9199), .ZN(n9864) );
  NAND3_X1 U8792 ( .A1(n9866), .A2(n9864), .A3(n9537), .ZN(n7112) );
  AOI22_X1 U8793 ( .A1(n9867), .A2(n9490), .B1(n7245), .B2(n9582), .ZN(n7111)
         );
  OAI211_X1 U8794 ( .C1(n7995), .C2(n9870), .A(n7112), .B(n7111), .ZN(n7113)
         );
  OR2_X1 U8795 ( .A1(n7114), .A2(n7113), .ZN(P1_U3283) );
  OAI21_X1 U8796 ( .B1(n7117), .B2(n7116), .A(n7115), .ZN(n7121) );
  XNOR2_X1 U8797 ( .A(n7119), .B(n7118), .ZN(n7120) );
  XNOR2_X1 U8798 ( .A(n7121), .B(n7120), .ZN(n7128) );
  NOR2_X1 U8799 ( .A1(n8988), .A2(n9851), .ZN(n7125) );
  NAND2_X1 U8800 ( .A1(n8984), .A2(n9281), .ZN(n7123) );
  OAI211_X1 U8801 ( .C1(n8986), .C2(n9080), .A(n7123), .B(n7122), .ZN(n7124)
         );
  AOI211_X1 U8802 ( .C1(n7126), .C2(n8991), .A(n7125), .B(n7124), .ZN(n7127)
         );
  OAI21_X1 U8803 ( .B1(n7128), .B2(n8993), .A(n7127), .ZN(P1_U3237) );
  XOR2_X1 U8804 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7297), .Z(n7251) );
  XNOR2_X1 U8805 ( .A(n7252), .B(n7251), .ZN(n7138) );
  NAND2_X1 U8806 ( .A1(n9375), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7131) );
  NAND2_X1 U8807 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7565) );
  OAI211_X1 U8808 ( .C1(n9791), .C2(n7250), .A(n7131), .B(n7565), .ZN(n7137)
         );
  XNOR2_X1 U8809 ( .A(n7297), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7135) );
  AOI211_X1 U8810 ( .C1(n7135), .C2(n7134), .A(n9799), .B(n7133), .ZN(n7136)
         );
  AOI211_X1 U8811 ( .C1(n9790), .C2(n7138), .A(n7137), .B(n7136), .ZN(n7139)
         );
  INV_X1 U8812 ( .A(n7139), .ZN(P1_U3253) );
  INV_X1 U8813 ( .A(n9986), .ZN(n9957) );
  AOI22_X1 U8814 ( .A1(n7140), .A2(n9957), .B1(n9956), .B2(n7378), .ZN(n7141)
         );
  OAI211_X1 U8815 ( .C1(n7143), .C2(n8751), .A(n7142), .B(n7141), .ZN(n7147)
         );
  NAND2_X1 U8816 ( .A1(n7147), .A2(n10004), .ZN(n7144) );
  OAI21_X1 U8817 ( .B1(n10004), .B2(n6670), .A(n7144), .ZN(P2_U3527) );
  INV_X1 U8818 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U8819 ( .A1(n7147), .A2(n9994), .ZN(n7148) );
  OAI21_X1 U8820 ( .B1(n9994), .B2(n7149), .A(n7148), .ZN(P2_U3472) );
  INV_X1 U8821 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7150) );
  INV_X1 U8822 ( .A(n8361), .ZN(n8350) );
  OAI222_X1 U8823 ( .A1(n8811), .A2(n7150), .B1(n8799), .B2(n7910), .C1(
        P2_U3152), .C2(n8350), .ZN(P2_U3340) );
  INV_X1 U8824 ( .A(n7733), .ZN(n7177) );
  OAI222_X1 U8825 ( .A1(n8811), .A2(n7151), .B1(n8799), .B2(n7177), .C1(n4954), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U8826 ( .A(n7239), .ZN(n9279) );
  NAND2_X1 U8827 ( .A1(n9867), .A2(n9279), .ZN(n7152) );
  NAND2_X1 U8828 ( .A1(n7153), .A2(n7087), .ZN(n7156) );
  AOI22_X1 U8829 ( .A1(n7734), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4438), .B2(
        n7154), .ZN(n7155) );
  OR2_X1 U8830 ( .A1(n9699), .A2(n7618), .ZN(n9092) );
  NAND2_X1 U8831 ( .A1(n9699), .A2(n7618), .ZN(n9090) );
  AND2_X1 U8832 ( .A1(n9092), .A2(n9090), .ZN(n9200) );
  XNOR2_X1 U8833 ( .A(n7327), .B(n9200), .ZN(n9698) );
  INV_X1 U8834 ( .A(n9601), .ZN(n7531) );
  NAND2_X1 U8835 ( .A1(n6743), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U8836 ( .A1(n6879), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7162) );
  OR2_X2 U8837 ( .A1(n7158), .A2(n7157), .ZN(n7291) );
  NAND2_X1 U8838 ( .A1(n7158), .A2(n7157), .ZN(n7159) );
  AND2_X1 U8839 ( .A1(n7291), .A2(n7159), .ZN(n7622) );
  NAND2_X1 U8840 ( .A1(n4264), .A2(n7622), .ZN(n7161) );
  NAND2_X1 U8841 ( .A1(n6532), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7160) );
  OAI22_X1 U8842 ( .A1(n7239), .A2(n9499), .B1(n7364), .B2(n9501), .ZN(n7170)
         );
  INV_X1 U8843 ( .A(n7164), .ZN(n7165) );
  INV_X1 U8844 ( .A(n7280), .ZN(n7168) );
  OAI21_X1 U8845 ( .B1(n7166), .B2(n9200), .A(n9577), .ZN(n7167) );
  AOI21_X1 U8846 ( .B1(n7168), .B2(n9092), .A(n7167), .ZN(n7169) );
  AOI211_X1 U8847 ( .C1(n9698), .C2(n7531), .A(n7170), .B(n7169), .ZN(n9702)
         );
  INV_X1 U8848 ( .A(n9699), .ZN(n7174) );
  AOI21_X1 U8849 ( .B1(n9699), .B2(n7171), .A(n7619), .ZN(n9700) );
  NAND2_X1 U8850 ( .A1(n9700), .A2(n9581), .ZN(n7173) );
  AOI22_X1 U8851 ( .A1(n9566), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7272), .B2(
        n9582), .ZN(n7172) );
  OAI211_X1 U8852 ( .C1(n7174), .C2(n9586), .A(n7173), .B(n7172), .ZN(n7175)
         );
  AOI21_X1 U8853 ( .B1(n7426), .B2(n9698), .A(n7175), .ZN(n7176) );
  OAI21_X1 U8854 ( .B1(n9702), .B2(n9566), .A(n7176), .ZN(P1_U3282) );
  OAI222_X1 U8855 ( .A1(n7178), .A2(n9743), .B1(P1_U3084), .B2(n9261), .C1(
        n4261), .C2(n7177), .ZN(P1_U3334) );
  XNOR2_X1 U8856 ( .A(n7179), .B(n7184), .ZN(n9976) );
  OAI22_X1 U8857 ( .A1(n9925), .A2(n9974), .B1(n9919), .B2(n7180), .ZN(n7189)
         );
  INV_X1 U8858 ( .A(n7181), .ZN(n7182) );
  OAI211_X1 U8859 ( .C1(n7182), .C2(n9974), .A(n7194), .B(n9957), .ZN(n9972)
         );
  INV_X1 U8860 ( .A(n6954), .ZN(n7183) );
  NAND2_X1 U8861 ( .A1(n7183), .A2(n9903), .ZN(n9896) );
  NAND2_X1 U8862 ( .A1(n9896), .A2(n4689), .ZN(n7202) );
  XNOR2_X1 U8863 ( .A(n7202), .B(n7184), .ZN(n7186) );
  AOI21_X1 U8864 ( .B1(n7186), .B2(n9913), .A(n7185), .ZN(n9973) );
  OAI21_X1 U8865 ( .B1(n8435), .B2(n9972), .A(n9973), .ZN(n7187) );
  MUX2_X1 U8866 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7187), .S(n8606), .Z(n7188)
         );
  AOI211_X1 U8867 ( .C1(n8611), .C2(n9976), .A(n7189), .B(n7188), .ZN(n7190)
         );
  INV_X1 U8868 ( .A(n7190), .ZN(P2_U3291) );
  XNOR2_X1 U8869 ( .A(n7192), .B(n7191), .ZN(n9982) );
  NAND2_X1 U8870 ( .A1(n7194), .A2(n7193), .ZN(n7195) );
  NAND2_X1 U8871 ( .A1(n7196), .A2(n7195), .ZN(n9978) );
  INV_X1 U8872 ( .A(n9978), .ZN(n7198) );
  AOI22_X1 U8873 ( .A1(n8629), .A2(n7198), .B1(n7197), .B2(n8649), .ZN(n7199)
         );
  OAI21_X1 U8874 ( .B1(n9925), .B2(n9977), .A(n7199), .ZN(n7208) );
  INV_X1 U8875 ( .A(n9910), .ZN(n8641) );
  OAI21_X1 U8876 ( .B1(n7202), .B2(n7201), .A(n7200), .ZN(n7204) );
  XNOR2_X1 U8877 ( .A(n7204), .B(n7203), .ZN(n7205) );
  OAI222_X1 U8878 ( .A1(n8641), .A2(n4631), .B1(n8640), .B2(n7206), .C1(n7205), 
        .C2(n9892), .ZN(n9979) );
  MUX2_X1 U8879 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9979), .S(n8606), .Z(n7207)
         );
  AOI211_X1 U8880 ( .C1(n8611), .C2(n9982), .A(n7208), .B(n7207), .ZN(n7209)
         );
  INV_X1 U8881 ( .A(n7209), .ZN(P2_U3290) );
  AOI21_X1 U8882 ( .B1(n7213), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8323), .ZN(
        n7224) );
  NOR2_X1 U8883 ( .A1(n7214), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7215) );
  AOI21_X1 U8884 ( .B1(n7217), .B2(n7216), .A(n7215), .ZN(n8331) );
  XOR2_X1 U8885 ( .A(n8330), .B(n8331), .Z(n7219) );
  AND2_X1 U8886 ( .A1(n7219), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8329) );
  INV_X1 U8887 ( .A(n8329), .ZN(n7218) );
  OAI211_X1 U8888 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n7219), .A(n7218), .B(
        n8359), .ZN(n7223) );
  INV_X1 U8889 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7220) );
  NAND2_X1 U8890 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8193) );
  OAI21_X1 U8891 ( .B1(n8375), .B2(n7220), .A(n8193), .ZN(n7221) );
  AOI21_X1 U8892 ( .B1(n8335), .B2(n8330), .A(n7221), .ZN(n7222) );
  OAI211_X1 U8893 ( .C1(n7224), .C2(n8370), .A(n7223), .B(n7222), .ZN(P2_U3260) );
  AOI21_X1 U8894 ( .B1(n7226), .B2(n7225), .A(n4366), .ZN(n7230) );
  NAND2_X1 U8895 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8298) );
  OAI21_X1 U8896 ( .B1(n8195), .B2(n7507), .A(n8298), .ZN(n7228) );
  OAI22_X1 U8897 ( .A1(n8166), .A2(n7375), .B1(n4982), .B2(n8115), .ZN(n7227)
         );
  AOI211_X1 U8898 ( .C1(n8192), .C2(n8211), .A(n7228), .B(n7227), .ZN(n7229)
         );
  OAI21_X1 U8899 ( .B1(n7230), .B2(n8202), .A(n7229), .ZN(P2_U3233) );
  NAND2_X1 U8900 ( .A1(n9867), .A2(n7893), .ZN(n7232) );
  OR2_X1 U8901 ( .A1(n7239), .A2(n7875), .ZN(n7231) );
  NAND2_X1 U8902 ( .A1(n7232), .A2(n7231), .ZN(n7233) );
  XNOR2_X1 U8903 ( .A(n7233), .B(n7890), .ZN(n7263) );
  INV_X1 U8904 ( .A(n7234), .ZN(n7236) );
  NAND2_X1 U8905 ( .A1(n7236), .A2(n7235), .ZN(n7237) );
  NOR2_X1 U8906 ( .A1(n7239), .A2(n7898), .ZN(n7240) );
  AOI21_X1 U8907 ( .B1(n9867), .B2(n7892), .A(n7240), .ZN(n7241) );
  NAND2_X1 U8908 ( .A1(n4367), .A2(n7264), .ZN(n7242) );
  XOR2_X1 U8909 ( .A(n7263), .B(n7242), .Z(n7248) );
  NAND2_X1 U8910 ( .A1(n8984), .A2(n9280), .ZN(n7243) );
  NAND2_X1 U8911 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9793) );
  OAI211_X1 U8912 ( .C1(n8986), .C2(n7618), .A(n7243), .B(n9793), .ZN(n7244)
         );
  AOI21_X1 U8913 ( .B1(n7245), .B2(n8991), .A(n7244), .ZN(n7247) );
  NAND2_X1 U8914 ( .A1(n9867), .A2(n8978), .ZN(n7246) );
  OAI211_X1 U8915 ( .C1(n7248), .C2(n8993), .A(n7247), .B(n7246), .ZN(P1_U3219) );
  XNOR2_X1 U8916 ( .A(n9293), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9286) );
  INV_X1 U8917 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7249) );
  XOR2_X1 U8918 ( .A(n9286), .B(n9287), .Z(n7262) );
  XNOR2_X1 U8919 ( .A(n9293), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7255) );
  AOI211_X1 U8920 ( .C1(n7256), .C2(n7255), .A(n9799), .B(n9292), .ZN(n7257)
         );
  INV_X1 U8921 ( .A(n7257), .ZN(n7261) );
  NOR2_X1 U8922 ( .A1(n7313), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8949) );
  NOR2_X1 U8923 ( .A1(n9791), .A2(n7258), .ZN(n7259) );
  AOI211_X1 U8924 ( .C1(n9375), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n8949), .B(
        n7259), .ZN(n7260) );
  OAI211_X1 U8925 ( .C1(n9807), .C2(n7262), .A(n7261), .B(n7260), .ZN(P1_U3254) );
  NAND2_X1 U8926 ( .A1(n9699), .A2(n7893), .ZN(n7266) );
  OR2_X1 U8927 ( .A1(n7618), .A2(n7875), .ZN(n7265) );
  NAND2_X1 U8928 ( .A1(n7266), .A2(n7265), .ZN(n7267) );
  XNOR2_X1 U8929 ( .A(n7267), .B(n7763), .ZN(n7343) );
  NOR2_X1 U8930 ( .A1(n7618), .A2(n7898), .ZN(n7268) );
  AOI21_X1 U8931 ( .B1(n9699), .B2(n7892), .A(n7268), .ZN(n7342) );
  XNOR2_X1 U8932 ( .A(n7343), .B(n7342), .ZN(n7345) );
  XOR2_X1 U8933 ( .A(n7346), .B(n7345), .Z(n7275) );
  NAND2_X1 U8934 ( .A1(n8984), .A2(n9279), .ZN(n7270) );
  OAI211_X1 U8935 ( .C1(n8986), .C2(n7364), .A(n7270), .B(n7269), .ZN(n7271)
         );
  AOI21_X1 U8936 ( .B1(n7272), .B2(n8991), .A(n7271), .ZN(n7274) );
  NAND2_X1 U8937 ( .A1(n9699), .A2(n8978), .ZN(n7273) );
  OAI211_X1 U8938 ( .C1(n7275), .C2(n8993), .A(n7274), .B(n7273), .ZN(P1_U3229) );
  INV_X1 U8939 ( .A(n7748), .ZN(n7277) );
  OAI222_X1 U8940 ( .A1(P1_U3084), .A2(n7276), .B1(n4261), .B2(n7277), .C1(
        n7749), .C2(n9743), .ZN(P1_U3333) );
  OAI222_X1 U8941 ( .A1(n8811), .A2(n7279), .B1(P2_U3152), .B2(n7278), .C1(
        n8799), .C2(n7277), .ZN(P2_U3338) );
  NAND2_X1 U8942 ( .A1(n7281), .A2(n7087), .ZN(n7284) );
  AOI22_X1 U8943 ( .A1(n7734), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4438), .B2(
        n7282), .ZN(n7283) );
  NAND2_X1 U8944 ( .A1(n9694), .A2(n7364), .ZN(n9093) );
  NAND2_X1 U8945 ( .A1(n7285), .A2(n7087), .ZN(n7288) );
  AOI22_X1 U8946 ( .A1(n7734), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4438), .B2(
        n7286), .ZN(n7287) );
  NAND2_X1 U8947 ( .A1(n6532), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7296) );
  NAND2_X1 U8948 ( .A1(n6743), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7295) );
  INV_X1 U8949 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7290) );
  NAND2_X1 U8950 ( .A1(n7291), .A2(n7290), .ZN(n7292) );
  AND2_X1 U8951 ( .A1(n7300), .A2(n7292), .ZN(n7463) );
  NAND2_X1 U8952 ( .A1(n4264), .A2(n7463), .ZN(n7294) );
  NAND2_X1 U8953 ( .A1(n6879), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7293) );
  NAND2_X1 U8954 ( .A1(n7455), .A2(n7615), .ZN(n8999) );
  NAND2_X1 U8955 ( .A1(n7362), .A2(n8999), .ZN(n7526) );
  NAND2_X1 U8956 ( .A1(n7526), .A2(n7525), .ZN(n7312) );
  NAND2_X1 U8957 ( .A1(n7308), .A2(n7087), .ZN(n7322) );
  AOI22_X1 U8958 ( .A1(n7734), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4438), .B2(
        n7297), .ZN(n7321) );
  NAND2_X1 U8959 ( .A1(n6743), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7305) );
  NAND2_X1 U8960 ( .A1(n6879), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7304) );
  INV_X1 U8961 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7299) );
  NAND2_X1 U8962 ( .A1(n7300), .A2(n7299), .ZN(n7301) );
  AND2_X1 U8963 ( .A1(n7314), .A2(n7301), .ZN(n7568) );
  NAND2_X1 U8964 ( .A1(n4264), .A2(n7568), .ZN(n7303) );
  NAND2_X1 U8965 ( .A1(n6532), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7302) );
  AND2_X1 U8966 ( .A1(n7321), .A2(n7309), .ZN(n7306) );
  NAND2_X1 U8967 ( .A1(n7322), .A2(n7306), .ZN(n9110) );
  AND2_X1 U8968 ( .A1(n7087), .A2(n8951), .ZN(n7307) );
  NAND2_X1 U8969 ( .A1(n7308), .A2(n7307), .ZN(n7311) );
  INV_X1 U8970 ( .A(n8951), .ZN(n7309) );
  OR2_X1 U8971 ( .A1(n7309), .A2(n7321), .ZN(n7310) );
  NAND2_X1 U8972 ( .A1(n7311), .A2(n7310), .ZN(n9016) );
  INV_X1 U8973 ( .A(n9016), .ZN(n9094) );
  NAND2_X1 U8974 ( .A1(n9110), .A2(n9094), .ZN(n9186) );
  XNOR2_X1 U8975 ( .A(n7312), .B(n9186), .ZN(n7320) );
  INV_X1 U8976 ( .A(n7615), .ZN(n9276) );
  NAND2_X1 U8977 ( .A1(n6532), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7319) );
  NAND2_X1 U8978 ( .A1(n6743), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7318) );
  NAND2_X1 U8979 ( .A1(n7314), .A2(n7313), .ZN(n7315) );
  AND2_X1 U8980 ( .A1(n7519), .A2(n7315), .ZN(n8953) );
  NAND2_X1 U8981 ( .A1(n4264), .A2(n8953), .ZN(n7317) );
  NAND2_X1 U8982 ( .A1(n6879), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7316) );
  INV_X1 U8983 ( .A(n8834), .ZN(n9275) );
  AOI222_X1 U8984 ( .A1(n9577), .A2(n7320), .B1(n9276), .B2(n9574), .C1(n9275), 
        .C2(n9572), .ZN(n9690) );
  INV_X1 U8985 ( .A(n9694), .ZN(n7624) );
  INV_X1 U8986 ( .A(n7533), .ZN(n7323) );
  AOI211_X1 U8987 ( .C1(n9688), .C2(n7361), .A(n9869), .B(n7323), .ZN(n9687)
         );
  INV_X1 U8988 ( .A(n7324), .ZN(n9564) );
  AOI22_X1 U8989 ( .A1(n9566), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7568), .B2(
        n9582), .ZN(n7325) );
  OAI21_X1 U8990 ( .B1(n4911), .B2(n9586), .A(n7325), .ZN(n7332) );
  INV_X1 U8991 ( .A(n7618), .ZN(n9278) );
  OR2_X1 U8992 ( .A1(n9699), .A2(n9278), .ZN(n7326) );
  NAND2_X1 U8993 ( .A1(n9699), .A2(n9278), .ZN(n7328) );
  NAND2_X1 U8994 ( .A1(n7525), .A2(n8999), .ZN(n7359) );
  INV_X1 U8995 ( .A(n7364), .ZN(n9277) );
  OR2_X1 U8996 ( .A1(n9694), .A2(n9277), .ZN(n7358) );
  AND2_X1 U8997 ( .A1(n7359), .A2(n7358), .ZN(n7329) );
  AOI22_X1 U8998 ( .A1(n7329), .A2(n9203), .B1(n9276), .B2(n7455), .ZN(n7330)
         );
  XNOR2_X1 U8999 ( .A(n7514), .B(n9186), .ZN(n9691) );
  NOR2_X1 U9000 ( .A1(n9691), .A2(n9592), .ZN(n7331) );
  AOI211_X1 U9001 ( .C1(n9687), .C2(n9564), .A(n7332), .B(n7331), .ZN(n7333)
         );
  OAI21_X1 U9002 ( .B1(n9690), .B2(n9566), .A(n7333), .ZN(P1_U3279) );
  XOR2_X1 U9003 ( .A(n7335), .B(n7334), .Z(n7340) );
  INV_X1 U9004 ( .A(n8759), .ZN(n7400) );
  AOI22_X1 U9005 ( .A1(n8191), .A2(n8208), .B1(n8192), .B2(n8210), .ZN(n7338)
         );
  AOI21_X1 U9006 ( .B1(n8186), .B2(n7398), .A(n7336), .ZN(n7337) );
  OAI211_X1 U9007 ( .C1(n7400), .C2(n8115), .A(n7338), .B(n7337), .ZN(n7339)
         );
  AOI21_X1 U9008 ( .B1(n7340), .B2(n8162), .A(n7339), .ZN(n7341) );
  INV_X1 U9009 ( .A(n7341), .ZN(P2_U3219) );
  NAND2_X1 U9010 ( .A1(n7343), .A2(n7342), .ZN(n7344) );
  NAND2_X1 U9011 ( .A1(n9694), .A2(n7893), .ZN(n7348) );
  OR2_X1 U9012 ( .A1(n7364), .A2(n7875), .ZN(n7347) );
  NAND2_X1 U9013 ( .A1(n7348), .A2(n7347), .ZN(n7349) );
  XNOR2_X1 U9014 ( .A(n7349), .B(n7890), .ZN(n7447) );
  NOR2_X1 U9015 ( .A1(n7364), .A2(n7898), .ZN(n7350) );
  AOI21_X1 U9016 ( .B1(n9694), .B2(n7892), .A(n7350), .ZN(n7448) );
  XNOR2_X1 U9017 ( .A(n7447), .B(n7448), .ZN(n7445) );
  XOR2_X1 U9018 ( .A(n7446), .B(n7445), .Z(n7356) );
  NAND2_X1 U9019 ( .A1(n8984), .A2(n9278), .ZN(n7352) );
  OAI211_X1 U9020 ( .C1(n8986), .C2(n7615), .A(n7352), .B(n7351), .ZN(n7354)
         );
  NOR2_X1 U9021 ( .A1(n7624), .A2(n8988), .ZN(n7353) );
  AOI211_X1 U9022 ( .C1(n7622), .C2(n8991), .A(n7354), .B(n7353), .ZN(n7355)
         );
  OAI21_X1 U9023 ( .B1(n7356), .B2(n8993), .A(n7355), .ZN(P1_U3215) );
  OR2_X1 U9024 ( .A1(n7357), .A2(n9203), .ZN(n7611) );
  NAND2_X1 U9025 ( .A1(n7611), .A2(n7358), .ZN(n7360) );
  INV_X1 U9026 ( .A(n7359), .ZN(n9102) );
  XNOR2_X1 U9027 ( .A(n7360), .B(n9102), .ZN(n7368) );
  INV_X1 U9028 ( .A(n7368), .ZN(n7425) );
  OAI21_X1 U9029 ( .B1(n7620), .B2(n7466), .A(n7361), .ZN(n7421) );
  OAI22_X1 U9030 ( .A1(n7421), .A2(n9869), .B1(n7466), .B2(n9868), .ZN(n7369)
         );
  XNOR2_X1 U9031 ( .A(n7362), .B(n7359), .ZN(n7363) );
  NAND2_X1 U9032 ( .A1(n7363), .A2(n9577), .ZN(n7367) );
  OAI22_X1 U9033 ( .A1(n7364), .A2(n9499), .B1(n8951), .B2(n9501), .ZN(n7365)
         );
  INV_X1 U9034 ( .A(n7365), .ZN(n7366) );
  OAI211_X1 U9035 ( .C1(n7368), .C2(n9601), .A(n7367), .B(n7366), .ZN(n7422)
         );
  AOI211_X1 U9036 ( .C1(n9856), .C2(n7425), .A(n7369), .B(n7422), .ZN(n7372)
         );
  NAND2_X1 U9037 ( .A1(n9874), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7370) );
  OAI21_X1 U9038 ( .B1(n7372), .B2(n9874), .A(n7370), .ZN(P1_U3487) );
  NAND2_X1 U9039 ( .A1(n9888), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7371) );
  OAI21_X1 U9040 ( .B1(n7372), .B2(n9888), .A(n7371), .ZN(P1_U3534) );
  XNOR2_X1 U9041 ( .A(n7373), .B(n7435), .ZN(n7374) );
  OAI222_X1 U9042 ( .A1(n8641), .A2(n7375), .B1(n8640), .B2(n8642), .C1(n9892), 
        .C2(n7374), .ZN(n7414) );
  INV_X1 U9043 ( .A(n7414), .ZN(n7388) );
  AND2_X1 U9044 ( .A1(n7471), .A2(n8211), .ZN(n7495) );
  NOR2_X1 U9045 ( .A1(n7499), .A2(n7495), .ZN(n7379) );
  NAND2_X1 U9046 ( .A1(n7468), .A2(n7379), .ZN(n7381) );
  INV_X1 U9047 ( .A(n7389), .ZN(n7391) );
  NAND2_X1 U9048 ( .A1(n8759), .A2(n8209), .ZN(n7382) );
  XNOR2_X1 U9049 ( .A(n7436), .B(n7383), .ZN(n7416) );
  INV_X1 U9050 ( .A(n7437), .ZN(n7412) );
  NAND2_X1 U9051 ( .A1(n7397), .A2(n7412), .ZN(n7438) );
  OAI21_X1 U9052 ( .B1(n7397), .B2(n7412), .A(n7438), .ZN(n7413) );
  AOI22_X1 U9053 ( .A1(n8651), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7406), .B2(
        n8649), .ZN(n7385) );
  NAND2_X1 U9054 ( .A1(n8653), .A2(n7437), .ZN(n7384) );
  OAI211_X1 U9055 ( .C1(n7413), .C2(n9921), .A(n7385), .B(n7384), .ZN(n7386)
         );
  AOI21_X1 U9056 ( .B1(n7416), .B2(n8611), .A(n7386), .ZN(n7387) );
  OAI21_X1 U9057 ( .B1(n7388), .B2(n8651), .A(n7387), .ZN(P2_U3285) );
  XNOR2_X1 U9058 ( .A(n7390), .B(n7389), .ZN(n7396) );
  INV_X1 U9059 ( .A(n7396), .ZN(n8763) );
  XNOR2_X1 U9060 ( .A(n7392), .B(n7391), .ZN(n7394) );
  AOI22_X1 U9061 ( .A1(n8596), .A2(n8208), .B1(n9910), .B2(n8210), .ZN(n7393)
         );
  OAI21_X1 U9062 ( .B1(n7394), .B2(n9892), .A(n7393), .ZN(n7395) );
  AOI21_X1 U9063 ( .B1(n7396), .B2(n8645), .A(n7395), .ZN(n8762) );
  MUX2_X1 U9064 ( .A(n6656), .B(n8762), .S(n8606), .Z(n7403) );
  AOI21_X1 U9065 ( .B1(n8759), .B2(n4984), .A(n7397), .ZN(n8760) );
  INV_X1 U9066 ( .A(n7398), .ZN(n7399) );
  OAI22_X1 U9067 ( .A1(n9925), .A2(n7400), .B1(n9919), .B2(n7399), .ZN(n7401)
         );
  AOI21_X1 U9068 ( .B1(n8760), .B2(n8629), .A(n7401), .ZN(n7402) );
  OAI211_X1 U9069 ( .C1(n8763), .C2(n8588), .A(n7403), .B(n7402), .ZN(P2_U3286) );
  XOR2_X1 U9070 ( .A(n7405), .B(n7404), .Z(n7410) );
  AOI22_X1 U9071 ( .A1(n8191), .A2(n8207), .B1(n8192), .B2(n8209), .ZN(n7408)
         );
  AOI22_X1 U9072 ( .A1(n8186), .A2(n7406), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n7407) );
  OAI211_X1 U9073 ( .C1(n7412), .C2(n8115), .A(n7408), .B(n7407), .ZN(n7409)
         );
  AOI21_X1 U9074 ( .B1(n7410), .B2(n8162), .A(n7409), .ZN(n7411) );
  INV_X1 U9075 ( .A(n7411), .ZN(P2_U3238) );
  INV_X1 U9076 ( .A(n7773), .ZN(n7553) );
  OAI222_X1 U9077 ( .A1(n9743), .A2(n7774), .B1(n4261), .B2(n7553), .C1(n9224), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  OAI22_X1 U9078 ( .A1(n7413), .A2(n9986), .B1(n7412), .B2(n9985), .ZN(n7415)
         );
  AOI211_X1 U9079 ( .C1(n7416), .C2(n9981), .A(n7415), .B(n7414), .ZN(n7419)
         );
  NAND2_X1 U9080 ( .A1(n9992), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7417) );
  OAI21_X1 U9081 ( .B1(n7419), .B2(n9992), .A(n7417), .ZN(P2_U3484) );
  NAND2_X1 U9082 ( .A1(n10002), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7418) );
  OAI21_X1 U9083 ( .B1(n7419), .B2(n10002), .A(n7418), .ZN(P2_U3531) );
  AOI22_X1 U9084 ( .A1(n7455), .A2(n9490), .B1(n7463), .B2(n9582), .ZN(n7420)
         );
  OAI21_X1 U9085 ( .B1(n7421), .B2(n7995), .A(n7420), .ZN(n7424) );
  MUX2_X1 U9086 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7422), .S(n9589), .Z(n7423)
         );
  AOI211_X1 U9087 ( .C1(n7426), .C2(n7425), .A(n7424), .B(n7423), .ZN(n7427)
         );
  INV_X1 U9088 ( .A(n7427), .ZN(P1_U3280) );
  NAND2_X1 U9089 ( .A1(n7429), .A2(n7428), .ZN(n7431) );
  XNOR2_X1 U9090 ( .A(n7431), .B(n7430), .ZN(n7432) );
  OAI222_X1 U9091 ( .A1(n8641), .A2(n7434), .B1(n8640), .B2(n7433), .C1(n7432), 
        .C2(n9892), .ZN(n7545) );
  INV_X1 U9092 ( .A(n7545), .ZN(n7444) );
  XNOR2_X1 U9093 ( .A(n8004), .B(n8003), .ZN(n7547) );
  INV_X1 U9094 ( .A(n8034), .ZN(n8646) );
  NAND2_X1 U9095 ( .A1(n7438), .A2(n8002), .ZN(n7439) );
  NAND2_X1 U9096 ( .A1(n8646), .A2(n7439), .ZN(n7544) );
  AOI22_X1 U9097 ( .A1(n8651), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7490), .B2(
        n8649), .ZN(n7441) );
  NAND2_X1 U9098 ( .A1(n8653), .A2(n8002), .ZN(n7440) );
  OAI211_X1 U9099 ( .C1(n7544), .C2(n9921), .A(n7441), .B(n7440), .ZN(n7442)
         );
  AOI21_X1 U9100 ( .B1(n7547), .B2(n8611), .A(n7442), .ZN(n7443) );
  OAI21_X1 U9101 ( .B1(n7444), .B2(n8651), .A(n7443), .ZN(P2_U3284) );
  INV_X1 U9102 ( .A(n7447), .ZN(n7449) );
  NAND2_X1 U9103 ( .A1(n7449), .A2(n7448), .ZN(n7450) );
  NAND2_X1 U9104 ( .A1(n7455), .A2(n7893), .ZN(n7452) );
  OR2_X1 U9105 ( .A1(n7615), .A2(n7875), .ZN(n7451) );
  NAND2_X1 U9106 ( .A1(n7452), .A2(n7451), .ZN(n7453) );
  XNOR2_X1 U9107 ( .A(n7453), .B(n7763), .ZN(n7557) );
  NOR2_X1 U9108 ( .A1(n7615), .A2(n7898), .ZN(n7454) );
  AOI21_X1 U9109 ( .B1(n7455), .B2(n7892), .A(n7454), .ZN(n7556) );
  XNOR2_X1 U9110 ( .A(n7557), .B(n7556), .ZN(n7457) );
  AOI21_X1 U9111 ( .B1(n7456), .B2(n7457), .A(n8993), .ZN(n7459) );
  INV_X1 U9112 ( .A(n7457), .ZN(n7458) );
  NAND2_X1 U9113 ( .A1(n7459), .A2(n7559), .ZN(n7465) );
  NAND2_X1 U9114 ( .A1(n8984), .A2(n9277), .ZN(n7461) );
  OAI211_X1 U9115 ( .C1(n8986), .C2(n8951), .A(n7461), .B(n7460), .ZN(n7462)
         );
  AOI21_X1 U9116 ( .B1(n7463), .B2(n8991), .A(n7462), .ZN(n7464) );
  OAI211_X1 U9117 ( .C1(n7466), .C2(n8988), .A(n7465), .B(n7464), .ZN(P1_U3234) );
  INV_X1 U9118 ( .A(n7792), .ZN(n7963) );
  OAI222_X1 U9119 ( .A1(n9743), .A2(n7793), .B1(n4261), .B2(n7963), .C1(
        P1_U3084), .C2(n9227), .ZN(P1_U3331) );
  AND2_X1 U9120 ( .A1(n7468), .A2(n7467), .ZN(n7469) );
  NOR2_X1 U9121 ( .A1(n7468), .A2(n7467), .ZN(n7496) );
  OR2_X1 U9122 ( .A1(n7469), .A2(n7496), .ZN(n7481) );
  INV_X1 U9123 ( .A(n7481), .ZN(n9990) );
  INV_X1 U9124 ( .A(n8588), .ZN(n8657) );
  OAI21_X1 U9125 ( .B1(n4360), .B2(n4983), .A(n7506), .ZN(n9987) );
  AOI22_X1 U9126 ( .A1(n8653), .A2(n7471), .B1(n8649), .B2(n7470), .ZN(n7472)
         );
  OAI21_X1 U9127 ( .B1(n9921), .B2(n9987), .A(n7472), .ZN(n7483) );
  AOI22_X1 U9128 ( .A1(n9910), .A2(n8212), .B1(n8596), .B2(n8210), .ZN(n7480)
         );
  NAND2_X1 U9129 ( .A1(n7475), .A2(n7474), .ZN(n7476) );
  NAND2_X1 U9130 ( .A1(n7477), .A2(n7476), .ZN(n7478) );
  NAND2_X1 U9131 ( .A1(n7478), .A2(n9913), .ZN(n7479) );
  OAI211_X1 U9132 ( .C1(n7481), .C2(n8581), .A(n7480), .B(n7479), .ZN(n9988)
         );
  MUX2_X1 U9133 ( .A(n9988), .B(P2_REG2_REG_8__SCAN_IN), .S(n8651), .Z(n7482)
         );
  AOI211_X1 U9134 ( .C1(n9990), .C2(n8657), .A(n7483), .B(n7482), .ZN(n7484)
         );
  INV_X1 U9135 ( .A(n7484), .ZN(P2_U3288) );
  NAND2_X1 U9136 ( .A1(n7486), .A2(n7485), .ZN(n7487) );
  AOI21_X1 U9137 ( .B1(n7488), .B2(n7487), .A(n8202), .ZN(n7494) );
  INV_X1 U9138 ( .A(n8002), .ZN(n7543) );
  AOI22_X1 U9139 ( .A1(n8191), .A2(n8619), .B1(n8192), .B2(n8208), .ZN(n7492)
         );
  AOI21_X1 U9140 ( .B1(n8186), .B2(n7490), .A(n7489), .ZN(n7491) );
  OAI211_X1 U9141 ( .C1(n7543), .C2(n8115), .A(n7492), .B(n7491), .ZN(n7493)
         );
  OR2_X1 U9142 ( .A1(n7494), .A2(n7493), .ZN(P2_U3226) );
  NOR2_X1 U9143 ( .A1(n7496), .A2(n7495), .ZN(n7497) );
  XOR2_X1 U9144 ( .A(n7499), .B(n7497), .Z(n7503) );
  INV_X1 U9145 ( .A(n7503), .ZN(n8768) );
  XOR2_X1 U9146 ( .A(n7499), .B(n7498), .Z(n7501) );
  AOI22_X1 U9147 ( .A1(n9910), .A2(n8211), .B1(n8596), .B2(n8209), .ZN(n7500)
         );
  OAI21_X1 U9148 ( .B1(n7501), .B2(n9892), .A(n7500), .ZN(n7502) );
  AOI21_X1 U9149 ( .B1(n7503), .B2(n8645), .A(n7502), .ZN(n8767) );
  MUX2_X1 U9150 ( .A(n7504), .B(n8767), .S(n8606), .Z(n7510) );
  AOI21_X1 U9151 ( .B1(n8764), .B2(n7506), .A(n7505), .ZN(n8765) );
  OAI22_X1 U9152 ( .A1(n9925), .A2(n4982), .B1(n9919), .B2(n7507), .ZN(n7508)
         );
  AOI21_X1 U9153 ( .B1(n8629), .B2(n8765), .A(n7508), .ZN(n7509) );
  OAI211_X1 U9154 ( .C1(n8768), .C2(n8588), .A(n7510), .B(n7509), .ZN(P2_U3287) );
  NAND2_X1 U9155 ( .A1(n7511), .A2(n7087), .ZN(n7513) );
  AOI22_X1 U9156 ( .A1(n7734), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4438), .B2(
        n9293), .ZN(n7512) );
  OR2_X1 U9157 ( .A1(n9682), .A2(n8834), .ZN(n9105) );
  NAND2_X1 U9158 ( .A1(n9682), .A2(n8834), .ZN(n9106) );
  NAND2_X1 U9159 ( .A1(n9105), .A2(n9106), .ZN(n9206) );
  NAND2_X1 U9160 ( .A1(n9688), .A2(n7309), .ZN(n7515) );
  XOR2_X1 U9161 ( .A(n9206), .B(n7581), .Z(n7535) );
  INV_X1 U9162 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U9163 ( .A1(n7519), .A2(n7518), .ZN(n7520) );
  NAND2_X1 U9164 ( .A1(n7592), .A2(n7520), .ZN(n8835) );
  OR2_X1 U9165 ( .A1(n7868), .A2(n8835), .ZN(n7524) );
  NAND2_X1 U9166 ( .A1(n6743), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U9167 ( .A1(n6879), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U9168 ( .A1(n6532), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7521) );
  OAI22_X1 U9169 ( .A1(n7662), .A2(n9501), .B1(n8951), .B2(n9499), .ZN(n7530)
         );
  AND2_X1 U9170 ( .A1(n9110), .A2(n7525), .ZN(n9017) );
  AOI21_X1 U9171 ( .B1(n7527), .B2(n9206), .A(n7590), .ZN(n7528) );
  NOR2_X1 U9172 ( .A1(n7528), .A2(n9496), .ZN(n7529) );
  AOI211_X1 U9173 ( .C1(n7535), .C2(n7531), .A(n7530), .B(n7529), .ZN(n9685)
         );
  INV_X1 U9174 ( .A(n7585), .ZN(n7532) );
  AOI21_X1 U9175 ( .B1(n9682), .B2(n7533), .A(n7532), .ZN(n9683) );
  AOI22_X1 U9176 ( .A1(n9566), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8953), .B2(
        n9582), .ZN(n7534) );
  OAI21_X1 U9177 ( .B1(n4910), .B2(n9586), .A(n7534), .ZN(n7538) );
  INV_X1 U9178 ( .A(n7535), .ZN(n9686) );
  NOR2_X1 U9179 ( .A1(n9686), .A2(n7536), .ZN(n7537) );
  AOI211_X1 U9180 ( .C1(n9683), .C2(n9581), .A(n7538), .B(n7537), .ZN(n7539)
         );
  OAI21_X1 U9181 ( .B1(n9685), .B2(n9566), .A(n7539), .ZN(P1_U3278) );
  INV_X1 U9182 ( .A(n7821), .ZN(n7542) );
  AOI21_X1 U9183 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8805), .A(n7540), .ZN(
        n7541) );
  OAI21_X1 U9184 ( .B1(n7542), .B2(n8799), .A(n7541), .ZN(P2_U3335) );
  OAI22_X1 U9185 ( .A1(n7544), .A2(n9986), .B1(n7543), .B2(n9985), .ZN(n7546)
         );
  AOI211_X1 U9186 ( .C1(n7547), .C2(n9981), .A(n7546), .B(n7545), .ZN(n7550)
         );
  NAND2_X1 U9187 ( .A1(n10002), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7548) );
  OAI21_X1 U9188 ( .B1(n7550), .B2(n10002), .A(n7548), .ZN(P2_U3532) );
  NAND2_X1 U9189 ( .A1(n9992), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7549) );
  OAI21_X1 U9190 ( .B1(n7550), .B2(n9992), .A(n7549), .ZN(P2_U3487) );
  NAND2_X1 U9191 ( .A1(n7821), .A2(n9735), .ZN(n7552) );
  OR2_X1 U9192 ( .A1(n7551), .A2(P1_U3084), .ZN(n9265) );
  OAI211_X1 U9193 ( .C1(n7822), .C2(n9743), .A(n7552), .B(n9265), .ZN(P1_U3330) );
  OAI222_X1 U9194 ( .A1(n8811), .A2(n7555), .B1(P2_U3152), .B2(n7554), .C1(
        n8799), .C2(n7553), .ZN(P2_U3337) );
  OR2_X1 U9195 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  NAND2_X1 U9196 ( .A1(n7559), .A2(n7558), .ZN(n7654) );
  NAND2_X1 U9197 ( .A1(n9688), .A2(n7893), .ZN(n7561) );
  OR2_X1 U9198 ( .A1(n8951), .A2(n7875), .ZN(n7560) );
  NAND2_X1 U9199 ( .A1(n7561), .A2(n7560), .ZN(n7562) );
  XNOR2_X1 U9200 ( .A(n7562), .B(n7763), .ZN(n7655) );
  NOR2_X1 U9201 ( .A1(n8951), .A2(n7898), .ZN(n7563) );
  AOI21_X1 U9202 ( .B1(n9688), .B2(n7892), .A(n7563), .ZN(n7652) );
  INV_X1 U9203 ( .A(n7652), .ZN(n7656) );
  XNOR2_X1 U9204 ( .A(n7655), .B(n7656), .ZN(n7564) );
  XNOR2_X1 U9205 ( .A(n7654), .B(n7564), .ZN(n7571) );
  NAND2_X1 U9206 ( .A1(n8984), .A2(n9276), .ZN(n7566) );
  OAI211_X1 U9207 ( .C1(n8986), .C2(n8834), .A(n7566), .B(n7565), .ZN(n7567)
         );
  AOI21_X1 U9208 ( .B1(n7568), .B2(n8991), .A(n7567), .ZN(n7570) );
  NAND2_X1 U9209 ( .A1(n9688), .A2(n8978), .ZN(n7569) );
  OAI211_X1 U9210 ( .C1(n7571), .C2(n8993), .A(n7570), .B(n7569), .ZN(P1_U3222) );
  XOR2_X1 U9211 ( .A(n7573), .B(n7572), .Z(n7578) );
  INV_X1 U9212 ( .A(n8652), .ZN(n8753) );
  AOI22_X1 U9213 ( .A1(n8192), .A2(n8207), .B1(n8191), .B2(n8595), .ZN(n7576)
         );
  AOI21_X1 U9214 ( .B1(n8186), .B2(n8650), .A(n7574), .ZN(n7575) );
  OAI211_X1 U9215 ( .C1(n8753), .C2(n8115), .A(n7576), .B(n7575), .ZN(n7577)
         );
  AOI21_X1 U9216 ( .B1(n7578), .B2(n8162), .A(n7577), .ZN(n7579) );
  INV_X1 U9217 ( .A(n7579), .ZN(P2_U3236) );
  AND2_X1 U9218 ( .A1(n9682), .A2(n9275), .ZN(n7580) );
  NAND2_X1 U9219 ( .A1(n7582), .A2(n7087), .ZN(n7584) );
  AOI22_X1 U9220 ( .A1(n7734), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4438), .B2(
        n9311), .ZN(n7583) );
  INV_X1 U9221 ( .A(n7588), .ZN(n9208) );
  XNOR2_X1 U9222 ( .A(n7922), .B(n9208), .ZN(n9681) );
  AOI211_X1 U9223 ( .C1(n9678), .C2(n7585), .A(n9578), .B(n9869), .ZN(n9677)
         );
  INV_X1 U9224 ( .A(n9678), .ZN(n8840) );
  INV_X1 U9225 ( .A(n8835), .ZN(n7586) );
  AOI22_X1 U9226 ( .A1(n9566), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7586), .B2(
        n9582), .ZN(n7587) );
  OAI21_X1 U9227 ( .B1(n8840), .B2(n9586), .A(n7587), .ZN(n7601) );
  INV_X1 U9228 ( .A(n9106), .ZN(n7589) );
  NOR2_X1 U9229 ( .A1(n7951), .A2(n9496), .ZN(n7599) );
  OAI21_X1 U9230 ( .B1(n7590), .B2(n7589), .A(n7588), .ZN(n7598) );
  INV_X1 U9231 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7591) );
  NAND2_X1 U9232 ( .A1(n7592), .A2(n7591), .ZN(n7593) );
  AND2_X1 U9233 ( .A1(n7670), .A2(n7593), .ZN(n9583) );
  NAND2_X1 U9234 ( .A1(n9583), .A2(n4264), .ZN(n7596) );
  AOI22_X1 U9235 ( .A1(n6532), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n6743), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U9236 ( .A1(n7986), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7594) );
  OAI22_X1 U9237 ( .A1(n7952), .A2(n9501), .B1(n8834), .B2(n9499), .ZN(n7597)
         );
  AOI21_X1 U9238 ( .B1(n7599), .B2(n7598), .A(n7597), .ZN(n9680) );
  NOR2_X1 U9239 ( .A1(n9680), .A2(n9566), .ZN(n7600) );
  AOI211_X1 U9240 ( .C1(n9677), .C2(n9564), .A(n7601), .B(n7600), .ZN(n7602)
         );
  OAI21_X1 U9241 ( .B1(n9681), .B2(n9592), .A(n7602), .ZN(P1_U3277) );
  INV_X1 U9242 ( .A(n7603), .ZN(n7604) );
  INV_X1 U9243 ( .A(n7807), .ZN(n7605) );
  OAI222_X1 U9244 ( .A1(n7604), .A2(P2_U3152), .B1(n8799), .B2(n7605), .C1(
        n10169), .C2(n8811), .ZN(P2_U3334) );
  OAI222_X1 U9245 ( .A1(P1_U3084), .A2(n7606), .B1(n4261), .B2(n7605), .C1(
        n7808), .C2(n9743), .ZN(P1_U3329) );
  INV_X1 U9246 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10160) );
  INV_X1 U9247 ( .A(n9044), .ZN(n8001) );
  OAI222_X1 U9248 ( .A1(n8811), .A2(n10160), .B1(n8799), .B2(n8001), .C1(n7607), .C2(P2_U3152), .ZN(P2_U3328) );
  OAI222_X1 U9249 ( .A1(n7610), .A2(P1_U3084), .B1(n4261), .B2(n7609), .C1(
        n7608), .C2(n9743), .ZN(P1_U3352) );
  INV_X1 U9250 ( .A(n7611), .ZN(n7612) );
  AOI21_X1 U9251 ( .B1(n9203), .B2(n7357), .A(n7612), .ZN(n9696) );
  OAI211_X1 U9252 ( .C1(n7614), .C2(n9203), .A(n7613), .B(n9577), .ZN(n7617)
         );
  OR2_X1 U9253 ( .A1(n7615), .A2(n9501), .ZN(n7616) );
  OAI211_X1 U9254 ( .C1(n7618), .C2(n9499), .A(n7617), .B(n7616), .ZN(n9692)
         );
  NAND2_X1 U9255 ( .A1(n9692), .A2(n9589), .ZN(n7627) );
  INV_X1 U9256 ( .A(n7619), .ZN(n7621) );
  AOI211_X1 U9257 ( .C1(n9694), .C2(n7621), .A(n9869), .B(n7620), .ZN(n9693)
         );
  AOI22_X1 U9258 ( .A1(n9566), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7622), .B2(
        n9582), .ZN(n7623) );
  OAI21_X1 U9259 ( .B1(n7624), .B2(n9586), .A(n7623), .ZN(n7625) );
  AOI21_X1 U9260 ( .B1(n9693), .B2(n9564), .A(n7625), .ZN(n7626) );
  OAI211_X1 U9261 ( .C1(n9592), .C2(n9696), .A(n7627), .B(n7626), .ZN(P1_U3281) );
  INV_X1 U9262 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7702) );
  OR2_X2 U9263 ( .A1(n7703), .A2(n7702), .ZN(n7720) );
  NAND2_X1 U9264 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n7629) );
  INV_X1 U9265 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8967) );
  INV_X1 U9266 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8846) );
  INV_X1 U9267 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7640) );
  OR2_X2 U9268 ( .A1(n7848), .A2(n7640), .ZN(n7866) );
  INV_X1 U9269 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7881) );
  INV_X1 U9270 ( .A(n7994), .ZN(n7636) );
  INV_X1 U9271 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7634) );
  NAND2_X1 U9272 ( .A1(n7986), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7633) );
  NAND2_X1 U9273 ( .A1(n6743), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7632) );
  OAI211_X1 U9274 ( .C1(n7990), .C2(n7634), .A(n7633), .B(n7632), .ZN(n7635)
         );
  NAND2_X1 U9275 ( .A1(n9274), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7637) );
  OAI21_X1 U9276 ( .B1(n9391), .B2(n9274), .A(n7637), .ZN(P1_U3584) );
  OR2_X1 U9277 ( .A1(n4635), .A2(n9744), .ZN(n7638) );
  NAND2_X1 U9278 ( .A1(n7848), .A2(n7640), .ZN(n7641) );
  AND2_X2 U9279 ( .A1(n7866), .A2(n7641), .ZN(n9424) );
  NAND2_X1 U9280 ( .A1(n9424), .A2(n4264), .ZN(n7647) );
  INV_X1 U9281 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U9282 ( .A1(n7986), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7643) );
  NAND2_X1 U9283 ( .A1(n6743), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7642) );
  OAI211_X1 U9284 ( .C1(n7990), .C2(n7644), .A(n7643), .B(n7642), .ZN(n7645)
         );
  INV_X1 U9285 ( .A(n7645), .ZN(n7646) );
  NOR2_X1 U9286 ( .A1(n9412), .A2(n7898), .ZN(n7648) );
  AOI21_X1 U9287 ( .B1(n9616), .B2(n7900), .A(n7648), .ZN(n7859) );
  INV_X1 U9288 ( .A(n7859), .ZN(n7861) );
  NAND2_X1 U9289 ( .A1(n9616), .A2(n7893), .ZN(n7650) );
  NAND2_X1 U9290 ( .A1(n9433), .A2(n7892), .ZN(n7649) );
  NAND2_X1 U9291 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  XNOR2_X1 U9292 ( .A(n7651), .B(n7890), .ZN(n7860) );
  NAND2_X1 U9293 ( .A1(n7655), .A2(n7652), .ZN(n7653) );
  INV_X1 U9294 ( .A(n7655), .ZN(n7657) );
  NAND2_X1 U9295 ( .A1(n7657), .A2(n7656), .ZN(n7658) );
  NAND2_X1 U9296 ( .A1(n9678), .A2(n7893), .ZN(n7660) );
  NAND2_X1 U9297 ( .A1(n9575), .A2(n7900), .ZN(n7659) );
  NAND2_X1 U9298 ( .A1(n7660), .A2(n7659), .ZN(n7661) );
  XNOR2_X1 U9299 ( .A(n7661), .B(n7763), .ZN(n8826) );
  NOR2_X1 U9300 ( .A1(n7662), .A2(n7898), .ZN(n7663) );
  AOI21_X1 U9301 ( .B1(n9678), .B2(n7892), .A(n7663), .ZN(n8830) );
  NOR2_X1 U9302 ( .A1(n8834), .A2(n7898), .ZN(n7664) );
  AOI21_X1 U9303 ( .B1(n9682), .B2(n7892), .A(n7664), .ZN(n7687) );
  AOI21_X1 U9304 ( .B1(n8826), .B2(n8830), .A(n8946), .ZN(n7665) );
  NAND2_X1 U9305 ( .A1(n7666), .A2(n7087), .ZN(n7668) );
  AOI22_X1 U9306 ( .A1(n7734), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9340), .B2(
        n4438), .ZN(n7667) );
  INV_X1 U9307 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7674) );
  INV_X1 U9308 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U9309 ( .A1(n7670), .A2(n7669), .ZN(n7671) );
  NAND2_X1 U9310 ( .A1(n7703), .A2(n7671), .ZN(n9556) );
  OR2_X1 U9311 ( .A1(n9556), .A2(n7868), .ZN(n7673) );
  AOI22_X1 U9312 ( .A1(n6743), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n6879), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n7672) );
  OAI211_X1 U9313 ( .C1(n7990), .C2(n7674), .A(n7673), .B(n7672), .ZN(n9573)
         );
  OAI22_X1 U9314 ( .A1(n9559), .A2(n6524), .B1(n8987), .B2(n7875), .ZN(n7675)
         );
  XNOR2_X1 U9315 ( .A(n7675), .B(n7890), .ZN(n8893) );
  OAI22_X1 U9316 ( .A1(n9559), .A2(n7875), .B1(n8987), .B2(n7898), .ZN(n8892)
         );
  NAND2_X1 U9317 ( .A1(n7676), .A2(n7087), .ZN(n7681) );
  OAI22_X1 U9318 ( .A1(n9323), .A2(n7678), .B1(n4635), .B2(n7677), .ZN(n7679)
         );
  INV_X1 U9319 ( .A(n7679), .ZN(n7680) );
  NAND2_X1 U9320 ( .A1(n9672), .A2(n7893), .ZN(n7683) );
  INV_X1 U9321 ( .A(n7952), .ZN(n9552) );
  NAND2_X1 U9322 ( .A1(n9552), .A2(n7900), .ZN(n7682) );
  NAND2_X1 U9323 ( .A1(n7683), .A2(n7682), .ZN(n7684) );
  XNOR2_X1 U9324 ( .A(n7684), .B(n7763), .ZN(n8888) );
  NOR2_X1 U9325 ( .A1(n7952), .A2(n7898), .ZN(n7685) );
  AOI21_X1 U9326 ( .B1(n9672), .B2(n7892), .A(n7685), .ZN(n8982) );
  INV_X1 U9327 ( .A(n7686), .ZN(n7689) );
  INV_X1 U9328 ( .A(n7687), .ZN(n7688) );
  NAND2_X1 U9329 ( .A1(n7689), .A2(n7688), .ZN(n8824) );
  NAND2_X1 U9330 ( .A1(n8824), .A2(n8830), .ZN(n7692) );
  INV_X1 U9331 ( .A(n8826), .ZN(n7691) );
  INV_X1 U9332 ( .A(n8830), .ZN(n8828) );
  AND2_X1 U9333 ( .A1(n8828), .A2(n7688), .ZN(n7690) );
  INV_X1 U9334 ( .A(n8893), .ZN(n7697) );
  NAND2_X1 U9335 ( .A1(n8888), .A2(n8982), .ZN(n7694) );
  NAND2_X1 U9336 ( .A1(n8892), .A2(n7694), .ZN(n7696) );
  INV_X1 U9337 ( .A(n8982), .ZN(n8891) );
  NOR2_X1 U9338 ( .A1(n8892), .A2(n8891), .ZN(n7695) );
  NAND2_X1 U9339 ( .A1(n7699), .A2(n7087), .ZN(n7701) );
  AOI22_X1 U9340 ( .A1(n7734), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4438), .B2(
        n9355), .ZN(n7700) );
  NAND2_X1 U9341 ( .A1(n9663), .A2(n7893), .ZN(n7709) );
  NAND2_X1 U9342 ( .A1(n7703), .A2(n7702), .ZN(n7704) );
  AND2_X1 U9343 ( .A1(n7720), .A2(n7704), .ZN(n9543) );
  NAND2_X1 U9344 ( .A1(n9543), .A2(n4264), .ZN(n7707) );
  AOI22_X1 U9345 ( .A1(n6532), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n6743), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n7706) );
  NAND2_X1 U9346 ( .A1(n7986), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7705) );
  OR2_X1 U9347 ( .A1(n8896), .A2(n7875), .ZN(n7708) );
  NAND2_X1 U9348 ( .A1(n7709), .A2(n7708), .ZN(n7710) );
  XNOR2_X1 U9349 ( .A(n7710), .B(n7890), .ZN(n7712) );
  NOR2_X1 U9350 ( .A1(n8896), .A2(n7898), .ZN(n7711) );
  AOI21_X1 U9351 ( .B1(n9663), .B2(n7892), .A(n7711), .ZN(n7713) );
  XNOR2_X1 U9352 ( .A(n7712), .B(n7713), .ZN(n8902) );
  INV_X1 U9353 ( .A(n7712), .ZN(n7714) );
  NAND2_X1 U9354 ( .A1(n7930), .A2(n7087), .ZN(n7928) );
  INV_X1 U9355 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U9356 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  NAND2_X1 U9357 ( .A1(n7717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7718) );
  XNOR2_X1 U9358 ( .A(n7718), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9367) );
  AOI22_X1 U9359 ( .A1(n7734), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4438), .B2(
        n9367), .ZN(n7931) );
  NAND2_X1 U9360 ( .A1(n7928), .A2(n7931), .ZN(n9656) );
  NAND2_X1 U9361 ( .A1(n9656), .A2(n7893), .ZN(n7728) );
  INV_X1 U9362 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7719) );
  NAND2_X1 U9363 ( .A1(n7720), .A2(n7719), .ZN(n7721) );
  NAND2_X1 U9364 ( .A1(n7753), .A2(n7721), .ZN(n9531) );
  OR2_X1 U9365 ( .A1(n9531), .A2(n7868), .ZN(n7726) );
  INV_X1 U9366 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U9367 ( .A1(n6743), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U9368 ( .A1(n7986), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7722) );
  OAI211_X1 U9369 ( .C1(n10095), .C2(n7990), .A(n7723), .B(n7722), .ZN(n7724)
         );
  INV_X1 U9370 ( .A(n7724), .ZN(n7725) );
  NAND2_X1 U9371 ( .A1(n7932), .A2(n7900), .ZN(n7727) );
  NAND2_X1 U9372 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  XNOR2_X1 U9373 ( .A(n7729), .B(n7763), .ZN(n7732) );
  NAND2_X1 U9374 ( .A1(n9656), .A2(n7900), .ZN(n7731) );
  NAND2_X1 U9375 ( .A1(n7731), .A2(n7730), .ZN(n7911) );
  NAND2_X1 U9376 ( .A1(n7733), .A2(n7087), .ZN(n7736) );
  AOI22_X1 U9377 ( .A1(n7734), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4438), .B2(
        n4259), .ZN(n7735) );
  NAND2_X1 U9378 ( .A1(n9651), .A2(n7900), .ZN(n7744) );
  XNOR2_X1 U9379 ( .A(n7753), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U9380 ( .A1(n9515), .A2(n4264), .ZN(n7742) );
  INV_X1 U9381 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U9382 ( .A1(n6743), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U9383 ( .A1(n7986), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7737) );
  OAI211_X1 U9384 ( .C1(n7739), .C2(n7990), .A(n7738), .B(n7737), .ZN(n7740)
         );
  INV_X1 U9385 ( .A(n7740), .ZN(n7741) );
  OR2_X1 U9386 ( .A1(n9498), .A2(n7898), .ZN(n7743) );
  NAND2_X1 U9387 ( .A1(n7744), .A2(n7743), .ZN(n7768) );
  INV_X1 U9388 ( .A(n7768), .ZN(n8860) );
  NAND2_X1 U9389 ( .A1(n9651), .A2(n7893), .ZN(n7746) );
  OR2_X1 U9390 ( .A1(n9498), .A2(n7875), .ZN(n7745) );
  NAND2_X1 U9391 ( .A1(n7746), .A2(n7745), .ZN(n7747) );
  XNOR2_X1 U9392 ( .A(n7747), .B(n7890), .ZN(n8864) );
  INV_X1 U9393 ( .A(n8864), .ZN(n8861) );
  NAND2_X1 U9394 ( .A1(n7748), .A2(n7087), .ZN(n7751) );
  OR2_X1 U9395 ( .A1(n4635), .A2(n7749), .ZN(n7750) );
  NAND2_X1 U9396 ( .A1(n9648), .A2(n4262), .ZN(n7762) );
  INV_X1 U9397 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8854) );
  INV_X1 U9398 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n7752) );
  OAI21_X1 U9399 ( .B1(n7753), .B2(n8854), .A(n7752), .ZN(n7754) );
  NAND2_X1 U9400 ( .A1(n7754), .A2(n7776), .ZN(n9503) );
  OR2_X1 U9401 ( .A1(n9503), .A2(n7868), .ZN(n7760) );
  INV_X1 U9402 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U9403 ( .A1(n6743), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U9404 ( .A1(n7986), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7755) );
  OAI211_X1 U9405 ( .C1(n7757), .C2(n7990), .A(n7756), .B(n7755), .ZN(n7758)
         );
  INV_X1 U9406 ( .A(n7758), .ZN(n7759) );
  NAND2_X1 U9407 ( .A1(n9511), .A2(n7900), .ZN(n7761) );
  NAND2_X1 U9408 ( .A1(n7762), .A2(n7761), .ZN(n7764) );
  XNOR2_X1 U9409 ( .A(n7764), .B(n7763), .ZN(n8870) );
  INV_X1 U9410 ( .A(n8870), .ZN(n7767) );
  NAND2_X1 U9411 ( .A1(n9648), .A2(n7900), .ZN(n7766) );
  NAND2_X1 U9412 ( .A1(n7766), .A2(n7765), .ZN(n8868) );
  NAND2_X1 U9413 ( .A1(n7767), .A2(n8868), .ZN(n8935) );
  OAI21_X1 U9414 ( .B1(n8860), .B2(n8861), .A(n8935), .ZN(n7772) );
  OAI21_X1 U9415 ( .B1(n8864), .B2(n7768), .A(n8868), .ZN(n7770) );
  NOR2_X1 U9416 ( .A1(n8868), .A2(n7768), .ZN(n7769) );
  AOI22_X1 U9417 ( .A1(n8870), .A2(n7770), .B1(n7769), .B2(n8861), .ZN(n7771)
         );
  NAND2_X1 U9418 ( .A1(n7773), .A2(n7087), .ZN(n7944) );
  OR2_X1 U9419 ( .A1(n4635), .A2(n7774), .ZN(n7941) );
  NAND2_X1 U9420 ( .A1(n9643), .A2(n7893), .ZN(n7785) );
  INV_X1 U9421 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U9422 ( .A1(n7776), .A2(n7775), .ZN(n7777) );
  NAND2_X1 U9423 ( .A1(n7794), .A2(n7777), .ZN(n9487) );
  OR2_X1 U9424 ( .A1(n9487), .A2(n7868), .ZN(n7783) );
  INV_X1 U9425 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U9426 ( .A1(n6879), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U9427 ( .A1(n6743), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7778) );
  OAI211_X1 U9428 ( .C1(n7990), .C2(n7780), .A(n7779), .B(n7778), .ZN(n7781)
         );
  INV_X1 U9429 ( .A(n7781), .ZN(n7782) );
  NAND2_X1 U9430 ( .A1(n7942), .A2(n7900), .ZN(n7784) );
  NAND2_X1 U9431 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  XNOR2_X1 U9432 ( .A(n7786), .B(n7890), .ZN(n7788) );
  NOR2_X1 U9433 ( .A1(n9500), .A2(n7898), .ZN(n7787) );
  AOI21_X1 U9434 ( .B1(n9643), .B2(n7892), .A(n7787), .ZN(n7789) );
  XNOR2_X1 U9435 ( .A(n7788), .B(n7789), .ZN(n8872) );
  INV_X1 U9436 ( .A(n7788), .ZN(n7790) );
  NAND2_X1 U9437 ( .A1(n7790), .A2(n7789), .ZN(n7791) );
  NAND2_X1 U9438 ( .A1(n7792), .A2(n7087), .ZN(n7948) );
  OR2_X1 U9439 ( .A1(n4635), .A2(n7793), .ZN(n7947) );
  OR2_X1 U9440 ( .A1(n9468), .A2(n7875), .ZN(n7803) );
  NAND2_X1 U9441 ( .A1(n7794), .A2(n8967), .ZN(n7795) );
  NAND2_X1 U9442 ( .A1(n7825), .A2(n7795), .ZN(n9465) );
  OR2_X1 U9443 ( .A1(n9465), .A2(n7868), .ZN(n7801) );
  INV_X1 U9444 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U9445 ( .A1(n7986), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U9446 ( .A1(n6743), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7796) );
  OAI211_X1 U9447 ( .C1(n7990), .C2(n7798), .A(n7797), .B(n7796), .ZN(n7799)
         );
  INV_X1 U9448 ( .A(n7799), .ZN(n7800) );
  NAND2_X1 U9449 ( .A1(n7801), .A2(n7800), .ZN(n9447) );
  AND2_X1 U9450 ( .A1(n7803), .A2(n7802), .ZN(n7805) );
  INV_X1 U9451 ( .A(n9447), .ZN(n9482) );
  OAI22_X1 U9452 ( .A1(n9468), .A2(n6524), .B1(n9482), .B2(n7875), .ZN(n7804)
         );
  XOR2_X1 U9453 ( .A(n7890), .B(n7804), .Z(n8960) );
  NAND2_X1 U9454 ( .A1(n7807), .A2(n7087), .ZN(n7810) );
  OR2_X1 U9455 ( .A1(n4635), .A2(n7808), .ZN(n7809) );
  INV_X1 U9456 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n7811) );
  NAND2_X1 U9457 ( .A1(n7827), .A2(n7811), .ZN(n7812) );
  NAND2_X1 U9458 ( .A1(n7846), .A2(n7812), .ZN(n8917) );
  OR2_X1 U9459 ( .A1(n8917), .A2(n7868), .ZN(n7818) );
  INV_X1 U9460 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U9461 ( .A1(n7986), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U9462 ( .A1(n6743), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7813) );
  OAI211_X1 U9463 ( .C1(n7990), .C2(n7815), .A(n7814), .B(n7813), .ZN(n7816)
         );
  INV_X1 U9464 ( .A(n7816), .ZN(n7817) );
  NAND2_X1 U9465 ( .A1(n9628), .A2(n7900), .ZN(n7820) );
  NAND2_X1 U9466 ( .A1(n7820), .A2(n7819), .ZN(n8913) );
  NAND2_X1 U9467 ( .A1(n7821), .A2(n7087), .ZN(n7824) );
  OR2_X1 U9468 ( .A1(n4635), .A2(n7822), .ZN(n7823) );
  NAND2_X1 U9469 ( .A1(n9631), .A2(n7900), .ZN(n7835) );
  NAND2_X1 U9470 ( .A1(n7825), .A2(n8846), .ZN(n7826) );
  AND2_X1 U9471 ( .A1(n7827), .A2(n7826), .ZN(n9453) );
  NAND2_X1 U9472 ( .A1(n9453), .A2(n4264), .ZN(n7833) );
  INV_X1 U9473 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U9474 ( .A1(n6743), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U9475 ( .A1(n7986), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7828) );
  OAI211_X1 U9476 ( .C1(n7990), .C2(n7830), .A(n7829), .B(n7828), .ZN(n7831)
         );
  INV_X1 U9477 ( .A(n7831), .ZN(n7832) );
  NAND2_X1 U9478 ( .A1(n7835), .A2(n7834), .ZN(n8912) );
  NAND2_X1 U9479 ( .A1(n9631), .A2(n4262), .ZN(n7837) );
  NAND2_X1 U9480 ( .A1(n9462), .A2(n7900), .ZN(n7836) );
  NAND2_X1 U9481 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  XNOR2_X1 U9482 ( .A(n7838), .B(n7890), .ZN(n7841) );
  AOI22_X1 U9483 ( .A1(n8914), .A2(n8913), .B1(n8912), .B2(n7841), .ZN(n7844)
         );
  INV_X1 U9484 ( .A(n7841), .ZN(n8841) );
  INV_X1 U9485 ( .A(n8912), .ZN(n8843) );
  INV_X1 U9486 ( .A(n8913), .ZN(n7839) );
  AOI21_X1 U9487 ( .B1(n8841), .B2(n8843), .A(n7839), .ZN(n7842) );
  NAND2_X1 U9488 ( .A1(n7839), .A2(n8843), .ZN(n7840) );
  OAI22_X1 U9489 ( .A1(n8914), .A2(n7842), .B1(n7841), .B2(n7840), .ZN(n7843)
         );
  OR2_X1 U9490 ( .A1(n4635), .A2(n7966), .ZN(n7973) );
  NAND2_X1 U9491 ( .A1(n9622), .A2(n4262), .ZN(n7855) );
  INV_X1 U9492 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U9493 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  NAND2_X1 U9494 ( .A1(n7848), .A2(n7847), .ZN(n8882) );
  INV_X1 U9495 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U9496 ( .A1(n6743), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U9497 ( .A1(n7986), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7849) );
  OAI211_X1 U9498 ( .C1(n10132), .C2(n7990), .A(n7850), .B(n7849), .ZN(n7851)
         );
  INV_X1 U9499 ( .A(n7851), .ZN(n7852) );
  NAND2_X1 U9500 ( .A1(n7972), .A2(n7900), .ZN(n7854) );
  NAND2_X1 U9501 ( .A1(n7855), .A2(n7854), .ZN(n7856) );
  XNOR2_X1 U9502 ( .A(n7856), .B(n7890), .ZN(n7858) );
  OAI22_X1 U9503 ( .A1(n9441), .A2(n7875), .B1(n8921), .B2(n7898), .ZN(n7857)
         );
  XNOR2_X1 U9504 ( .A(n7858), .B(n7857), .ZN(n8881) );
  XOR2_X1 U9505 ( .A(n7860), .B(n7859), .Z(n8976) );
  NAND2_X1 U9506 ( .A1(n8801), .A2(n7087), .ZN(n7864) );
  OR2_X1 U9507 ( .A1(n4635), .A2(n7862), .ZN(n7863) );
  INV_X1 U9508 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U9509 ( .A1(n7866), .A2(n7865), .ZN(n7867) );
  NAND2_X1 U9510 ( .A1(n7882), .A2(n7867), .ZN(n8817) );
  INV_X1 U9511 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U9512 ( .A1(n6743), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U9513 ( .A1(n7986), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7869) );
  OAI211_X1 U9514 ( .C1(n7990), .C2(n7871), .A(n7870), .B(n7869), .ZN(n7872)
         );
  INV_X1 U9515 ( .A(n7872), .ZN(n7873) );
  OAI22_X1 U9516 ( .A1(n9409), .A2(n6524), .B1(n9390), .B2(n7875), .ZN(n7876)
         );
  XOR2_X1 U9517 ( .A(n7890), .B(n7876), .Z(n8814) );
  INV_X1 U9518 ( .A(n8814), .ZN(n7877) );
  NAND2_X1 U9519 ( .A1(n7878), .A2(n7877), .ZN(n7908) );
  OR2_X1 U9520 ( .A1(n4635), .A2(n10133), .ZN(n7879) );
  NAND2_X1 U9521 ( .A1(n9606), .A2(n7900), .ZN(n7889) );
  NAND2_X1 U9522 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  INV_X1 U9523 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U9524 ( .A1(n6743), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U9525 ( .A1(n6879), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7884) );
  OAI211_X1 U9526 ( .C1(n7886), .C2(n7990), .A(n7885), .B(n7884), .ZN(n7887)
         );
  AOI21_X2 U9527 ( .B1(n9395), .B2(n4264), .A(n7887), .ZN(n9413) );
  OR2_X1 U9528 ( .A1(n9413), .A2(n7898), .ZN(n7888) );
  NAND2_X1 U9529 ( .A1(n7889), .A2(n7888), .ZN(n7891) );
  XNOR2_X1 U9530 ( .A(n7890), .B(n7891), .ZN(n7895) );
  INV_X1 U9531 ( .A(n9413), .ZN(n9273) );
  AOI22_X1 U9532 ( .A1(n9606), .A2(n7893), .B1(n7892), .B2(n9273), .ZN(n7894)
         );
  XNOR2_X1 U9533 ( .A(n7895), .B(n7894), .ZN(n7897) );
  INV_X1 U9534 ( .A(n7897), .ZN(n7896) );
  NAND2_X1 U9535 ( .A1(n7896), .A2(n8964), .ZN(n7907) );
  NOR2_X1 U9536 ( .A1(n9390), .A2(n7898), .ZN(n7899) );
  AOI21_X1 U9537 ( .B1(n9612), .B2(n7900), .A(n7899), .ZN(n8813) );
  AOI21_X1 U9538 ( .B1(n8816), .B2(n8814), .A(n8813), .ZN(n7901) );
  NAND2_X1 U9539 ( .A1(n9422), .A2(n8984), .ZN(n7903) );
  AOI22_X1 U9540 ( .A1(n9395), .A2(n8991), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7902) );
  OAI211_X1 U9541 ( .C1(n9391), .C2(n8986), .A(n7903), .B(n7902), .ZN(n7904)
         );
  AOI21_X1 U9542 ( .B1(n9606), .B2(n8978), .A(n7904), .ZN(n7905) );
  OAI211_X1 U9543 ( .C1(n7908), .C2(n7907), .A(n7906), .B(n7905), .ZN(P1_U3218) );
  AOI22_X1 U9544 ( .A1(n9367), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9740), .ZN(n7909) );
  OAI21_X1 U9545 ( .B1(n7910), .B2(n4261), .A(n7909), .ZN(P1_U3335) );
  INV_X1 U9546 ( .A(n7913), .ZN(n7917) );
  AOI21_X1 U9547 ( .B1(n7913), .B2(n7912), .A(n7911), .ZN(n7914) );
  NOR2_X1 U9548 ( .A1(n7914), .A2(n8993), .ZN(n7915) );
  OAI21_X1 U9549 ( .B1(n7917), .B2(n7916), .A(n7915), .ZN(n7921) );
  NAND2_X1 U9550 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9358) );
  OAI21_X1 U9551 ( .B1(n8896), .B2(n8968), .A(n9358), .ZN(n7919) );
  NOR2_X1 U9552 ( .A1(n8966), .A2(n9531), .ZN(n7918) );
  AOI211_X1 U9553 ( .C1(n8971), .C2(n9524), .A(n7919), .B(n7918), .ZN(n7920)
         );
  OAI211_X1 U9554 ( .C1(n9528), .C2(n8988), .A(n7921), .B(n7920), .ZN(P1_U3236) );
  NAND2_X1 U9555 ( .A1(n9672), .A2(n9552), .ZN(n7923) );
  NAND2_X1 U9556 ( .A1(n9559), .A2(n9573), .ZN(n9130) );
  NAND2_X1 U9557 ( .A1(n9130), .A2(n7953), .ZN(n9561) );
  NAND2_X1 U9558 ( .A1(n9668), .A2(n9573), .ZN(n7924) );
  INV_X1 U9559 ( .A(n8896), .ZN(n9553) );
  OR2_X1 U9560 ( .A1(n9663), .A2(n9553), .ZN(n7926) );
  INV_X1 U9561 ( .A(n8905), .ZN(n7932) );
  AND2_X1 U9562 ( .A1(n7931), .A2(n7932), .ZN(n7927) );
  NAND2_X1 U9563 ( .A1(n7928), .A2(n7927), .ZN(n9134) );
  AND2_X1 U9564 ( .A1(n7087), .A2(n8905), .ZN(n7929) );
  NAND2_X1 U9565 ( .A1(n7930), .A2(n7929), .ZN(n7934) );
  OR2_X1 U9566 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  AND2_X2 U9567 ( .A1(n7934), .A2(n7933), .ZN(n9030) );
  AND2_X2 U9568 ( .A1(n9134), .A2(n9030), .ZN(n9535) );
  NAND2_X1 U9569 ( .A1(n9656), .A2(n7932), .ZN(n7936) );
  OR2_X1 U9570 ( .A1(n9651), .A2(n9524), .ZN(n7937) );
  NAND2_X1 U9571 ( .A1(n9519), .A2(n7937), .ZN(n7939) );
  NAND2_X1 U9572 ( .A1(n9651), .A2(n9524), .ZN(n7938) );
  OR2_X1 U9573 ( .A1(n9648), .A2(n9511), .ZN(n7940) );
  INV_X1 U9574 ( .A(n9500), .ZN(n7942) );
  AND2_X1 U9575 ( .A1(n7942), .A2(n7941), .ZN(n7943) );
  NAND2_X1 U9576 ( .A1(n7944), .A2(n7943), .ZN(n9148) );
  NAND2_X1 U9577 ( .A1(n9643), .A2(n9500), .ZN(n9144) );
  NAND2_X1 U9578 ( .A1(n9148), .A2(n9144), .ZN(n9475) );
  NAND2_X1 U9579 ( .A1(n9643), .A2(n7942), .ZN(n7945) );
  OR2_X1 U9580 ( .A1(n9636), .A2(n9447), .ZN(n7949) );
  INV_X1 U9581 ( .A(n7970), .ZN(n7950) );
  XOR2_X1 U9582 ( .A(n7967), .B(n9216), .Z(n9630) );
  INV_X1 U9583 ( .A(n9021), .ZN(n9107) );
  OR2_X1 U9584 ( .A1(n9672), .A2(n7952), .ZN(n9123) );
  NAND2_X1 U9585 ( .A1(n9672), .A2(n7952), .ZN(n9122) );
  INV_X1 U9586 ( .A(n7953), .ZN(n9129) );
  NOR2_X1 U9587 ( .A1(n9663), .A2(n8896), .ZN(n9128) );
  NAND2_X1 U9588 ( .A1(n9663), .A2(n8896), .ZN(n9126) );
  INV_X1 U9589 ( .A(n9030), .ZN(n7954) );
  OR2_X1 U9590 ( .A1(n9651), .A2(n9498), .ZN(n9133) );
  NAND2_X1 U9591 ( .A1(n9651), .A2(n9498), .ZN(n9135) );
  NAND2_X1 U9592 ( .A1(n9133), .A2(n9135), .ZN(n9518) );
  NAND2_X1 U9593 ( .A1(n9648), .A2(n9483), .ZN(n9184) );
  INV_X1 U9594 ( .A(n9144), .ZN(n7955) );
  NAND2_X1 U9595 ( .A1(n9636), .A2(n9482), .ZN(n9155) );
  NAND2_X1 U9596 ( .A1(n9631), .A2(n7957), .ZN(n9156) );
  XOR2_X1 U9597 ( .A(n9216), .B(n7982), .Z(n7956) );
  OAI222_X1 U9598 ( .A1(n9501), .A2(n8921), .B1(n9499), .B2(n7957), .C1(n9496), 
        .C2(n7956), .ZN(n9626) );
  INV_X1 U9599 ( .A(n9631), .ZN(n9455) );
  INV_X1 U9600 ( .A(n9672), .ZN(n9587) );
  NAND2_X1 U9601 ( .A1(n9578), .A2(n9587), .ZN(n9579) );
  INV_X1 U9602 ( .A(n9651), .ZN(n9517) );
  INV_X1 U9603 ( .A(n9643), .ZN(n8879) );
  NAND2_X1 U9604 ( .A1(n9455), .A2(n9464), .ZN(n9450) );
  AOI211_X1 U9605 ( .C1(n9628), .C2(n9450), .A(n9869), .B(n9435), .ZN(n9627)
         );
  INV_X1 U9606 ( .A(n9627), .ZN(n7958) );
  OAI22_X1 U9607 ( .A1(n7958), .A2(n4259), .B1(n8917), .B2(n9530), .ZN(n7959)
         );
  OAI21_X1 U9608 ( .B1(n9626), .B2(n7959), .A(n9589), .ZN(n7961) );
  AOI22_X1 U9609 ( .A1(n9628), .A2(n9490), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9566), .ZN(n7960) );
  OAI211_X1 U9610 ( .C1(n9630), .C2(n9592), .A(n7961), .B(n7960), .ZN(P1_U3267) );
  OAI222_X1 U9611 ( .A1(n8811), .A2(n7964), .B1(n8799), .B2(n7963), .C1(n7962), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9612 ( .A(n7965), .ZN(n8809) );
  OAI222_X1 U9613 ( .A1(n9743), .A2(n7966), .B1(n4261), .B2(n8809), .C1(
        P1_U3084), .C2(n6150), .ZN(P1_U3328) );
  INV_X1 U9614 ( .A(n7968), .ZN(n7969) );
  INV_X1 U9615 ( .A(n8921), .ZN(n7972) );
  AND2_X1 U9616 ( .A1(n7973), .A2(n7972), .ZN(n7974) );
  NAND2_X1 U9617 ( .A1(n7975), .A2(n7974), .ZN(n9419) );
  NAND2_X1 U9618 ( .A1(n9622), .A2(n8921), .ZN(n9160) );
  NAND2_X1 U9619 ( .A1(n9419), .A2(n9160), .ZN(n9431) );
  OR2_X1 U9620 ( .A1(n9622), .A2(n7972), .ZN(n7976) );
  NAND2_X1 U9621 ( .A1(n9612), .A2(n9390), .ZN(n9163) );
  NAND2_X1 U9622 ( .A1(n9606), .A2(n9273), .ZN(n7978) );
  NAND2_X1 U9623 ( .A1(n8793), .A2(n7087), .ZN(n7980) );
  OR2_X1 U9624 ( .A1(n4635), .A2(n9734), .ZN(n7979) );
  NAND2_X1 U9625 ( .A1(n7998), .A2(n9391), .ZN(n9253) );
  NAND2_X1 U9626 ( .A1(n9420), .A2(n9040), .ZN(n7983) );
  NAND2_X1 U9627 ( .A1(n9616), .A2(n9412), .ZN(n9162) );
  XNOR2_X1 U9628 ( .A(n7984), .B(n9061), .ZN(n7992) );
  AND2_X1 U9629 ( .A1(n9778), .A2(P1_B_REG_SCAN_IN), .ZN(n7985) );
  NOR2_X1 U9630 ( .A1(n9501), .A2(n7985), .ZN(n9377) );
  INV_X1 U9631 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U9632 ( .A1(n6743), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U9633 ( .A1(n7986), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7987) );
  OAI211_X1 U9634 ( .C1(n7990), .C2(n7989), .A(n7988), .B(n7987), .ZN(n9272)
         );
  AOI22_X1 U9635 ( .A1(n9273), .A2(n9574), .B1(n9377), .B2(n9272), .ZN(n7991)
         );
  OAI21_X1 U9636 ( .B1(n7992), .B2(n9496), .A(n7991), .ZN(n9600) );
  NAND2_X1 U9637 ( .A1(n9600), .A2(n9589), .ZN(n8000) );
  INV_X1 U9638 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7993) );
  OAI22_X1 U9639 ( .A1(n7994), .A2(n9530), .B1(n7993), .B2(n9589), .ZN(n7997)
         );
  XNOR2_X1 U9640 ( .A(n9394), .B(n9603), .ZN(n9604) );
  NOR2_X1 U9641 ( .A1(n9604), .A2(n7995), .ZN(n7996) );
  AOI211_X1 U9642 ( .C1(n9490), .C2(n7998), .A(n7997), .B(n7996), .ZN(n7999)
         );
  OAI211_X1 U9643 ( .C1(n9602), .C2(n9592), .A(n8000), .B(n7999), .ZN(P1_U3355) );
  INV_X1 U9644 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U9645 ( .A1(n8652), .A2(n8619), .ZN(n8614) );
  INV_X1 U9646 ( .A(n8614), .ZN(n8005) );
  NOR2_X1 U9647 ( .A1(n8635), .A2(n8005), .ZN(n8006) );
  INV_X1 U9648 ( .A(n8746), .ZN(n8618) );
  AOI22_X1 U9649 ( .A1(n8623), .A2(n8006), .B1(n8618), .B2(n8639), .ZN(n8007)
         );
  OR2_X1 U9650 ( .A1(n8608), .A2(n8626), .ZN(n8008) );
  NAND2_X1 U9651 ( .A1(n8735), .A2(n8597), .ZN(n8559) );
  NAND2_X1 U9652 ( .A1(n8575), .A2(n8559), .ZN(n8009) );
  OAI22_X1 U9653 ( .A1(n8010), .A2(n8009), .B1(n8731), .B2(n8579), .ZN(n8011)
         );
  INV_X1 U9654 ( .A(n8011), .ZN(n8012) );
  NAND2_X1 U9655 ( .A1(n8725), .A2(n8563), .ZN(n8013) );
  NOR2_X1 U9656 ( .A1(n8721), .A2(n8547), .ZN(n8015) );
  NAND2_X1 U9657 ( .A1(n8721), .A2(n8547), .ZN(n8014) );
  NOR2_X1 U9658 ( .A1(n8703), .A2(n8505), .ZN(n8016) );
  NAND2_X1 U9659 ( .A1(n8696), .A2(n8492), .ZN(n8017) );
  NOR2_X1 U9660 ( .A1(n8691), .A2(n8474), .ZN(n8448) );
  NOR2_X1 U9661 ( .A1(n8688), .A2(n8459), .ZN(n8020) );
  AOI21_X1 U9662 ( .B1(n8021), .B2(n8448), .A(n8020), .ZN(n8420) );
  OR2_X1 U9663 ( .A1(n8680), .A2(n8206), .ZN(n8022) );
  INV_X1 U9664 ( .A(n8022), .ZN(n8023) );
  OR2_X1 U9665 ( .A1(n8675), .A2(n8398), .ZN(n8024) );
  NAND2_X1 U9666 ( .A1(n8025), .A2(n8024), .ZN(n8390) );
  NOR2_X1 U9667 ( .A1(n8670), .A2(n8205), .ZN(n8026) );
  NAND2_X1 U9668 ( .A1(n8366), .A2(P2_B_REG_SCAN_IN), .ZN(n8029) );
  NAND2_X1 U9669 ( .A1(n8596), .A2(n8029), .ZN(n8378) );
  NOR2_X1 U9670 ( .A1(n8378), .A2(n8030), .ZN(n8031) );
  AOI21_X1 U9671 ( .B1(n8205), .B2(n9910), .A(n8031), .ZN(n8032) );
  NAND2_X1 U9672 ( .A1(n8033), .A2(n8032), .ZN(n8665) );
  NAND2_X1 U9673 ( .A1(n8665), .A2(n8606), .ZN(n8042) );
  INV_X1 U9674 ( .A(n8666), .ZN(n8039) );
  INV_X1 U9675 ( .A(n8675), .ZN(n8409) );
  INV_X1 U9676 ( .A(n8721), .ZN(n8081) );
  INV_X1 U9677 ( .A(n8608), .ZN(n8740) );
  NOR2_X2 U9678 ( .A1(n8584), .A2(n8731), .ZN(n8567) );
  AND2_X2 U9679 ( .A1(n8567), .A2(n5013), .ZN(n8549) );
  INV_X1 U9680 ( .A(n8703), .ZN(n8500) );
  OR2_X2 U9681 ( .A1(n8496), .A2(n8696), .ZN(n8477) );
  INV_X1 U9682 ( .A(n8688), .ZN(n8452) );
  NOR2_X2 U9683 ( .A1(n8404), .A2(n8670), .ZN(n8391) );
  NAND2_X1 U9684 ( .A1(n8039), .A2(n8391), .ZN(n8382) );
  INV_X1 U9685 ( .A(n8391), .ZN(n8035) );
  NAND2_X1 U9686 ( .A1(n8666), .A2(n8035), .ZN(n8036) );
  AND2_X1 U9687 ( .A1(n8382), .A2(n8036), .ZN(n8667) );
  AOI22_X1 U9688 ( .A1(n8037), .A2(n8649), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8651), .ZN(n8038) );
  OAI21_X1 U9689 ( .B1(n8039), .B2(n9925), .A(n8038), .ZN(n8040) );
  AOI21_X1 U9690 ( .B1(n8667), .B2(n8629), .A(n8040), .ZN(n8041) );
  OAI211_X1 U9691 ( .C1(n8669), .C2(n9924), .A(n8042), .B(n8041), .ZN(P2_U3267) );
  OAI22_X1 U9692 ( .A1(n8406), .A2(n8195), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8044), .ZN(n8046) );
  OAI22_X1 U9693 ( .A1(n8413), .A2(n8166), .B1(n8412), .B2(n8167), .ZN(n8045)
         );
  AOI211_X1 U9694 ( .C1(n8675), .C2(n8197), .A(n8046), .B(n8045), .ZN(n8047)
         );
  OAI21_X1 U9695 ( .B1(n8048), .B2(n8202), .A(n8047), .ZN(P2_U3216) );
  OAI21_X1 U9696 ( .B1(n8051), .B2(n8050), .A(n8049), .ZN(n8056) );
  AOI21_X1 U9697 ( .B1(n8186), .B2(n8616), .A(n8052), .ZN(n8054) );
  AOI22_X1 U9698 ( .A1(n8192), .A2(n8619), .B1(n8191), .B2(n8626), .ZN(n8053)
         );
  OAI211_X1 U9699 ( .C1(n8618), .C2(n8115), .A(n8054), .B(n8053), .ZN(n8055)
         );
  AOI21_X1 U9700 ( .B1(n8056), .B2(n8162), .A(n8055), .ZN(n8057) );
  INV_X1 U9701 ( .A(n8057), .ZN(P2_U3217) );
  INV_X1 U9702 ( .A(n8058), .ZN(n8125) );
  XNOR2_X1 U9703 ( .A(n8126), .B(n8125), .ZN(n8065) );
  INV_X1 U9704 ( .A(n8478), .ZN(n8060) );
  OAI22_X1 U9705 ( .A1(n8195), .A2(n8060), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8059), .ZN(n8063) );
  OAI22_X1 U9706 ( .A1(n8061), .A2(n8166), .B1(n8167), .B2(n8086), .ZN(n8062)
         );
  AOI211_X1 U9707 ( .C1(n8696), .C2(n8197), .A(n8063), .B(n8062), .ZN(n8064)
         );
  OAI21_X1 U9708 ( .B1(n8065), .B2(n8202), .A(n8064), .ZN(P2_U3218) );
  MUX2_X1 U9709 ( .A(n8195), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n8071) );
  XOR2_X1 U9710 ( .A(n8067), .B(n8066), .Z(n8068) );
  AOI22_X1 U9711 ( .A1(n8197), .A2(n9955), .B1(n8162), .B2(n8068), .ZN(n8070)
         );
  AOI22_X1 U9712 ( .A1(n8192), .A2(n8216), .B1(n8191), .B2(n8215), .ZN(n8069)
         );
  NAND3_X1 U9713 ( .A1(n8071), .A2(n8070), .A3(n8069), .ZN(P2_U3220) );
  OAI21_X1 U9714 ( .B1(n8074), .B2(n8073), .A(n8072), .ZN(n8075) );
  NAND2_X1 U9715 ( .A1(n8075), .A2(n8162), .ZN(n8080) );
  INV_X1 U9716 ( .A(n8076), .ZN(n8540) );
  NAND2_X1 U9717 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8374) );
  INV_X1 U9718 ( .A(n8374), .ZN(n8078) );
  OAI22_X1 U9719 ( .A1(n8085), .A2(n8166), .B1(n8167), .B2(n8118), .ZN(n8077)
         );
  AOI211_X1 U9720 ( .C1(n8186), .C2(n8540), .A(n8078), .B(n8077), .ZN(n8079)
         );
  OAI211_X1 U9721 ( .C1(n8081), .C2(n8115), .A(n8080), .B(n8079), .ZN(P2_U3221) );
  XNOR2_X1 U9722 ( .A(n8082), .B(n8083), .ZN(n8090) );
  INV_X1 U9723 ( .A(n8507), .ZN(n8084) );
  OAI22_X1 U9724 ( .A1(n8195), .A2(n8084), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10083), .ZN(n8088) );
  OAI22_X1 U9725 ( .A1(n8086), .A2(n8166), .B1(n8167), .B2(n8085), .ZN(n8087)
         );
  AOI211_X1 U9726 ( .C1(n8709), .C2(n8197), .A(n8088), .B(n8087), .ZN(n8089)
         );
  OAI21_X1 U9727 ( .B1(n8090), .B2(n8202), .A(n8089), .ZN(P2_U3225) );
  XNOR2_X1 U9728 ( .A(n8092), .B(n8091), .ZN(n8098) );
  AND2_X1 U9729 ( .A1(n8474), .A2(n9910), .ZN(n8093) );
  AOI21_X1 U9730 ( .B1(n8206), .B2(n8596), .A(n8093), .ZN(n8446) );
  INV_X1 U9731 ( .A(n8143), .ZN(n8184) );
  OAI22_X1 U9732 ( .A1(n8446), .A2(n8184), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8094), .ZN(n8096) );
  NOR2_X1 U9733 ( .A1(n8452), .A2(n8115), .ZN(n8095) );
  AOI211_X1 U9734 ( .C1(n8186), .C2(n8450), .A(n8096), .B(n8095), .ZN(n8097)
         );
  OAI21_X1 U9735 ( .B1(n8098), .B2(n8202), .A(n8097), .ZN(P2_U3227) );
  NAND2_X1 U9736 ( .A1(n8101), .A2(n8100), .ZN(n8103) );
  OAI21_X1 U9737 ( .B1(n8101), .B2(n8100), .A(n8103), .ZN(n8199) );
  NOR2_X1 U9738 ( .A1(n8199), .A2(n8102), .ZN(n8190) );
  INV_X1 U9739 ( .A(n8103), .ZN(n8105) );
  NOR3_X1 U9740 ( .A1(n8190), .A2(n8105), .A3(n8104), .ZN(n8108) );
  INV_X1 U9741 ( .A(n8106), .ZN(n8107) );
  OAI21_X1 U9742 ( .B1(n8108), .B2(n8107), .A(n8162), .ZN(n8114) );
  INV_X1 U9743 ( .A(n8109), .ZN(n8586) );
  AND2_X1 U9744 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8328) );
  OAI22_X1 U9745 ( .A1(n8111), .A2(n8166), .B1(n8167), .B2(n8110), .ZN(n8112)
         );
  AOI211_X1 U9746 ( .C1(n8186), .C2(n8586), .A(n8328), .B(n8112), .ZN(n8113)
         );
  OAI211_X1 U9747 ( .C1(n4985), .C2(n8115), .A(n8114), .B(n8113), .ZN(P2_U3228) );
  XNOR2_X1 U9748 ( .A(n8117), .B(n8116), .ZN(n8123) );
  OAI22_X1 U9749 ( .A1(n8195), .A2(n8569), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10193), .ZN(n8121) );
  OAI22_X1 U9750 ( .A1(n8119), .A2(n8167), .B1(n8166), .B2(n8118), .ZN(n8120)
         );
  AOI211_X1 U9751 ( .C1(n8731), .C2(n8197), .A(n8121), .B(n8120), .ZN(n8122)
         );
  OAI21_X1 U9752 ( .B1(n8123), .B2(n8202), .A(n8122), .ZN(P2_U3230) );
  AOI21_X1 U9753 ( .B1(n8126), .B2(n8125), .A(n8124), .ZN(n8130) );
  XNOR2_X1 U9754 ( .A(n8128), .B(n8127), .ZN(n8129) );
  XNOR2_X1 U9755 ( .A(n8130), .B(n8129), .ZN(n8136) );
  OAI22_X1 U9756 ( .A1(n8195), .A2(n8465), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8131), .ZN(n8134) );
  OAI22_X1 U9757 ( .A1(n8132), .A2(n8166), .B1(n8165), .B2(n8167), .ZN(n8133)
         );
  AOI211_X1 U9758 ( .C1(n8691), .C2(n8197), .A(n8134), .B(n8133), .ZN(n8135)
         );
  OAI21_X1 U9759 ( .B1(n8136), .B2(n8202), .A(n8135), .ZN(P2_U3231) );
  AOI22_X1 U9760 ( .A1(n8197), .A2(n9898), .B1(n8186), .B2(n9900), .ZN(n8147)
         );
  OAI21_X1 U9761 ( .B1(n8139), .B2(n8138), .A(n8137), .ZN(n8140) );
  NAND2_X1 U9762 ( .A1(n8162), .A2(n8140), .ZN(n8145) );
  NAND2_X1 U9763 ( .A1(n8596), .A2(n8214), .ZN(n8142) );
  NAND2_X1 U9764 ( .A1(n9910), .A2(n9909), .ZN(n8141) );
  NAND2_X1 U9765 ( .A1(n8142), .A2(n8141), .ZN(n9894) );
  NAND2_X1 U9766 ( .A1(n8143), .A2(n9894), .ZN(n8144) );
  NAND4_X1 U9767 ( .A1(n8147), .A2(n8146), .A3(n8145), .A4(n8144), .ZN(
        P2_U3232) );
  XNOR2_X1 U9768 ( .A(n8149), .B(n8148), .ZN(n8155) );
  OAI22_X1 U9769 ( .A1(n8195), .A2(n8525), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8150), .ZN(n8153) );
  OAI22_X1 U9770 ( .A1(n8168), .A2(n8166), .B1(n8167), .B2(n8151), .ZN(n8152)
         );
  AOI211_X1 U9771 ( .C1(n8714), .C2(n8197), .A(n8153), .B(n8152), .ZN(n8154)
         );
  OAI21_X1 U9772 ( .B1(n8155), .B2(n8202), .A(n8154), .ZN(P2_U3235) );
  NAND2_X1 U9773 ( .A1(n8157), .A2(n8156), .ZN(n8159) );
  XNOR2_X1 U9774 ( .A(n8159), .B(n8158), .ZN(n8160) );
  NAND3_X1 U9775 ( .A1(n8160), .A2(n8198), .A3(n8505), .ZN(n8173) );
  INV_X1 U9776 ( .A(n8160), .ZN(n8163) );
  NAND3_X1 U9777 ( .A1(n8163), .A2(n8162), .A3(n8161), .ZN(n8172) );
  OAI22_X1 U9778 ( .A1(n8195), .A2(n8497), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8164), .ZN(n8170) );
  OAI22_X1 U9779 ( .A1(n8168), .A2(n8167), .B1(n8166), .B2(n8165), .ZN(n8169)
         );
  AOI211_X1 U9780 ( .C1(n8703), .C2(n8197), .A(n8170), .B(n8169), .ZN(n8171)
         );
  NAND3_X1 U9781 ( .A1(n8173), .A2(n8172), .A3(n8171), .ZN(P2_U3237) );
  XNOR2_X1 U9782 ( .A(n8175), .B(n8174), .ZN(n8179) );
  AOI22_X1 U9783 ( .A1(n8191), .A2(n8547), .B1(n8192), .B2(n8579), .ZN(n8176)
         );
  NAND2_X1 U9784 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8351) );
  OAI211_X1 U9785 ( .C1(n8195), .C2(n8551), .A(n8176), .B(n8351), .ZN(n8177)
         );
  AOI21_X1 U9786 ( .B1(n8725), .B2(n8197), .A(n8177), .ZN(n8178) );
  OAI21_X1 U9787 ( .B1(n8179), .B2(n8202), .A(n8178), .ZN(P2_U3240) );
  XNOR2_X1 U9788 ( .A(n8180), .B(n8181), .ZN(n8189) );
  AND2_X1 U9789 ( .A1(n8459), .A2(n9910), .ZN(n8182) );
  AOI21_X1 U9790 ( .B1(n8398), .B2(n8596), .A(n8182), .ZN(n8429) );
  OAI22_X1 U9791 ( .A1(n8429), .A2(n8184), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8183), .ZN(n8185) );
  AOI21_X1 U9792 ( .B1(n8433), .B2(n8186), .A(n8185), .ZN(n8188) );
  NAND2_X1 U9793 ( .A1(n8680), .A2(n8197), .ZN(n8187) );
  OAI211_X1 U9794 ( .C1(n8189), .C2(n8202), .A(n8188), .B(n8187), .ZN(P2_U3242) );
  INV_X1 U9795 ( .A(n8190), .ZN(n8203) );
  AOI22_X1 U9796 ( .A1(n8192), .A2(n8595), .B1(n8191), .B2(n8597), .ZN(n8194)
         );
  OAI211_X1 U9797 ( .C1(n8195), .C2(n8604), .A(n8194), .B(n8193), .ZN(n8196)
         );
  AOI21_X1 U9798 ( .B1(n8608), .B2(n8197), .A(n8196), .ZN(n8201) );
  NAND3_X1 U9799 ( .A1(n8199), .A2(n8198), .A3(n8626), .ZN(n8200) );
  OAI211_X1 U9800 ( .C1(n8203), .C2(n8202), .A(n8201), .B(n8200), .ZN(P2_U3243) );
  MUX2_X1 U9801 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8204), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9802 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8399), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9803 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8205), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9804 ( .A(n8398), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8217), .Z(
        P2_U3579) );
  MUX2_X1 U9805 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8206), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9806 ( .A(n8459), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8217), .Z(
        P2_U3577) );
  MUX2_X1 U9807 ( .A(n8474), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8217), .Z(
        P2_U3576) );
  MUX2_X1 U9808 ( .A(n8492), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8217), .Z(
        P2_U3575) );
  MUX2_X1 U9809 ( .A(n8505), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8217), .Z(
        P2_U3574) );
  MUX2_X1 U9810 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8520), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9811 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8535), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9812 ( .A(n8547), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8217), .Z(
        P2_U3571) );
  MUX2_X1 U9813 ( .A(n8563), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8217), .Z(
        P2_U3570) );
  MUX2_X1 U9814 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8579), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9815 ( .A(n8597), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8217), .Z(
        P2_U3568) );
  MUX2_X1 U9816 ( .A(n8626), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8217), .Z(
        P2_U3567) );
  MUX2_X1 U9817 ( .A(n8595), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8217), .Z(
        P2_U3566) );
  MUX2_X1 U9818 ( .A(n8619), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8217), .Z(
        P2_U3565) );
  MUX2_X1 U9819 ( .A(n8207), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8217), .Z(
        P2_U3564) );
  MUX2_X1 U9820 ( .A(n8208), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8217), .Z(
        P2_U3563) );
  MUX2_X1 U9821 ( .A(n8209), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8217), .Z(
        P2_U3562) );
  MUX2_X1 U9822 ( .A(n8210), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8217), .Z(
        P2_U3561) );
  MUX2_X1 U9823 ( .A(n8211), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8217), .Z(
        P2_U3560) );
  MUX2_X1 U9824 ( .A(n8212), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8217), .Z(
        P2_U3559) );
  MUX2_X1 U9825 ( .A(n8213), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8217), .Z(
        P2_U3558) );
  MUX2_X1 U9826 ( .A(n8214), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8217), .Z(
        P2_U3557) );
  MUX2_X1 U9827 ( .A(n8215), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8217), .Z(
        P2_U3556) );
  MUX2_X1 U9828 ( .A(n9909), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8217), .Z(
        P2_U3555) );
  MUX2_X1 U9829 ( .A(n8216), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8217), .Z(
        P2_U3554) );
  MUX2_X1 U9830 ( .A(n9911), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8217), .Z(
        P2_U3553) );
  MUX2_X1 U9831 ( .A(n8218), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8217), .Z(
        P2_U3552) );
  INV_X1 U9832 ( .A(n8219), .ZN(n8221) );
  MUX2_X1 U9833 ( .A(n7064), .B(P2_REG2_REG_3__SCAN_IN), .S(n8225), .Z(n8220)
         );
  NAND2_X1 U9834 ( .A1(n8221), .A2(n8220), .ZN(n8223) );
  OAI211_X1 U9835 ( .C1(n8224), .C2(n8223), .A(n10190), .B(n8222), .ZN(n8232)
         );
  AOI22_X1 U9836 ( .A1(n10200), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n8231) );
  NAND2_X1 U9837 ( .A1(n8335), .A2(n8225), .ZN(n8230) );
  OAI211_X1 U9838 ( .C1(n8228), .C2(n8227), .A(n8359), .B(n8226), .ZN(n8229)
         );
  NAND4_X1 U9839 ( .A1(n8232), .A2(n8231), .A3(n8230), .A4(n8229), .ZN(
        P2_U3248) );
  INV_X1 U9840 ( .A(n8233), .ZN(n8236) );
  MUX2_X1 U9841 ( .A(n8234), .B(P2_REG2_REG_5__SCAN_IN), .S(n8239), .Z(n8235)
         );
  NAND3_X1 U9842 ( .A1(n8237), .A2(n8236), .A3(n8235), .ZN(n8238) );
  NAND3_X1 U9843 ( .A1(n10190), .A2(n8251), .A3(n8238), .ZN(n8247) );
  NAND2_X1 U9844 ( .A1(n8335), .A2(n8239), .ZN(n8246) );
  AOI21_X1 U9845 ( .B1(n10200), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8240), .ZN(
        n8245) );
  OAI211_X1 U9846 ( .C1(n8243), .C2(n8242), .A(n8359), .B(n8241), .ZN(n8244)
         );
  NAND4_X1 U9847 ( .A1(n8247), .A2(n8246), .A3(n8245), .A4(n8244), .ZN(
        P2_U3250) );
  INV_X1 U9848 ( .A(n8248), .ZN(n8266) );
  NAND3_X1 U9849 ( .A1(n8251), .A2(n8250), .A3(n8249), .ZN(n8252) );
  NAND3_X1 U9850 ( .A1(n10190), .A2(n8266), .A3(n8252), .ZN(n8262) );
  NAND2_X1 U9851 ( .A1(n8335), .A2(n8253), .ZN(n8261) );
  INV_X1 U9852 ( .A(n8254), .ZN(n8255) );
  AOI21_X1 U9853 ( .B1(n10200), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8255), .ZN(
        n8260) );
  OAI211_X1 U9854 ( .C1(n8258), .C2(n8257), .A(n8359), .B(n8256), .ZN(n8259)
         );
  NAND4_X1 U9855 ( .A1(n8262), .A2(n8261), .A3(n8260), .A4(n8259), .ZN(
        P2_U3251) );
  INV_X1 U9856 ( .A(n8263), .ZN(n8265) );
  MUX2_X1 U9857 ( .A(n6965), .B(P2_REG2_REG_7__SCAN_IN), .S(n8268), .Z(n8264)
         );
  NAND3_X1 U9858 ( .A1(n8266), .A2(n8265), .A3(n8264), .ZN(n8267) );
  NAND3_X1 U9859 ( .A1(n10190), .A2(n8286), .A3(n8267), .ZN(n8276) );
  NAND2_X1 U9860 ( .A1(n8335), .A2(n8268), .ZN(n8275) );
  AOI21_X1 U9861 ( .B1(n10200), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8269), .ZN(
        n8274) );
  OAI211_X1 U9862 ( .C1(n8272), .C2(n8271), .A(n8359), .B(n8270), .ZN(n8273)
         );
  NAND4_X1 U9863 ( .A1(n8276), .A2(n8275), .A3(n8274), .A4(n8273), .ZN(
        P2_U3252) );
  INV_X1 U9864 ( .A(n8277), .ZN(n8280) );
  NOR2_X1 U9865 ( .A1(n10204), .A2(n8278), .ZN(n8279) );
  AOI211_X1 U9866 ( .C1(n10200), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n8280), .B(
        n8279), .ZN(n8291) );
  OAI211_X1 U9867 ( .C1(n8283), .C2(n8282), .A(n8359), .B(n8281), .ZN(n8290)
         );
  INV_X1 U9868 ( .A(n8297), .ZN(n8288) );
  NAND3_X1 U9869 ( .A1(n8286), .A2(n8285), .A3(n8284), .ZN(n8287) );
  NAND3_X1 U9870 ( .A1(n8288), .A2(n10190), .A3(n8287), .ZN(n8289) );
  NAND3_X1 U9871 ( .A1(n8291), .A2(n8290), .A3(n8289), .ZN(P2_U3253) );
  MUX2_X1 U9872 ( .A(n7504), .B(P2_REG2_REG_9__SCAN_IN), .S(n8303), .Z(n8294)
         );
  INV_X1 U9873 ( .A(n8292), .ZN(n8293) );
  NAND2_X1 U9874 ( .A1(n8294), .A2(n8293), .ZN(n8296) );
  OAI211_X1 U9875 ( .C1(n8297), .C2(n8296), .A(n8295), .B(n10190), .ZN(n8307)
         );
  INV_X1 U9876 ( .A(n8298), .ZN(n8299) );
  AOI21_X1 U9877 ( .B1(n10200), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8299), .ZN(
        n8306) );
  OAI211_X1 U9878 ( .C1(n8302), .C2(n8301), .A(n8359), .B(n8300), .ZN(n8305)
         );
  NAND2_X1 U9879 ( .A1(n8335), .A2(n8303), .ZN(n8304) );
  NAND4_X1 U9880 ( .A1(n8307), .A2(n8306), .A3(n8305), .A4(n8304), .ZN(
        P2_U3254) );
  NOR2_X1 U9881 ( .A1(n8309), .A2(n8308), .ZN(n8311) );
  OAI21_X1 U9882 ( .B1(n8311), .B2(n8310), .A(n10190), .ZN(n8321) );
  NOR2_X1 U9883 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8312), .ZN(n8315) );
  NOR2_X1 U9884 ( .A1(n10204), .A2(n8313), .ZN(n8314) );
  AOI211_X1 U9885 ( .C1(n10200), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n8315), .B(
        n8314), .ZN(n8320) );
  OAI211_X1 U9886 ( .C1(n8318), .C2(n8317), .A(n8316), .B(n8359), .ZN(n8319)
         );
  NAND3_X1 U9887 ( .A1(n8321), .A2(n8320), .A3(n8319), .ZN(P2_U3256) );
  NOR2_X1 U9888 ( .A1(n8330), .A2(n8322), .ZN(n8324) );
  MUX2_X1 U9889 ( .A(n5543), .B(P2_REG2_REG_16__SCAN_IN), .S(n8346), .Z(n8325)
         );
  INV_X1 U9890 ( .A(n8325), .ZN(n8326) );
  NAND2_X1 U9891 ( .A1(n8326), .A2(n8327), .ZN(n8341) );
  OAI211_X1 U9892 ( .C1(n8327), .C2(n8326), .A(n10190), .B(n8341), .ZN(n8339)
         );
  AOI21_X1 U9893 ( .B1(n10200), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8328), .ZN(
        n8338) );
  AOI21_X1 U9894 ( .B1(n8331), .B2(n8330), .A(n8329), .ZN(n8333) );
  XOR2_X1 U9895 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8346), .Z(n8332) );
  NAND2_X1 U9896 ( .A1(n8332), .A2(n8333), .ZN(n8345) );
  OAI21_X1 U9897 ( .B1(n8333), .B2(n8332), .A(n8345), .ZN(n8334) );
  NAND2_X1 U9898 ( .A1(n8334), .A2(n8359), .ZN(n8337) );
  NAND2_X1 U9899 ( .A1(n8335), .A2(n8346), .ZN(n8336) );
  NAND4_X1 U9900 ( .A1(n8339), .A2(n8338), .A3(n8337), .A4(n8336), .ZN(
        P2_U3261) );
  NAND2_X1 U9901 ( .A1(n8347), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8343) );
  NOR2_X1 U9902 ( .A1(n8347), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8340) );
  AOI21_X1 U9903 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8347), .A(n8340), .ZN(
        n10191) );
  NAND2_X1 U9904 ( .A1(n8346), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U9905 ( .A1(n8342), .A2(n8341), .ZN(n10192) );
  NAND2_X1 U9906 ( .A1(n10191), .A2(n10192), .ZN(n10189) );
  NAND2_X1 U9907 ( .A1(n8343), .A2(n10189), .ZN(n8360) );
  OAI21_X1 U9908 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8344), .A(n8363), .ZN(
        n8356) );
  XNOR2_X1 U9909 ( .A(n8347), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n10196) );
  OAI21_X1 U9910 ( .B1(n8346), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8345), .ZN(
        n10197) );
  NOR2_X1 U9911 ( .A1(n10196), .A2(n10197), .ZN(n10195) );
  AOI21_X1 U9912 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8347), .A(n10195), .ZN(
        n8349) );
  INV_X1 U9913 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10068) );
  AOI22_X1 U9914 ( .A1(n8361), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n10068), .B2(
        n8350), .ZN(n8348) );
  NAND2_X1 U9915 ( .A1(n8349), .A2(n8348), .ZN(n8357) );
  OAI21_X1 U9916 ( .B1(n8349), .B2(n8348), .A(n8357), .ZN(n8354) );
  NOR2_X1 U9917 ( .A1(n10204), .A2(n8350), .ZN(n8353) );
  INV_X1 U9918 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10213) );
  OAI21_X1 U9919 ( .B1(n8375), .B2(n10213), .A(n8351), .ZN(n8352) );
  AOI211_X1 U9920 ( .C1(n8354), .C2(n8359), .A(n8353), .B(n8352), .ZN(n8355)
         );
  OAI21_X1 U9921 ( .B1(n8356), .B2(n8370), .A(n8355), .ZN(P2_U3263) );
  OAI21_X1 U9922 ( .B1(n8361), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8357), .ZN(
        n8358) );
  XOR2_X1 U9923 ( .A(n8358), .B(P2_REG1_REG_19__SCAN_IN), .Z(n8369) );
  NAND2_X1 U9924 ( .A1(n8369), .A2(n8359), .ZN(n8368) );
  NAND2_X1 U9925 ( .A1(n8361), .A2(n8360), .ZN(n8362) );
  XNOR2_X1 U9926 ( .A(n8364), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8371) );
  NAND3_X1 U9927 ( .A1(n8371), .A2(n8366), .A3(n8365), .ZN(n8367) );
  NAND3_X1 U9928 ( .A1(n8368), .A2(n10204), .A3(n8367), .ZN(n8373) );
  OAI22_X1 U9929 ( .A1(n8371), .A2(n8370), .B1(n8369), .B2(n10194), .ZN(n8372)
         );
  OAI21_X1 U9930 ( .B1(n8375), .B2(n5005), .A(n8374), .ZN(n8376) );
  NOR2_X1 U9931 ( .A1(n8378), .A2(n8377), .ZN(n8662) );
  INV_X1 U9932 ( .A(n8662), .ZN(n8379) );
  NOR2_X1 U9933 ( .A1(n8651), .A2(n8379), .ZN(n8387) );
  AOI21_X1 U9934 ( .B1(n8651), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8387), .ZN(
        n8381) );
  NAND2_X1 U9935 ( .A1(n8659), .A2(n8653), .ZN(n8380) );
  OAI211_X1 U9936 ( .C1(n8661), .C2(n9921), .A(n8381), .B(n8380), .ZN(P2_U3265) );
  INV_X1 U9937 ( .A(n8382), .ZN(n8385) );
  INV_X1 U9938 ( .A(n5030), .ZN(n8384) );
  AND2_X1 U9939 ( .A1(n8651), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8386) );
  NOR2_X1 U9940 ( .A1(n8387), .A2(n8386), .ZN(n8389) );
  NAND2_X1 U9941 ( .A1(n5030), .A2(n8653), .ZN(n8388) );
  OAI211_X1 U9942 ( .C1(n8664), .C2(n9921), .A(n8389), .B(n8388), .ZN(P2_U3266) );
  XNOR2_X1 U9943 ( .A(n8390), .B(n8396), .ZN(n8674) );
  AOI21_X1 U9944 ( .B1(n8670), .B2(n8404), .A(n8391), .ZN(n8671) );
  AOI22_X1 U9945 ( .A1(n8392), .A2(n8649), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8651), .ZN(n8393) );
  OAI21_X1 U9946 ( .B1(n8394), .B2(n9925), .A(n8393), .ZN(n8402) );
  OAI211_X1 U9947 ( .C1(n8397), .C2(n8396), .A(n8395), .B(n9913), .ZN(n8401)
         );
  AOI22_X1 U9948 ( .A1(n8399), .A2(n8596), .B1(n8398), .B2(n9910), .ZN(n8400)
         );
  OAI21_X1 U9949 ( .B1(n8674), .B2(n9924), .A(n4356), .ZN(P2_U3268) );
  XNOR2_X1 U9950 ( .A(n8403), .B(n4890), .ZN(n8679) );
  INV_X1 U9951 ( .A(n8404), .ZN(n8405) );
  AOI21_X1 U9952 ( .B1(n8675), .B2(n8432), .A(n8405), .ZN(n8676) );
  INV_X1 U9953 ( .A(n8406), .ZN(n8407) );
  AOI22_X1 U9954 ( .A1(n8407), .A2(n8649), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8651), .ZN(n8408) );
  OAI21_X1 U9955 ( .B1(n8409), .B2(n9925), .A(n8408), .ZN(n8418) );
  AOI21_X1 U9956 ( .B1(n8411), .B2(n8410), .A(n9892), .ZN(n8416) );
  OAI22_X1 U9957 ( .A1(n8413), .A2(n8640), .B1(n8412), .B2(n8641), .ZN(n8414)
         );
  AOI21_X1 U9958 ( .B1(n8416), .B2(n8415), .A(n8414), .ZN(n8678) );
  NOR2_X1 U9959 ( .A1(n8678), .A2(n8651), .ZN(n8417) );
  AOI211_X1 U9960 ( .C1(n8676), .C2(n8629), .A(n8418), .B(n8417), .ZN(n8419)
         );
  OAI21_X1 U9961 ( .B1(n8679), .B2(n9924), .A(n8419), .ZN(P2_U3269) );
  INV_X1 U9962 ( .A(n8426), .ZN(n8421) );
  XNOR2_X1 U9963 ( .A(n8422), .B(n8421), .ZN(n8683) );
  NAND2_X1 U9964 ( .A1(n8457), .A2(n8424), .ZN(n8445) );
  NAND2_X1 U9965 ( .A1(n8445), .A2(n8444), .ZN(n8443) );
  NAND2_X1 U9966 ( .A1(n8443), .A2(n8425), .ZN(n8427) );
  XNOR2_X1 U9967 ( .A(n8427), .B(n8426), .ZN(n8428) );
  NAND2_X1 U9968 ( .A1(n8428), .A2(n9913), .ZN(n8430) );
  NAND2_X1 U9969 ( .A1(n8430), .A2(n8429), .ZN(n8685) );
  NAND2_X1 U9970 ( .A1(n8440), .A2(n8680), .ZN(n8431) );
  NAND3_X1 U9971 ( .A1(n8432), .A2(n9957), .A3(n8431), .ZN(n8681) );
  INV_X1 U9972 ( .A(n8433), .ZN(n8434) );
  OAI22_X1 U9973 ( .A1(n8681), .A2(n8435), .B1(n8434), .B2(n9919), .ZN(n8436)
         );
  OAI21_X1 U9974 ( .B1(n8685), .B2(n8436), .A(n8606), .ZN(n8438) );
  AOI22_X1 U9975 ( .A1(n8680), .A2(n8653), .B1(n8651), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8437) );
  OAI211_X1 U9976 ( .C1(n8683), .C2(n9924), .A(n8438), .B(n8437), .ZN(P2_U3270) );
  INV_X1 U9977 ( .A(n8439), .ZN(n8442) );
  INV_X1 U9978 ( .A(n8440), .ZN(n8441) );
  AOI211_X1 U9979 ( .C1(n8688), .C2(n8442), .A(n9986), .B(n8441), .ZN(n8687)
         );
  OAI211_X1 U9980 ( .C1(n8445), .C2(n8444), .A(n8443), .B(n9913), .ZN(n8447)
         );
  AOI21_X1 U9981 ( .B1(n8687), .B2(n4954), .A(n8686), .ZN(n8456) );
  NOR2_X1 U9982 ( .A1(n8463), .A2(n8464), .ZN(n8462) );
  NOR2_X1 U9983 ( .A1(n8462), .A2(n8448), .ZN(n8449) );
  XNOR2_X1 U9984 ( .A(n8449), .B(n8021), .ZN(n8690) );
  INV_X1 U9985 ( .A(n8690), .ZN(n8454) );
  AOI22_X1 U9986 ( .A1(n8450), .A2(n8649), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8651), .ZN(n8451) );
  OAI21_X1 U9987 ( .B1(n8452), .B2(n9925), .A(n8451), .ZN(n8453) );
  AOI21_X1 U9988 ( .B1(n8454), .B2(n8611), .A(n8453), .ZN(n8455) );
  OAI21_X1 U9989 ( .B1(n8456), .B2(n8651), .A(n8455), .ZN(P2_U3271) );
  OAI211_X1 U9990 ( .C1(n8464), .C2(n8458), .A(n8457), .B(n9913), .ZN(n8461)
         );
  AOI22_X1 U9991 ( .A1(n8459), .A2(n8596), .B1(n9910), .B2(n8492), .ZN(n8460)
         );
  AOI21_X1 U9992 ( .B1(n8464), .B2(n8463), .A(n8462), .ZN(n8695) );
  INV_X1 U9993 ( .A(n8695), .ZN(n8471) );
  INV_X1 U9994 ( .A(n8691), .ZN(n8469) );
  XOR2_X1 U9995 ( .A(n8477), .B(n8691), .Z(n8692) );
  NAND2_X1 U9996 ( .A1(n8692), .A2(n8629), .ZN(n8468) );
  INV_X1 U9997 ( .A(n8465), .ZN(n8466) );
  AOI22_X1 U9998 ( .A1(n8466), .A2(n8649), .B1(n8651), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8467) );
  OAI211_X1 U9999 ( .C1(n8469), .C2(n9925), .A(n8468), .B(n8467), .ZN(n8470)
         );
  AOI21_X1 U10000 ( .B1(n8471), .B2(n8611), .A(n8470), .ZN(n8472) );
  OAI21_X1 U10001 ( .B1(n8651), .B2(n8694), .A(n8472), .ZN(P2_U3272) );
  XNOR2_X1 U10002 ( .A(n8473), .B(n8482), .ZN(n8475) );
  AOI222_X1 U10003 ( .A1(n9913), .A2(n8475), .B1(n8505), .B2(n9910), .C1(n8474), .C2(n8596), .ZN(n8702) );
  NAND2_X1 U10004 ( .A1(n8696), .A2(n8496), .ZN(n8476) );
  AND2_X1 U10005 ( .A1(n8477), .A2(n8476), .ZN(n8697) );
  NAND2_X1 U10006 ( .A1(n8696), .A2(n8653), .ZN(n8480) );
  AOI22_X1 U10007 ( .A1(n8651), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8478), .B2(
        n8649), .ZN(n8479) );
  NAND2_X1 U10008 ( .A1(n8480), .A2(n8479), .ZN(n8481) );
  AOI21_X1 U10009 ( .B1(n8697), .B2(n8629), .A(n8481), .ZN(n8485) );
  OR2_X1 U10010 ( .A1(n8483), .A2(n8482), .ZN(n8698) );
  NAND3_X1 U10011 ( .A1(n8698), .A2(n8699), .A3(n8611), .ZN(n8484) );
  OAI211_X1 U10012 ( .C1(n8702), .C2(n8651), .A(n8485), .B(n8484), .ZN(
        P2_U3273) );
  XNOR2_X1 U10013 ( .A(n8487), .B(n8486), .ZN(n8706) );
  NAND2_X1 U10014 ( .A1(n8489), .A2(n8488), .ZN(n8490) );
  NAND3_X1 U10015 ( .A1(n8491), .A2(n9913), .A3(n8490), .ZN(n8494) );
  AOI22_X1 U10016 ( .A1(n8492), .A2(n8596), .B1(n9910), .B2(n8520), .ZN(n8493)
         );
  NAND2_X1 U10017 ( .A1(n8494), .A2(n8493), .ZN(n8708) );
  NAND2_X1 U10018 ( .A1(n8708), .A2(n8606), .ZN(n8503) );
  OR2_X1 U10019 ( .A1(n8500), .A2(n4349), .ZN(n8495) );
  AND2_X1 U10020 ( .A1(n8496), .A2(n8495), .ZN(n8704) );
  INV_X1 U10021 ( .A(n8497), .ZN(n8498) );
  AOI22_X1 U10022 ( .A1(n8651), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8498), .B2(
        n8649), .ZN(n8499) );
  OAI21_X1 U10023 ( .B1(n8500), .B2(n9925), .A(n8499), .ZN(n8501) );
  AOI21_X1 U10024 ( .B1(n8704), .B2(n8629), .A(n8501), .ZN(n8502) );
  OAI211_X1 U10025 ( .C1(n8706), .C2(n9924), .A(n8503), .B(n8502), .ZN(
        P2_U3274) );
  XNOR2_X1 U10026 ( .A(n8504), .B(n8510), .ZN(n8506) );
  AOI222_X1 U10027 ( .A1(n9913), .A2(n8506), .B1(n8535), .B2(n9910), .C1(n8505), .C2(n8596), .ZN(n8712) );
  XOR2_X1 U10028 ( .A(n8524), .B(n8709), .Z(n8710) );
  INV_X1 U10029 ( .A(n8709), .ZN(n8509) );
  AOI22_X1 U10030 ( .A1(n8651), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8507), .B2(
        n8649), .ZN(n8508) );
  OAI21_X1 U10031 ( .B1(n8509), .B2(n9925), .A(n8508), .ZN(n8513) );
  XOR2_X1 U10032 ( .A(n8511), .B(n8510), .Z(n8713) );
  NOR2_X1 U10033 ( .A1(n8713), .A2(n9924), .ZN(n8512) );
  AOI211_X1 U10034 ( .C1(n8710), .C2(n8629), .A(n8513), .B(n8512), .ZN(n8514)
         );
  OAI21_X1 U10035 ( .B1(n8651), .B2(n8712), .A(n8514), .ZN(P2_U3275) );
  XNOR2_X1 U10036 ( .A(n8515), .B(n8517), .ZN(n8717) );
  INV_X1 U10037 ( .A(n8517), .ZN(n8518) );
  XNOR2_X1 U10038 ( .A(n8516), .B(n8518), .ZN(n8519) );
  NAND2_X1 U10039 ( .A1(n8519), .A2(n9913), .ZN(n8522) );
  AOI22_X1 U10040 ( .A1(n8520), .A2(n8596), .B1(n9910), .B2(n8547), .ZN(n8521)
         );
  NAND2_X1 U10041 ( .A1(n8522), .A2(n8521), .ZN(n8719) );
  NAND2_X1 U10042 ( .A1(n8719), .A2(n8606), .ZN(n8531) );
  NAND2_X1 U10043 ( .A1(n8537), .A2(n8714), .ZN(n8523) );
  AND2_X1 U10044 ( .A1(n8524), .A2(n8523), .ZN(n8715) );
  INV_X1 U10045 ( .A(n8714), .ZN(n8528) );
  INV_X1 U10046 ( .A(n8525), .ZN(n8526) );
  AOI22_X1 U10047 ( .A1(n8651), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8526), .B2(
        n8649), .ZN(n8527) );
  OAI21_X1 U10048 ( .B1(n8528), .B2(n9925), .A(n8527), .ZN(n8529) );
  AOI21_X1 U10049 ( .B1(n8629), .B2(n8715), .A(n8529), .ZN(n8530) );
  OAI211_X1 U10050 ( .C1(n8717), .C2(n9924), .A(n8531), .B(n8530), .ZN(
        P2_U3276) );
  XOR2_X1 U10051 ( .A(n8533), .B(n8532), .Z(n8724) );
  OAI21_X1 U10052 ( .B1(n5887), .B2(n5129), .A(n8534), .ZN(n8536) );
  AOI222_X1 U10053 ( .A1(n9913), .A2(n8536), .B1(n8563), .B2(n9910), .C1(n8535), .C2(n8596), .ZN(n8723) );
  INV_X1 U10054 ( .A(n8549), .ZN(n8539) );
  INV_X1 U10055 ( .A(n8537), .ZN(n8538) );
  AOI211_X1 U10056 ( .C1(n8721), .C2(n8539), .A(n9986), .B(n8538), .ZN(n8720)
         );
  AOI22_X1 U10057 ( .A1(n8720), .A2(n4954), .B1(n8649), .B2(n8540), .ZN(n8541)
         );
  AOI21_X1 U10058 ( .B1(n8723), .B2(n8541), .A(n8651), .ZN(n8542) );
  INV_X1 U10059 ( .A(n8542), .ZN(n8544) );
  AOI22_X1 U10060 ( .A1(n8721), .A2(n8653), .B1(n8651), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8543) );
  OAI211_X1 U10061 ( .C1(n8724), .C2(n9924), .A(n8544), .B(n8543), .ZN(
        P2_U3277) );
  XNOR2_X1 U10062 ( .A(n8546), .B(n8545), .ZN(n8548) );
  AOI222_X1 U10063 ( .A1(n9913), .A2(n8548), .B1(n8579), .B2(n9910), .C1(n8547), .C2(n8596), .ZN(n8728) );
  INV_X1 U10064 ( .A(n8567), .ZN(n8550) );
  AOI21_X1 U10065 ( .B1(n8725), .B2(n8550), .A(n8549), .ZN(n8726) );
  INV_X1 U10066 ( .A(n8551), .ZN(n8552) );
  AOI22_X1 U10067 ( .A1(n8651), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8552), .B2(
        n8649), .ZN(n8553) );
  OAI21_X1 U10068 ( .B1(n5013), .B2(n9925), .A(n8553), .ZN(n8557) );
  XNOR2_X1 U10069 ( .A(n8555), .B(n8554), .ZN(n8729) );
  NOR2_X1 U10070 ( .A1(n8729), .A2(n9924), .ZN(n8556) );
  AOI211_X1 U10071 ( .C1(n8726), .C2(n8629), .A(n8557), .B(n8556), .ZN(n8558)
         );
  OAI21_X1 U10072 ( .B1(n8728), .B2(n8651), .A(n8558), .ZN(P2_U3278) );
  NAND2_X1 U10073 ( .A1(n8578), .A2(n8559), .ZN(n8560) );
  XNOR2_X1 U10074 ( .A(n8560), .B(n8561), .ZN(n8734) );
  XNOR2_X1 U10075 ( .A(n8562), .B(n8561), .ZN(n8564) );
  AOI222_X1 U10076 ( .A1(n9913), .A2(n8564), .B1(n8563), .B2(n8596), .C1(n8597), .C2(n9910), .ZN(n8733) );
  NAND2_X1 U10077 ( .A1(n8584), .A2(n8731), .ZN(n8565) );
  NAND2_X1 U10078 ( .A1(n8565), .A2(n9957), .ZN(n8566) );
  NOR2_X1 U10079 ( .A1(n8567), .A2(n8566), .ZN(n8730) );
  NAND2_X1 U10080 ( .A1(n8730), .A2(n4954), .ZN(n8568) );
  OAI211_X1 U10081 ( .C1(n9919), .C2(n8569), .A(n8733), .B(n8568), .ZN(n8570)
         );
  NAND2_X1 U10082 ( .A1(n8570), .A2(n8606), .ZN(n8572) );
  AOI22_X1 U10083 ( .A1(n8731), .A2(n8653), .B1(n8651), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8571) );
  OAI211_X1 U10084 ( .C1(n8734), .C2(n9924), .A(n8572), .B(n8571), .ZN(
        P2_U3279) );
  XNOR2_X1 U10085 ( .A(n8574), .B(n8573), .ZN(n8583) );
  NAND2_X1 U10086 ( .A1(n8576), .A2(n8575), .ZN(n8577) );
  NAND2_X1 U10087 ( .A1(n8578), .A2(n8577), .ZN(n8739) );
  AOI22_X1 U10088 ( .A1(n8579), .A2(n8596), .B1(n9910), .B2(n8626), .ZN(n8580)
         );
  OAI21_X1 U10089 ( .B1(n8739), .B2(n8581), .A(n8580), .ZN(n8582) );
  AOI21_X1 U10090 ( .B1(n9913), .B2(n8583), .A(n8582), .ZN(n8738) );
  INV_X1 U10091 ( .A(n8584), .ZN(n8585) );
  AOI21_X1 U10092 ( .B1(n8735), .B2(n8603), .A(n8585), .ZN(n8736) );
  AOI22_X1 U10093 ( .A1(n8651), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8586), .B2(
        n8649), .ZN(n8587) );
  OAI21_X1 U10094 ( .B1(n4985), .B2(n9925), .A(n8587), .ZN(n8590) );
  NOR2_X1 U10095 ( .A1(n8739), .A2(n8588), .ZN(n8589) );
  AOI211_X1 U10096 ( .C1(n8736), .C2(n8629), .A(n8590), .B(n8589), .ZN(n8591)
         );
  OAI21_X1 U10097 ( .B1(n8651), .B2(n8738), .A(n8591), .ZN(P2_U3280) );
  OAI211_X1 U10098 ( .C1(n8594), .C2(n8593), .A(n8592), .B(n9913), .ZN(n8599)
         );
  AOI22_X1 U10099 ( .A1(n8597), .A2(n8596), .B1(n9910), .B2(n8595), .ZN(n8598)
         );
  NAND2_X1 U10100 ( .A1(n8599), .A2(n8598), .ZN(n8742) );
  INV_X1 U10101 ( .A(n8742), .ZN(n8613) );
  OAI21_X1 U10102 ( .B1(n8602), .B2(n8601), .A(n8600), .ZN(n8744) );
  OAI21_X1 U10103 ( .B1(n4361), .B2(n8740), .A(n8603), .ZN(n8741) );
  INV_X1 U10104 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8605) );
  OAI22_X1 U10105 ( .A1(n8606), .A2(n8605), .B1(n8604), .B2(n9919), .ZN(n8607)
         );
  AOI21_X1 U10106 ( .B1(n8608), .B2(n8653), .A(n8607), .ZN(n8609) );
  OAI21_X1 U10107 ( .B1(n8741), .B2(n9921), .A(n8609), .ZN(n8610) );
  AOI21_X1 U10108 ( .B1(n8744), .B2(n8611), .A(n8610), .ZN(n8612) );
  OAI21_X1 U10109 ( .B1(n8613), .B2(n8651), .A(n8612), .ZN(P2_U3281) );
  OR2_X1 U10110 ( .A1(n8632), .A2(n8631), .ZN(n8634) );
  NAND2_X1 U10111 ( .A1(n8634), .A2(n8614), .ZN(n8615) );
  XNOR2_X1 U10112 ( .A(n8615), .B(n8623), .ZN(n8750) );
  AOI21_X1 U10113 ( .B1(n8746), .B2(n8648), .A(n4361), .ZN(n8747) );
  AOI22_X1 U10114 ( .A1(n8651), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8616), .B2(
        n8649), .ZN(n8617) );
  OAI21_X1 U10115 ( .B1(n8618), .B2(n9925), .A(n8617), .ZN(n8628) );
  AND2_X1 U10116 ( .A1(n9910), .A2(n8619), .ZN(n8625) );
  INV_X1 U10117 ( .A(n8620), .ZN(n8621) );
  AOI211_X1 U10118 ( .C1(n8623), .C2(n8622), .A(n9892), .B(n8621), .ZN(n8624)
         );
  AOI211_X1 U10119 ( .C1(n8596), .C2(n8626), .A(n8625), .B(n8624), .ZN(n8749)
         );
  NOR2_X1 U10120 ( .A1(n8749), .A2(n8651), .ZN(n8627) );
  AOI211_X1 U10121 ( .C1(n8747), .C2(n8629), .A(n8628), .B(n8627), .ZN(n8630)
         );
  OAI21_X1 U10122 ( .B1(n9924), .B2(n8750), .A(n8630), .ZN(P2_U3282) );
  NAND2_X1 U10123 ( .A1(n8632), .A2(n8631), .ZN(n8633) );
  NAND2_X1 U10124 ( .A1(n8636), .A2(n8635), .ZN(n8637) );
  AOI21_X1 U10125 ( .B1(n8638), .B2(n8637), .A(n9892), .ZN(n8644) );
  OAI22_X1 U10126 ( .A1(n8642), .A2(n8641), .B1(n8640), .B2(n8639), .ZN(n8643)
         );
  AOI211_X1 U10127 ( .C1(n8752), .C2(n8645), .A(n8644), .B(n8643), .ZN(n8757)
         );
  NAND2_X1 U10128 ( .A1(n8646), .A2(n8652), .ZN(n8647) );
  NAND2_X1 U10129 ( .A1(n8648), .A2(n8647), .ZN(n8754) );
  AOI22_X1 U10130 ( .A1(n8651), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8650), .B2(
        n8649), .ZN(n8655) );
  NAND2_X1 U10131 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  OAI211_X1 U10132 ( .C1(n8754), .C2(n9921), .A(n8655), .B(n8654), .ZN(n8656)
         );
  AOI21_X1 U10133 ( .B1(n8752), .B2(n8657), .A(n8656), .ZN(n8658) );
  OAI21_X1 U10134 ( .B1(n8757), .B2(n8651), .A(n8658), .ZN(P2_U3283) );
  AOI21_X1 U10135 ( .B1(n8659), .B2(n9956), .A(n8662), .ZN(n8660) );
  OAI21_X1 U10136 ( .B1(n8661), .B2(n9986), .A(n8660), .ZN(n8769) );
  MUX2_X1 U10137 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8769), .S(n10004), .Z(
        P2_U3551) );
  AOI21_X1 U10138 ( .B1(n5030), .B2(n9956), .A(n8662), .ZN(n8663) );
  OAI21_X1 U10139 ( .B1(n8664), .B2(n9986), .A(n8663), .ZN(n8770) );
  MUX2_X1 U10140 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8770), .S(n10004), .Z(
        P2_U3550) );
  AOI22_X1 U10141 ( .A1(n8667), .A2(n9957), .B1(n9956), .B2(n8666), .ZN(n8668)
         );
  AOI22_X1 U10142 ( .A1(n8671), .A2(n9957), .B1(n9956), .B2(n8670), .ZN(n8672)
         );
  OAI211_X1 U10143 ( .C1(n8751), .C2(n8674), .A(n8673), .B(n8672), .ZN(n8772)
         );
  MUX2_X1 U10144 ( .A(n8772), .B(P2_REG1_REG_28__SCAN_IN), .S(n10002), .Z(
        P2_U3548) );
  AOI22_X1 U10145 ( .A1(n8676), .A2(n9957), .B1(n9956), .B2(n8675), .ZN(n8677)
         );
  OAI211_X1 U10146 ( .C1(n8679), .C2(n8751), .A(n8678), .B(n8677), .ZN(n8773)
         );
  MUX2_X1 U10147 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8773), .S(n10004), .Z(
        P2_U3547) );
  NAND2_X1 U10148 ( .A1(n8680), .A2(n9956), .ZN(n8682) );
  OAI211_X1 U10149 ( .C1(n8683), .C2(n8751), .A(n8682), .B(n8681), .ZN(n8684)
         );
  OR2_X2 U10150 ( .A1(n8685), .A2(n8684), .ZN(n8774) );
  MUX2_X1 U10151 ( .A(n8774), .B(P2_REG1_REG_26__SCAN_IN), .S(n10002), .Z(
        P2_U3546) );
  OAI21_X1 U10152 ( .B1(n8751), .B2(n8690), .A(n8689), .ZN(n8775) );
  MUX2_X1 U10153 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8775), .S(n10004), .Z(
        P2_U3545) );
  AOI22_X1 U10154 ( .A1(n8692), .A2(n9957), .B1(n9956), .B2(n8691), .ZN(n8693)
         );
  OAI211_X1 U10155 ( .C1(n8695), .C2(n8751), .A(n8694), .B(n8693), .ZN(n8776)
         );
  MUX2_X1 U10156 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8776), .S(n10004), .Z(
        P2_U3544) );
  AOI22_X1 U10157 ( .A1(n8697), .A2(n9957), .B1(n9956), .B2(n8696), .ZN(n8701)
         );
  NAND3_X1 U10158 ( .A1(n8699), .A2(n8698), .A3(n9981), .ZN(n8700) );
  NAND3_X1 U10159 ( .A1(n8702), .A2(n8701), .A3(n8700), .ZN(n8777) );
  MUX2_X1 U10160 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8777), .S(n10004), .Z(
        P2_U3543) );
  AOI22_X1 U10161 ( .A1(n8704), .A2(n9957), .B1(n9956), .B2(n8703), .ZN(n8705)
         );
  OAI21_X1 U10162 ( .B1(n8706), .B2(n8751), .A(n8705), .ZN(n8707) );
  MUX2_X1 U10163 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8778), .S(n10004), .Z(
        P2_U3542) );
  AOI22_X1 U10164 ( .A1(n8710), .A2(n9957), .B1(n9956), .B2(n8709), .ZN(n8711)
         );
  OAI211_X1 U10165 ( .C1(n8751), .C2(n8713), .A(n8712), .B(n8711), .ZN(n8779)
         );
  MUX2_X1 U10166 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8779), .S(n10004), .Z(
        P2_U3541) );
  AOI22_X1 U10167 ( .A1(n8715), .A2(n9957), .B1(n9956), .B2(n8714), .ZN(n8716)
         );
  OAI21_X1 U10168 ( .B1(n8717), .B2(n8751), .A(n8716), .ZN(n8718) );
  MUX2_X1 U10169 ( .A(n8780), .B(P2_REG1_REG_20__SCAN_IN), .S(n10002), .Z(
        P2_U3540) );
  AOI21_X1 U10170 ( .B1(n9956), .B2(n8721), .A(n8720), .ZN(n8722) );
  OAI211_X1 U10171 ( .C1(n8751), .C2(n8724), .A(n8723), .B(n8722), .ZN(n8781)
         );
  MUX2_X1 U10172 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8781), .S(n10004), .Z(
        P2_U3539) );
  AOI22_X1 U10173 ( .A1(n8726), .A2(n9957), .B1(n9956), .B2(n8725), .ZN(n8727)
         );
  OAI211_X1 U10174 ( .C1(n8751), .C2(n8729), .A(n8728), .B(n8727), .ZN(n8782)
         );
  MUX2_X1 U10175 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8782), .S(n10004), .Z(
        P2_U3538) );
  AOI21_X1 U10176 ( .B1(n9956), .B2(n8731), .A(n8730), .ZN(n8732) );
  OAI211_X1 U10177 ( .C1(n8751), .C2(n8734), .A(n8733), .B(n8732), .ZN(n8783)
         );
  MUX2_X1 U10178 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8783), .S(n10004), .Z(
        P2_U3537) );
  AOI22_X1 U10179 ( .A1(n8736), .A2(n9957), .B1(n9956), .B2(n8735), .ZN(n8737)
         );
  OAI211_X1 U10180 ( .C1(n9984), .C2(n8739), .A(n8738), .B(n8737), .ZN(n8784)
         );
  MUX2_X1 U10181 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8784), .S(n10004), .Z(
        P2_U3536) );
  OAI22_X1 U10182 ( .A1(n8741), .A2(n9986), .B1(n8740), .B2(n9985), .ZN(n8743)
         );
  AOI211_X1 U10183 ( .C1(n9981), .C2(n8744), .A(n8743), .B(n8742), .ZN(n8745)
         );
  INV_X1 U10184 ( .A(n8745), .ZN(n8785) );
  MUX2_X1 U10185 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8785), .S(n10004), .Z(
        P2_U3535) );
  AOI22_X1 U10186 ( .A1(n8747), .A2(n9957), .B1(n9956), .B2(n8746), .ZN(n8748)
         );
  OAI211_X1 U10187 ( .C1(n8751), .C2(n8750), .A(n8749), .B(n8748), .ZN(n8786)
         );
  MUX2_X1 U10188 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8786), .S(n10004), .Z(
        P2_U3534) );
  INV_X1 U10189 ( .A(n8752), .ZN(n8758) );
  OAI22_X1 U10190 ( .A1(n8754), .A2(n9986), .B1(n8753), .B2(n9985), .ZN(n8755)
         );
  INV_X1 U10191 ( .A(n8755), .ZN(n8756) );
  OAI211_X1 U10192 ( .C1(n9984), .C2(n8758), .A(n8757), .B(n8756), .ZN(n8787)
         );
  MUX2_X1 U10193 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8787), .S(n10004), .Z(
        P2_U3533) );
  AOI22_X1 U10194 ( .A1(n8760), .A2(n9957), .B1(n9956), .B2(n8759), .ZN(n8761)
         );
  OAI211_X1 U10195 ( .C1(n8763), .C2(n9984), .A(n8762), .B(n8761), .ZN(n8788)
         );
  MUX2_X1 U10196 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8788), .S(n10004), .Z(
        P2_U3530) );
  AOI22_X1 U10197 ( .A1(n8765), .A2(n9957), .B1(n9956), .B2(n8764), .ZN(n8766)
         );
  OAI211_X1 U10198 ( .C1(n9984), .C2(n8768), .A(n8767), .B(n8766), .ZN(n8789)
         );
  MUX2_X1 U10199 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8789), .S(n10004), .Z(
        P2_U3529) );
  MUX2_X1 U10200 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8769), .S(n9994), .Z(
        P2_U3519) );
  MUX2_X1 U10201 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8770), .S(n9994), .Z(
        P2_U3518) );
  MUX2_X1 U10202 ( .A(n8772), .B(P2_REG0_REG_28__SCAN_IN), .S(n9992), .Z(
        P2_U3516) );
  MUX2_X1 U10203 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8773), .S(n9994), .Z(
        P2_U3515) );
  MUX2_X1 U10204 ( .A(n8774), .B(P2_REG0_REG_26__SCAN_IN), .S(n9992), .Z(
        P2_U3514) );
  MUX2_X1 U10205 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8775), .S(n9994), .Z(
        P2_U3513) );
  MUX2_X1 U10206 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8776), .S(n9994), .Z(
        P2_U3512) );
  MUX2_X1 U10207 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8777), .S(n9994), .Z(
        P2_U3511) );
  MUX2_X1 U10208 ( .A(n8778), .B(P2_REG0_REG_22__SCAN_IN), .S(n9992), .Z(
        P2_U3510) );
  MUX2_X1 U10209 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8779), .S(n9994), .Z(
        P2_U3509) );
  MUX2_X1 U10210 ( .A(n8780), .B(P2_REG0_REG_20__SCAN_IN), .S(n9992), .Z(
        P2_U3508) );
  MUX2_X1 U10211 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8781), .S(n9994), .Z(
        P2_U3507) );
  MUX2_X1 U10212 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8782), .S(n9994), .Z(
        P2_U3505) );
  MUX2_X1 U10213 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8783), .S(n9994), .Z(
        P2_U3502) );
  MUX2_X1 U10214 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8784), .S(n9994), .Z(
        P2_U3499) );
  MUX2_X1 U10215 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8785), .S(n9994), .Z(
        P2_U3496) );
  MUX2_X1 U10216 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8786), .S(n9994), .Z(
        P2_U3493) );
  MUX2_X1 U10217 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8787), .S(n9994), .Z(
        P2_U3490) );
  MUX2_X1 U10218 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n8788), .S(n9994), .Z(
        P2_U3481) );
  MUX2_X1 U10219 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n8789), .S(n9994), .Z(
        P2_U3478) );
  INV_X1 U10220 ( .A(n9048), .ZN(n9731) );
  NOR4_X1 U10221 ( .A1(n8790), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5168), .A4(
        P2_U3152), .ZN(n8791) );
  AOI21_X1 U10222 ( .B1(n8805), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8791), .ZN(
        n8792) );
  OAI21_X1 U10223 ( .B1(n9731), .B2(n8799), .A(n8792), .ZN(P2_U3327) );
  INV_X1 U10224 ( .A(n8793), .ZN(n9733) );
  OAI222_X1 U10225 ( .A1(n8811), .A2(n8796), .B1(P2_U3152), .B2(n8794), .C1(
        n8799), .C2(n9733), .ZN(P2_U3329) );
  INV_X1 U10226 ( .A(n9736), .ZN(n8800) );
  NAND2_X1 U10227 ( .A1(n8805), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U10228 ( .C1(n8800), .C2(n8799), .A(n8798), .B(n8797), .ZN(
        P2_U3330) );
  INV_X1 U10229 ( .A(n8801), .ZN(n9742) );
  AOI21_X1 U10230 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8805), .A(n8802), .ZN(
        n8803) );
  OAI21_X1 U10231 ( .B1(n9742), .B2(n8799), .A(n8803), .ZN(P2_U3331) );
  INV_X1 U10232 ( .A(n8804), .ZN(n9745) );
  AOI22_X1 U10233 ( .A1(n8806), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8805), .ZN(n8807) );
  OAI21_X1 U10234 ( .B1(n9745), .B2(n8799), .A(n8807), .ZN(P2_U3332) );
  OAI222_X1 U10235 ( .A1(n8811), .A2(n8810), .B1(n8799), .B2(n8809), .C1(n8808), .C2(P2_U3152), .ZN(P2_U3333) );
  MUX2_X1 U10236 ( .A(n8812), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10237 ( .A(n8814), .B(n8813), .ZN(n8815) );
  XNOR2_X1 U10238 ( .A(n8816), .B(n8815), .ZN(n8822) );
  INV_X1 U10239 ( .A(n8817), .ZN(n9407) );
  AOI22_X1 U10240 ( .A1(n9407), .A2(n8991), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8819) );
  NAND2_X1 U10241 ( .A1(n9433), .A2(n8984), .ZN(n8818) );
  OAI211_X1 U10242 ( .C1(n9413), .C2(n8986), .A(n8819), .B(n8818), .ZN(n8820)
         );
  AOI21_X1 U10243 ( .B1(n9612), .B2(n8978), .A(n8820), .ZN(n8821) );
  OAI21_X1 U10244 ( .B1(n8822), .B2(n8993), .A(n8821), .ZN(P1_U3212) );
  INV_X1 U10245 ( .A(n8824), .ZN(n8944) );
  INV_X1 U10246 ( .A(n8946), .ZN(n8825) );
  NAND2_X1 U10247 ( .A1(n8947), .A2(n8825), .ZN(n8827) );
  INV_X1 U10248 ( .A(n8889), .ZN(n8833) );
  NAND2_X1 U10249 ( .A1(n8827), .A2(n8826), .ZN(n8829) );
  NAND2_X1 U10250 ( .A1(n8829), .A2(n8828), .ZN(n8890) );
  INV_X1 U10251 ( .A(n8829), .ZN(n8831) );
  OAI21_X1 U10252 ( .B1(n8833), .B2(n8831), .A(n8830), .ZN(n8832) );
  OAI211_X1 U10253 ( .C1(n8833), .C2(n8890), .A(n8832), .B(n8964), .ZN(n8839)
         );
  NAND2_X1 U10254 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9290) );
  OAI21_X1 U10255 ( .B1(n8968), .B2(n8834), .A(n9290), .ZN(n8837) );
  NOR2_X1 U10256 ( .A1(n8966), .A2(n8835), .ZN(n8836) );
  AOI211_X1 U10257 ( .C1(n8971), .C2(n9552), .A(n8837), .B(n8836), .ZN(n8838)
         );
  OAI211_X1 U10258 ( .C1(n8840), .C2(n8988), .A(n8839), .B(n8838), .ZN(
        P1_U3213) );
  NOR2_X1 U10259 ( .A1(n8956), .A2(n8841), .ZN(n8910) );
  INV_X1 U10260 ( .A(n8910), .ZN(n8842) );
  NAND2_X1 U10261 ( .A1(n8956), .A2(n8841), .ZN(n8911) );
  NAND2_X1 U10262 ( .A1(n8842), .A2(n8911), .ZN(n8844) );
  XNOR2_X1 U10263 ( .A(n8844), .B(n8843), .ZN(n8852) );
  NAND2_X1 U10264 ( .A1(n9447), .A2(n8984), .ZN(n8845) );
  OAI21_X1 U10265 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n8846), .A(n8845), .ZN(
        n8847) );
  AOI21_X1 U10266 ( .B1(n9453), .B2(n8991), .A(n8847), .ZN(n8848) );
  OAI21_X1 U10267 ( .B1(n8849), .B2(n8986), .A(n8848), .ZN(n8850) );
  AOI21_X1 U10268 ( .B1(n9631), .B2(n8978), .A(n8850), .ZN(n8851) );
  OAI21_X1 U10269 ( .B1(n8852), .B2(n8993), .A(n8851), .ZN(P1_U3214) );
  XNOR2_X1 U10270 ( .A(n8864), .B(n8860), .ZN(n8853) );
  XNOR2_X1 U10271 ( .A(n8865), .B(n8853), .ZN(n8859) );
  NOR2_X1 U10272 ( .A1(n8854), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9374) );
  AOI21_X1 U10273 ( .B1(n7932), .B2(n8984), .A(n9374), .ZN(n8856) );
  NAND2_X1 U10274 ( .A1(n9515), .A2(n8991), .ZN(n8855) );
  OAI211_X1 U10275 ( .C1(n9483), .C2(n8986), .A(n8856), .B(n8855), .ZN(n8857)
         );
  AOI21_X1 U10276 ( .B1(n9651), .B2(n8978), .A(n8857), .ZN(n8858) );
  OAI21_X1 U10277 ( .B1(n8859), .B2(n8993), .A(n8858), .ZN(P1_U3217) );
  INV_X1 U10278 ( .A(n8865), .ZN(n8862) );
  AOI21_X1 U10279 ( .B1(n8862), .B2(n8861), .A(n8860), .ZN(n8863) );
  AOI21_X1 U10280 ( .B1(n8865), .B2(n8864), .A(n8863), .ZN(n8934) );
  INV_X1 U10281 ( .A(n8934), .ZN(n8867) );
  INV_X1 U10282 ( .A(n8935), .ZN(n8866) );
  NOR2_X1 U10283 ( .A1(n8867), .A2(n8866), .ZN(n8938) );
  INV_X1 U10284 ( .A(n8868), .ZN(n8869) );
  NAND2_X1 U10285 ( .A1(n8870), .A2(n8869), .ZN(n8937) );
  INV_X1 U10286 ( .A(n8937), .ZN(n8871) );
  NOR3_X1 U10287 ( .A1(n8938), .A2(n8872), .A3(n8871), .ZN(n8873) );
  OAI21_X1 U10288 ( .B1(n8873), .B2(n4336), .A(n8964), .ZN(n8878) );
  INV_X1 U10289 ( .A(n9487), .ZN(n8876) );
  AOI22_X1 U10290 ( .A1(n9511), .A2(n8984), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8874) );
  OAI21_X1 U10291 ( .B1(n9482), .B2(n8986), .A(n8874), .ZN(n8875) );
  AOI21_X1 U10292 ( .B1(n8876), .B2(n8991), .A(n8875), .ZN(n8877) );
  OAI211_X1 U10293 ( .C1(n8879), .C2(n8988), .A(n8878), .B(n8877), .ZN(
        P1_U3221) );
  XOR2_X1 U10294 ( .A(n8880), .B(n8881), .Z(n8887) );
  INV_X1 U10295 ( .A(n8882), .ZN(n9439) );
  AOI22_X1 U10296 ( .A1(n9439), .A2(n8991), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8884) );
  NAND2_X1 U10297 ( .A1(n9448), .A2(n8984), .ZN(n8883) );
  OAI211_X1 U10298 ( .C1(n9412), .C2(n8986), .A(n8884), .B(n8883), .ZN(n8885)
         );
  AOI21_X1 U10299 ( .B1(n9622), .B2(n8978), .A(n8885), .ZN(n8886) );
  OAI21_X1 U10300 ( .B1(n8887), .B2(n8993), .A(n8886), .ZN(P1_U3223) );
  NAND3_X1 U10301 ( .A1(n8890), .A2(n8888), .A3(n8889), .ZN(n8980) );
  AOI21_X1 U10302 ( .B1(n8890), .B2(n8889), .A(n8888), .ZN(n8979) );
  AOI21_X1 U10303 ( .B1(n8891), .B2(n8980), .A(n8979), .ZN(n8895) );
  XNOR2_X1 U10304 ( .A(n8893), .B(n8892), .ZN(n8894) );
  XNOR2_X1 U10305 ( .A(n8895), .B(n8894), .ZN(n8901) );
  NAND2_X1 U10306 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9328) );
  OAI21_X1 U10307 ( .B1(n8896), .B2(n8986), .A(n9328), .ZN(n8897) );
  AOI21_X1 U10308 ( .B1(n8984), .B2(n9552), .A(n8897), .ZN(n8898) );
  OAI21_X1 U10309 ( .B1(n8966), .B2(n9556), .A(n8898), .ZN(n8899) );
  AOI21_X1 U10310 ( .B1(n9668), .B2(n8978), .A(n8899), .ZN(n8900) );
  OAI21_X1 U10311 ( .B1(n8901), .B2(n8993), .A(n8900), .ZN(P1_U3224) );
  XOR2_X1 U10312 ( .A(n8903), .B(n8902), .Z(n8909) );
  NAND2_X1 U10313 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U10314 ( .A1(n8984), .A2(n9573), .ZN(n8904) );
  OAI211_X1 U10315 ( .C1(n8905), .C2(n8986), .A(n9343), .B(n8904), .ZN(n8906)
         );
  AOI21_X1 U10316 ( .B1(n9543), .B2(n8991), .A(n8906), .ZN(n8908) );
  NAND2_X1 U10317 ( .A1(n9663), .A2(n8978), .ZN(n8907) );
  OAI211_X1 U10318 ( .C1(n8909), .C2(n8993), .A(n8908), .B(n8907), .ZN(
        P1_U3226) );
  AOI21_X1 U10319 ( .B1(n8912), .B2(n8911), .A(n8910), .ZN(n8916) );
  XNOR2_X1 U10320 ( .A(n8914), .B(n8913), .ZN(n8915) );
  XNOR2_X1 U10321 ( .A(n8916), .B(n8915), .ZN(n8924) );
  INV_X1 U10322 ( .A(n8917), .ZN(n8918) );
  AOI22_X1 U10323 ( .A1(n8918), .A2(n8991), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8920) );
  NAND2_X1 U10324 ( .A1(n9462), .A2(n8984), .ZN(n8919) );
  OAI211_X1 U10325 ( .C1(n8921), .C2(n8986), .A(n8920), .B(n8919), .ZN(n8922)
         );
  AOI21_X1 U10326 ( .B1(n9628), .B2(n8978), .A(n8922), .ZN(n8923) );
  OAI21_X1 U10327 ( .B1(n8924), .B2(n8993), .A(n8923), .ZN(P1_U3227) );
  OAI211_X1 U10328 ( .C1(n8927), .C2(n8926), .A(n8925), .B(n8964), .ZN(n8933)
         );
  AOI21_X1 U10329 ( .B1(n8984), .B2(n9283), .A(n8928), .ZN(n8932) );
  AOI22_X1 U10330 ( .A1(n8971), .A2(n9281), .B1(n9833), .B2(n8978), .ZN(n8931)
         );
  NAND2_X1 U10331 ( .A1(n8991), .A2(n8929), .ZN(n8930) );
  NAND4_X1 U10332 ( .A1(n8933), .A2(n8932), .A3(n8931), .A4(n8930), .ZN(
        P1_U3228) );
  AOI21_X1 U10333 ( .B1(n8935), .B2(n8937), .A(n8934), .ZN(n8936) );
  AOI21_X1 U10334 ( .B1(n8938), .B2(n8937), .A(n8936), .ZN(n8943) );
  AOI22_X1 U10335 ( .A1(n7942), .A2(n8971), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8940) );
  NAND2_X1 U10336 ( .A1(n9524), .A2(n8984), .ZN(n8939) );
  OAI211_X1 U10337 ( .C1(n8966), .C2(n9503), .A(n8940), .B(n8939), .ZN(n8941)
         );
  AOI21_X1 U10338 ( .B1(n9648), .B2(n8978), .A(n8941), .ZN(n8942) );
  OAI21_X1 U10339 ( .B1(n8943), .B2(n8993), .A(n8942), .ZN(P1_U3231) );
  OAI21_X1 U10340 ( .B1(n8946), .B2(n8944), .A(n8823), .ZN(n8945) );
  OAI21_X1 U10341 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8948) );
  NAND2_X1 U10342 ( .A1(n8948), .A2(n8964), .ZN(n8955) );
  AOI21_X1 U10343 ( .B1(n8971), .B2(n9575), .A(n8949), .ZN(n8950) );
  OAI21_X1 U10344 ( .B1(n8951), .B2(n8968), .A(n8950), .ZN(n8952) );
  AOI21_X1 U10345 ( .B1(n8953), .B2(n8991), .A(n8952), .ZN(n8954) );
  OAI211_X1 U10346 ( .C1(n4910), .C2(n8988), .A(n8955), .B(n8954), .ZN(
        P1_U3232) );
  INV_X1 U10347 ( .A(n8956), .ZN(n8963) );
  NOR2_X1 U10348 ( .A1(n8959), .A2(n8958), .ZN(n8961) );
  OAI22_X1 U10349 ( .A1(n8963), .A2(n8962), .B1(n8961), .B2(n8960), .ZN(n8965)
         );
  NAND2_X1 U10350 ( .A1(n8965), .A2(n8964), .ZN(n8973) );
  NOR2_X1 U10351 ( .A1(n9465), .A2(n8966), .ZN(n8970) );
  OAI22_X1 U10352 ( .A1(n9500), .A2(n8968), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8967), .ZN(n8969) );
  AOI211_X1 U10353 ( .C1(n9462), .C2(n8971), .A(n8970), .B(n8969), .ZN(n8972)
         );
  OAI211_X1 U10354 ( .C1(n9468), .C2(n8988), .A(n8973), .B(n8972), .ZN(
        P1_U3233) );
  AOI22_X1 U10355 ( .A1(n9424), .A2(n8991), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8975) );
  NAND2_X1 U10356 ( .A1(n7972), .A2(n8984), .ZN(n8974) );
  OAI211_X1 U10357 ( .C1(n9390), .C2(n8986), .A(n8975), .B(n8974), .ZN(n8977)
         );
  INV_X1 U10358 ( .A(n8979), .ZN(n8981) );
  NAND2_X1 U10359 ( .A1(n8981), .A2(n8980), .ZN(n8983) );
  XNOR2_X1 U10360 ( .A(n8983), .B(n8982), .ZN(n8994) );
  NAND2_X1 U10361 ( .A1(n8984), .A2(n9575), .ZN(n8985) );
  NAND2_X1 U10362 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9304) );
  OAI211_X1 U10363 ( .C1(n8987), .C2(n8986), .A(n8985), .B(n9304), .ZN(n8990)
         );
  NOR2_X1 U10364 ( .A1(n9587), .A2(n8988), .ZN(n8989) );
  AOI211_X1 U10365 ( .C1(n9583), .C2(n8991), .A(n8990), .B(n8989), .ZN(n8992)
         );
  OAI21_X1 U10366 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(P1_U3239) );
  INV_X1 U10367 ( .A(n9184), .ZN(n9476) );
  NAND2_X1 U10368 ( .A1(n9148), .A2(n9476), .ZN(n8995) );
  AND2_X1 U10369 ( .A1(n9144), .A2(n8995), .ZN(n8996) );
  NAND2_X1 U10370 ( .A1(n8996), .A2(n9155), .ZN(n9149) );
  NOR2_X1 U10371 ( .A1(n9149), .A2(n4563), .ZN(n8997) );
  NAND2_X1 U10372 ( .A1(n8997), .A2(n9156), .ZN(n9028) );
  NAND2_X1 U10373 ( .A1(n9030), .A2(n9126), .ZN(n9071) );
  OR2_X1 U10374 ( .A1(n9071), .A2(n9129), .ZN(n9026) );
  NAND2_X1 U10375 ( .A1(n9122), .A2(n9114), .ZN(n9023) );
  INV_X1 U10376 ( .A(n8998), .ZN(n9001) );
  AND2_X1 U10377 ( .A1(n9093), .A2(n9090), .ZN(n9099) );
  INV_X1 U10378 ( .A(n8999), .ZN(n9000) );
  NOR2_X1 U10379 ( .A1(n9016), .A2(n9000), .ZN(n9112) );
  OAI211_X1 U10380 ( .C1(n5093), .C2(n9099), .A(n9112), .B(n9106), .ZN(n9020)
         );
  OR3_X1 U10381 ( .A1(n9023), .A2(n9001), .A3(n9020), .ZN(n9002) );
  OR3_X1 U10382 ( .A1(n9028), .A2(n9026), .A3(n9002), .ZN(n9245) );
  INV_X1 U10383 ( .A(n9245), .ZN(n9037) );
  AOI211_X1 U10384 ( .C1(n9821), .C2(n9285), .A(n9224), .B(n9003), .ZN(n9005)
         );
  OAI21_X1 U10385 ( .B1(n9006), .B2(n9005), .A(n9004), .ZN(n9008) );
  NAND3_X1 U10386 ( .A1(n9008), .A2(n9230), .A3(n9007), .ZN(n9010) );
  AND2_X1 U10387 ( .A1(n9009), .A2(n9231), .ZN(n9237) );
  NAND2_X1 U10388 ( .A1(n9010), .A2(n9237), .ZN(n9013) );
  NAND4_X1 U10389 ( .A1(n9013), .A2(n9012), .A3(n9239), .A4(n9011), .ZN(n9014)
         );
  NAND3_X1 U10390 ( .A1(n9014), .A2(n9242), .A3(n9236), .ZN(n9036) );
  AND2_X1 U10391 ( .A1(n9092), .A2(n9015), .ZN(n9096) );
  AND2_X1 U10392 ( .A1(n9096), .A2(n9101), .ZN(n9019) );
  NOR2_X1 U10393 ( .A1(n9017), .A2(n9016), .ZN(n9103) );
  NAND2_X1 U10394 ( .A1(n9103), .A2(n9106), .ZN(n9018) );
  OAI21_X1 U10395 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(n9022) );
  NAND2_X1 U10396 ( .A1(n9021), .A2(n9105), .ZN(n9115) );
  NOR2_X1 U10397 ( .A1(n9022), .A2(n9115), .ZN(n9024) );
  OAI211_X1 U10398 ( .C1(n9024), .C2(n9023), .A(n9130), .B(n9123), .ZN(n9025)
         );
  INV_X1 U10399 ( .A(n9025), .ZN(n9027) );
  OR3_X1 U10400 ( .A1(n9028), .A2(n9027), .A3(n9026), .ZN(n9035) );
  INV_X1 U10401 ( .A(n9128), .ZN(n9029) );
  AND2_X1 U10402 ( .A1(n9134), .A2(n9029), .ZN(n9069) );
  NAND2_X1 U10403 ( .A1(n9135), .A2(n9030), .ZN(n9137) );
  AND2_X1 U10404 ( .A1(n9185), .A2(n9133), .ZN(n9141) );
  OAI211_X1 U10405 ( .C1(n9069), .C2(n9137), .A(n9148), .B(n9141), .ZN(n9031)
         );
  INV_X1 U10406 ( .A(n9031), .ZN(n9032) );
  INV_X1 U10407 ( .A(n9183), .ZN(n9153) );
  OAI21_X1 U10408 ( .B1(n9149), .B2(n9032), .A(n9153), .ZN(n9033) );
  NAND2_X1 U10409 ( .A1(n9033), .A2(n9156), .ZN(n9034) );
  NAND4_X1 U10410 ( .A1(n9035), .A2(n9159), .A3(n9157), .A4(n9034), .ZN(n9246)
         );
  AOI21_X1 U10411 ( .B1(n9037), .B2(n9036), .A(n9246), .ZN(n9043) );
  NAND2_X1 U10412 ( .A1(n9062), .A2(n9163), .ZN(n9065) );
  INV_X1 U10413 ( .A(n9162), .ZN(n9038) );
  AND2_X1 U10414 ( .A1(n9249), .A2(n9038), .ZN(n9039) );
  INV_X1 U10415 ( .A(n9248), .ZN(n9041) );
  INV_X1 U10416 ( .A(n9068), .ZN(n9158) );
  AND2_X1 U10417 ( .A1(n9160), .A2(n9158), .ZN(n9146) );
  NAND2_X1 U10418 ( .A1(n9041), .A2(n9146), .ZN(n9251) );
  AOI21_X1 U10419 ( .B1(n9041), .B2(n9410), .A(n9254), .ZN(n9042) );
  NAND2_X1 U10420 ( .A1(n9044), .A2(n7087), .ZN(n9047) );
  OR2_X1 U10421 ( .A1(n4635), .A2(n9045), .ZN(n9046) );
  INV_X1 U10422 ( .A(n9272), .ZN(n9053) );
  NAND2_X1 U10423 ( .A1(n9383), .A2(n9053), .ZN(n9219) );
  NAND2_X1 U10424 ( .A1(n9048), .A2(n7087), .ZN(n9051) );
  OR2_X1 U10425 ( .A1(n4635), .A2(n6183), .ZN(n9050) );
  NAND2_X1 U10426 ( .A1(n9376), .A2(n9052), .ZN(n9179) );
  AND2_X1 U10427 ( .A1(n9179), .A2(n9175), .ZN(n9223) );
  AOI21_X1 U10428 ( .B1(n9054), .B2(n9223), .A(n9180), .ZN(n9268) );
  NOR2_X1 U10429 ( .A1(n9056), .A2(n9055), .ZN(n9059) );
  OAI21_X1 U10430 ( .B1(n9057), .B2(n9265), .A(P1_B_REG_SCAN_IN), .ZN(n9058)
         );
  AOI21_X1 U10431 ( .B1(n9060), .B2(n9059), .A(n9058), .ZN(n9269) );
  NOR4_X1 U10432 ( .A1(n9268), .A2(n9261), .A3(n9263), .A4(n9269), .ZN(n9271)
         );
  INV_X1 U10433 ( .A(n9170), .ZN(n9177) );
  INV_X1 U10434 ( .A(n9061), .ZN(n9221) );
  NAND2_X1 U10435 ( .A1(n9064), .A2(n9249), .ZN(n9063) );
  NAND2_X1 U10436 ( .A1(n9063), .A2(n9062), .ZN(n9067) );
  NAND2_X1 U10437 ( .A1(n9065), .A2(n9064), .ZN(n9066) );
  MUX2_X1 U10438 ( .A(n9067), .B(n9066), .S(n9177), .Z(n9169) );
  OAI211_X1 U10439 ( .C1(n9068), .C2(n9157), .A(n9419), .B(n9159), .ZN(n9147)
         );
  INV_X1 U10440 ( .A(n9069), .ZN(n9070) );
  MUX2_X1 U10441 ( .A(n9071), .B(n9070), .S(n9177), .Z(n9072) );
  INV_X1 U10442 ( .A(n9072), .ZN(n9132) );
  NAND3_X1 U10443 ( .A1(n9073), .A2(n9177), .A3(n9239), .ZN(n9074) );
  AOI21_X1 U10444 ( .B1(n9075), .B2(n9232), .A(n9074), .ZN(n9089) );
  NAND2_X1 U10445 ( .A1(n9079), .A2(n9170), .ZN(n9078) );
  INV_X1 U10446 ( .A(n9078), .ZN(n9076) );
  AOI22_X1 U10447 ( .A1(n9076), .A2(n9081), .B1(n9170), .B2(n9080), .ZN(n9088)
         );
  OAI21_X1 U10448 ( .B1(n9078), .B2(n9280), .A(n9081), .ZN(n9085) );
  OR2_X1 U10449 ( .A1(n9079), .A2(n9170), .ZN(n9082) );
  OAI21_X1 U10450 ( .B1(n9082), .B2(n9080), .A(n9851), .ZN(n9084) );
  OAI22_X1 U10451 ( .A1(n9082), .A2(n9081), .B1(n9170), .B2(n9080), .ZN(n9083)
         );
  AOI22_X1 U10452 ( .A1(n9085), .A2(n9084), .B1(n9083), .B2(n9859), .ZN(n9086)
         );
  INV_X1 U10453 ( .A(n9095), .ZN(n9097) );
  OAI21_X1 U10454 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(n9100) );
  INV_X1 U10455 ( .A(n9103), .ZN(n9104) );
  AND2_X1 U10456 ( .A1(n9114), .A2(n9106), .ZN(n9111) );
  AOI21_X1 U10457 ( .B1(n9108), .B2(n9111), .A(n9107), .ZN(n9121) );
  INV_X1 U10458 ( .A(n9109), .ZN(n9119) );
  INV_X1 U10459 ( .A(n9110), .ZN(n9113) );
  OAI21_X1 U10460 ( .B1(n9113), .B2(n9112), .A(n9111), .ZN(n9118) );
  INV_X1 U10461 ( .A(n9114), .ZN(n9117) );
  INV_X1 U10462 ( .A(n9115), .ZN(n9116) );
  OAI22_X1 U10463 ( .A1(n9119), .A2(n9118), .B1(n9117), .B2(n9116), .ZN(n9120)
         );
  MUX2_X1 U10464 ( .A(n9121), .B(n9120), .S(n9170), .Z(n9125) );
  INV_X1 U10465 ( .A(n9571), .ZN(n9567) );
  MUX2_X1 U10466 ( .A(n9123), .B(n9122), .S(n9170), .Z(n9124) );
  INV_X1 U10467 ( .A(n9126), .ZN(n9127) );
  INV_X1 U10468 ( .A(n9546), .ZN(n9211) );
  MUX2_X1 U10469 ( .A(n7953), .B(n9130), .S(n9170), .Z(n9131) );
  NAND3_X1 U10470 ( .A1(n9136), .A2(n9135), .A3(n9184), .ZN(n9143) );
  INV_X1 U10471 ( .A(n9137), .ZN(n9138) );
  NAND2_X1 U10472 ( .A1(n9139), .A2(n9138), .ZN(n9140) );
  NAND2_X1 U10473 ( .A1(n9141), .A2(n9140), .ZN(n9142) );
  NAND3_X1 U10474 ( .A1(n9152), .A2(n9185), .A3(n9148), .ZN(n9145) );
  INV_X1 U10475 ( .A(n9148), .ZN(n9151) );
  INV_X1 U10476 ( .A(n9149), .ZN(n9150) );
  OAI21_X1 U10477 ( .B1(n9152), .B2(n9151), .A(n9150), .ZN(n9154) );
  NAND2_X1 U10478 ( .A1(n9157), .A2(n9156), .ZN(n9214) );
  MUX2_X1 U10479 ( .A(n9160), .B(n9419), .S(n9170), .Z(n9161) );
  AND2_X1 U10480 ( .A1(n9163), .A2(n9162), .ZN(n9164) );
  MUX2_X1 U10481 ( .A(n9165), .B(n9164), .S(n9170), .Z(n9166) );
  NAND3_X1 U10482 ( .A1(n9221), .A2(n9169), .A3(n9168), .ZN(n9174) );
  MUX2_X1 U10483 ( .A(n9171), .B(n9253), .S(n9170), .Z(n9173) );
  NAND2_X1 U10484 ( .A1(n9378), .A2(n9272), .ZN(n9172) );
  NAND2_X1 U10485 ( .A1(n9383), .A2(n9172), .ZN(n9252) );
  NAND2_X1 U10486 ( .A1(n9175), .A2(n9378), .ZN(n9176) );
  NAND2_X1 U10487 ( .A1(n9176), .A2(n9376), .ZN(n9256) );
  INV_X1 U10488 ( .A(n9252), .ZN(n9178) );
  NAND3_X1 U10489 ( .A1(n9179), .A2(n9178), .A3(n9177), .ZN(n9181) );
  AND2_X1 U10490 ( .A1(n9181), .A2(n9258), .ZN(n9182) );
  NOR2_X1 U10491 ( .A1(n9183), .A2(n5103), .ZN(n9469) );
  INV_X1 U10492 ( .A(n9475), .ZN(n9477) );
  INV_X1 U10493 ( .A(n9186), .ZN(n9204) );
  INV_X1 U10494 ( .A(n9187), .ZN(n9198) );
  NOR2_X1 U10495 ( .A1(n9189), .A2(n9188), .ZN(n9193) );
  NAND4_X1 U10496 ( .A1(n9193), .A2(n9192), .A3(n9191), .A4(n9190), .ZN(n9196)
         );
  NOR3_X1 U10497 ( .A1(n9196), .A2(n9195), .A3(n9194), .ZN(n9197) );
  NAND4_X1 U10498 ( .A1(n9200), .A2(n9199), .A3(n9198), .A4(n9197), .ZN(n9201)
         );
  NOR2_X1 U10499 ( .A1(n7359), .A2(n9201), .ZN(n9202) );
  NAND3_X1 U10500 ( .A1(n9204), .A2(n9203), .A3(n9202), .ZN(n9205) );
  NOR2_X1 U10501 ( .A1(n9206), .A2(n9205), .ZN(n9207) );
  NAND3_X1 U10502 ( .A1(n9571), .A2(n9208), .A3(n9207), .ZN(n9209) );
  NOR2_X1 U10503 ( .A1(n9561), .A2(n9209), .ZN(n9210) );
  NAND3_X1 U10504 ( .A1(n9535), .A2(n9211), .A3(n9210), .ZN(n9212) );
  NOR2_X1 U10505 ( .A1(n9518), .A2(n9212), .ZN(n9213) );
  NAND4_X1 U10506 ( .A1(n9469), .A2(n9477), .A3(n9495), .A4(n9213), .ZN(n9215)
         );
  NOR2_X1 U10507 ( .A1(n9215), .A2(n9214), .ZN(n9217) );
  NAND4_X1 U10508 ( .A1(n9426), .A2(n4941), .A3(n9217), .A4(n9216), .ZN(n9218)
         );
  NOR2_X1 U10509 ( .A1(n9410), .A2(n9218), .ZN(n9220) );
  AND4_X1 U10510 ( .A1(n9221), .A2(n9388), .A3(n9220), .A4(n9219), .ZN(n9222)
         );
  NAND3_X1 U10511 ( .A1(n9223), .A2(n9222), .A3(n9258), .ZN(n9225) );
  NAND2_X1 U10512 ( .A1(n9225), .A2(n9224), .ZN(n9260) );
  AND3_X1 U10513 ( .A1(n9258), .A2(n9259), .A3(n9227), .ZN(n9228) );
  INV_X1 U10514 ( .A(n9230), .ZN(n9233) );
  AND3_X1 U10515 ( .A1(n9233), .A2(n9232), .A3(n9231), .ZN(n9234) );
  NAND3_X1 U10516 ( .A1(n9238), .A2(n9237), .A3(n9236), .ZN(n9240) );
  NAND3_X1 U10517 ( .A1(n9241), .A2(n9240), .A3(n9239), .ZN(n9243) );
  AND2_X1 U10518 ( .A1(n9243), .A2(n9242), .ZN(n9244) );
  NOR2_X1 U10519 ( .A1(n9245), .A2(n9244), .ZN(n9247) );
  NOR2_X1 U10520 ( .A1(n9247), .A2(n9246), .ZN(n9250) );
  OAI22_X1 U10521 ( .A1(n9251), .A2(n9250), .B1(n9249), .B2(n9248), .ZN(n9255)
         );
  OAI211_X1 U10522 ( .C1(n9255), .C2(n9254), .A(n9253), .B(n9252), .ZN(n9257)
         );
  NAND3_X1 U10523 ( .A1(n9262), .A2(n9261), .A3(n9260), .ZN(n9264) );
  INV_X1 U10524 ( .A(n9269), .ZN(n9266) );
  MUX2_X1 U10525 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9272), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10526 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9273), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10527 ( .A(n9422), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9274), .Z(
        P1_U3582) );
  MUX2_X1 U10528 ( .A(n9433), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9274), .Z(
        P1_U3581) );
  MUX2_X1 U10529 ( .A(n7972), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9274), .Z(
        P1_U3580) );
  MUX2_X1 U10530 ( .A(n9448), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9274), .Z(
        P1_U3579) );
  MUX2_X1 U10531 ( .A(n9462), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9274), .Z(
        P1_U3578) );
  MUX2_X1 U10532 ( .A(n9447), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9274), .Z(
        P1_U3577) );
  MUX2_X1 U10533 ( .A(n7942), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9274), .Z(
        P1_U3576) );
  MUX2_X1 U10534 ( .A(n9511), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9274), .Z(
        P1_U3575) );
  MUX2_X1 U10535 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9524), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10536 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n7932), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10537 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9553), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10538 ( .A(n9573), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9274), .Z(
        P1_U3571) );
  MUX2_X1 U10539 ( .A(n9552), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9274), .Z(
        P1_U3570) );
  MUX2_X1 U10540 ( .A(n9575), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9274), .Z(
        P1_U3569) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9275), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10542 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n7309), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10543 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9276), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9277), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9278), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10546 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9279), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9280), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10548 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n4928), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10549 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9281), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10550 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9282), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10551 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9283), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10552 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9284), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10553 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9285), .S(P1_U4006), .Z(
        P1_U3556) );
  XNOR2_X1 U10554 ( .A(n9294), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9289) );
  OAI21_X1 U10555 ( .B1(n9289), .B2(n9288), .A(n9310), .ZN(n9302) );
  NAND2_X1 U10556 ( .A1(n9375), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n9291) );
  OAI211_X1 U10557 ( .C1(n9791), .C2(n9294), .A(n9291), .B(n9290), .ZN(n9301)
         );
  INV_X1 U10558 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9299) );
  AOI211_X1 U10559 ( .C1(n9299), .C2(n9298), .A(n9799), .B(n9306), .ZN(n9300)
         );
  AOI211_X1 U10560 ( .C1(n9790), .C2(n9302), .A(n9301), .B(n9300), .ZN(n9303)
         );
  INV_X1 U10561 ( .A(n9303), .ZN(P1_U3255) );
  NAND2_X1 U10562 ( .A1(n9375), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n9305) );
  OAI211_X1 U10563 ( .C1(n9791), .C2(n9323), .A(n9305), .B(n9304), .ZN(n9316)
         );
  INV_X1 U10564 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9308) );
  AOI211_X1 U10565 ( .C1(n9309), .C2(n9308), .A(n9318), .B(n9799), .ZN(n9315)
         );
  INV_X1 U10566 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9312) );
  NOR2_X1 U10567 ( .A1(n9312), .A2(n9313), .ZN(n9324) );
  AOI211_X1 U10568 ( .C1(n9313), .C2(n9312), .A(n9324), .B(n9807), .ZN(n9314)
         );
  OR3_X1 U10569 ( .A1(n9316), .A2(n9315), .A3(n9314), .ZN(P1_U3256) );
  NAND2_X1 U10570 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9340), .ZN(n9320) );
  OAI21_X1 U10571 ( .B1(n9340), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9320), .ZN(
        n9321) );
  AOI211_X1 U10572 ( .C1(n4305), .C2(n9321), .A(n9334), .B(n9799), .ZN(n9333)
         );
  NOR2_X1 U10573 ( .A1(n9323), .A2(n9322), .ZN(n9325) );
  XNOR2_X1 U10574 ( .A(n9340), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9326) );
  AOI211_X1 U10575 ( .C1(n9327), .C2(n9326), .A(n9339), .B(n9807), .ZN(n9332)
         );
  NAND2_X1 U10576 ( .A1(n9375), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9329) );
  OAI211_X1 U10577 ( .C1(n9791), .C2(n9330), .A(n9329), .B(n9328), .ZN(n9331)
         );
  OR3_X1 U10578 ( .A1(n9333), .A2(n9332), .A3(n9331), .ZN(P1_U3257) );
  INV_X1 U10579 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U10580 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9355), .ZN(n9335) );
  OAI21_X1 U10581 ( .B1(n9355), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9335), .ZN(
        n9336) );
  AOI211_X1 U10582 ( .C1(n9337), .C2(n9336), .A(n9349), .B(n9799), .ZN(n9338)
         );
  AOI21_X1 U10583 ( .B1(n9369), .B2(n9355), .A(n9338), .ZN(n9347) );
  XNOR2_X1 U10584 ( .A(n9355), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9341) );
  AOI211_X1 U10585 ( .C1(n9342), .C2(n9341), .A(n9354), .B(n9807), .ZN(n9345)
         );
  INV_X1 U10586 ( .A(n9343), .ZN(n9344) );
  NOR2_X1 U10587 ( .A1(n9345), .A2(n9344), .ZN(n9346) );
  OAI211_X1 U10588 ( .C1(n9813), .C2(n9348), .A(n9347), .B(n9346), .ZN(
        P1_U3258) );
  INV_X1 U10589 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U10590 ( .A1(n9367), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9350) );
  OAI21_X1 U10591 ( .B1(n9367), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9350), .ZN(
        n9351) );
  AOI211_X1 U10592 ( .C1(n9352), .C2(n9351), .A(n9364), .B(n9799), .ZN(n9353)
         );
  AOI21_X1 U10593 ( .B1(n9369), .B2(n9367), .A(n9353), .ZN(n9362) );
  XOR2_X1 U10594 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9367), .Z(n9357) );
  NAND2_X1 U10595 ( .A1(n9357), .A2(n9356), .ZN(n9366) );
  OAI21_X1 U10596 ( .B1(n9357), .B2(n9356), .A(n9366), .ZN(n9360) );
  INV_X1 U10597 ( .A(n9358), .ZN(n9359) );
  AOI21_X1 U10598 ( .B1(n9790), .B2(n9360), .A(n9359), .ZN(n9361) );
  OAI211_X1 U10599 ( .C1(n9813), .C2(n9363), .A(n9362), .B(n9361), .ZN(
        P1_U3259) );
  INV_X1 U10600 ( .A(n9368), .ZN(n9372) );
  AOI21_X1 U10601 ( .B1(n9370), .B2(n9790), .A(n9369), .ZN(n9371) );
  NOR2_X2 U10602 ( .A1(n9382), .A2(n9383), .ZN(n9381) );
  XNOR2_X1 U10603 ( .A(n9376), .B(n9381), .ZN(n9593) );
  NAND2_X1 U10604 ( .A1(n9593), .A2(n9581), .ZN(n9380) );
  NAND2_X1 U10605 ( .A1(n9378), .A2(n9377), .ZN(n9597) );
  NOR2_X1 U10606 ( .A1(n9566), .A2(n9597), .ZN(n9384) );
  AOI21_X1 U10607 ( .B1(n9566), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9384), .ZN(
        n9379) );
  OAI211_X1 U10608 ( .C1(n9595), .C2(n9586), .A(n9380), .B(n9379), .ZN(
        P1_U3261) );
  INV_X1 U10609 ( .A(n9383), .ZN(n9599) );
  AOI21_X1 U10610 ( .B1(n9383), .B2(n9382), .A(n9381), .ZN(n9596) );
  NAND2_X1 U10611 ( .A1(n9596), .A2(n9581), .ZN(n9386) );
  AOI21_X1 U10612 ( .B1(n9566), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9384), .ZN(
        n9385) );
  OAI211_X1 U10613 ( .C1(n9599), .C2(n9586), .A(n9386), .B(n9385), .ZN(
        P1_U3262) );
  OAI21_X1 U10614 ( .B1(n9389), .B2(n9388), .A(n9387), .ZN(n9393) );
  OAI22_X1 U10615 ( .A1(n9391), .A2(n9501), .B1(n9390), .B2(n9499), .ZN(n9392)
         );
  AOI21_X1 U10616 ( .B1(n9606), .B2(n9404), .A(n9394), .ZN(n9607) );
  INV_X1 U10617 ( .A(n9606), .ZN(n9397) );
  AOI22_X1 U10618 ( .A1(n9395), .A2(n9582), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9566), .ZN(n9396) );
  OAI21_X1 U10619 ( .B1(n9397), .B2(n9586), .A(n9396), .ZN(n9401) );
  NOR2_X1 U10620 ( .A1(n9610), .A2(n9592), .ZN(n9400) );
  OAI21_X1 U10621 ( .B1(n9609), .B2(n9566), .A(n9402), .ZN(P1_U3263) );
  XNOR2_X1 U10622 ( .A(n9403), .B(n9410), .ZN(n9615) );
  INV_X1 U10623 ( .A(n9423), .ZN(n9406) );
  INV_X1 U10624 ( .A(n9404), .ZN(n9405) );
  AOI211_X1 U10625 ( .C1(n9612), .C2(n9406), .A(n9869), .B(n9405), .ZN(n9611)
         );
  AOI22_X1 U10626 ( .A1(n9407), .A2(n9582), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9566), .ZN(n9408) );
  OAI21_X1 U10627 ( .B1(n9409), .B2(n9586), .A(n9408), .ZN(n9417) );
  AOI21_X1 U10628 ( .B1(n9411), .B2(n9410), .A(n9496), .ZN(n9416) );
  OAI22_X1 U10629 ( .A1(n9413), .A2(n9501), .B1(n9412), .B2(n9499), .ZN(n9414)
         );
  OAI21_X1 U10630 ( .B1(n9592), .B2(n9615), .A(n9418), .ZN(P1_U3264) );
  NAND2_X1 U10631 ( .A1(n9420), .A2(n9419), .ZN(n9421) );
  AOI21_X1 U10632 ( .B1(n9616), .B2(n9436), .A(n9423), .ZN(n9617) );
  AOI22_X1 U10633 ( .A1(n9424), .A2(n9582), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9566), .ZN(n9425) );
  OAI21_X1 U10634 ( .B1(n4925), .B2(n9586), .A(n9425), .ZN(n9429) );
  XNOR2_X1 U10635 ( .A(n9427), .B(n9426), .ZN(n9620) );
  NOR2_X1 U10636 ( .A1(n9620), .A2(n9592), .ZN(n9428) );
  AOI211_X1 U10637 ( .C1(n9617), .C2(n9581), .A(n9429), .B(n9428), .ZN(n9430)
         );
  OAI21_X1 U10638 ( .B1(n9619), .B2(n9566), .A(n9430), .ZN(P1_U3265) );
  XNOR2_X1 U10639 ( .A(n9432), .B(n9431), .ZN(n9434) );
  AOI222_X1 U10640 ( .A1(n9577), .A2(n9434), .B1(n9448), .B2(n9574), .C1(n9433), .C2(n9572), .ZN(n9624) );
  INV_X1 U10641 ( .A(n9435), .ZN(n9438) );
  INV_X1 U10642 ( .A(n9436), .ZN(n9437) );
  AOI211_X1 U10643 ( .C1(n9622), .C2(n9438), .A(n9869), .B(n9437), .ZN(n9621)
         );
  AOI22_X1 U10644 ( .A1(n9439), .A2(n9582), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9566), .ZN(n9440) );
  OAI21_X1 U10645 ( .B1(n9441), .B2(n9586), .A(n9440), .ZN(n9444) );
  XNOR2_X1 U10646 ( .A(n9442), .B(n4941), .ZN(n9625) );
  NOR2_X1 U10647 ( .A1(n9625), .A2(n9592), .ZN(n9443) );
  AOI211_X1 U10648 ( .C1(n9621), .C2(n9564), .A(n9444), .B(n9443), .ZN(n9445)
         );
  OAI21_X1 U10649 ( .B1(n9624), .B2(n9566), .A(n9445), .ZN(P1_U3266) );
  XNOR2_X1 U10650 ( .A(n9446), .B(n9456), .ZN(n9449) );
  AOI222_X1 U10651 ( .A1(n9577), .A2(n9449), .B1(n9448), .B2(n9572), .C1(n9447), .C2(n9574), .ZN(n9634) );
  INV_X1 U10652 ( .A(n9464), .ZN(n9452) );
  INV_X1 U10653 ( .A(n9450), .ZN(n9451) );
  AOI21_X1 U10654 ( .B1(n9631), .B2(n9452), .A(n9451), .ZN(n9632) );
  AOI22_X1 U10655 ( .A1(n9453), .A2(n9582), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9566), .ZN(n9454) );
  OAI21_X1 U10656 ( .B1(n9455), .B2(n9586), .A(n9454), .ZN(n9459) );
  XNOR2_X1 U10657 ( .A(n9457), .B(n9456), .ZN(n9635) );
  NOR2_X1 U10658 ( .A1(n9635), .A2(n9592), .ZN(n9458) );
  AOI211_X1 U10659 ( .C1(n9632), .C2(n9581), .A(n9459), .B(n9458), .ZN(n9460)
         );
  OAI21_X1 U10660 ( .B1(n9634), .B2(n9566), .A(n9460), .ZN(P1_U3268) );
  XOR2_X1 U10661 ( .A(n9461), .B(n9469), .Z(n9463) );
  AOI222_X1 U10662 ( .A1(n9577), .A2(n9463), .B1(n9462), .B2(n9572), .C1(n7942), .C2(n9574), .ZN(n9639) );
  AOI21_X1 U10663 ( .B1(n9636), .B2(n9484), .A(n9464), .ZN(n9637) );
  INV_X1 U10664 ( .A(n9465), .ZN(n9466) );
  AOI22_X1 U10665 ( .A1(n9466), .A2(n9582), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9566), .ZN(n9467) );
  OAI21_X1 U10666 ( .B1(n9468), .B2(n9586), .A(n9467), .ZN(n9472) );
  XOR2_X1 U10667 ( .A(n9470), .B(n9469), .Z(n9640) );
  NOR2_X1 U10668 ( .A1(n9640), .A2(n9592), .ZN(n9471) );
  AOI211_X1 U10669 ( .C1(n9637), .C2(n9581), .A(n9472), .B(n9471), .ZN(n9473)
         );
  OAI21_X1 U10670 ( .B1(n9639), .B2(n9566), .A(n9473), .ZN(P1_U3269) );
  XNOR2_X1 U10671 ( .A(n9475), .B(n9474), .ZN(n9645) );
  NOR2_X1 U10672 ( .A1(n9477), .A2(n9476), .ZN(n9480) );
  AOI21_X1 U10673 ( .B1(n9480), .B2(n9479), .A(n9478), .ZN(n9481) );
  OAI222_X1 U10674 ( .A1(n9499), .A2(n9483), .B1(n9501), .B2(n9482), .C1(n9496), .C2(n9481), .ZN(n9641) );
  INV_X1 U10675 ( .A(n9502), .ZN(n9486) );
  INV_X1 U10676 ( .A(n9484), .ZN(n9485) );
  AOI211_X1 U10677 ( .C1(n9643), .C2(n9486), .A(n9869), .B(n9485), .ZN(n9642)
         );
  INV_X1 U10678 ( .A(n9642), .ZN(n9488) );
  OAI22_X1 U10679 ( .A1(n9488), .A2(n4259), .B1(n9487), .B2(n9530), .ZN(n9489)
         );
  OAI21_X1 U10680 ( .B1(n9641), .B2(n9489), .A(n9589), .ZN(n9492) );
  AOI22_X1 U10681 ( .A1(n9643), .A2(n9490), .B1(n9566), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9491) );
  OAI211_X1 U10682 ( .C1(n9645), .C2(n9592), .A(n9492), .B(n9491), .ZN(
        P1_U3270) );
  XOR2_X1 U10683 ( .A(n9493), .B(n9495), .Z(n9650) );
  XOR2_X1 U10684 ( .A(n9495), .B(n9494), .Z(n9497) );
  OAI222_X1 U10685 ( .A1(n9501), .A2(n9500), .B1(n9499), .B2(n9498), .C1(n9497), .C2(n9496), .ZN(n9646) );
  NAND2_X1 U10686 ( .A1(n9646), .A2(n9589), .ZN(n9509) );
  AOI211_X1 U10687 ( .C1(n9648), .C2(n9513), .A(n9869), .B(n9502), .ZN(n9647)
         );
  INV_X1 U10688 ( .A(n9648), .ZN(n9506) );
  INV_X1 U10689 ( .A(n9503), .ZN(n9504) );
  AOI22_X1 U10690 ( .A1(n9504), .A2(n9582), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9566), .ZN(n9505) );
  OAI21_X1 U10691 ( .B1(n9506), .B2(n9586), .A(n9505), .ZN(n9507) );
  AOI21_X1 U10692 ( .B1(n9647), .B2(n9564), .A(n9507), .ZN(n9508) );
  OAI211_X1 U10693 ( .C1(n9650), .C2(n9592), .A(n9509), .B(n9508), .ZN(
        P1_U3271) );
  XNOR2_X1 U10694 ( .A(n9510), .B(n9518), .ZN(n9512) );
  AOI222_X1 U10695 ( .A1(n9577), .A2(n9512), .B1(n7932), .B2(n9574), .C1(n9511), .C2(n9572), .ZN(n9654) );
  INV_X1 U10696 ( .A(n9526), .ZN(n9514) );
  AOI21_X1 U10697 ( .B1(n9651), .B2(n9514), .A(n4917), .ZN(n9652) );
  AOI22_X1 U10698 ( .A1(n9515), .A2(n9582), .B1(P1_REG2_REG_19__SCAN_IN), .B2(
        n9566), .ZN(n9516) );
  OAI21_X1 U10699 ( .B1(n9517), .B2(n9586), .A(n9516), .ZN(n9521) );
  XNOR2_X1 U10700 ( .A(n9519), .B(n9518), .ZN(n9655) );
  NOR2_X1 U10701 ( .A1(n9655), .A2(n9592), .ZN(n9520) );
  AOI211_X1 U10702 ( .C1(n9652), .C2(n9581), .A(n9521), .B(n9520), .ZN(n9522)
         );
  OAI21_X1 U10703 ( .B1(n9654), .B2(n9566), .A(n9522), .ZN(P1_U3272) );
  XNOR2_X1 U10704 ( .A(n9523), .B(n9535), .ZN(n9525) );
  AOI222_X1 U10705 ( .A1(n9577), .A2(n9525), .B1(n9553), .B2(n9574), .C1(n9524), .C2(n9572), .ZN(n9661) );
  NOR2_X1 U10706 ( .A1(n9528), .A2(n9542), .ZN(n9527) );
  NOR2_X1 U10707 ( .A1(n9527), .A2(n9526), .ZN(n9657) );
  NOR2_X1 U10708 ( .A1(n9528), .A2(n9586), .ZN(n9533) );
  INV_X1 U10709 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9529) );
  OAI22_X1 U10710 ( .A1(n9531), .A2(n9530), .B1(n9529), .B2(n9589), .ZN(n9532)
         );
  AOI211_X1 U10711 ( .C1(n9657), .C2(n9581), .A(n9533), .B(n9532), .ZN(n9539)
         );
  NAND2_X1 U10712 ( .A1(n9536), .A2(n9535), .ZN(n9658) );
  NAND3_X1 U10713 ( .A1(n9534), .A2(n9658), .A3(n9537), .ZN(n9538) );
  OAI211_X1 U10714 ( .C1(n9661), .C2(n9566), .A(n9539), .B(n9538), .ZN(
        P1_U3273) );
  XNOR2_X1 U10715 ( .A(n9540), .B(n9546), .ZN(n9541) );
  AOI222_X1 U10716 ( .A1(n9577), .A2(n9541), .B1(n7932), .B2(n9572), .C1(n9573), .C2(n9574), .ZN(n9665) );
  AOI211_X1 U10717 ( .C1(n9663), .C2(n5125), .A(n9869), .B(n9542), .ZN(n9662)
         );
  INV_X1 U10718 ( .A(n9663), .ZN(n9545) );
  AOI22_X1 U10719 ( .A1(n9566), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9543), .B2(
        n9582), .ZN(n9544) );
  OAI21_X1 U10720 ( .B1(n9545), .B2(n9586), .A(n9544), .ZN(n9549) );
  XNOR2_X1 U10721 ( .A(n9547), .B(n9546), .ZN(n9666) );
  NOR2_X1 U10722 ( .A1(n9666), .A2(n9592), .ZN(n9548) );
  AOI211_X1 U10723 ( .C1(n9662), .C2(n9564), .A(n9549), .B(n9548), .ZN(n9550)
         );
  OAI21_X1 U10724 ( .B1(n9665), .B2(n9566), .A(n9550), .ZN(P1_U3274) );
  XNOR2_X1 U10725 ( .A(n9551), .B(n4426), .ZN(n9554) );
  AOI222_X1 U10726 ( .A1(n9577), .A2(n9554), .B1(n9553), .B2(n9572), .C1(n9552), .C2(n9574), .ZN(n9670) );
  INV_X1 U10727 ( .A(n5125), .ZN(n9555) );
  AOI211_X1 U10728 ( .C1(n9668), .C2(n9579), .A(n9869), .B(n9555), .ZN(n9667)
         );
  INV_X1 U10729 ( .A(n9556), .ZN(n9557) );
  AOI22_X1 U10730 ( .A1(n9566), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9557), .B2(
        n9582), .ZN(n9558) );
  OAI21_X1 U10731 ( .B1(n9559), .B2(n9586), .A(n9558), .ZN(n9563) );
  XNOR2_X1 U10732 ( .A(n9560), .B(n9561), .ZN(n9671) );
  NOR2_X1 U10733 ( .A1(n9671), .A2(n9592), .ZN(n9562) );
  AOI211_X1 U10734 ( .C1(n9667), .C2(n9564), .A(n9563), .B(n9562), .ZN(n9565)
         );
  OAI21_X1 U10735 ( .B1(n9670), .B2(n9566), .A(n9565), .ZN(P1_U3275) );
  XNOR2_X1 U10736 ( .A(n9568), .B(n9567), .ZN(n9676) );
  OAI21_X1 U10737 ( .B1(n9571), .B2(n9570), .A(n9569), .ZN(n9576) );
  AOI222_X1 U10738 ( .A1(n9577), .A2(n9576), .B1(n9575), .B2(n9574), .C1(n9573), .C2(n9572), .ZN(n9675) );
  INV_X1 U10739 ( .A(n9675), .ZN(n9590) );
  OR2_X1 U10740 ( .A1(n9578), .A2(n9587), .ZN(n9580) );
  AND2_X1 U10741 ( .A1(n9580), .A2(n9579), .ZN(n9673) );
  NAND2_X1 U10742 ( .A1(n9673), .A2(n9581), .ZN(n9585) );
  AOI22_X1 U10743 ( .A1(n9566), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9583), .B2(
        n9582), .ZN(n9584) );
  OAI211_X1 U10744 ( .C1(n9587), .C2(n9586), .A(n9585), .B(n9584), .ZN(n9588)
         );
  AOI21_X1 U10745 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9591) );
  OAI21_X1 U10746 ( .B1(n9592), .B2(n9676), .A(n9591), .ZN(P1_U3276) );
  NAND2_X1 U10747 ( .A1(n9593), .A2(n9835), .ZN(n9594) );
  OAI211_X1 U10748 ( .C1(n9595), .C2(n9868), .A(n9594), .B(n9597), .ZN(n9705)
         );
  MUX2_X1 U10749 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9705), .S(n9891), .Z(
        P1_U3554) );
  NAND2_X1 U10750 ( .A1(n9596), .A2(n9835), .ZN(n9598) );
  OAI211_X1 U10751 ( .C1(n9599), .C2(n9868), .A(n9598), .B(n9597), .ZN(n9706)
         );
  MUX2_X1 U10752 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9706), .S(n9891), .Z(
        P1_U3553) );
  INV_X1 U10753 ( .A(n9856), .ZN(n9839) );
  OAI22_X1 U10754 ( .A1(n9604), .A2(n9869), .B1(n9603), .B2(n9868), .ZN(n9605)
         );
  AOI22_X1 U10755 ( .A1(n9607), .A2(n9835), .B1(n9834), .B2(n9606), .ZN(n9608)
         );
  MUX2_X1 U10756 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9708), .S(n9891), .Z(
        P1_U3551) );
  AOI21_X1 U10757 ( .B1(n9834), .B2(n9612), .A(n9611), .ZN(n9613) );
  OAI211_X1 U10758 ( .C1(n9697), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9709)
         );
  MUX2_X1 U10759 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9709), .S(n9891), .Z(
        P1_U3550) );
  AOI22_X1 U10760 ( .A1(n9617), .A2(n9835), .B1(n9834), .B2(n9616), .ZN(n9618)
         );
  OAI211_X1 U10761 ( .C1(n9697), .C2(n9620), .A(n9619), .B(n9618), .ZN(n9710)
         );
  MUX2_X1 U10762 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9710), .S(n9891), .Z(
        P1_U3549) );
  AOI21_X1 U10763 ( .B1(n9834), .B2(n9622), .A(n9621), .ZN(n9623) );
  OAI211_X1 U10764 ( .C1(n9697), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9711)
         );
  MUX2_X1 U10765 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9711), .S(n9891), .Z(
        P1_U3548) );
  OAI21_X1 U10766 ( .B1(n9697), .B2(n9630), .A(n9629), .ZN(n9712) );
  MUX2_X1 U10767 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9712), .S(n9891), .Z(
        P1_U3547) );
  AOI22_X1 U10768 ( .A1(n9632), .A2(n9835), .B1(n9834), .B2(n9631), .ZN(n9633)
         );
  OAI211_X1 U10769 ( .C1(n9697), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9713)
         );
  MUX2_X1 U10770 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9713), .S(n9891), .Z(
        P1_U3546) );
  AOI22_X1 U10771 ( .A1(n9637), .A2(n9835), .B1(n9834), .B2(n9636), .ZN(n9638)
         );
  OAI211_X1 U10772 ( .C1(n9697), .C2(n9640), .A(n9639), .B(n9638), .ZN(n9714)
         );
  MUX2_X1 U10773 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9714), .S(n9891), .Z(
        P1_U3545) );
  AOI211_X1 U10774 ( .C1(n9834), .C2(n9643), .A(n9642), .B(n9641), .ZN(n9644)
         );
  OAI21_X1 U10775 ( .B1(n9697), .B2(n9645), .A(n9644), .ZN(n9715) );
  MUX2_X1 U10776 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9715), .S(n9891), .Z(
        P1_U3544) );
  AOI211_X1 U10777 ( .C1(n9834), .C2(n9648), .A(n9647), .B(n9646), .ZN(n9649)
         );
  OAI21_X1 U10778 ( .B1(n9697), .B2(n9650), .A(n9649), .ZN(n9716) );
  MUX2_X1 U10779 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9716), .S(n9891), .Z(
        P1_U3543) );
  AOI22_X1 U10780 ( .A1(n9652), .A2(n9835), .B1(n9834), .B2(n9651), .ZN(n9653)
         );
  OAI211_X1 U10781 ( .C1(n9697), .C2(n9655), .A(n9654), .B(n9653), .ZN(n9717)
         );
  MUX2_X1 U10782 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9717), .S(n9891), .Z(
        P1_U3542) );
  AOI22_X1 U10783 ( .A1(n9657), .A2(n9835), .B1(n9834), .B2(n9656), .ZN(n9660)
         );
  INV_X1 U10784 ( .A(n9697), .ZN(n9865) );
  NAND3_X1 U10785 ( .A1(n9534), .A2(n9658), .A3(n9865), .ZN(n9659) );
  NAND3_X1 U10786 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n9718) );
  MUX2_X1 U10787 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9718), .S(n9891), .Z(
        P1_U3541) );
  AOI21_X1 U10788 ( .B1(n9834), .B2(n9663), .A(n9662), .ZN(n9664) );
  OAI211_X1 U10789 ( .C1(n9697), .C2(n9666), .A(n9665), .B(n9664), .ZN(n9719)
         );
  MUX2_X1 U10790 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9719), .S(n9891), .Z(
        P1_U3540) );
  AOI21_X1 U10791 ( .B1(n9834), .B2(n9668), .A(n9667), .ZN(n9669) );
  OAI211_X1 U10792 ( .C1(n9697), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9720)
         );
  MUX2_X1 U10793 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9720), .S(n9891), .Z(
        P1_U3539) );
  AOI22_X1 U10794 ( .A1(n9673), .A2(n9835), .B1(n9834), .B2(n9672), .ZN(n9674)
         );
  OAI211_X1 U10795 ( .C1(n9697), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9721)
         );
  MUX2_X1 U10796 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9721), .S(n9891), .Z(
        P1_U3538) );
  AOI21_X1 U10797 ( .B1(n9834), .B2(n9678), .A(n9677), .ZN(n9679) );
  OAI211_X1 U10798 ( .C1(n9697), .C2(n9681), .A(n9680), .B(n9679), .ZN(n9722)
         );
  MUX2_X1 U10799 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9722), .S(n9891), .Z(
        P1_U3537) );
  AOI22_X1 U10800 ( .A1(n9683), .A2(n9835), .B1(n9834), .B2(n9682), .ZN(n9684)
         );
  OAI211_X1 U10801 ( .C1(n9839), .C2(n9686), .A(n9685), .B(n9684), .ZN(n9723)
         );
  MUX2_X1 U10802 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9723), .S(n9891), .Z(
        P1_U3536) );
  AOI21_X1 U10803 ( .B1(n9834), .B2(n9688), .A(n9687), .ZN(n9689) );
  OAI211_X1 U10804 ( .C1(n9697), .C2(n9691), .A(n9690), .B(n9689), .ZN(n9724)
         );
  MUX2_X1 U10805 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9724), .S(n9891), .Z(
        P1_U3535) );
  AOI211_X1 U10806 ( .C1(n9834), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9695)
         );
  OAI21_X1 U10807 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n9725) );
  MUX2_X1 U10808 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9725), .S(n9891), .Z(
        P1_U3533) );
  INV_X1 U10809 ( .A(n9698), .ZN(n9703) );
  AOI22_X1 U10810 ( .A1(n9700), .A2(n9835), .B1(n9834), .B2(n9699), .ZN(n9701)
         );
  OAI211_X1 U10811 ( .C1(n9839), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9726)
         );
  MUX2_X1 U10812 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9726), .S(n9891), .Z(
        P1_U3532) );
  MUX2_X1 U10813 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9704), .S(n9891), .Z(
        P1_U3523) );
  MUX2_X1 U10814 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9705), .S(n9876), .Z(
        P1_U3522) );
  MUX2_X1 U10815 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9706), .S(n9876), .Z(
        P1_U3521) );
  MUX2_X1 U10816 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9708), .S(n9876), .Z(
        P1_U3519) );
  MUX2_X1 U10817 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9709), .S(n9876), .Z(
        P1_U3518) );
  MUX2_X1 U10818 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9710), .S(n9876), .Z(
        P1_U3517) );
  MUX2_X1 U10819 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9711), .S(n9876), .Z(
        P1_U3516) );
  MUX2_X1 U10820 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9712), .S(n9876), .Z(
        P1_U3515) );
  MUX2_X1 U10821 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9713), .S(n9876), .Z(
        P1_U3514) );
  MUX2_X1 U10822 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9714), .S(n9876), .Z(
        P1_U3513) );
  MUX2_X1 U10823 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9715), .S(n9876), .Z(
        P1_U3512) );
  MUX2_X1 U10824 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9716), .S(n9876), .Z(
        P1_U3511) );
  MUX2_X1 U10825 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9717), .S(n9876), .Z(
        P1_U3510) );
  MUX2_X1 U10826 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9718), .S(n9876), .Z(
        P1_U3508) );
  MUX2_X1 U10827 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9719), .S(n9876), .Z(
        P1_U3505) );
  MUX2_X1 U10828 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9720), .S(n9876), .Z(
        P1_U3502) );
  MUX2_X1 U10829 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9721), .S(n9876), .Z(
        P1_U3499) );
  MUX2_X1 U10830 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9722), .S(n9876), .Z(
        P1_U3496) );
  MUX2_X1 U10831 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9723), .S(n9876), .Z(
        P1_U3493) );
  MUX2_X1 U10832 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9724), .S(n9876), .Z(
        P1_U3490) );
  MUX2_X1 U10833 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n9725), .S(n9876), .Z(
        P1_U3484) );
  MUX2_X1 U10834 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n9726), .S(n9876), .Z(
        P1_U3481) );
  NOR4_X1 U10835 ( .A1(n9728), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9727), .A4(
        P1_U3084), .ZN(n9729) );
  AOI21_X1 U10836 ( .B1(n9740), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9729), .ZN(
        n9730) );
  OAI21_X1 U10837 ( .B1(n9731), .B2(n4261), .A(n9730), .ZN(P1_U3322) );
  OAI222_X1 U10838 ( .A1(n9743), .A2(n9734), .B1(n4261), .B2(n9733), .C1(n9732), .C2(P1_U3084), .ZN(P1_U3324) );
  NAND2_X1 U10839 ( .A1(n9736), .A2(n9735), .ZN(n9738) );
  OAI211_X1 U10840 ( .C1(n9743), .C2(n10133), .A(n9738), .B(n9737), .ZN(
        P1_U3325) );
  AOI21_X1 U10841 ( .B1(n9740), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9739), .ZN(
        n9741) );
  OAI21_X1 U10842 ( .B1(n9742), .B2(n4261), .A(n9741), .ZN(P1_U3326) );
  OAI222_X1 U10843 ( .A1(P1_U3084), .A2(n9746), .B1(n4261), .B2(n9745), .C1(
        n9744), .C2(n9743), .ZN(P1_U3327) );
  INV_X1 U10844 ( .A(n9747), .ZN(n9748) );
  MUX2_X1 U10845 ( .A(n9748), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U10846 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9749) );
  AOI21_X1 U10847 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9749), .ZN(n10012) );
  NOR2_X1 U10848 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9750) );
  AOI21_X1 U10849 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9750), .ZN(n10015) );
  NOR2_X1 U10850 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9751) );
  AOI21_X1 U10851 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9751), .ZN(n10018) );
  NOR2_X1 U10852 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9752) );
  AOI21_X1 U10853 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9752), .ZN(n10021) );
  NOR2_X1 U10854 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9753) );
  AOI21_X1 U10855 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9753), .ZN(n10024) );
  NOR2_X1 U10856 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9760) );
  XNOR2_X1 U10857 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10225) );
  NAND2_X1 U10858 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9758) );
  XOR2_X1 U10859 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10223) );
  NAND2_X1 U10860 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9756) );
  XOR2_X1 U10861 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10219) );
  AOI21_X1 U10862 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10005) );
  INV_X1 U10863 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9754) );
  NAND3_X1 U10864 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U10865 ( .A1(n10219), .A2(n10218), .ZN(n9755) );
  NAND2_X1 U10866 ( .A1(n9756), .A2(n9755), .ZN(n10222) );
  NAND2_X1 U10867 ( .A1(n10223), .A2(n10222), .ZN(n9757) );
  NAND2_X1 U10868 ( .A1(n9758), .A2(n9757), .ZN(n10224) );
  NOR2_X1 U10869 ( .A1(n10225), .A2(n10224), .ZN(n9759) );
  NOR2_X1 U10870 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9761), .ZN(n10208) );
  NAND2_X1 U10871 ( .A1(n9763), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9764) );
  XOR2_X1 U10872 ( .A(n9763), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10210) );
  NAND2_X1 U10873 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9765), .ZN(n9766) );
  XOR2_X1 U10874 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9765), .Z(n10221) );
  NAND2_X1 U10875 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9767), .ZN(n9769) );
  XOR2_X1 U10876 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9767), .Z(n10220) );
  NAND2_X1 U10877 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10220), .ZN(n9768) );
  NAND2_X1 U10878 ( .A1(n9769), .A2(n9768), .ZN(n9770) );
  AND2_X1 U10879 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9770), .ZN(n9771) );
  XNOR2_X1 U10880 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9770), .ZN(n10216) );
  NAND2_X1 U10881 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9772) );
  OAI21_X1 U10882 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9772), .ZN(n10032) );
  NAND2_X1 U10883 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9773) );
  OAI21_X1 U10884 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9773), .ZN(n10029) );
  NOR2_X1 U10885 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9774) );
  AOI21_X1 U10886 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9774), .ZN(n10026) );
  NAND2_X1 U10887 ( .A1(n10021), .A2(n10020), .ZN(n10019) );
  NAND2_X1 U10888 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  OAI21_X1 U10889 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10013), .ZN(n10011) );
  NAND2_X1 U10890 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  NOR2_X1 U10891 ( .A1(n10213), .A2(n10212), .ZN(n9775) );
  NAND2_X1 U10892 ( .A1(n10213), .A2(n10212), .ZN(n10211) );
  XOR2_X1 U10893 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9776) );
  XNOR2_X1 U10894 ( .A(n9777), .B(n9776), .ZN(ADD_1071_U4) );
  XNOR2_X1 U10895 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10896 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10897 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10009) );
  INV_X1 U10898 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9785) );
  OAI22_X1 U10899 ( .A1(n9779), .A2(n9786), .B1(n9778), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U10900 ( .A1(n9781), .A2(n9780), .ZN(n9783) );
  AOI21_X1 U10901 ( .B1(n9783), .B2(n9782), .A(P1_U3084), .ZN(n9784) );
  AOI21_X1 U10902 ( .B1(n9785), .B2(P1_U3084), .A(n9784), .ZN(n9788) );
  NOR3_X1 U10903 ( .A1(n9807), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9786), .ZN(
        n9787) );
  AOI21_X1 U10904 ( .B1(n9788), .B2(P1_U3083), .A(n9787), .ZN(n9789) );
  OAI21_X1 U10905 ( .B1(n9813), .B2(n10009), .A(n9789), .ZN(P1_U3241) );
  INV_X1 U10906 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9814) );
  NAND2_X1 U10907 ( .A1(n9790), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9792) );
  OAI21_X1 U10908 ( .B1(n9808), .B2(n9792), .A(n9791), .ZN(n9804) );
  INV_X1 U10909 ( .A(n9793), .ZN(n9803) );
  INV_X1 U10910 ( .A(n9795), .ZN(n9797) );
  MUX2_X1 U10911 ( .A(n6343), .B(P1_REG2_REG_8__SCAN_IN), .S(n9805), .Z(n9796)
         );
  NAND3_X1 U10912 ( .A1(n9798), .A2(n9797), .A3(n9796), .ZN(n9800) );
  AOI21_X1 U10913 ( .B1(n9801), .B2(n9800), .A(n9799), .ZN(n9802) );
  AOI211_X1 U10914 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9812)
         );
  AOI211_X1 U10915 ( .C1(n9809), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9810)
         );
  INV_X1 U10916 ( .A(n9810), .ZN(n9811) );
  OAI211_X1 U10917 ( .C1(n9814), .C2(n9813), .A(n9812), .B(n9811), .ZN(
        P1_U3249) );
  AND2_X1 U10918 ( .A1(n9816), .A2(n9815), .ZN(n9817) );
  AND2_X1 U10919 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9818), .ZN(P1_U3292) );
  AND2_X1 U10920 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9818), .ZN(P1_U3293) );
  AND2_X1 U10921 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9818), .ZN(P1_U3294) );
  AND2_X1 U10922 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9818), .ZN(P1_U3295) );
  AND2_X1 U10923 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9818), .ZN(P1_U3296) );
  AND2_X1 U10924 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9818), .ZN(P1_U3297) );
  AND2_X1 U10925 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9818), .ZN(P1_U3298) );
  AND2_X1 U10926 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9818), .ZN(P1_U3299) );
  AND2_X1 U10927 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9818), .ZN(P1_U3300) );
  AND2_X1 U10928 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9818), .ZN(P1_U3301) );
  AND2_X1 U10929 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9818), .ZN(P1_U3302) );
  AND2_X1 U10930 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9818), .ZN(P1_U3303) );
  NOR2_X1 U10931 ( .A1(n9817), .A2(n10109), .ZN(P1_U3304) );
  AND2_X1 U10932 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9818), .ZN(P1_U3305) );
  NOR2_X1 U10933 ( .A1(n9817), .A2(n10155), .ZN(P1_U3306) );
  NOR2_X1 U10934 ( .A1(n9817), .A2(n10147), .ZN(P1_U3307) );
  AND2_X1 U10935 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9818), .ZN(P1_U3308) );
  AND2_X1 U10936 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9818), .ZN(P1_U3309) );
  AND2_X1 U10937 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9818), .ZN(P1_U3310) );
  AND2_X1 U10938 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9818), .ZN(P1_U3311) );
  AND2_X1 U10939 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9818), .ZN(P1_U3312) );
  AND2_X1 U10940 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9818), .ZN(P1_U3313) );
  AND2_X1 U10941 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9818), .ZN(P1_U3314) );
  AND2_X1 U10942 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9818), .ZN(P1_U3315) );
  AND2_X1 U10943 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9818), .ZN(P1_U3316) );
  NOR2_X1 U10944 ( .A1(n9817), .A2(n10172), .ZN(P1_U3317) );
  AND2_X1 U10945 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9818), .ZN(P1_U3318) );
  AND2_X1 U10946 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9818), .ZN(P1_U3319) );
  AND2_X1 U10947 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9818), .ZN(P1_U3320) );
  AND2_X1 U10948 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9818), .ZN(P1_U3321) );
  INV_X1 U10949 ( .A(n9819), .ZN(n9824) );
  OAI21_X1 U10950 ( .B1(n9821), .B2(n9868), .A(n9820), .ZN(n9823) );
  AOI211_X1 U10951 ( .C1(n9856), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9878)
         );
  INV_X1 U10952 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9825) );
  AOI22_X1 U10953 ( .A1(n9876), .A2(n9878), .B1(n9825), .B2(n9874), .ZN(
        P1_U3457) );
  INV_X1 U10954 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10108) );
  AOI22_X1 U10955 ( .A1(n9876), .A2(n9826), .B1(n10108), .B2(n9874), .ZN(
        P1_U3460) );
  OAI22_X1 U10956 ( .A1(n9828), .A2(n9869), .B1(n9827), .B2(n9868), .ZN(n9830)
         );
  AOI211_X1 U10957 ( .C1(n9856), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9879)
         );
  INV_X1 U10958 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9832) );
  AOI22_X1 U10959 ( .A1(n9876), .A2(n9879), .B1(n9832), .B2(n9874), .ZN(
        P1_U3463) );
  AOI22_X1 U10960 ( .A1(n9836), .A2(n9835), .B1(n9834), .B2(n9833), .ZN(n9837)
         );
  OAI211_X1 U10961 ( .C1(n9840), .C2(n9839), .A(n9838), .B(n9837), .ZN(n9841)
         );
  INV_X1 U10962 ( .A(n9841), .ZN(n9881) );
  INV_X1 U10963 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9842) );
  AOI22_X1 U10964 ( .A1(n9876), .A2(n9881), .B1(n9842), .B2(n9874), .ZN(
        P1_U3466) );
  AND3_X1 U10965 ( .A1(n9844), .A2(n9865), .A3(n9843), .ZN(n9848) );
  NOR2_X1 U10966 ( .A1(n9845), .A2(n9868), .ZN(n9846) );
  NOR4_X1 U10967 ( .A1(n9849), .A2(n9848), .A3(n9847), .A4(n9846), .ZN(n9883)
         );
  INV_X1 U10968 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10969 ( .A1(n9876), .A2(n9883), .B1(n9850), .B2(n9874), .ZN(
        P1_U3469) );
  OAI22_X1 U10970 ( .A1(n9852), .A2(n9869), .B1(n9851), .B2(n9868), .ZN(n9854)
         );
  AOI211_X1 U10971 ( .C1(n9856), .C2(n9855), .A(n9854), .B(n9853), .ZN(n9885)
         );
  INV_X1 U10972 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U10973 ( .A1(n9876), .A2(n9885), .B1(n9857), .B2(n9874), .ZN(
        P1_U3472) );
  OAI21_X1 U10974 ( .B1(n9859), .B2(n9868), .A(n9858), .ZN(n9861) );
  AOI211_X1 U10975 ( .C1(n9865), .C2(n9862), .A(n9861), .B(n9860), .ZN(n9887)
         );
  INV_X1 U10976 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9863) );
  AOI22_X1 U10977 ( .A1(n9876), .A2(n9887), .B1(n9863), .B2(n9874), .ZN(
        P1_U3475) );
  AND3_X1 U10978 ( .A1(n9866), .A2(n9865), .A3(n9864), .ZN(n9872) );
  OAI22_X1 U10979 ( .A1(n9870), .A2(n9869), .B1(n4913), .B2(n9868), .ZN(n9871)
         );
  NOR3_X1 U10980 ( .A1(n9873), .A2(n9872), .A3(n9871), .ZN(n9890) );
  INV_X1 U10981 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9875) );
  AOI22_X1 U10982 ( .A1(n9876), .A2(n9890), .B1(n9875), .B2(n9874), .ZN(
        P1_U3478) );
  AOI22_X1 U10983 ( .A1(n9891), .A2(n9878), .B1(n9877), .B2(n9888), .ZN(
        P1_U3524) );
  AOI22_X1 U10984 ( .A1(n9891), .A2(n9879), .B1(n6192), .B2(n9888), .ZN(
        P1_U3526) );
  AOI22_X1 U10985 ( .A1(n9891), .A2(n9881), .B1(n9880), .B2(n9888), .ZN(
        P1_U3527) );
  AOI22_X1 U10986 ( .A1(n9891), .A2(n9883), .B1(n9882), .B2(n9888), .ZN(
        P1_U3528) );
  AOI22_X1 U10987 ( .A1(n9891), .A2(n9885), .B1(n9884), .B2(n9888), .ZN(
        P1_U3529) );
  AOI22_X1 U10988 ( .A1(n9891), .A2(n9887), .B1(n9886), .B2(n9888), .ZN(
        P1_U3530) );
  INV_X1 U10989 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U10990 ( .A1(n9891), .A2(n9890), .B1(n9889), .B2(n9888), .ZN(
        P1_U3531) );
  AOI21_X1 U10991 ( .B1(n6954), .B2(n9893), .A(n9892), .ZN(n9895) );
  AOI21_X1 U10992 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n9967) );
  XNOR2_X1 U10993 ( .A(n9899), .B(n9898), .ZN(n9966) );
  INV_X1 U10994 ( .A(n9900), .ZN(n9901) );
  OAI22_X1 U10995 ( .A1(n9921), .A2(n9966), .B1(n9901), .B2(n9919), .ZN(n9905)
         );
  XNOR2_X1 U10996 ( .A(n9902), .B(n9903), .ZN(n9964) );
  OAI22_X1 U10997 ( .A1(n9965), .A2(n9925), .B1(n9924), .B2(n9964), .ZN(n9904)
         );
  AOI211_X1 U10998 ( .C1(n8651), .C2(P2_REG2_REG_4__SCAN_IN), .A(n9905), .B(
        n9904), .ZN(n9906) );
  OAI21_X1 U10999 ( .B1(n8651), .B2(n9967), .A(n9906), .ZN(P2_U3292) );
  OAI21_X1 U11000 ( .B1(n9922), .B2(n9908), .A(n9907), .ZN(n9912) );
  AOI222_X1 U11001 ( .A1(n9913), .A2(n9912), .B1(n9911), .B2(n9910), .C1(n9909), .C2(n8596), .ZN(n9950) );
  AND2_X1 U11002 ( .A1(n9916), .A2(n9915), .ZN(n9918) );
  OR2_X1 U11003 ( .A1(n9918), .A2(n9917), .ZN(n9949) );
  INV_X1 U11004 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9920) );
  OAI22_X1 U11005 ( .A1(n9921), .A2(n9949), .B1(n9920), .B2(n9919), .ZN(n9927)
         );
  XNOR2_X1 U11006 ( .A(n9923), .B(n9922), .ZN(n9947) );
  OAI22_X1 U11007 ( .A1(n9948), .A2(n9925), .B1(n9924), .B2(n9947), .ZN(n9926)
         );
  AOI211_X1 U11008 ( .C1(n8651), .C2(P2_REG2_REG_2__SCAN_IN), .A(n9927), .B(
        n9926), .ZN(n9928) );
  OAI21_X1 U11009 ( .B1(n8651), .B2(n9950), .A(n9928), .ZN(P2_U3294) );
  NOR2_X1 U11010 ( .A1(n9930), .A2(n9929), .ZN(n9931) );
  AND2_X1 U11011 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9935), .ZN(P2_U3297) );
  INV_X1 U11012 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10178) );
  NOR2_X1 U11013 ( .A1(n9931), .A2(n10178), .ZN(P2_U3298) );
  AND2_X1 U11014 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9935), .ZN(P2_U3299) );
  AND2_X1 U11015 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9935), .ZN(P2_U3300) );
  AND2_X1 U11016 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9935), .ZN(P2_U3301) );
  AND2_X1 U11017 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9935), .ZN(P2_U3302) );
  AND2_X1 U11018 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9935), .ZN(P2_U3303) );
  AND2_X1 U11019 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9935), .ZN(P2_U3304) );
  AND2_X1 U11020 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9935), .ZN(P2_U3305) );
  AND2_X1 U11021 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9935), .ZN(P2_U3306) );
  AND2_X1 U11022 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9935), .ZN(P2_U3307) );
  INV_X1 U11023 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10073) );
  NOR2_X1 U11024 ( .A1(n9931), .A2(n10073), .ZN(P2_U3308) );
  AND2_X1 U11025 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9935), .ZN(P2_U3309) );
  AND2_X1 U11026 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9935), .ZN(P2_U3310) );
  AND2_X1 U11027 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9935), .ZN(P2_U3311) );
  AND2_X1 U11028 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9935), .ZN(P2_U3312) );
  AND2_X1 U11029 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9935), .ZN(P2_U3313) );
  AND2_X1 U11030 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9935), .ZN(P2_U3314) );
  AND2_X1 U11031 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9935), .ZN(P2_U3315) );
  AND2_X1 U11032 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9935), .ZN(P2_U3316) );
  AND2_X1 U11033 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9935), .ZN(P2_U3317) );
  AND2_X1 U11034 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9935), .ZN(P2_U3318) );
  AND2_X1 U11035 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9935), .ZN(P2_U3319) );
  AND2_X1 U11036 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9935), .ZN(P2_U3320) );
  AND2_X1 U11037 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9935), .ZN(P2_U3321) );
  AND2_X1 U11038 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9935), .ZN(P2_U3322) );
  AND2_X1 U11039 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9935), .ZN(P2_U3323) );
  AND2_X1 U11040 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9935), .ZN(P2_U3324) );
  AND2_X1 U11041 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9935), .ZN(P2_U3325) );
  AND2_X1 U11042 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9935), .ZN(P2_U3326) );
  INV_X1 U11043 ( .A(n9932), .ZN(n9934) );
  AOI22_X1 U11044 ( .A1(n9938), .A2(n9934), .B1(n9933), .B2(n9935), .ZN(
        P2_U3437) );
  AOI22_X1 U11045 ( .A1(n9938), .A2(n9937), .B1(n9936), .B2(n9935), .ZN(
        P2_U3438) );
  INV_X1 U11046 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9939) );
  AOI22_X1 U11047 ( .A1(n9994), .A2(n9940), .B1(n9939), .B2(n9992), .ZN(
        P2_U3451) );
  OAI22_X1 U11048 ( .A1(n9942), .A2(n9986), .B1(n9941), .B2(n9985), .ZN(n9945)
         );
  INV_X1 U11049 ( .A(n9943), .ZN(n9944) );
  AOI211_X1 U11050 ( .C1(n9981), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9996)
         );
  AOI22_X1 U11051 ( .A1(n9994), .A2(n9996), .B1(n5039), .B2(n9992), .ZN(
        P2_U3454) );
  INV_X1 U11052 ( .A(n9947), .ZN(n9953) );
  OAI22_X1 U11053 ( .A1(n9949), .A2(n9986), .B1(n9948), .B2(n9985), .ZN(n9952)
         );
  INV_X1 U11054 ( .A(n9950), .ZN(n9951) );
  AOI211_X1 U11055 ( .C1(n9981), .C2(n9953), .A(n9952), .B(n9951), .ZN(n9997)
         );
  INV_X1 U11056 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U11057 ( .A1(n9994), .A2(n9997), .B1(n9954), .B2(n9992), .ZN(
        P2_U3457) );
  AOI22_X1 U11058 ( .A1(n9958), .A2(n9957), .B1(n9956), .B2(n9955), .ZN(n9959)
         );
  OAI211_X1 U11059 ( .C1(n9961), .C2(n9984), .A(n9960), .B(n9959), .ZN(n9962)
         );
  INV_X1 U11060 ( .A(n9962), .ZN(n9998) );
  INV_X1 U11061 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U11062 ( .A1(n9994), .A2(n9998), .B1(n9963), .B2(n9992), .ZN(
        P2_U3460) );
  INV_X1 U11063 ( .A(n9964), .ZN(n9970) );
  OAI22_X1 U11064 ( .A1(n9966), .A2(n9986), .B1(n9965), .B2(n9985), .ZN(n9969)
         );
  INV_X1 U11065 ( .A(n9967), .ZN(n9968) );
  AOI211_X1 U11066 ( .C1(n9981), .C2(n9970), .A(n9969), .B(n9968), .ZN(n9999)
         );
  INV_X1 U11067 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U11068 ( .A1(n9994), .A2(n9999), .B1(n9971), .B2(n9992), .ZN(
        P2_U3463) );
  OAI211_X1 U11069 ( .C1(n9974), .C2(n9985), .A(n9973), .B(n9972), .ZN(n9975)
         );
  AOI21_X1 U11070 ( .B1(n9981), .B2(n9976), .A(n9975), .ZN(n10000) );
  INV_X1 U11071 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U11072 ( .A1(n9994), .A2(n10000), .B1(n10177), .B2(n9992), .ZN(
        P2_U3466) );
  OAI22_X1 U11073 ( .A1(n9978), .A2(n9986), .B1(n9977), .B2(n9985), .ZN(n9980)
         );
  AOI211_X1 U11074 ( .C1(n9982), .C2(n9981), .A(n9980), .B(n9979), .ZN(n10001)
         );
  INV_X1 U11075 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U11076 ( .A1(n9994), .A2(n10001), .B1(n9983), .B2(n9992), .ZN(
        P2_U3469) );
  INV_X1 U11077 ( .A(n9984), .ZN(n9991) );
  OAI22_X1 U11078 ( .A1(n9987), .A2(n9986), .B1(n4983), .B2(n9985), .ZN(n9989)
         );
  AOI211_X1 U11079 ( .C1(n9991), .C2(n9990), .A(n9989), .B(n9988), .ZN(n10003)
         );
  INV_X1 U11080 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U11081 ( .A1(n9994), .A2(n10003), .B1(n9993), .B2(n9992), .ZN(
        P2_U3475) );
  INV_X1 U11082 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9995) );
  AOI22_X1 U11083 ( .A1(n10004), .A2(n9996), .B1(n9995), .B2(n10002), .ZN(
        P2_U3521) );
  AOI22_X1 U11084 ( .A1(n10004), .A2(n9997), .B1(n6426), .B2(n10002), .ZN(
        P2_U3522) );
  AOI22_X1 U11085 ( .A1(n10004), .A2(n9998), .B1(n6560), .B2(n10002), .ZN(
        P2_U3523) );
  AOI22_X1 U11086 ( .A1(n10004), .A2(n9999), .B1(n10130), .B2(n10002), .ZN(
        P2_U3524) );
  AOI22_X1 U11087 ( .A1(n10004), .A2(n10000), .B1(n6666), .B2(n10002), .ZN(
        P2_U3525) );
  AOI22_X1 U11088 ( .A1(n10004), .A2(n10001), .B1(n6668), .B2(n10002), .ZN(
        P2_U3526) );
  AOI22_X1 U11089 ( .A1(n10004), .A2(n10003), .B1(n10141), .B2(n10002), .ZN(
        P2_U3528) );
  INV_X1 U11090 ( .A(n10005), .ZN(n10006) );
  NAND2_X1 U11091 ( .A1(n10007), .A2(n10006), .ZN(n10008) );
  XNOR2_X1 U11092 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10008), .ZN(ADD_1071_U5)
         );
  AOI22_X1 U11093 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n6627), .B2(n10009), .ZN(ADD_1071_U46) );
  OAI21_X1 U11094 ( .B1(n10012), .B2(n10011), .A(n10010), .ZN(ADD_1071_U56) );
  OAI21_X1 U11095 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(ADD_1071_U57) );
  OAI21_X1 U11096 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(ADD_1071_U58) );
  OAI21_X1 U11097 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(ADD_1071_U59) );
  OAI21_X1 U11098 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(ADD_1071_U60) );
  OAI21_X1 U11099 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(ADD_1071_U61) );
  AOI21_X1 U11100 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(ADD_1071_U62) );
  AOI21_X1 U11101 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(ADD_1071_U63) );
  NAND3_X1 U11102 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .A3(
        P2_IR_REG_10__SCAN_IN), .ZN(n10035) );
  NAND3_X1 U11103 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(P2_REG2_REG_27__SCAN_IN), .A3(SI_31_), .ZN(n10034) );
  NOR4_X1 U11104 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        n10035), .A4(n10034), .ZN(n10065) );
  NOR3_X1 U11105 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(P2_REG2_REG_28__SCAN_IN), 
        .A3(n7640), .ZN(n10062) );
  NOR3_X1 U11106 ( .A1(n10036), .A2(P1_DATAO_REG_30__SCAN_IN), .A3(
        P1_ADDR_REG_15__SCAN_IN), .ZN(n10050) );
  AND4_X1 U11107 ( .A1(n10037), .A2(n10129), .A3(n10085), .A4(n10084), .ZN(
        n10049) );
  OR4_X1 U11108 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n10141), .A3(n6965), .A4(
        n10130), .ZN(n10039) );
  NOR2_X1 U11109 ( .A1(n10039), .A2(n10038), .ZN(n10046) );
  INV_X1 U11110 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10115) );
  NOR4_X1 U11111 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(SI_23_), .A3(
        P2_REG2_REG_18__SCAN_IN), .A4(n10115), .ZN(n10045) );
  NAND4_X1 U11112 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(P2_DATAO_REG_28__SCAN_IN), .A3(n10169), .A4(n10132), .ZN(n10040) );
  NOR2_X1 U11113 ( .A1(n6343), .A2(n10040), .ZN(n10044) );
  INV_X1 U11114 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10041) );
  INV_X1 U11115 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10097) );
  NAND4_X1 U11116 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(n10041), .A3(n10095), .A4(
        n10097), .ZN(n10042) );
  INV_X1 U11117 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10168) );
  NOR2_X1 U11118 ( .A1(n10042), .A2(n10168), .ZN(n10043) );
  NAND4_X1 U11119 ( .A1(n10046), .A2(n10045), .A3(n10044), .A4(n10043), .ZN(
        n10047) );
  NOR2_X1 U11120 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(n10047), .ZN(n10048) );
  AND4_X1 U11121 ( .A1(n10050), .A2(n10049), .A3(P2_D_REG_30__SCAN_IN), .A4(
        n10048), .ZN(n10061) );
  NAND4_X1 U11122 ( .A1(n5141), .A2(n10051), .A3(n10083), .A4(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n10054) );
  INV_X1 U11123 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10052) );
  NAND4_X1 U11124 ( .A1(n10052), .A2(P1_REG0_REG_2__SCAN_IN), .A3(
        P1_REG1_REG_2__SCAN_IN), .A4(P1_REG2_REG_1__SCAN_IN), .ZN(n10053) );
  NOR2_X1 U11125 ( .A1(n10054), .A2(n10053), .ZN(n10060) );
  NAND4_X1 U11126 ( .A1(n10055), .A2(n10177), .A3(P1_DATAO_REG_6__SCAN_IN), 
        .A4(P1_DATAO_REG_3__SCAN_IN), .ZN(n10058) );
  NAND4_X1 U11127 ( .A1(n10056), .A2(n10171), .A3(P2_REG1_REG_18__SCAN_IN), 
        .A4(P2_REG0_REG_25__SCAN_IN), .ZN(n10057) );
  NOR2_X1 U11128 ( .A1(n10058), .A2(n10057), .ZN(n10059) );
  AND4_X1 U11129 ( .A1(n10062), .A2(n10061), .A3(n10060), .A4(n10059), .ZN(
        n10064) );
  INV_X1 U11130 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10082) );
  INV_X1 U11131 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n10154) );
  INV_X1 U11132 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10162) );
  NOR4_X1 U11133 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10082), .A3(n10154), 
        .A4(n10162), .ZN(n10063) );
  NAND3_X1 U11134 ( .A1(n10065), .A2(n10064), .A3(n10063), .ZN(n10066) );
  NAND2_X1 U11135 ( .A1(n10066), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U11136 ( .A1(n5785), .A2(keyinput45), .B1(keyinput16), .B2(n10068), 
        .ZN(n10067) );
  OAI221_X1 U11137 ( .B1(n5785), .B2(keyinput45), .C1(n10068), .C2(keyinput16), 
        .A(n10067), .ZN(n10080) );
  AOI22_X1 U11138 ( .A1(n10071), .A2(keyinput18), .B1(keyinput4), .B2(n10070), 
        .ZN(n10069) );
  OAI221_X1 U11139 ( .B1(n10071), .B2(keyinput18), .C1(n10070), .C2(keyinput4), 
        .A(n10069), .ZN(n10079) );
  XNOR2_X1 U11140 ( .A(P1_REG1_REG_13__SCAN_IN), .B(keyinput30), .ZN(n10072)
         );
  OAI21_X1 U11141 ( .B1(n10073), .B2(keyinput36), .A(n10072), .ZN(n10078) );
  XNOR2_X1 U11142 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput41), .ZN(n10075) );
  NAND2_X1 U11143 ( .A1(n10073), .A2(keyinput36), .ZN(n10074) );
  OAI211_X1 U11144 ( .C1(keyinput31), .C2(n10076), .A(n10075), .B(n10074), 
        .ZN(n10077) );
  NOR4_X1 U11145 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10125) );
  AOI22_X1 U11146 ( .A1(n10083), .A2(keyinput6), .B1(keyinput58), .B2(n10082), 
        .ZN(n10081) );
  OAI221_X1 U11147 ( .B1(n10083), .B2(keyinput6), .C1(n10082), .C2(keyinput58), 
        .A(n10081), .ZN(n10093) );
  XNOR2_X1 U11148 ( .A(n10084), .B(keyinput48), .ZN(n10092) );
  XNOR2_X1 U11149 ( .A(n10085), .B(keyinput5), .ZN(n10091) );
  XNOR2_X1 U11150 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput2), .ZN(n10089) );
  XNOR2_X1 U11151 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput37), .ZN(n10088)
         );
  XNOR2_X1 U11152 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput0), .ZN(n10087) );
  XNOR2_X1 U11153 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput55), .ZN(n10086) );
  NAND4_X1 U11154 ( .A1(n10089), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        n10090) );
  NOR4_X1 U11155 ( .A1(n10093), .A2(n10092), .A3(n10091), .A4(n10090), .ZN(
        n10124) );
  AOI22_X1 U11156 ( .A1(n10095), .A2(keyinput62), .B1(keyinput23), .B2(n5532), 
        .ZN(n10094) );
  OAI221_X1 U11157 ( .B1(n10095), .B2(keyinput62), .C1(n5532), .C2(keyinput23), 
        .A(n10094), .ZN(n10106) );
  INV_X1 U11158 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10098) );
  AOI22_X1 U11159 ( .A1(n10098), .A2(keyinput53), .B1(n10097), .B2(keyinput22), 
        .ZN(n10096) );
  OAI221_X1 U11160 ( .B1(n10098), .B2(keyinput53), .C1(n10097), .C2(keyinput22), .A(n10096), .ZN(n10105) );
  INV_X1 U11161 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U11162 ( .A1(n5798), .A2(keyinput51), .B1(n10100), .B2(keyinput14), 
        .ZN(n10099) );
  OAI221_X1 U11163 ( .B1(n5798), .B2(keyinput51), .C1(n10100), .C2(keyinput14), 
        .A(n10099), .ZN(n10104) );
  XNOR2_X1 U11164 ( .A(P1_REG0_REG_14__SCAN_IN), .B(keyinput42), .ZN(n10102)
         );
  XNOR2_X1 U11165 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput26), .ZN(n10101) );
  NAND2_X1 U11166 ( .A1(n10102), .A2(n10101), .ZN(n10103) );
  NOR4_X1 U11167 ( .A1(n10106), .A2(n10105), .A3(n10104), .A4(n10103), .ZN(
        n10123) );
  AOI22_X1 U11168 ( .A1(n10108), .A2(keyinput9), .B1(keyinput46), .B2(n5436), 
        .ZN(n10107) );
  OAI221_X1 U11169 ( .B1(n10108), .B2(keyinput9), .C1(n5436), .C2(keyinput46), 
        .A(n10107), .ZN(n10111) );
  XNOR2_X1 U11170 ( .A(n10109), .B(keyinput43), .ZN(n10110) );
  NOR2_X1 U11171 ( .A1(n10111), .A2(n10110), .ZN(n10121) );
  AOI22_X1 U11172 ( .A1(n10051), .A2(keyinput39), .B1(n7640), .B2(keyinput60), 
        .ZN(n10112) );
  OAI221_X1 U11173 ( .B1(n10051), .B2(keyinput39), .C1(n7640), .C2(keyinput60), 
        .A(n10112), .ZN(n10113) );
  INV_X1 U11174 ( .A(n10113), .ZN(n10120) );
  INV_X1 U11175 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U11176 ( .A1(n10116), .A2(keyinput50), .B1(n10115), .B2(keyinput38), 
        .ZN(n10114) );
  OAI221_X1 U11177 ( .B1(n10116), .B2(keyinput50), .C1(n10115), .C2(keyinput38), .A(n10114), .ZN(n10117) );
  INV_X1 U11178 ( .A(n10117), .ZN(n10119) );
  XNOR2_X1 U11179 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput3), .ZN(n10118) );
  AND4_X1 U11180 ( .A1(n10121), .A2(n10120), .A3(n10119), .A4(n10118), .ZN(
        n10122) );
  NAND4_X1 U11181 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10187) );
  AOI22_X1 U11182 ( .A1(n6965), .A2(keyinput56), .B1(n10127), .B2(keyinput33), 
        .ZN(n10126) );
  OAI221_X1 U11183 ( .B1(n6965), .B2(keyinput56), .C1(n10127), .C2(keyinput33), 
        .A(n10126), .ZN(n10139) );
  AOI22_X1 U11184 ( .A1(n10130), .A2(keyinput44), .B1(n10129), .B2(keyinput8), 
        .ZN(n10128) );
  OAI221_X1 U11185 ( .B1(n10130), .B2(keyinput44), .C1(n10129), .C2(keyinput8), 
        .A(n10128), .ZN(n10138) );
  AOI22_X1 U11186 ( .A1(n10133), .A2(keyinput17), .B1(keyinput47), .B2(n10132), 
        .ZN(n10131) );
  OAI221_X1 U11187 ( .B1(n10133), .B2(keyinput17), .C1(n10132), .C2(keyinput47), .A(n10131), .ZN(n10137) );
  XNOR2_X1 U11188 ( .A(P2_REG1_REG_19__SCAN_IN), .B(keyinput32), .ZN(n10135)
         );
  XNOR2_X1 U11189 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput34), .ZN(n10134) );
  NAND2_X1 U11190 ( .A1(n10135), .A2(n10134), .ZN(n10136) );
  NOR4_X1 U11191 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n10185) );
  AOI22_X1 U11192 ( .A1(n10142), .A2(keyinput27), .B1(keyinput13), .B2(n10141), 
        .ZN(n10140) );
  OAI221_X1 U11193 ( .B1(n10142), .B2(keyinput27), .C1(n10141), .C2(keyinput13), .A(n10140), .ZN(n10151) );
  AOI22_X1 U11194 ( .A1(n5141), .A2(keyinput24), .B1(keyinput61), .B2(n5583), 
        .ZN(n10143) );
  OAI221_X1 U11195 ( .B1(n5141), .B2(keyinput24), .C1(n5583), .C2(keyinput61), 
        .A(n10143), .ZN(n10150) );
  XOR2_X1 U11196 ( .A(n5340), .B(keyinput11), .Z(n10146) );
  XNOR2_X1 U11197 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput29), .ZN(n10145) );
  XNOR2_X1 U11198 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput1), .ZN(n10144) );
  NAND3_X1 U11199 ( .A1(n10146), .A2(n10145), .A3(n10144), .ZN(n10149) );
  XNOR2_X1 U11200 ( .A(n10147), .B(keyinput49), .ZN(n10148) );
  NOR4_X1 U11201 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10184) );
  INV_X1 U11202 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U11203 ( .A1(n10154), .A2(keyinput25), .B1(keyinput40), .B2(n10153), 
        .ZN(n10152) );
  OAI221_X1 U11204 ( .B1(n10154), .B2(keyinput25), .C1(n10153), .C2(keyinput40), .A(n10152), .ZN(n10158) );
  XOR2_X1 U11205 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput7), .Z(n10157) );
  XNOR2_X1 U11206 ( .A(n10155), .B(keyinput20), .ZN(n10156) );
  OR3_X1 U11207 ( .A1(n10158), .A2(n10157), .A3(n10156), .ZN(n10166) );
  AOI22_X1 U11208 ( .A1(n10160), .A2(keyinput52), .B1(n6343), .B2(keyinput54), 
        .ZN(n10159) );
  OAI221_X1 U11209 ( .B1(n10160), .B2(keyinput52), .C1(n6343), .C2(keyinput54), 
        .A(n10159), .ZN(n10165) );
  AOI22_X1 U11210 ( .A1(n10163), .A2(keyinput10), .B1(keyinput57), .B2(n10162), 
        .ZN(n10161) );
  OAI221_X1 U11211 ( .B1(n10163), .B2(keyinput10), .C1(n10162), .C2(keyinput57), .A(n10161), .ZN(n10164) );
  NOR3_X1 U11212 ( .A1(n10166), .A2(n10165), .A3(n10164), .ZN(n10183) );
  AOI22_X1 U11213 ( .A1(n10169), .A2(keyinput19), .B1(keyinput63), .B2(n10168), 
        .ZN(n10167) );
  OAI221_X1 U11214 ( .B1(n10169), .B2(keyinput19), .C1(n10168), .C2(keyinput63), .A(n10167), .ZN(n10181) );
  AOI22_X1 U11215 ( .A1(n10055), .A2(keyinput59), .B1(n10171), .B2(keyinput12), 
        .ZN(n10170) );
  OAI221_X1 U11216 ( .B1(n10055), .B2(keyinput59), .C1(n10171), .C2(keyinput12), .A(n10170), .ZN(n10175) );
  XNOR2_X1 U11217 ( .A(n10172), .B(keyinput35), .ZN(n10174) );
  XOR2_X1 U11218 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput21), .Z(n10173) );
  OR3_X1 U11219 ( .A1(n10175), .A2(n10174), .A3(n10173), .ZN(n10180) );
  AOI22_X1 U11220 ( .A1(n10178), .A2(keyinput15), .B1(keyinput28), .B2(n10177), 
        .ZN(n10176) );
  OAI221_X1 U11221 ( .B1(n10178), .B2(keyinput15), .C1(n10177), .C2(keyinput28), .A(n10176), .ZN(n10179) );
  NOR3_X1 U11222 ( .A1(n10181), .A2(n10180), .A3(n10179), .ZN(n10182) );
  NAND4_X1 U11223 ( .A1(n10185), .A2(n10184), .A3(n10183), .A4(n10182), .ZN(
        n10186) );
  AOI211_X1 U11224 ( .C1(keyinput31), .C2(n10188), .A(n10187), .B(n10186), 
        .ZN(n10206) );
  OAI211_X1 U11225 ( .C1(n10192), .C2(n10191), .A(n10190), .B(n10189), .ZN(
        n10202) );
  NOR2_X1 U11226 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10193), .ZN(n10199) );
  AOI211_X1 U11227 ( .C1(n10197), .C2(n10196), .A(n10195), .B(n10194), .ZN(
        n10198) );
  AOI211_X1 U11228 ( .C1(n10200), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n10199), 
        .B(n10198), .ZN(n10201) );
  OAI211_X1 U11229 ( .C1(n10204), .C2(n10203), .A(n10202), .B(n10201), .ZN(
        n10205) );
  XOR2_X1 U11230 ( .A(n10206), .B(n10205), .Z(P2_U3262) );
  NOR2_X1 U11231 ( .A1(n10208), .A2(n10207), .ZN(n10209) );
  XOR2_X1 U11232 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10209), .Z(ADD_1071_U51) );
  XOR2_X1 U11233 ( .A(n10210), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  OAI21_X1 U11234 ( .B1(n10213), .B2(n10212), .A(n10211), .ZN(n10214) );
  XNOR2_X1 U11235 ( .A(n10214), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11236 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(ADD_1071_U47) );
  XOR2_X1 U11237 ( .A(n10219), .B(n10218), .Z(ADD_1071_U54) );
  XOR2_X1 U11238 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10220), .Z(ADD_1071_U48) );
  XOR2_X1 U11239 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10221), .Z(ADD_1071_U49) );
  XOR2_X1 U11240 ( .A(n10222), .B(n10223), .Z(ADD_1071_U53) );
  XNOR2_X1 U11241 ( .A(n10225), .B(n10224), .ZN(ADD_1071_U52) );
  NAND2_X1 U4770 ( .A1(n5972), .A2(n7278), .ZN(n6923) );
  AND4_X2 U4799 ( .A1(n5135), .A2(n5435), .A3(n5532), .A4(n5464), .ZN(n5136)
         );
  NAND2_X1 U4801 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5294) );
  NAND2_X1 U4902 ( .A1(n5997), .A2(n5996), .ZN(n7377) );
  CLKBUF_X2 U6830 ( .A(n6320), .Z(n4259) );
  NAND4_X1 U6845 ( .A1(n5234), .A2(n5233), .A3(n5232), .A4(n5231), .ZN(n9909)
         );
endmodule

