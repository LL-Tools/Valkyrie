

module b17_C_SARLock_k_64_7 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886;

  OR2_X1 U11036 ( .A1(n17303), .A2(n10225), .ZN(n10226) );
  AND2_X1 U11037 ( .A1(n14651), .A2(n14668), .ZN(n9669) );
  NOR2_X1 U11038 ( .A1(n18402), .A2(n17200), .ZN(n18634) );
  NAND2_X1 U11039 ( .A1(n15441), .A2(n15438), .ZN(n9827) );
  XNOR2_X1 U11040 ( .A(n12309), .B(n12460), .ZN(n15429) );
  OR2_X1 U11041 ( .A1(n12400), .A2(n12399), .ZN(n12406) );
  CLKBUF_X2 U11042 ( .A(n10661), .Z(n10774) );
  NAND2_X1 U11043 ( .A1(n9957), .A2(n12403), .ZN(n12411) );
  CLKBUF_X1 U11044 ( .A(n12604), .Z(n9633) );
  CLKBUF_X2 U11045 ( .A(n9626), .Z(n14238) );
  CLKBUF_X2 U11046 ( .A(n10171), .Z(n15537) );
  BUF_X2 U11047 ( .A(n10144), .Z(n9600) );
  NAND4_X1 U11048 ( .A1(n10654), .A2(n10653), .A3(n10648), .A4(n10652), .ZN(
        n12159) );
  AND2_X1 U11049 ( .A1(n13446), .A2(n10814), .ZN(n10856) );
  CLKBUF_X2 U11050 ( .A(n10270), .Z(n9604) );
  CLKBUF_X1 U11051 ( .A(n16697), .Z(n16876) );
  CLKBUF_X1 U11052 ( .A(n10171), .Z(n9605) );
  NOR2_X1 U11053 ( .A1(n10104), .A2(n18429), .ZN(n10150) );
  CLKBUF_X2 U11054 ( .A(n11271), .Z(n14146) );
  NOR2_X2 U11055 ( .A1(n18429), .A2(n10105), .ZN(n10188) );
  CLKBUF_X2 U11056 ( .A(n11264), .Z(n12058) );
  INV_X1 U11057 ( .A(n10627), .ZN(n12774) );
  CLKBUF_X2 U11058 ( .A(n14139), .Z(n12052) );
  CLKBUF_X2 U11059 ( .A(n11503), .Z(n12057) );
  CLKBUF_X2 U11060 ( .A(n11376), .Z(n11497) );
  NAND3_X1 U11061 ( .A1(n9996), .A2(n10575), .A3(n10576), .ZN(n12821) );
  CLKBUF_X1 U11062 ( .A(n11305), .Z(n20029) );
  CLKBUF_X1 U11063 ( .A(n11308), .Z(n20044) );
  NAND2_X1 U11064 ( .A1(n10533), .A2(n10547), .ZN(n10534) );
  AND4_X1 U11065 ( .A1(n11263), .A2(n11262), .A3(n11261), .A4(n11260), .ZN(
        n11270) );
  AND2_X1 U11066 ( .A1(n10827), .A2(n10785), .ZN(n13141) );
  AND2_X1 U11067 ( .A1(n10827), .A2(n10785), .ZN(n9601) );
  AND2_X1 U11068 ( .A1(n11194), .A2(n11193), .ZN(n11376) );
  AND2_X1 U11069 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n11183), .ZN(
        n11195) );
  CLKBUF_X1 U11070 ( .A(n16660), .Z(n9591) );
  NOR2_X1 U11071 ( .A1(n16676), .A2(n18566), .ZN(n16660) );
  CLKBUF_X1 U11072 ( .A(n18187), .Z(n9592) );
  NOR2_X1 U11073 ( .A1(n18109), .A2(n18108), .ZN(n18187) );
  INV_X1 U11074 ( .A(n18473), .ZN(n9593) );
  INV_X1 U11075 ( .A(n9593), .ZN(n9594) );
  INV_X1 U11076 ( .A(n9593), .ZN(n9595) );
  INV_X1 U11077 ( .A(n19617), .ZN(n9596) );
  INV_X1 U11078 ( .A(n9596), .ZN(n9597) );
  INV_X1 U11079 ( .A(n9596), .ZN(n9598) );
  OR2_X1 U11080 ( .A1(n11321), .A2(n12623), .ZN(n13467) );
  AND2_X1 U11081 ( .A1(n10622), .A2(n12814), .ZN(n10649) );
  AND2_X1 U11082 ( .A1(n12462), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12467) );
  NOR2_X1 U11083 ( .A1(n17988), .A2(n17993), .ZN(n10338) );
  AND2_X1 U11084 ( .A1(n11193), .A2(n11191), .ZN(n11264) );
  AND4_X1 U11085 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(
        n11255) );
  AND2_X1 U11086 ( .A1(n10827), .A2(n10785), .ZN(n9602) );
  INV_X1 U11087 ( .A(n12601), .ZN(n12605) );
  NAND2_X1 U11088 ( .A1(n11563), .A2(n11562), .ZN(n11591) );
  AND2_X1 U11089 ( .A1(n19930), .A2(n9962), .ZN(n9961) );
  NAND2_X1 U11090 ( .A1(n19940), .A2(n11415), .ZN(n11466) );
  AND4_X1 U11091 ( .A1(n11208), .A2(n11207), .A3(n11206), .A4(n11205), .ZN(
        n9639) );
  NAND2_X1 U11092 ( .A1(n19071), .A2(n19700), .ZN(n11140) );
  AOI21_X1 U11093 ( .B1(n12535), .B2(n9891), .A(n9888), .ZN(n9895) );
  INV_X1 U11094 ( .A(n9615), .ZN(n10689) );
  INV_X2 U11095 ( .A(n9622), .ZN(n12555) );
  AND4_X1 U11096 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .ZN(
        n10654) );
  CLKBUF_X2 U11098 ( .A(n11361), .Z(n13481) );
  INV_X2 U11099 ( .A(n12403), .ZN(n19061) );
  AND2_X1 U11100 ( .A1(n12411), .A2(n12418), .ZN(n12547) );
  NAND2_X1 U11101 ( .A1(n12331), .A2(n12339), .ZN(n12368) );
  INV_X2 U11102 ( .A(n13231), .ZN(n12750) );
  NAND2_X1 U11103 ( .A1(n15013), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15001) );
  NAND2_X1 U11104 ( .A1(n12446), .A2(n12290), .ZN(n13894) );
  INV_X2 U11105 ( .A(n13945), .ZN(n10466) );
  INV_X1 U11106 ( .A(n13639), .ZN(n12747) );
  NAND2_X2 U11107 ( .A1(n9657), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17818) );
  INV_X1 U11108 ( .A(n16804), .ZN(n16921) );
  OR2_X1 U11109 ( .A1(n9782), .A2(n9781), .ZN(n14277) );
  NAND2_X1 U11110 ( .A1(n13835), .A2(n13834), .ZN(n13833) );
  NAND2_X1 U11111 ( .A1(n13510), .A2(n13509), .ZN(n13511) );
  INV_X1 U11113 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19700) );
  CLKBUF_X2 U11114 ( .A(n10806), .Z(n13231) );
  NOR2_X1 U11115 ( .A1(n10459), .A2(n18794), .ZN(n10461) );
  INV_X1 U11116 ( .A(n16646), .ZN(n16666) );
  AOI21_X1 U11117 ( .B1(n17531), .B2(n15572), .A(n10229), .ZN(n15612) );
  NOR2_X1 U11118 ( .A1(n10227), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17271) );
  AND2_X1 U11119 ( .A1(n11595), .A2(n9654), .ZN(n9599) );
  INV_X2 U11120 ( .A(n20040), .ZN(n14239) );
  NAND2_X4 U11121 ( .A1(n11270), .A2(n11269), .ZN(n20040) );
  OR2_X2 U11122 ( .A1(n17536), .A2(n10210), .ZN(n9657) );
  NAND2_X2 U11123 ( .A1(n12313), .A2(n9643), .ZN(n10063) );
  INV_X4 U11124 ( .A(n10094), .ZN(n15538) );
  NOR2_X2 U11125 ( .A1(n10106), .A2(n10107), .ZN(n10144) );
  NOR3_X2 U11126 ( .A1(n12198), .A2(n12197), .A3(n12196), .ZN(n12208) );
  NAND2_X2 U11127 ( .A1(n9655), .A2(n11237), .ZN(n11308) );
  NAND2_X4 U11128 ( .A1(n10535), .A2(n10534), .ZN(n12808) );
  XNOR2_X1 U11129 ( .A(n11466), .B(n9764), .ZN(n13510) );
  AOI221_X1 U11130 ( .B1(n16973), .B2(n16985), .C1(n17032), .C2(n16985), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n16975) );
  XNOR2_X2 U11132 ( .A(n10679), .B(n10680), .ZN(n12156) );
  AND2_X4 U11133 ( .A1(n10472), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13619) );
  NOR2_X2 U11134 ( .A1(n16135), .A2(n14179), .ZN(n15413) );
  AND2_X4 U11135 ( .A1(n10821), .A2(n10785), .ZN(n9603) );
  AND2_X2 U11136 ( .A1(n10821), .A2(n10785), .ZN(n10820) );
  NOR2_X1 U11137 ( .A1(n10103), .A2(n10106), .ZN(n10270) );
  AND2_X4 U11138 ( .A1(n11591), .A2(n11590), .ZN(n9634) );
  NOR2_X1 U11139 ( .A1(n10102), .A2(n10107), .ZN(n10171) );
  XNOR2_X2 U11140 ( .A(n10371), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17613) );
  AND2_X2 U11141 ( .A1(n9659), .A2(n10149), .ZN(n10371) );
  AND2_X1 U11142 ( .A1(n14303), .A2(n12096), .ZN(n14286) );
  INV_X1 U11143 ( .A(n15001), .ZN(n9606) );
  AND2_X2 U11144 ( .A1(n12478), .A2(n9716), .ZN(n15013) );
  AOI21_X1 U11145 ( .B1(n14843), .B2(n14837), .A(n14839), .ZN(n14832) );
  NAND2_X1 U11146 ( .A1(n19929), .A2(n11518), .ZN(n13835) );
  NAND2_X1 U11147 ( .A1(n12924), .A2(n12923), .ZN(n14878) );
  AND2_X1 U11148 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16743), .ZN(n16737) );
  NAND2_X1 U11149 ( .A1(n11487), .A2(n11488), .ZN(n11538) );
  OAI21_X1 U11150 ( .B1(n13381), .B2(n13382), .A(n13383), .ZN(n19320) );
  NAND2_X1 U11152 ( .A1(n10215), .A2(n10214), .ZN(n17409) );
  AND2_X1 U11153 ( .A1(n12413), .A2(n11162), .ZN(n12415) );
  AND2_X1 U11154 ( .A1(n14111), .A2(n14110), .ZN(n14389) );
  NAND2_X1 U11155 ( .A1(n12199), .A2(n12168), .ZN(n19114) );
  INV_X2 U11157 ( .A(n16603), .ZN(n10414) );
  OAI21_X1 U11158 ( .B1(n9984), .B2(n10206), .A(n9981), .ZN(n10209) );
  NAND2_X1 U11159 ( .A1(n9907), .A2(n9906), .ZN(n10352) );
  NAND2_X1 U11160 ( .A1(n10207), .A2(n17103), .ZN(n17428) );
  NAND2_X1 U11161 ( .A1(n12774), .A2(n10637), .ZN(n10760) );
  NOR2_X2 U11162 ( .A1(n17999), .A2(n17979), .ZN(n10360) );
  NAND2_X1 U11163 ( .A1(n12605), .A2(n12623), .ZN(n12694) );
  INV_X1 U11164 ( .A(n16992), .ZN(n17988) );
  INV_X1 U11165 ( .A(n17971), .ZN(n18619) );
  NAND2_X2 U11166 ( .A1(n10623), .A2(n19045), .ZN(n12768) );
  INV_X2 U11167 ( .A(n10847), .ZN(n10838) );
  AND2_X1 U11168 ( .A1(n14239), .A2(n11310), .ZN(n13489) );
  INV_X2 U11169 ( .A(n20025), .ZN(n12599) );
  NAND2_X2 U11170 ( .A1(n10096), .A2(n9639), .ZN(n11340) );
  AND4_X2 U11171 ( .A1(n11228), .A2(n11227), .A3(n11226), .A4(n11225), .ZN(
        n20012) );
  AND4_X1 U11172 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n11256) );
  AND4_X1 U11173 ( .A1(n11236), .A2(n11235), .A3(n11234), .A4(n11233), .ZN(
        n11237) );
  AND4_X1 U11174 ( .A1(n11199), .A2(n11198), .A3(n11197), .A4(n11196), .ZN(
        n11200) );
  CLKBUF_X2 U11175 ( .A(n11250), .Z(n11988) );
  CLKBUF_X2 U11176 ( .A(n10280), .Z(n16914) );
  CLKBUF_X2 U11177 ( .A(n10552), .Z(n10813) );
  CLKBUF_X2 U11178 ( .A(n11523), .Z(n12038) );
  BUF_X2 U11179 ( .A(n11766), .Z(n12130) );
  BUF_X2 U11180 ( .A(n11283), .Z(n14144) );
  CLKBUF_X3 U11181 ( .A(n10138), .Z(n9609) );
  AND2_X2 U11182 ( .A1(n11184), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13479) );
  AND2_X1 U11183 ( .A1(n13475), .A2(n11192), .ZN(n11361) );
  NOR2_X1 U11184 ( .A1(n10473), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10826) );
  INV_X2 U11185 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10472) );
  AND2_X1 U11186 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11192) );
  INV_X1 U11187 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10547) );
  NOR2_X1 U11188 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13443) );
  XNOR2_X1 U11189 ( .A(n14271), .B(n14165), .ZN(n14452) );
  AOI211_X1 U11190 ( .C1(n16108), .C2(n18669), .A(n15080), .B(n15079), .ZN(
        n15081) );
  AOI21_X1 U11191 ( .B1(n14305), .B2(n14496), .A(n14286), .ZN(n14488) );
  AND2_X1 U11192 ( .A1(n14303), .A2(n10046), .ZN(n12143) );
  INV_X1 U11193 ( .A(n14414), .ZN(n15680) );
  AND2_X1 U11194 ( .A1(n12852), .A2(n9855), .ZN(n9854) );
  AND2_X1 U11195 ( .A1(n14460), .A2(n9774), .ZN(n9675) );
  AOI211_X1 U11196 ( .C1(n16108), .C2(n15004), .A(n15003), .B(n15002), .ZN(
        n15005) );
  OAI21_X1 U11197 ( .B1(n15160), .B2(n9843), .A(n9672), .ZN(n9840) );
  AND2_X1 U11198 ( .A1(n9740), .A2(n9738), .ZN(n15302) );
  AOI21_X1 U11199 ( .B1(n15097), .B2(n15071), .A(n15089), .ZN(n15249) );
  AND2_X1 U11200 ( .A1(n9606), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12479) );
  AND2_X1 U11201 ( .A1(n15001), .A2(n20763), .ZN(n15160) );
  AND2_X1 U11202 ( .A1(n14501), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11618) );
  NAND2_X1 U11203 ( .A1(n11608), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14521) );
  INV_X2 U11204 ( .A(n9745), .ZN(n15358) );
  NAND2_X1 U11205 ( .A1(n15353), .A2(n12343), .ZN(n9793) );
  NOR2_X1 U11206 ( .A1(n14853), .A2(n14852), .ZN(n14851) );
  XNOR2_X1 U11207 ( .A(n13081), .B(n10090), .ZN(n14853) );
  NAND2_X1 U11208 ( .A1(n15867), .A2(n11573), .ZN(n15860) );
  NAND2_X1 U11209 ( .A1(n14921), .A2(n14920), .ZN(n14919) );
  XNOR2_X1 U11210 ( .A(n14856), .B(n13063), .ZN(n14921) );
  AOI21_X1 U11211 ( .B1(n9599), .B2(n11596), .A(n9673), .ZN(n9968) );
  XNOR2_X1 U11212 ( .A(n12311), .B(n12828), .ZN(n15119) );
  NAND2_X1 U11213 ( .A1(n10001), .A2(n10004), .ZN(n14856) );
  NAND2_X1 U11214 ( .A1(n9791), .A2(n12310), .ZN(n15120) );
  NOR3_X1 U11215 ( .A1(n17270), .A2(n17271), .A3(n17428), .ZN(n17269) );
  OR2_X1 U11216 ( .A1(n14868), .A2(n10005), .ZN(n10001) );
  NOR2_X1 U11217 ( .A1(n15864), .A2(n9975), .ZN(n9974) );
  AND2_X1 U11218 ( .A1(n14559), .A2(n14557), .ZN(n14535) );
  NOR2_X2 U11219 ( .A1(n14878), .A2(n10015), .ZN(n13020) );
  INV_X2 U11220 ( .A(n9634), .ZN(n14539) );
  INV_X2 U11221 ( .A(n9634), .ZN(n14705) );
  XNOR2_X1 U11222 ( .A(n11591), .B(n11576), .ZN(n11725) );
  NAND2_X1 U11223 ( .A1(n10067), .A2(n12278), .ZN(n12274) );
  NAND2_X1 U11224 ( .A1(n13511), .A2(n11467), .ZN(n11494) );
  NAND2_X1 U11225 ( .A1(n17483), .A2(n10214), .ZN(n17422) );
  AND2_X1 U11226 ( .A1(n11565), .A2(n11539), .ZN(n11706) );
  INV_X1 U11227 ( .A(n13521), .ZN(n13590) );
  OAI21_X1 U11228 ( .B1(n11701), .B2(n11811), .A(n11700), .ZN(n13586) );
  NAND2_X1 U11229 ( .A1(n11538), .A2(n11490), .ZN(n11701) );
  NAND2_X1 U11230 ( .A1(n12271), .A2(n12270), .ZN(n12465) );
  INV_X1 U11231 ( .A(n17529), .ZN(n17494) );
  CLKBUF_X1 U11232 ( .A(n13521), .Z(n9625) );
  XNOR2_X1 U11233 ( .A(n11538), .B(n11534), .ZN(n11716) );
  AND2_X1 U11234 ( .A1(n9807), .A2(n9644), .ZN(n14782) );
  AND2_X1 U11235 ( .A1(n12247), .A2(n12246), .ZN(n12278) );
  OR3_X1 U11236 ( .A1(n12268), .A2(n12267), .A3(n12266), .ZN(n12271) );
  NOR2_X1 U11237 ( .A1(n16681), .A2(n16762), .ZN(n16744) );
  NAND2_X1 U11238 ( .A1(n13415), .A2(n13414), .ZN(n13413) );
  NAND2_X1 U11239 ( .A1(n11680), .A2(n11679), .ZN(n13415) );
  INV_X1 U11240 ( .A(n19174), .ZN(n12201) );
  INV_X1 U11241 ( .A(n12256), .ZN(n12205) );
  AND2_X1 U11242 ( .A1(n12882), .A2(n12880), .ZN(n10000) );
  OAI21_X1 U11243 ( .B1(n13391), .B2(n13392), .A(n12869), .ZN(n13381) );
  NOR2_X2 U11244 ( .A1(n12204), .A2(n13653), .ZN(n12248) );
  INV_X1 U11245 ( .A(n19114), .ZN(n19110) );
  AND2_X1 U11246 ( .A1(n12199), .A2(n19007), .ZN(n12202) );
  NAND2_X1 U11247 ( .A1(n12179), .A2(n14238), .ZN(n19382) );
  AND2_X1 U11248 ( .A1(n12188), .A2(n14238), .ZN(n12253) );
  NAND2_X1 U11249 ( .A1(n17897), .A2(n17971), .ZN(n17801) );
  NOR2_X2 U11250 ( .A1(n17922), .A2(n18438), .ZN(n17897) );
  AND2_X1 U11251 ( .A1(n14238), .A2(n12203), .ZN(n12168) );
  AND2_X1 U11252 ( .A1(n19007), .A2(n12191), .ZN(n12192) );
  OR2_X1 U11253 ( .A1(n14073), .A2(n14089), .ZN(n14091) );
  AND2_X1 U11254 ( .A1(n12590), .A2(n14260), .ZN(n12723) );
  NAND2_X1 U11255 ( .A1(n11425), .A2(n11426), .ZN(n11468) );
  BUF_X2 U11256 ( .A(n12857), .Z(n9626) );
  NAND2_X1 U11257 ( .A1(n9772), .A2(n9670), .ZN(n11681) );
  OAI21_X1 U11258 ( .B1(n18871), .B2(n12874), .A(n12864), .ZN(n13345) );
  AOI21_X2 U11259 ( .B1(n14128), .B2(n15457), .A(n10352), .ZN(n18427) );
  XNOR2_X1 U11260 ( .A(n9973), .B(n11389), .ZN(n11684) );
  NAND2_X1 U11261 ( .A1(n12411), .A2(n12340), .ZN(n12331) );
  OR2_X1 U11262 ( .A1(n12764), .A2(n12763), .ZN(n13631) );
  OR2_X1 U11263 ( .A1(n9728), .A2(n9727), .ZN(n10423) );
  OR2_X1 U11264 ( .A1(n14126), .A2(n9678), .ZN(n9907) );
  NOR2_X1 U11265 ( .A1(n12315), .A2(n9953), .ZN(n12330) );
  NAND2_X1 U11266 ( .A1(n10648), .A2(n10626), .ZN(n9614) );
  AND2_X1 U11267 ( .A1(n12608), .A2(n12607), .ZN(n13500) );
  OR2_X1 U11268 ( .A1(n10660), .A2(n16155), .ZN(n10677) );
  AND2_X1 U11269 ( .A1(n9988), .A2(n9983), .ZN(n9982) );
  NAND2_X1 U11270 ( .A1(n10601), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10660) );
  OR2_X1 U11271 ( .A1(n12505), .A2(n17199), .ZN(n9758) );
  NAND2_X1 U11272 ( .A1(n11326), .A2(n13409), .ZN(n12586) );
  NOR2_X1 U11273 ( .A1(n17598), .A2(n10195), .ZN(n17591) );
  AOI21_X1 U11274 ( .B1(n11444), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10027), 
        .ZN(n10026) );
  NOR2_X1 U11275 ( .A1(n10347), .A2(n9759), .ZN(n17199) );
  CLKBUF_X2 U11276 ( .A(n10760), .Z(n9621) );
  CLKBUF_X3 U11277 ( .A(n10760), .Z(n9622) );
  MUX2_X1 U11278 ( .A(n12435), .B(P2_EBX_REG_2__SCAN_IN), .S(n19061), .Z(
        n12293) );
  NAND2_X1 U11279 ( .A1(n10621), .A2(n12769), .ZN(n12811) );
  NAND2_X1 U11280 ( .A1(n9761), .A2(n9760), .ZN(n9759) );
  MUX2_X1 U11281 ( .A(n12210), .B(n11147), .S(n19731), .Z(n12435) );
  NAND2_X1 U11282 ( .A1(n11343), .A2(n11324), .ZN(n12704) );
  INV_X1 U11283 ( .A(n12821), .ZN(n15557) );
  INV_X2 U11284 ( .A(n12280), .ZN(n12548) );
  NAND2_X1 U11285 ( .A1(n19731), .A2(n13639), .ZN(n12776) );
  NAND2_X1 U11286 ( .A1(n17993), .A2(n17983), .ZN(n10346) );
  NOR2_X1 U11287 ( .A1(n17115), .A2(n10199), .ZN(n10203) );
  INV_X1 U11288 ( .A(n10332), .ZN(n17993) );
  INV_X1 U11289 ( .A(n10345), .ZN(n17975) );
  OR2_X1 U11290 ( .A1(n11390), .A2(n20012), .ZN(n11652) );
  NAND3_X1 U11291 ( .A1(n10330), .A2(n10329), .A3(n10328), .ZN(n16992) );
  AND2_X1 U11292 ( .A1(n10806), .A2(n12743), .ZN(n10637) );
  AND2_X1 U11293 ( .A1(n20044), .A2(n11310), .ZN(n13425) );
  NAND2_X1 U11294 ( .A1(n10577), .A2(n10841), .ZN(n13639) );
  OR2_X1 U11295 ( .A1(n10594), .A2(n10593), .ZN(n10595) );
  NOR2_X2 U11296 ( .A1(n20029), .A2(n11340), .ZN(n13557) );
  AND2_X1 U11297 ( .A1(n10578), .A2(n13188), .ZN(n9736) );
  INV_X1 U11298 ( .A(n10841), .ZN(n10806) );
  NAND2_X1 U11299 ( .A1(n10578), .A2(n10612), .ZN(n10620) );
  NAND2_X1 U11300 ( .A1(n9656), .A2(n10087), .ZN(n17620) );
  CLKBUF_X2 U11301 ( .A(n10612), .Z(n13165) );
  NAND4_X1 U11302 ( .A1(n9660), .A2(n9908), .A3(n10288), .A4(n10287), .ZN(
        n17032) );
  INV_X1 U11303 ( .A(n11305), .ZN(n12580) );
  CLKBUF_X1 U11304 ( .A(n11325), .Z(n20036) );
  OR2_X1 U11305 ( .A1(n11382), .A2(n11381), .ZN(n11409) );
  OR2_X1 U11306 ( .A1(n11402), .A2(n11401), .ZN(n11581) );
  INV_X1 U11307 ( .A(n10614), .ZN(n19045) );
  NOR2_X2 U11308 ( .A1(n10134), .A2(n10133), .ZN(n17124) );
  INV_X1 U11310 ( .A(n10611), .ZN(n19071) );
  AND4_X1 U11311 ( .A1(n10148), .A2(n10147), .A3(n10146), .A4(n10145), .ZN(
        n10149) );
  NAND2_X2 U11312 ( .A1(n10493), .A2(n10492), .ZN(n12785) );
  NAND2_X1 U11313 ( .A1(n10097), .A2(n11200), .ZN(n11305) );
  NAND2_X1 U11314 ( .A1(n10049), .A2(n10047), .ZN(n10614) );
  INV_X1 U11315 ( .A(n10963), .ZN(n9620) );
  AND2_X1 U11316 ( .A1(n13645), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12743) );
  INV_X1 U11317 ( .A(n10963), .ZN(n9619) );
  NOR2_X2 U11319 ( .A1(n20007), .A2(n20006), .ZN(n20008) );
  AND4_X1 U11320 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11228) );
  AND4_X1 U11321 ( .A1(n11299), .A2(n11298), .A3(n11297), .A4(n11296), .ZN(
        n11300) );
  AND4_X1 U11322 ( .A1(n11295), .A2(n11294), .A3(n11293), .A4(n11292), .ZN(
        n11301) );
  INV_X2 U11323 ( .A(n10240), .ZN(n16903) );
  AND4_X1 U11324 ( .A1(n11204), .A2(n11203), .A3(n11202), .A4(n11201), .ZN(
        n10096) );
  AND4_X1 U11325 ( .A1(n11241), .A2(n11240), .A3(n11239), .A4(n11238), .ZN(
        n11258) );
  AND4_X1 U11326 ( .A1(n11245), .A2(n11244), .A3(n11243), .A4(n11242), .ZN(
        n11257) );
  AND4_X1 U11327 ( .A1(n11268), .A2(n11267), .A3(n11266), .A4(n11265), .ZN(
        n11269) );
  AND4_X1 U11328 ( .A1(n11216), .A2(n11215), .A3(n11214), .A4(n11213), .ZN(
        n11227) );
  AND4_X1 U11329 ( .A1(n11220), .A2(n11219), .A3(n11218), .A4(n11217), .ZN(
        n11226) );
  AND4_X1 U11330 ( .A1(n11224), .A2(n11223), .A3(n11222), .A4(n11221), .ZN(
        n11225) );
  AND4_X1 U11331 ( .A1(n11287), .A2(n11286), .A3(n11285), .A4(n11284), .ZN(
        n11303) );
  NAND2_X1 U11332 ( .A1(n10813), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10963) );
  BUF_X2 U11333 ( .A(n11502), .Z(n11355) );
  AND2_X2 U11334 ( .A1(n13146), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10904) );
  BUF_X2 U11335 ( .A(n11392), .Z(n11370) );
  INV_X1 U11336 ( .A(n19689), .ZN(n19617) );
  CLKBUF_X2 U11337 ( .A(n10135), .Z(n16913) );
  CLKBUF_X3 U11338 ( .A(n10150), .Z(n16932) );
  CLKBUF_X2 U11339 ( .A(n10135), .Z(n10299) );
  NAND2_X2 U11340 ( .A1(n19761), .A2(n19634), .ZN(n19678) );
  INV_X1 U11341 ( .A(n10143), .ZN(n10235) );
  BUF_X2 U11342 ( .A(n10311), .Z(n16938) );
  INV_X1 U11343 ( .A(n10136), .ZN(n10240) );
  BUF_X2 U11344 ( .A(n11360), .Z(n12131) );
  NAND2_X2 U11345 ( .A1(n18610), .A2(n18490), .ZN(n18538) );
  AND2_X2 U11346 ( .A1(n13149), .A2(n10547), .ZN(n10851) );
  INV_X1 U11347 ( .A(n18563), .ZN(n18473) );
  INV_X2 U11348 ( .A(n16302), .ZN(n16304) );
  AND2_X2 U11349 ( .A1(n10821), .A2(n13443), .ZN(n10875) );
  INV_X2 U11350 ( .A(n19758), .ZN(n19761) );
  OR2_X1 U11351 ( .A1(n10107), .A2(n16663), .ZN(n10094) );
  BUF_X2 U11352 ( .A(n16697), .Z(n16920) );
  INV_X2 U11353 ( .A(n16622), .ZN(n9607) );
  BUF_X2 U11354 ( .A(n11272), .Z(n14138) );
  BUF_X4 U11355 ( .A(n10114), .Z(n9608) );
  NOR2_X1 U11356 ( .A1(n10102), .A2(n10104), .ZN(n10280) );
  AND2_X2 U11357 ( .A1(n11191), .A2(n11192), .ZN(n14139) );
  NAND2_X1 U11358 ( .A1(n18572), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10107) );
  NAND2_X1 U11359 ( .A1(n18592), .A2(n18598), .ZN(n16663) );
  NAND2_X1 U11360 ( .A1(n10822), .A2(n10785), .ZN(n13027) );
  AND2_X2 U11361 ( .A1(n10827), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10815) );
  NAND2_X2 U11362 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18429) );
  INV_X1 U11363 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18572) );
  OR2_X1 U11364 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10103) );
  INV_X1 U11365 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18592) );
  NOR2_X2 U11366 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11193) );
  NOR2_X2 U11368 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11191) );
  INV_X1 U11369 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19719) );
  INV_X2 U11370 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10785) );
  AND2_X1 U11372 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n12565), .ZN(
        n9611) );
  OAI21_X2 U11373 ( .B1(n9617), .B2(n11811), .A(n11671), .ZN(n11672) );
  AOI21_X1 U11374 ( .B1(n11706), .B2(n11856), .A(n11705), .ZN(n13751) );
  NAND2_X1 U11376 ( .A1(n12471), .A2(n12275), .ZN(n9613) );
  NAND2_X1 U11377 ( .A1(n12393), .A2(n12392), .ZN(n15049) );
  NAND2_X1 U11378 ( .A1(n12471), .A2(n12275), .ZN(n12463) );
  NAND2_X1 U11379 ( .A1(n10648), .A2(n10626), .ZN(n10672) );
  AND2_X1 U11380 ( .A1(n10574), .A2(n10610), .ZN(n10513) );
  OR2_X1 U11381 ( .A1(n10657), .A2(n10656), .ZN(n10658) );
  INV_X1 U11382 ( .A(n10660), .ZN(n9615) );
  INV_X1 U11383 ( .A(n10660), .ZN(n9616) );
  AND2_X4 U11384 ( .A1(n10826), .A2(n10785), .ZN(n10552) );
  XNOR2_X1 U11385 ( .A(n11468), .B(n20159), .ZN(n20666) );
  INV_X2 U11386 ( .A(n11325), .ZN(n11309) );
  NAND3_X2 U11387 ( .A1(n11719), .A2(n11718), .A3(n11717), .ZN(n13750) );
  NAND2_X2 U11388 ( .A1(n12158), .A2(n12159), .ZN(n12166) );
  BUF_X2 U11389 ( .A(n20009), .Z(n9617) );
  INV_X1 U11390 ( .A(n10963), .ZN(n9618) );
  OAI211_X2 U11391 ( .C1(n11327), .C2(n11316), .A(n11315), .B(n11314), .ZN(
        n11317) );
  NOR2_X2 U11392 ( .A1(n11341), .A2(n11309), .ZN(n11327) );
  AND2_X2 U11393 ( .A1(n13479), .A2(n11191), .ZN(n11503) );
  NAND2_X1 U11394 ( .A1(n10616), .A2(n9996), .ZN(n19737) );
  NAND2_X2 U11395 ( .A1(n14337), .A2(n14338), .ZN(n14336) );
  NAND2_X1 U11396 ( .A1(n12286), .A2(n12287), .ZN(n12446) );
  NOR2_X2 U11397 ( .A1(n14561), .A2(n11599), .ZN(n14702) );
  AND2_X1 U11398 ( .A1(n13475), .A2(n11192), .ZN(n9623) );
  AND2_X1 U11399 ( .A1(n13475), .A2(n11192), .ZN(n9624) );
  NAND2_X1 U11400 ( .A1(n11682), .A2(n20040), .ZN(n11341) );
  XNOR2_X1 U11401 ( .A(n11413), .B(n11412), .ZN(n19941) );
  AND2_X2 U11402 ( .A1(n14314), .A2(n15720), .ZN(n14364) );
  NAND2_X2 U11404 ( .A1(n11588), .A2(n11587), .ZN(n14010) );
  XNOR2_X2 U11405 ( .A(n12434), .B(n12433), .ZN(n15142) );
  NOR2_X2 U11406 ( .A1(n15165), .A2(n12428), .ZN(n12434) );
  NOR2_X2 U11407 ( .A1(n12875), .A2(n12177), .ZN(n12200) );
  NAND2_X2 U11408 ( .A1(n12583), .A2(n14251), .ZN(n12592) );
  AND2_X2 U11409 ( .A1(n12713), .A2(n12593), .ZN(n12583) );
  NOR2_X2 U11410 ( .A1(n14998), .A2(n20763), .ZN(n15165) );
  NAND2_X2 U11411 ( .A1(n12426), .A2(n10095), .ZN(n14998) );
  OAI21_X1 U11412 ( .B1(n12875), .B2(n12874), .A(n12873), .ZN(n12881) );
  AND2_X1 U11413 ( .A1(n12875), .A2(n18871), .ZN(n12199) );
  NAND2_X2 U11414 ( .A1(n11335), .A2(n11331), .ZN(n11419) );
  NAND2_X2 U11415 ( .A1(n11319), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11335) );
  NAND3_X2 U11416 ( .A1(n11617), .A2(n9770), .A3(n11616), .ZN(n14455) );
  OR2_X4 U11417 ( .A1(n11282), .A2(n11281), .ZN(n11310) );
  AOI21_X2 U11418 ( .B1(n14287), .B2(n14304), .A(n12143), .ZN(n14479) );
  NOR2_X2 U11419 ( .A1(n14470), .A2(n9719), .ZN(n14469) );
  NAND2_X2 U11420 ( .A1(n11614), .A2(n15811), .ZN(n14470) );
  AND2_X1 U11421 ( .A1(n11193), .A2(n11191), .ZN(n9627) );
  AND2_X1 U11422 ( .A1(n11194), .A2(n11193), .ZN(n9628) );
  NOR2_X1 U11423 ( .A1(n14127), .A2(n18430), .ZN(n18419) );
  BUF_X2 U11424 ( .A(n11391), .Z(n9630) );
  BUF_X4 U11425 ( .A(n11391), .Z(n9631) );
  NOR2_X4 U11426 ( .A1(n14336), .A2(n14494), .ZN(n14303) );
  NAND2_X2 U11427 ( .A1(n11429), .A2(n20057), .ZN(n13829) );
  NAND2_X2 U11428 ( .A1(n20120), .A2(n11354), .ZN(n20057) );
  OR2_X1 U11429 ( .A1(n11340), .A2(n20012), .ZN(n12604) );
  NOR2_X1 U11430 ( .A1(n19855), .A2(n20709), .ZN(n19883) );
  AND4_X1 U11431 ( .A1(n10971), .A2(n10970), .A3(n10969), .A4(n10968), .ZN(
        n10978) );
  AND4_X1 U11432 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n10976) );
  AOI21_X1 U11433 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20778), .A(
        n10250), .ZN(n10356) );
  NOR2_X1 U11434 ( .A1(n10352), .A2(n9905), .ZN(n18411) );
  AND2_X1 U11435 ( .A1(n15457), .A2(n10351), .ZN(n9905) );
  NAND2_X1 U11436 ( .A1(n12788), .A2(n13460), .ZN(n12850) );
  CLKBUF_X1 U11437 ( .A(n9631), .Z(n14145) );
  AND4_X1 U11438 ( .A1(n10967), .A2(n10966), .A3(n10965), .A4(n10964), .ZN(
        n10979) );
  OAI21_X1 U11439 ( .B1(n9830), .B2(n9829), .A(n12821), .ZN(n9828) );
  AND2_X1 U11440 ( .A1(n12123), .A2(n12096), .ZN(n10046) );
  INV_X1 U11441 ( .A(n14287), .ZN(n12123) );
  NAND2_X1 U11442 ( .A1(n14612), .A2(n9708), .ZN(n9782) );
  INV_X1 U11443 ( .A(n14297), .ZN(n9778) );
  NAND2_X1 U11444 ( .A1(n11445), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9773) );
  AND2_X1 U11445 ( .A1(n9689), .A2(n11159), .ZN(n9951) );
  OR2_X1 U11446 ( .A1(n12315), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n9960) );
  OR2_X1 U11447 ( .A1(n11151), .A2(n9947), .ZN(n9945) );
  NOR2_X1 U11448 ( .A1(n11150), .A2(n9948), .ZN(n9947) );
  INV_X1 U11449 ( .A(n12298), .ZN(n9948) );
  NOR2_X1 U11450 ( .A1(n12296), .A2(n12291), .ZN(n11149) );
  INV_X1 U11451 ( .A(n10620), .ZN(n9832) );
  NAND2_X1 U11452 ( .A1(n15557), .A2(n19028), .ZN(n12765) );
  INV_X1 U11453 ( .A(n9896), .ZN(n9890) );
  INV_X1 U11454 ( .A(n14989), .ZN(n9904) );
  NAND2_X1 U11455 ( .A1(n9792), .A2(n15066), .ZN(n15068) );
  NAND2_X1 U11456 ( .A1(n9793), .A2(n15354), .ZN(n9792) );
  INV_X1 U11457 ( .A(n9845), .ZN(n9844) );
  AOI21_X1 U11458 ( .B1(n15044), .B2(n10055), .A(n9694), .ZN(n10054) );
  INV_X1 U11459 ( .A(n15047), .ZN(n10055) );
  NAND2_X1 U11460 ( .A1(n15120), .A2(n15119), .ZN(n12313) );
  NAND2_X1 U11461 ( .A1(n12472), .A2(n12548), .ZN(n12474) );
  INV_X1 U11462 ( .A(n12471), .ZN(n12472) );
  BUF_X1 U11463 ( .A(n12808), .Z(n12403) );
  INV_X1 U11464 ( .A(n10349), .ZN(n9757) );
  AOI211_X1 U11465 ( .C1(n17979), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        n12506) );
  AOI21_X1 U11466 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n15628) );
  OR2_X1 U11467 ( .A1(n16311), .A2(n18620), .ZN(n9916) );
  NAND2_X1 U11468 ( .A1(n17199), .A2(n18619), .ZN(n9917) );
  INV_X1 U11469 ( .A(n19763), .ZN(n14260) );
  NAND2_X1 U11470 ( .A1(n9974), .A2(n13833), .ZN(n15867) );
  INV_X1 U11471 ( .A(n11549), .ZN(n9975) );
  INV_X1 U11472 ( .A(n9945), .ZN(n12307) );
  NAND2_X1 U11473 ( .A1(n11149), .A2(n11148), .ZN(n12308) );
  NAND2_X1 U11474 ( .A1(n13020), .A2(n10002), .ZN(n10004) );
  NOR2_X1 U11475 ( .A1(n14857), .A2(n10003), .ZN(n10002) );
  AND2_X1 U11476 ( .A1(n10841), .A2(n19700), .ZN(n13342) );
  NAND2_X1 U11477 ( .A1(n15097), .A2(n9800), .ZN(n9797) );
  NOR2_X1 U11478 ( .A1(n15073), .A2(n9801), .ZN(n9800) );
  INV_X1 U11479 ( .A(n15071), .ZN(n9801) );
  AOI21_X1 U11480 ( .B1(n12535), .B2(n9900), .A(n9901), .ZN(n9899) );
  NAND2_X1 U11481 ( .A1(n9797), .A2(n9796), .ZN(n15229) );
  NOR2_X1 U11482 ( .A1(n9798), .A2(n9802), .ZN(n9796) );
  NAND2_X1 U11483 ( .A1(n15077), .A2(n15230), .ZN(n9802) );
  NOR2_X1 U11484 ( .A1(n15333), .A2(n9739), .ZN(n9738) );
  NAND2_X1 U11485 ( .A1(n9742), .A2(n9741), .ZN(n9740) );
  AND2_X1 U11486 ( .A1(n19002), .A2(n15315), .ZN(n9739) );
  INV_X1 U11487 ( .A(n13361), .ZN(n9928) );
  NAND2_X1 U11488 ( .A1(n12447), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9746) );
  NAND2_X1 U11489 ( .A1(n13894), .A2(n13955), .ZN(n9878) );
  CLKBUF_X1 U11490 ( .A(n10780), .Z(n13632) );
  AOI21_X1 U11491 ( .B1(n12872), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12863), .ZN(n12864) );
  INV_X1 U11492 ( .A(n16167), .ZN(n13460) );
  INV_X1 U11493 ( .A(n19416), .ZN(n19690) );
  NOR3_X1 U11494 ( .A1(n17199), .A2(n14126), .A3(n18433), .ZN(n18402) );
  AOI211_X1 U11495 ( .C1(n9604), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n10327), .B(n10326), .ZN(n10328) );
  NAND2_X1 U11496 ( .A1(n17362), .A2(n9995), .ZN(n17304) );
  AND2_X1 U11497 ( .A1(n10221), .A2(n17676), .ZN(n9995) );
  AND2_X2 U11498 ( .A1(n20012), .A2(n12599), .ZN(n14251) );
  NAND2_X2 U11499 ( .A1(n10806), .A2(n13645), .ZN(n19731) );
  NOR2_X1 U11500 ( .A1(n9842), .A2(n20763), .ZN(n9841) );
  INV_X1 U11501 ( .A(n15162), .ZN(n9842) );
  INV_X1 U11502 ( .A(n11636), .ZN(n11632) );
  NAND2_X1 U11503 ( .A1(n19033), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12174) );
  AOI22_X1 U11504 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10518) );
  NAND2_X1 U11505 ( .A1(n12694), .A2(n9786), .ZN(n9785) );
  NAND2_X1 U11506 ( .A1(n11533), .A2(n11532), .ZN(n11565) );
  AND2_X1 U11507 ( .A1(n11534), .A2(n11535), .ZN(n11532) );
  AND2_X1 U11508 ( .A1(n11561), .A2(n11560), .ZN(n11564) );
  NOR2_X1 U11509 ( .A1(n11440), .A2(n11439), .ZN(n11491) );
  OR2_X1 U11510 ( .A1(n20036), .A2(n20702), .ZN(n11473) );
  AOI21_X1 U11511 ( .B1(n20673), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11625), .ZN(n11624) );
  INV_X1 U11512 ( .A(n11652), .ZN(n11656) );
  AOI21_X1 U11513 ( .B1(n10661), .B2(P2_EBX_REG_1__SCAN_IN), .A(n10632), .ZN(
        n10635) );
  NOR2_X1 U11514 ( .A1(n15633), .A2(n9934), .ZN(n9933) );
  INV_X1 U11515 ( .A(n14962), .ZN(n9934) );
  INV_X1 U11516 ( .A(n12279), .ZN(n10067) );
  NAND2_X1 U11517 ( .A1(n9886), .A2(n9882), .ZN(n9881) );
  INV_X1 U11518 ( .A(n13955), .ZN(n9882) );
  OAI211_X1 U11519 ( .C1(n10675), .C2(n13394), .A(n10663), .B(n10662), .ZN(
        n10664) );
  INV_X1 U11520 ( .A(n14160), .ZN(n12140) );
  NOR2_X1 U11521 ( .A1(n14363), .A2(n10042), .ZN(n10041) );
  INV_X1 U11522 ( .A(n14365), .ZN(n10042) );
  NOR2_X1 U11523 ( .A1(n9966), .A2(n11607), .ZN(n9965) );
  INV_X1 U11524 ( .A(n9968), .ZN(n9966) );
  INV_X1 U11525 ( .A(n14377), .ZN(n11915) );
  OR2_X1 U11526 ( .A1(n14742), .A2(n20702), .ZN(n14160) );
  NAND2_X1 U11527 ( .A1(n10034), .A2(n11863), .ZN(n10033) );
  INV_X1 U11528 ( .A(n14386), .ZN(n10034) );
  NAND2_X1 U11529 ( .A1(n14166), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12112) );
  NAND2_X1 U11530 ( .A1(n11387), .A2(n11386), .ZN(n11413) );
  NAND2_X1 U11531 ( .A1(n9976), .A2(n14705), .ZN(n14501) );
  NOR2_X1 U11532 ( .A1(n9979), .A2(n14663), .ZN(n9977) );
  OR2_X1 U11533 ( .A1(n11446), .A2(n20702), .ZN(n11589) );
  INV_X1 U11535 ( .A(n12694), .ZN(n12686) );
  OR2_X1 U11536 ( .A1(n11484), .A2(n11483), .ZN(n11542) );
  INV_X1 U11537 ( .A(n9788), .ZN(n9787) );
  NOR2_X2 U11538 ( .A1(n12601), .A2(n12623), .ZN(n12696) );
  NAND2_X1 U11539 ( .A1(n20036), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11390) );
  INV_X1 U11540 ( .A(n20059), .ZN(n20164) );
  AND2_X1 U11541 ( .A1(n13571), .A2(n13570), .ZN(n13574) );
  NOR2_X2 U11542 ( .A1(n12406), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12413) );
  NOR2_X1 U11543 ( .A1(n9955), .A2(n9954), .ZN(n9953) );
  NOR2_X1 U11544 ( .A1(n9956), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n9954) );
  AND2_X1 U11545 ( .A1(n12403), .A2(n9958), .ZN(n9955) );
  INV_X1 U11546 ( .A(n13101), .ZN(n10013) );
  OAI21_X1 U11547 ( .B1(n14853), .B2(n10011), .A(n10010), .ZN(n13104) );
  NAND2_X1 U11548 ( .A1(n10013), .A2(n10012), .ZN(n10011) );
  NAND2_X1 U11549 ( .A1(n10082), .A2(n10013), .ZN(n10010) );
  INV_X1 U11550 ( .A(n14852), .ZN(n10012) );
  NOR2_X1 U11551 ( .A1(n10958), .A2(n10957), .ZN(n12269) );
  AND2_X1 U11552 ( .A1(n13340), .A2(n13231), .ZN(n13099) );
  NAND2_X1 U11553 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9806) );
  OR2_X1 U11554 ( .A1(n10444), .A2(n15000), .ZN(n10443) );
  NAND2_X1 U11555 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U11556 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9825) );
  OR2_X1 U11557 ( .A1(n9871), .A2(n13903), .ZN(n9870) );
  INV_X1 U11558 ( .A(n13763), .ZN(n9871) );
  NOR2_X1 U11559 ( .A1(n15113), .A2(n9823), .ZN(n9822) );
  NOR2_X1 U11560 ( .A1(n9927), .A2(n9926), .ZN(n9925) );
  INV_X1 U11561 ( .A(n14776), .ZN(n9926) );
  INV_X1 U11562 ( .A(n14909), .ZN(n9927) );
  NAND2_X1 U11563 ( .A1(n15977), .A2(n12548), .ZN(n12420) );
  OR2_X1 U11564 ( .A1(n15996), .A2(n12280), .ZN(n15008) );
  NAND2_X1 U11565 ( .A1(n9861), .A2(n14818), .ZN(n9860) );
  INV_X1 U11566 ( .A(n15061), .ZN(n9861) );
  AND2_X1 U11567 ( .A1(n12378), .A2(n9874), .ZN(n9873) );
  NAND2_X1 U11568 ( .A1(n12343), .A2(n15378), .ZN(n9874) );
  OR2_X1 U11569 ( .A1(n15323), .A2(n15318), .ZN(n15065) );
  OAI21_X1 U11570 ( .B1(n15073), .B2(n9799), .A(n15072), .ZN(n9798) );
  INV_X1 U11571 ( .A(n15089), .ZN(n9799) );
  NAND2_X1 U11572 ( .A1(n15292), .A2(n18996), .ZN(n9741) );
  OR2_X1 U11573 ( .A1(n9938), .A2(n15304), .ZN(n9937) );
  OR2_X1 U11574 ( .A1(n16118), .A2(n9939), .ZN(n9938) );
  INV_X1 U11575 ( .A(n13811), .ZN(n9939) );
  NAND2_X1 U11576 ( .A1(n12323), .A2(n10062), .ZN(n10061) );
  INV_X1 U11577 ( .A(n15405), .ZN(n10062) );
  NOR2_X1 U11578 ( .A1(n9851), .A2(n9849), .ZN(n9848) );
  INV_X1 U11579 ( .A(n13539), .ZN(n9849) );
  NAND2_X1 U11580 ( .A1(n13545), .A2(n13597), .ZN(n9851) );
  NAND2_X1 U11581 ( .A1(n9880), .A2(n9885), .ZN(n9877) );
  NAND2_X1 U11582 ( .A1(n10649), .A2(n9828), .ZN(n10615) );
  NAND2_X1 U11583 ( .A1(n12776), .A2(n10599), .ZN(n13437) );
  AND3_X1 U11584 ( .A1(n10598), .A2(n19045), .A3(n10578), .ZN(n10599) );
  NAND2_X1 U11585 ( .A1(n12182), .A2(n12200), .ZN(n12212) );
  NAND2_X1 U11586 ( .A1(n12200), .A2(n19007), .ZN(n12204) );
  AND4_X1 U11587 ( .A1(n12781), .A2(n12812), .A3(n12780), .A4(n12779), .ZN(
        n13454) );
  AOI221_X1 U11588 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10799), 
        .C1(n15561), .C2(n10799), .A(n10798), .ZN(n12762) );
  NOR2_X1 U11589 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13672) );
  NAND2_X1 U11590 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10105) );
  NOR3_X1 U11591 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18572), .A3(
        n18432), .ZN(n10138) );
  NOR2_X1 U11592 ( .A1(n10102), .A2(n10103), .ZN(n10114) );
  NOR2_X1 U11593 ( .A1(n17124), .A2(n10371), .ZN(n10197) );
  NOR3_X1 U11594 ( .A1(n15456), .A2(n10362), .A3(n10361), .ZN(n12507) );
  INV_X1 U11595 ( .A(n20706), .ZN(n13803) );
  OR2_X1 U11596 ( .A1(n15801), .A2(n13428), .ZN(n14123) );
  AND2_X1 U11597 ( .A1(n20700), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14163) );
  CLKBUF_X1 U11598 ( .A(n11685), .Z(n14164) );
  AND2_X1 U11599 ( .A1(n13789), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14137) );
  AND2_X1 U11600 ( .A1(n14303), .A2(n10043), .ZN(n14271) );
  AND2_X1 U11601 ( .A1(n10045), .A2(n10044), .ZN(n10043) );
  INV_X1 U11602 ( .A(n14273), .ZN(n10044) );
  INV_X1 U11603 ( .A(n14055), .ZN(n11845) );
  NAND2_X1 U11604 ( .A1(n11720), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11726) );
  AOI21_X1 U11605 ( .B1(n11716), .B2(n11856), .A(n11715), .ZN(n13752) );
  AND2_X1 U11606 ( .A1(n14252), .A2(n11667), .ZN(n15590) );
  NAND2_X1 U11607 ( .A1(n9611), .A2(n12566), .ZN(n14460) );
  INV_X1 U11608 ( .A(n14481), .ZN(n11617) );
  NOR2_X2 U11609 ( .A1(n14355), .A2(n14348), .ZN(n14347) );
  NAND2_X1 U11610 ( .A1(n14656), .A2(n9709), .ZN(n14361) );
  AND2_X1 U11611 ( .A1(n14654), .A2(n14653), .ZN(n14656) );
  NOR2_X2 U11612 ( .A1(n14091), .A2(n14057), .ZN(n14111) );
  AND2_X1 U11613 ( .A1(n12650), .A2(n12642), .ZN(n9783) );
  NAND2_X1 U11614 ( .A1(n9971), .A2(n9970), .ZN(n9969) );
  INV_X1 U11615 ( .A(n14010), .ZN(n9971) );
  NAND2_X1 U11616 ( .A1(n9777), .A2(n9642), .ZN(n13754) );
  NAND2_X1 U11617 ( .A1(n9674), .A2(n9773), .ZN(n9771) );
  AND2_X1 U11618 ( .A1(n20164), .A2(n20352), .ZN(n20478) );
  INV_X1 U11619 ( .A(n20443), .ZN(n20470) );
  OAI221_X2 U11620 ( .B1(n20703), .B2(n14753), .C1(n13578), .C2(n14753), .A(
        n20702), .ZN(n20059) );
  NAND2_X1 U11621 ( .A1(n9819), .A2(n13945), .ZN(n9818) );
  INV_X1 U11622 ( .A(n14993), .ZN(n9817) );
  OR2_X1 U11623 ( .A1(n15969), .A2(n15970), .ZN(n9819) );
  NAND2_X1 U11624 ( .A1(n9808), .A2(n9711), .ZN(n9807) );
  INV_X1 U11625 ( .A(n16031), .ZN(n9810) );
  NAND2_X1 U11626 ( .A1(n10466), .A2(n15019), .ZN(n9809) );
  AND2_X1 U11627 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  NAND2_X1 U11628 ( .A1(n13945), .A2(n16040), .ZN(n9814) );
  NAND2_X1 U11629 ( .A1(n12373), .A2(n9951), .ZN(n12354) );
  INV_X1 U11630 ( .A(n12315), .ZN(n9957) );
  NOR2_X1 U11631 ( .A1(n12308), .A2(n9696), .ZN(n12284) );
  INV_X1 U11632 ( .A(n12281), .ZN(n9946) );
  AND2_X1 U11633 ( .A1(n10724), .A2(n10723), .ZN(n13994) );
  NAND2_X1 U11634 ( .A1(n13926), .A2(n15101), .ZN(n15100) );
  AND2_X1 U11635 ( .A1(n12885), .A2(n13589), .ZN(n12886) );
  INV_X1 U11636 ( .A(n12978), .ZN(n13013) );
  INV_X1 U11637 ( .A(n11140), .ZN(n12803) );
  OR2_X1 U11638 ( .A1(n14868), .A2(n14867), .ZN(n10007) );
  NAND2_X1 U11639 ( .A1(n10017), .A2(n10016), .ZN(n10015) );
  INV_X1 U11640 ( .A(n14945), .ZN(n10016) );
  AND4_X1 U11641 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n13387) );
  NOR2_X1 U11642 ( .A1(n10622), .A2(n12768), .ZN(n13162) );
  NAND2_X1 U11643 ( .A1(n10840), .A2(n10886), .ZN(n13337) );
  AND2_X1 U11644 ( .A1(n10836), .A2(n10835), .ZN(n10840) );
  AND2_X1 U11645 ( .A1(n13337), .A2(n13336), .ZN(n13339) );
  CLKBUF_X1 U11646 ( .A(n12765), .Z(n12766) );
  NAND2_X1 U11647 ( .A1(n13631), .A2(n13231), .ZN(n13319) );
  NAND2_X1 U11648 ( .A1(n12537), .A2(n9893), .ZN(n9887) );
  NOR2_X1 U11649 ( .A1(n9896), .A2(n9894), .ZN(n9893) );
  NOR2_X1 U11650 ( .A1(n9896), .A2(n9892), .ZN(n9891) );
  INV_X1 U11651 ( .A(n9889), .ZN(n9888) );
  INV_X1 U11652 ( .A(n9900), .ZN(n9892) );
  NAND2_X1 U11653 ( .A1(n10449), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10465) );
  INV_X1 U11654 ( .A(n9798), .ZN(n9795) );
  NAND2_X1 U11655 ( .A1(n15279), .A2(n14877), .ZN(n15060) );
  OR2_X1 U11656 ( .A1(n15100), .A2(n13994), .ZN(n15278) );
  AND2_X1 U11657 ( .A1(n10729), .A2(n10728), .ZN(n15277) );
  NOR2_X1 U11658 ( .A1(n15278), .A2(n15277), .ZN(n15279) );
  NAND2_X1 U11659 ( .A1(n10450), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10464) );
  INV_X1 U11660 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18703) );
  AND2_X1 U11661 ( .A1(n10708), .A2(n10707), .ZN(n13820) );
  NAND2_X1 U11662 ( .A1(n10461), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10460) );
  AND2_X1 U11663 ( .A1(n10698), .A2(n10697), .ZN(n15396) );
  NAND2_X1 U11664 ( .A1(n14789), .A2(n9923), .ZN(n14765) );
  AND2_X1 U11665 ( .A1(n9707), .A2(n14766), .ZN(n9923) );
  NOR2_X1 U11666 ( .A1(n14765), .A2(n11141), .ZN(n12806) );
  NAND2_X1 U11667 ( .A1(n10070), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10068) );
  AND2_X1 U11668 ( .A1(n14789), .A2(n9707), .ZN(n14894) );
  OR2_X1 U11669 ( .A1(n14814), .A2(n12398), .ZN(n15047) );
  NOR2_X1 U11670 ( .A1(n10066), .A2(n15636), .ZN(n10065) );
  NOR2_X2 U11671 ( .A1(n15272), .A2(n14970), .ZN(n15271) );
  NAND2_X1 U11672 ( .A1(n9794), .A2(n12334), .ZN(n15353) );
  INV_X1 U11673 ( .A(n15376), .ZN(n9794) );
  NAND2_X1 U11674 ( .A1(n13591), .A2(n13592), .ZN(n13902) );
  INV_X1 U11675 ( .A(n10061), .ZN(n10058) );
  AND4_X1 U11676 ( .A1(n11035), .A2(n11034), .A3(n11033), .A4(n11032), .ZN(
        n15390) );
  AOI21_X1 U11677 ( .B1(n9835), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n9834), .ZN(n9838) );
  INV_X1 U11678 ( .A(n15108), .ZN(n9834) );
  INV_X1 U11679 ( .A(n12470), .ZN(n9835) );
  OR2_X1 U11680 ( .A1(n10982), .A2(n10981), .ZN(n13361) );
  NAND2_X1 U11681 ( .A1(n15429), .A2(n15430), .ZN(n9791) );
  AOI21_X1 U11682 ( .B1(n13955), .B2(n12548), .A(n16155), .ZN(n9886) );
  NAND2_X1 U11683 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  AND2_X1 U11684 ( .A1(n9922), .A2(n13734), .ZN(n9919) );
  NAND2_X1 U11685 ( .A1(n12868), .A2(n12867), .ZN(n13392) );
  NAND2_X1 U11686 ( .A1(n19320), .A2(n19724), .ZN(n19232) );
  OR3_X1 U11687 ( .A1(n12238), .A2(n19293), .A3(n19549), .ZN(n19262) );
  AND2_X1 U11688 ( .A1(n19320), .A2(n19287), .ZN(n19258) );
  OR2_X1 U11689 ( .A1(n19177), .A2(n19715), .ZN(n19327) );
  NAND2_X1 U11690 ( .A1(n19549), .A2(n19700), .ZN(n19416) );
  AND2_X1 U11691 ( .A1(n12220), .A2(n19440), .ZN(n19447) );
  NAND2_X1 U11692 ( .A1(n19177), .A2(n19712), .ZN(n19451) );
  INV_X1 U11693 ( .A(n19554), .ZN(n19509) );
  OR2_X1 U11694 ( .A1(n19320), .A2(n19287), .ZN(n19504) );
  AND2_X1 U11695 ( .A1(n19177), .A2(n19715), .ZN(n19696) );
  NAND2_X1 U11696 ( .A1(n12487), .A2(n12486), .ZN(n19554) );
  NAND2_X1 U11697 ( .A1(n12764), .A2(n12485), .ZN(n12487) );
  INV_X1 U11698 ( .A(n17276), .ZN(n9734) );
  NOR2_X1 U11699 ( .A1(n16371), .A2(n9658), .ZN(n16370) );
  OAI21_X1 U11700 ( .B1(n16392), .B2(n9688), .A(n9730), .ZN(n16380) );
  NAND2_X1 U11701 ( .A1(n9733), .A2(n17297), .ZN(n9730) );
  NAND2_X1 U11702 ( .A1(n16454), .A2(n10081), .ZN(n16431) );
  AND2_X1 U11703 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n9909) );
  NOR2_X1 U11704 ( .A1(n17968), .A2(n16992), .ZN(n9760) );
  INV_X1 U11705 ( .A(n10346), .ZN(n9761) );
  NAND2_X1 U11706 ( .A1(n9724), .A2(n9722), .ZN(n17379) );
  NOR2_X1 U11707 ( .A1(n17414), .A2(n9723), .ZN(n9722) );
  INV_X1 U11708 ( .A(n17413), .ZN(n9724) );
  NOR2_X1 U11709 ( .A1(n17413), .A2(n17414), .ZN(n17398) );
  NAND2_X1 U11710 ( .A1(n10220), .A2(n10078), .ZN(n10221) );
  NAND2_X1 U11711 ( .A1(n10222), .A2(n10402), .ZN(n10220) );
  INV_X1 U11712 ( .A(n17304), .ZN(n17308) );
  NOR2_X1 U11713 ( .A1(n17408), .A2(n10218), .ZN(n17404) );
  NAND2_X1 U11714 ( .A1(n17409), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10217) );
  INV_X1 U11715 ( .A(n10350), .ZN(n9906) );
  NAND2_X1 U11716 ( .A1(n9989), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9988) );
  INV_X1 U11717 ( .A(n17565), .ZN(n9989) );
  NOR2_X1 U11718 ( .A1(n17552), .A2(n9985), .ZN(n9984) );
  INV_X1 U11719 ( .A(n9987), .ZN(n9985) );
  NAND2_X1 U11720 ( .A1(n17565), .A2(n9990), .ZN(n9987) );
  AND2_X1 U11721 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10200), .ZN(
        n10201) );
  OAI21_X1 U11722 ( .B1(n10357), .B2(n10359), .A(n10356), .ZN(n16311) );
  AND2_X1 U11723 ( .A1(n15659), .A2(n13806), .ZN(n19837) );
  AND2_X1 U11724 ( .A1(n14450), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13806) );
  AND2_X2 U11725 ( .A1(n13412), .A2(n14260), .ZN(n19854) );
  INV_X1 U11726 ( .A(n11310), .ZN(n14166) );
  OR2_X1 U11727 ( .A1(n12143), .A2(n12144), .ZN(n12145) );
  OR2_X1 U11728 ( .A1(n15801), .A2(n13468), .ZN(n14442) );
  INV_X1 U11729 ( .A(n14208), .ZN(n12153) );
  AND2_X1 U11730 ( .A1(n15823), .A2(n12148), .ZN(n15849) );
  AND2_X1 U11731 ( .A1(n15590), .A2(n14260), .ZN(n19935) );
  INV_X1 U11732 ( .A(n19935), .ZN(n19943) );
  INV_X1 U11733 ( .A(n14278), .ZN(n9790) );
  INV_X1 U11734 ( .A(n13836), .ZN(n19961) );
  AND2_X1 U11735 ( .A1(n12723), .A2(n12702), .ZN(n19979) );
  INV_X1 U11736 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20673) );
  OR2_X1 U11737 ( .A1(n10627), .A2(n10803), .ZN(n13233) );
  AND2_X1 U11738 ( .A1(n13632), .A2(n13222), .ZN(n18643) );
  AND2_X1 U11739 ( .A1(n9818), .A2(n9817), .ZN(n14770) );
  OAI21_X1 U11740 ( .B1(n9818), .B2(n9817), .A(n18827), .ZN(n9816) );
  NAND2_X1 U11741 ( .A1(n18974), .A2(n10805), .ZN(n18836) );
  AND2_X1 U11742 ( .A1(n18903), .A2(n13188), .ZN(n18899) );
  NOR2_X1 U11743 ( .A1(n14984), .A2(n18989), .ZN(n9868) );
  INV_X1 U11744 ( .A(n16108), .ZN(n18989) );
  NAND2_X1 U11745 ( .A1(n13230), .A2(n12488), .ZN(n16117) );
  XOR2_X1 U11746 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n14992), .Z(
        n14985) );
  NAND2_X1 U11747 ( .A1(n14990), .A2(n14988), .ZN(n14193) );
  XNOR2_X1 U11748 ( .A(n15233), .B(n10091), .ZN(n16043) );
  NAND2_X1 U11749 ( .A1(n15302), .A2(n9710), .ZN(n9737) );
  AND2_X1 U11750 ( .A1(n12790), .A2(n12789), .ZN(n18992) );
  OR2_X1 U11751 ( .A1(n12850), .A2(n12802), .ZN(n16146) );
  INV_X1 U11752 ( .A(n18996), .ZN(n16152) );
  INV_X1 U11753 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19710) );
  INV_X1 U11754 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19704) );
  AND2_X1 U11755 ( .A1(n19258), .A2(n19446), .ZN(n19249) );
  NOR2_X1 U11756 ( .A1(n17621), .A2(n18631), .ZN(n18617) );
  NOR2_X1 U11757 ( .A1(n17008), .A2(n17144), .ZN(n17003) );
  NOR2_X1 U11758 ( .A1(n17032), .A2(n17026), .ZN(n17023) );
  NOR2_X1 U11759 ( .A1(n17075), .A2(n17250), .ZN(n17070) );
  OR2_X1 U11760 ( .A1(n17261), .A2(n17260), .ZN(n17262) );
  AOI21_X1 U11761 ( .B1(n12524), .B2(n17258), .A(n17470), .ZN(n17263) );
  OAI21_X1 U11762 ( .B1(n17278), .B2(n9726), .A(n9750), .ZN(n9749) );
  AOI21_X1 U11763 ( .B1(n17475), .B2(n17276), .A(n17643), .ZN(n9750) );
  INV_X1 U11764 ( .A(n17277), .ZN(n9751) );
  NAND2_X1 U11765 ( .A1(n9755), .A2(n17627), .ZN(n9754) );
  NAND2_X1 U11766 ( .A1(n17328), .A2(n17268), .ZN(n9755) );
  INV_X1 U11767 ( .A(n17275), .ZN(n9753) );
  INV_X1 U11768 ( .A(n17475), .ZN(n17417) );
  NAND2_X1 U11769 ( .A1(n17614), .A2(n17103), .ZN(n17470) );
  NOR2_X1 U11770 ( .A1(n17269), .A2(n17273), .ZN(n17646) );
  INV_X1 U11771 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18631) );
  XNOR2_X1 U11772 ( .A(n11184), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11627) );
  NAND2_X1 U11773 ( .A1(n11621), .A2(n11620), .ZN(n11630) );
  AND2_X1 U11774 ( .A1(n13408), .A2(n11310), .ZN(n11343) );
  NAND2_X1 U11775 ( .A1(n11682), .A2(n11309), .ZN(n11311) );
  OR2_X1 U11776 ( .A1(n9621), .A2(n14224), .ZN(n10663) );
  OR2_X1 U11777 ( .A1(n10255), .A2(n10256), .ZN(n10248) );
  OR2_X1 U11778 ( .A1(n11529), .A2(n11528), .ZN(n11566) );
  INV_X1 U11779 ( .A(n11341), .ZN(n12584) );
  NAND2_X1 U11780 ( .A1(n12580), .A2(n11340), .ZN(n11320) );
  NAND2_X1 U11781 ( .A1(n9768), .A2(n11320), .ZN(n12709) );
  AOI22_X1 U11782 ( .A1(n11360), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9630), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U11783 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14139), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11229) );
  AND2_X2 U11784 ( .A1(n11186), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11194) );
  AND2_X1 U11785 ( .A1(n12324), .A2(n9959), .ZN(n9958) );
  INV_X1 U11786 ( .A(n9958), .ZN(n9956) );
  NOR2_X1 U11787 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10822) );
  INV_X1 U11788 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10814) );
  NOR2_X1 U11789 ( .A1(n10056), .A2(n10053), .ZN(n10052) );
  INV_X1 U11790 ( .A(n15048), .ZN(n10053) );
  INV_X1 U11791 ( .A(n15044), .ZN(n10056) );
  OR2_X1 U11792 ( .A1(n10943), .A2(n10942), .ZN(n12244) );
  NAND2_X1 U11793 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12173) );
  AOI22_X1 U11794 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12201), .B1(
        n12248), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12207) );
  AND2_X1 U11795 ( .A1(n12765), .A2(n10628), .ZN(n10600) );
  INV_X1 U11796 ( .A(n12768), .ZN(n12816) );
  CLKBUF_X1 U11797 ( .A(n10614), .Z(n12819) );
  NOR2_X1 U11798 ( .A1(n12875), .A2(n12178), .ZN(n12188) );
  AND2_X1 U11799 ( .A1(n10787), .A2(n10786), .ZN(n10793) );
  NAND2_X1 U11800 ( .A1(n9763), .A2(n9762), .ZN(n16705) );
  INV_X1 U11801 ( .A(n10105), .ZN(n9762) );
  INV_X1 U11802 ( .A(n16663), .ZN(n9763) );
  NOR2_X1 U11803 ( .A1(n10105), .A2(n10106), .ZN(n10137) );
  AOI21_X1 U11804 ( .B1(n18423), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10247), .ZN(n10256) );
  AND2_X1 U11805 ( .A1(n10354), .A2(n10355), .ZN(n10247) );
  NOR2_X1 U11806 ( .A1(n10107), .A2(n18429), .ZN(n10136) );
  XNOR2_X1 U11807 ( .A(n11336), .B(n11335), .ZN(n11352) );
  NOR2_X1 U11808 ( .A1(n14352), .A2(n10040), .ZN(n10039) );
  INV_X1 U11809 ( .A(n10041), .ZN(n10040) );
  NAND2_X1 U11810 ( .A1(n9785), .A2(n9784), .ZN(n12603) );
  AND2_X1 U11811 ( .A1(n10046), .A2(n12144), .ZN(n10045) );
  INV_X1 U11812 ( .A(n14305), .ZN(n12096) );
  AND2_X1 U11813 ( .A1(n13870), .A2(n11764), .ZN(n10038) );
  NOR2_X1 U11814 ( .A1(n14300), .A2(n9780), .ZN(n9779) );
  INV_X1 U11815 ( .A(n14611), .ZN(n9780) );
  NAND2_X1 U11816 ( .A1(n9980), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9979) );
  NAND2_X1 U11817 ( .A1(n14705), .A2(n11609), .ZN(n9980) );
  INV_X1 U11818 ( .A(n13768), .ZN(n9963) );
  INV_X1 U11819 ( .A(n11321), .ZN(n12593) );
  NAND2_X1 U11820 ( .A1(n10025), .A2(n10023), .ZN(n11455) );
  AOI21_X1 U11821 ( .B1(n10026), .B2(n10028), .A(n10024), .ZN(n10023) );
  INV_X1 U11822 ( .A(n11589), .ZN(n10024) );
  NAND2_X1 U11823 ( .A1(n11424), .A2(n11423), .ZN(n11426) );
  NAND2_X1 U11824 ( .A1(n20666), .A2(n20702), .ZN(n11486) );
  AOI221_X1 U11825 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11624), 
        .C1(n15947), .C2(n11624), .A(n11622), .ZN(n12573) );
  INV_X1 U11826 ( .A(n12297), .ZN(n10781) );
  NAND2_X1 U11827 ( .A1(n11165), .A2(n11164), .ZN(n12430) );
  INV_X1 U11828 ( .A(n12362), .ZN(n9952) );
  NOR2_X1 U11829 ( .A1(n12368), .A2(n11154), .ZN(n12346) );
  CLKBUF_X1 U11830 ( .A(n13149), .Z(n13137) );
  INV_X1 U11831 ( .A(n10071), .ZN(n10003) );
  OR2_X1 U11832 ( .A1(n14857), .A2(n14867), .ZN(n10005) );
  NAND2_X1 U11833 ( .A1(n10020), .A2(n16010), .ZN(n10019) );
  INV_X1 U11834 ( .A(n14880), .ZN(n10020) );
  NOR2_X1 U11835 ( .A1(n10019), .A2(n10018), .ZN(n10017) );
  INV_X1 U11836 ( .A(n14874), .ZN(n10018) );
  AND2_X1 U11837 ( .A1(n13099), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12876) );
  INV_X1 U11838 ( .A(n14194), .ZN(n9897) );
  NOR3_X1 U11839 ( .A1(n10443), .A2(n10442), .A3(n12489), .ZN(n10441) );
  NAND2_X1 U11840 ( .A1(n14811), .A2(n13213), .ZN(n9858) );
  NOR2_X1 U11841 ( .A1(n14775), .A2(n9865), .ZN(n9864) );
  INV_X1 U11842 ( .A(n14847), .ZN(n9865) );
  AOI21_X1 U11843 ( .B1(n12536), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9903), .ZN(n9902) );
  NOR2_X1 U11844 ( .A1(n12539), .A2(n20763), .ZN(n9900) );
  INV_X1 U11845 ( .A(n14892), .ZN(n9924) );
  NAND2_X1 U11846 ( .A1(n9651), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9845) );
  OR2_X1 U11847 ( .A1(n11118), .A2(n11117), .ZN(n14962) );
  NAND2_X1 U11848 ( .A1(n15271), .A2(n14962), .ZN(n15632) );
  NAND2_X1 U11849 ( .A1(n12477), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10066) );
  INV_X1 U11850 ( .A(n12465), .ZN(n12272) );
  OAI211_X1 U11851 ( .C1(n10675), .C2(n10678), .A(n10677), .B(n10676), .ZN(
        n10680) );
  NAND2_X1 U11852 ( .A1(n10674), .A2(n10673), .ZN(n10679) );
  NAND2_X1 U11853 ( .A1(n10625), .A2(n10624), .ZN(n10651) );
  NAND2_X1 U11854 ( .A1(n10623), .A2(n10622), .ZN(n10624) );
  OR2_X1 U11855 ( .A1(n10833), .A2(n10832), .ZN(n12449) );
  NOR2_X1 U11856 ( .A1(n12798), .A2(n12797), .ZN(n13650) );
  INV_X1 U11857 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U11858 ( .A1(n12853), .A2(n19700), .ZN(n12872) );
  AND2_X1 U11859 ( .A1(n13099), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12858) );
  AND2_X1 U11860 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12985) );
  AND2_X2 U11861 ( .A1(n13950), .A2(n12190), .ZN(n19084) );
  OR2_X1 U11862 ( .A1(n13319), .A2(n13229), .ZN(n13459) );
  NAND2_X1 U11863 ( .A1(n12484), .A2(n12483), .ZN(n12764) );
  NAND2_X1 U11864 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18592), .ZN(
        n10106) );
  NOR2_X1 U11865 ( .A1(n10104), .A2(n10106), .ZN(n10135) );
  INV_X1 U11866 ( .A(n10137), .ZN(n16804) );
  INV_X1 U11867 ( .A(n16622), .ZN(n16939) );
  NAND2_X1 U11868 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18584), .ZN(
        n10104) );
  NAND2_X1 U11869 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18598), .ZN(
        n10102) );
  NAND2_X1 U11870 ( .A1(n10360), .A2(n17975), .ZN(n10347) );
  NAND2_X1 U11871 ( .A1(n17253), .A2(n9725), .ZN(n9728) );
  NOR2_X1 U11872 ( .A1(n17617), .A2(n9726), .ZN(n9725) );
  AND2_X1 U11873 ( .A1(n17524), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17487) );
  NAND2_X1 U11874 ( .A1(n9994), .A2(n9993), .ZN(n10228) );
  AND2_X1 U11875 ( .A1(n12521), .A2(n17627), .ZN(n9993) );
  INV_X1 U11876 ( .A(n10227), .ZN(n9994) );
  OAI21_X1 U11877 ( .B1(n17979), .B2(n10343), .A(n12506), .ZN(n10350) );
  NOR2_X1 U11878 ( .A1(n10210), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9992) );
  NOR2_X1 U11879 ( .A1(n17539), .A2(n17542), .ZN(n10395) );
  NOR2_X1 U11880 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18598), .ZN(
        n10355) );
  XNOR2_X1 U11881 ( .A(n17124), .B(n10371), .ZN(n10194) );
  NOR2_X1 U11882 ( .A1(n10348), .A2(n10350), .ZN(n14127) );
  AND2_X1 U11883 ( .A1(n14246), .A2(n14245), .ZN(n14253) );
  INV_X1 U11884 ( .A(n13413), .ZN(n11690) );
  NAND2_X1 U11885 ( .A1(n11352), .A2(n11353), .ZN(n11429) );
  OR3_X1 U11886 ( .A1(n20706), .A2(n19977), .A3(n13787), .ZN(n15659) );
  NAND2_X1 U11887 ( .A1(n12695), .A2(n9769), .ZN(n14297) );
  AND2_X1 U11888 ( .A1(n13398), .A2(n13397), .ZN(n19855) );
  OR2_X1 U11889 ( .A1(n12122), .A2(n12121), .ZN(n14287) );
  OR2_X1 U11890 ( .A1(n12076), .A2(n12075), .ZN(n14494) );
  INV_X1 U11891 ( .A(n14303), .ZN(n14496) );
  AND2_X1 U11892 ( .A1(n15666), .A2(n14157), .ZN(n12047) );
  AND2_X1 U11893 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12027), .ZN(
        n12028) );
  NAND2_X1 U11894 ( .A1(n12028), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12070) );
  NAND2_X1 U11895 ( .A1(n11968), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12026) );
  AND2_X1 U11896 ( .A1(n11966), .A2(n11965), .ZN(n14365) );
  NOR2_X1 U11897 ( .A1(n11934), .A2(n11933), .ZN(n11935) );
  NOR2_X1 U11898 ( .A1(n11911), .A2(n14543), .ZN(n11912) );
  NAND2_X1 U11899 ( .A1(n9967), .A2(n9965), .ZN(n9972) );
  CLKBUF_X1 U11900 ( .A(n14312), .Z(n14313) );
  NOR2_X1 U11901 ( .A1(n10031), .A2(n10033), .ZN(n10030) );
  INV_X1 U11902 ( .A(n14121), .ZN(n10031) );
  NOR2_X1 U11903 ( .A1(n11865), .A2(n11864), .ZN(n11866) );
  AND2_X1 U11904 ( .A1(n11829), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11847) );
  AND2_X1 U11905 ( .A1(n11782), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11783) );
  AND2_X1 U11906 ( .A1(n11856), .A2(n11796), .ZN(n14078) );
  CLKBUF_X1 U11907 ( .A(n13982), .Z(n13983) );
  OR2_X1 U11908 ( .A1(n11748), .A2(n13879), .ZN(n11765) );
  AOI21_X1 U11909 ( .B1(n11724), .B2(n11856), .A(n11723), .ZN(n13844) );
  NOR2_X1 U11910 ( .A1(n11711), .A2(n19812), .ZN(n11720) );
  INV_X1 U11911 ( .A(n13752), .ZN(n11717) );
  AND2_X1 U11912 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11693), .ZN(
        n11712) );
  NAND2_X1 U11913 ( .A1(n13503), .A2(n11692), .ZN(n13587) );
  CLKBUF_X1 U11914 ( .A(n13584), .Z(n13585) );
  OAI21_X1 U11915 ( .B1(n12601), .B2(P1_EBX_REG_29__SCAN_IN), .A(n9766), .ZN(
        n14274) );
  NAND2_X1 U11916 ( .A1(n12566), .A2(n12565), .ZN(n14458) );
  INV_X1 U11917 ( .A(n14219), .ZN(n9781) );
  NAND2_X1 U11918 ( .A1(n14612), .A2(n9779), .ZN(n14302) );
  NAND2_X1 U11919 ( .A1(n14469), .A2(n11615), .ZN(n14481) );
  NAND2_X1 U11920 ( .A1(n14612), .A2(n14611), .ZN(n14614) );
  OR2_X1 U11921 ( .A1(n14470), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14502) );
  AND2_X1 U11922 ( .A1(n12679), .A2(n12678), .ZN(n14353) );
  INV_X1 U11923 ( .A(n9978), .ZN(n11614) );
  AOI21_X1 U11924 ( .B1(n14521), .B2(n14705), .A(n9979), .ZN(n9978) );
  AND2_X1 U11925 ( .A1(n14656), .A2(n14366), .ZN(n14368) );
  AND2_X1 U11926 ( .A1(n12670), .A2(n12669), .ZN(n14653) );
  AND2_X1 U11927 ( .A1(n12667), .A2(n12666), .ZN(n14316) );
  INV_X1 U11928 ( .A(n11608), .ZN(n14526) );
  AND2_X1 U11929 ( .A1(n12653), .A2(n12652), .ZN(n14089) );
  OR2_X1 U11930 ( .A1(n14728), .A2(n14727), .ZN(n14725) );
  AND2_X1 U11931 ( .A1(n13987), .A2(n12642), .ZN(n15781) );
  AND2_X1 U11932 ( .A1(n12639), .A2(n12638), .ZN(n13916) );
  OR2_X1 U11933 ( .A1(n15936), .A2(n12634), .ZN(n13917) );
  INV_X1 U11934 ( .A(n19986), .ZN(n15922) );
  NAND2_X1 U11935 ( .A1(n15934), .A2(n15933), .ZN(n15936) );
  NAND2_X1 U11936 ( .A1(n12615), .A2(n9787), .ZN(n12616) );
  NAND2_X1 U11937 ( .A1(n11465), .A2(n11464), .ZN(n13509) );
  OR2_X1 U11938 ( .A1(n20001), .A2(n19991), .ZN(n14661) );
  NAND2_X1 U11939 ( .A1(n11327), .A2(n11310), .ZN(n14742) );
  AND2_X1 U11940 ( .A1(n12583), .A2(n12703), .ZN(n13506) );
  AND2_X1 U11941 ( .A1(n11701), .A2(n9617), .ZN(n20118) );
  OR2_X1 U11942 ( .A1(n9617), .A2(n11488), .ZN(n20214) );
  NAND2_X1 U11943 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20164), .ZN(n20024) );
  OR2_X1 U11944 ( .A1(n20010), .A2(n20259), .ZN(n20404) );
  NOR2_X2 U11945 ( .A1(n20006), .A2(n20005), .ZN(n20048) );
  AND2_X1 U11946 ( .A1(n20010), .A2(n20259), .ZN(n20383) );
  OR2_X1 U11947 ( .A1(n9617), .A2(n20158), .ZN(n20443) );
  AOI21_X1 U11948 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20446), .A(n20059), 
        .ZN(n20527) );
  INV_X1 U11949 ( .A(n20024), .ZN(n20049) );
  AND2_X1 U11950 ( .A1(n14789), .A2(n14909), .ZN(n14911) );
  AND2_X1 U11951 ( .A1(n12406), .A2(n12401), .ZN(n13211) );
  NAND2_X1 U11952 ( .A1(n9636), .A2(n9814), .ZN(n9815) );
  NAND2_X1 U11953 ( .A1(n12367), .A2(n11156), .ZN(n9942) );
  NAND2_X1 U11954 ( .A1(n12314), .A2(n12324), .ZN(n12326) );
  INV_X1 U11955 ( .A(n11149), .ZN(n9943) );
  AND2_X1 U11956 ( .A1(n9641), .A2(n10022), .ZN(n10021) );
  OR2_X1 U11957 ( .A1(n13631), .A2(n13634), .ZN(n13455) );
  NOR2_X1 U11958 ( .A1(n14851), .A2(n10009), .ZN(n10008) );
  OR2_X1 U11959 ( .A1(n10082), .A2(n10013), .ZN(n10009) );
  NOR4_X1 U11960 ( .A1(n12983), .A2(n12982), .A3(n12981), .A4(n12980), .ZN(
        n14945) );
  NAND2_X1 U11961 ( .A1(n10014), .A2(n10017), .ZN(n14873) );
  OR2_X1 U11962 ( .A1(n12910), .A2(n12909), .ZN(n13993) );
  NOR2_X1 U11963 ( .A1(n15391), .A2(n15390), .ZN(n13537) );
  NAND2_X1 U11964 ( .A1(n15431), .A2(n10960), .ZN(n13360) );
  OR2_X1 U11965 ( .A1(n10962), .A2(n10961), .ZN(n13359) );
  NAND2_X1 U11966 ( .A1(n12881), .A2(n12876), .ZN(n13781) );
  OAI21_X1 U11967 ( .B1(n13174), .B2(n13173), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13272) );
  CLKBUF_X1 U11968 ( .A(n10837), .Z(n13334) );
  NOR2_X1 U11969 ( .A1(n18921), .A2(n19071), .ZN(n13335) );
  INV_X1 U11970 ( .A(n13272), .ZN(n19027) );
  OR3_X1 U11971 ( .A1(n10442), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A3(
        n9806), .ZN(n9805) );
  OAI21_X1 U11972 ( .B1(n10443), .B2(n9804), .A(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9803) );
  OR2_X1 U11973 ( .A1(n10442), .A2(n9806), .ZN(n9804) );
  NAND2_X1 U11974 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U11975 ( .A1(n9857), .A2(n14858), .ZN(n14861) );
  AND2_X1 U11976 ( .A1(n10736), .A2(n10735), .ZN(n15061) );
  OR2_X1 U11977 ( .A1(n9825), .A2(n18703), .ZN(n9824) );
  AND2_X1 U11978 ( .A1(n15320), .A2(n15338), .ZN(n15067) );
  NAND2_X1 U11979 ( .A1(n10452), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10463) );
  OR2_X1 U11980 ( .A1(n9870), .A2(n13820), .ZN(n9869) );
  OR2_X1 U11981 ( .A1(n13902), .A2(n9870), .ZN(n13819) );
  NAND2_X1 U11982 ( .A1(n10453), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10462) );
  AND2_X1 U11983 ( .A1(n10603), .A2(n10602), .ZN(n13903) );
  NOR2_X1 U11984 ( .A1(n13902), .A2(n13903), .ZN(n13904) );
  NAND2_X1 U11985 ( .A1(n10454), .A2(n9692), .ZN(n10459) );
  NAND2_X1 U11986 ( .A1(n10454), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10458) );
  NAND2_X1 U11987 ( .A1(n10455), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10457) );
  NAND2_X1 U11988 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10456) );
  INV_X1 U11989 ( .A(n12167), .ZN(n12171) );
  NOR2_X1 U11990 ( .A1(n20763), .A2(n14201), .ZN(n10069) );
  NOR2_X1 U11991 ( .A1(n15128), .A2(n12539), .ZN(n10070) );
  AND2_X1 U11992 ( .A1(n14848), .A2(n9862), .ZN(n14762) );
  NOR2_X1 U11993 ( .A1(n9863), .A2(n12481), .ZN(n9862) );
  INV_X1 U11994 ( .A(n9864), .ZN(n9863) );
  NAND2_X1 U11995 ( .A1(n14789), .A2(n9925), .ZN(n14893) );
  NOR2_X1 U11996 ( .A1(n14861), .A2(n14787), .ZN(n14848) );
  OAI21_X1 U11997 ( .B1(n15007), .B2(n12417), .A(n9941), .ZN(n9940) );
  INV_X1 U11998 ( .A(n12416), .ZN(n9941) );
  XNOR2_X1 U11999 ( .A(n12420), .B(n15166), .ZN(n15011) );
  OAI21_X1 U12000 ( .B1(n14793), .B2(n12280), .A(n15187), .ZN(n15177) );
  AND2_X1 U12001 ( .A1(n13214), .A2(n14932), .ZN(n14930) );
  AND2_X1 U12002 ( .A1(n15271), .A2(n9713), .ZN(n13216) );
  INV_X1 U12003 ( .A(n14808), .ZN(n9931) );
  NAND2_X1 U12004 ( .A1(n12478), .A2(n9651), .ZN(n15038) );
  NOR3_X1 U12005 ( .A1(n15060), .A2(n9860), .A3(n10741), .ZN(n14809) );
  AND2_X1 U12006 ( .A1(n12355), .A2(n15227), .ZN(n15231) );
  INV_X1 U12007 ( .A(n15082), .ZN(n10064) );
  AND3_X1 U12008 ( .A1(n10811), .A2(n10810), .A3(n10809), .ZN(n15272) );
  INV_X1 U12009 ( .A(n16119), .ZN(n9935) );
  INV_X1 U12010 ( .A(n14971), .ZN(n9936) );
  OR2_X1 U12011 ( .A1(n16119), .A2(n9938), .ZN(n15305) );
  INV_X1 U12012 ( .A(n9793), .ZN(n15337) );
  NAND2_X1 U12013 ( .A1(n13731), .A2(n13730), .ZN(n16119) );
  NOR2_X1 U12014 ( .A1(n13535), .A2(n13677), .ZN(n13731) );
  INV_X1 U12015 ( .A(n15396), .ZN(n9847) );
  NOR2_X1 U12016 ( .A1(n10061), .A2(n10060), .ZN(n10059) );
  INV_X1 U12017 ( .A(n15387), .ZN(n10060) );
  NAND2_X1 U12018 ( .A1(n13362), .A2(n9929), .ZN(n15391) );
  NOR2_X1 U12019 ( .A1(n13387), .A2(n9930), .ZN(n9929) );
  NAND2_X1 U12020 ( .A1(n13361), .A2(n13416), .ZN(n9930) );
  NOR2_X1 U12021 ( .A1(n9852), .A2(n9851), .ZN(n13547) );
  INV_X1 U12022 ( .A(n13597), .ZN(n9850) );
  OR2_X1 U12023 ( .A1(n15452), .A2(n13363), .ZN(n14178) );
  INV_X1 U12024 ( .A(n14178), .ZN(n15410) );
  NAND2_X1 U12025 ( .A1(n12461), .A2(n12460), .ZN(n15438) );
  NOR2_X1 U12026 ( .A1(n13732), .A2(n13775), .ZN(n15433) );
  NAND2_X1 U12027 ( .A1(n9876), .A2(n9875), .ZN(n13935) );
  AOI21_X1 U12028 ( .B1(n9879), .B2(n9883), .A(n9697), .ZN(n9875) );
  INV_X1 U12029 ( .A(n9886), .ZN(n9883) );
  OAI21_X1 U12030 ( .B1(n13894), .B2(n13893), .A(n12458), .ZN(n13933) );
  NOR2_X1 U12031 ( .A1(n16155), .A2(n16154), .ZN(n15435) );
  OAI22_X1 U12032 ( .A1(n10672), .A2(n10639), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10661), .ZN(n10641) );
  INV_X1 U12033 ( .A(n13437), .ZN(n12792) );
  NOR2_X1 U12034 ( .A1(n12850), .A2(n13441), .ZN(n19000) );
  XNOR2_X1 U12035 ( .A(n13339), .B(n10850), .ZN(n13431) );
  NAND2_X1 U12036 ( .A1(n9922), .A2(n9920), .ZN(n13604) );
  INV_X1 U12037 ( .A(n10890), .ZN(n9920) );
  XNOR2_X1 U12038 ( .A(n13345), .B(n12866), .ZN(n13374) );
  NOR2_X1 U12039 ( .A1(n10610), .A2(n10574), .ZN(n10576) );
  AND2_X1 U12040 ( .A1(n12985), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13446) );
  INV_X1 U12041 ( .A(n19382), .ZN(n19379) );
  INV_X1 U12042 ( .A(n12785), .ZN(n19055) );
  NAND2_X1 U12043 ( .A1(n19554), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19072) );
  OR2_X1 U12044 ( .A1(n19320), .A2(n19724), .ZN(n19452) );
  INV_X1 U12045 ( .A(n19452), .ZN(n19376) );
  NOR2_X2 U12046 ( .A1(n19027), .A2(n19026), .ZN(n19076) );
  NOR2_X2 U12047 ( .A1(n19025), .A2(n19026), .ZN(n19077) );
  OR2_X1 U12048 ( .A1(n12751), .A2(n12440), .ZN(n10800) );
  INV_X1 U12049 ( .A(n16311), .ZN(n18403) );
  NOR2_X1 U12050 ( .A1(n16342), .A2(n16343), .ZN(n16341) );
  NAND2_X1 U12051 ( .A1(n9732), .A2(n9731), .ZN(n16351) );
  OR2_X1 U12052 ( .A1(n9733), .A2(n9734), .ZN(n9731) );
  OR2_X1 U12053 ( .A1(n16370), .A2(n9733), .ZN(n9732) );
  NOR2_X1 U12055 ( .A1(n16421), .A2(n9733), .ZN(n16413) );
  NOR2_X1 U12056 ( .A1(n16413), .A2(n17334), .ZN(n16412) );
  NOR2_X1 U12057 ( .A1(n16431), .A2(n17371), .ZN(n16430) );
  NAND2_X1 U12058 ( .A1(n10414), .A2(n10093), .ZN(n16454) );
  INV_X1 U12059 ( .A(n10188), .ZN(n16622) );
  NAND2_X1 U12060 ( .A1(n17138), .A2(n18634), .ZN(n10429) );
  NOR2_X1 U12061 ( .A1(n17148), .A2(n20815), .ZN(n9910) );
  NAND2_X1 U12062 ( .A1(n9915), .A2(n9914), .ZN(n16987) );
  NAND2_X1 U12063 ( .A1(n15627), .A2(n15626), .ZN(n9914) );
  INV_X1 U12064 ( .A(n10334), .ZN(n18418) );
  AOI21_X1 U12065 ( .B1(n9756), .B2(n18453), .A(n18478), .ZN(n17137) );
  INV_X1 U12066 ( .A(n17196), .ZN(n17139) );
  INV_X1 U12067 ( .A(n17200), .ZN(n17198) );
  NOR2_X1 U12068 ( .A1(n10423), .A2(n16182), .ZN(n10422) );
  NAND2_X1 U12069 ( .A1(n17253), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17254) );
  NOR2_X1 U12070 ( .A1(n17332), .A2(n10408), .ZN(n17295) );
  NAND2_X1 U12071 ( .A1(n10407), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17332) );
  NOR2_X1 U12072 ( .A1(n17366), .A2(n17330), .ZN(n10417) );
  NAND2_X1 U12073 ( .A1(n10363), .A2(n10077), .ZN(n17413) );
  NOR2_X1 U12074 ( .A1(n17477), .A2(n17463), .ZN(n17437) );
  NAND2_X1 U12075 ( .A1(n16532), .A2(n17454), .ZN(n17458) );
  AND3_X1 U12076 ( .A1(n17487), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17454) );
  INV_X1 U12077 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16634) );
  NOR2_X1 U12078 ( .A1(n17608), .A2(n16634), .ZN(n17582) );
  NAND2_X1 U12079 ( .A1(n17581), .A2(n17622), .ZN(n17551) );
  OAI21_X1 U12080 ( .B1(n10228), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17428), .ZN(n10230) );
  OAI21_X1 U12081 ( .B1(n17257), .B2(n12501), .A(n12500), .ZN(n12502) );
  NOR2_X1 U12082 ( .A1(n17302), .A2(n12504), .ZN(n17628) );
  AOI21_X1 U12083 ( .B1(n17443), .B2(n10212), .A(n17531), .ZN(n17408) );
  NOR2_X1 U12084 ( .A1(n17471), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17443) );
  INV_X1 U12085 ( .A(n17818), .ZN(n17495) );
  NOR2_X1 U12086 ( .A1(n10345), .A2(n10344), .ZN(n15457) );
  AOI21_X1 U12087 ( .B1(n17988), .B2(n18411), .A(n14126), .ZN(n14128) );
  INV_X1 U12088 ( .A(n17493), .ZN(n17820) );
  NAND2_X1 U12089 ( .A1(n9991), .A2(n9992), .ZN(n10213) );
  NOR2_X1 U12090 ( .A1(n17541), .A2(n17540), .ZN(n17539) );
  OAI21_X1 U12091 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n10198), .A(
        n17590), .ZN(n17579) );
  NAND2_X1 U12092 ( .A1(n18419), .A2(n18427), .ZN(n17922) );
  INV_X1 U12093 ( .A(n14128), .ZN(n18430) );
  NAND2_X1 U12094 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18432) );
  INV_X1 U12095 ( .A(n10240), .ZN(n16819) );
  NOR2_X2 U12096 ( .A1(n18633), .A2(n15460), .ZN(n18438) );
  AND2_X1 U12097 ( .A1(n14127), .A2(n14128), .ZN(n18433) );
  NOR2_X1 U12098 ( .A1(n10268), .A2(n10267), .ZN(n17968) );
  NOR2_X2 U12099 ( .A1(n10246), .A2(n10245), .ZN(n17971) );
  INV_X1 U12100 ( .A(n10344), .ZN(n17979) );
  NOR2_X1 U12101 ( .A1(n10309), .A2(n10308), .ZN(n17983) );
  INV_X1 U12102 ( .A(n17991), .ZN(n18344) );
  NAND2_X1 U12103 ( .A1(n18622), .A2(n17966), .ZN(n18043) );
  OAI22_X1 U12104 ( .A1(n15458), .A2(n17801), .B1(n12510), .B2(n18405), .ZN(
        n18451) );
  CLKBUF_X1 U12105 ( .A(n13272), .Z(n19025) );
  NAND2_X1 U12106 ( .A1(n13695), .A2(n13298), .ZN(n20706) );
  INV_X1 U12107 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19812) );
  INV_X1 U12108 ( .A(n15770), .ZN(n19832) );
  AND2_X1 U12109 ( .A1(n13800), .A2(n13798), .ZN(n19833) );
  INV_X1 U12110 ( .A(n19837), .ZN(n19818) );
  AND2_X1 U12111 ( .A1(n15659), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19838) );
  INV_X1 U12112 ( .A(n14383), .ZN(n19849) );
  INV_X1 U12113 ( .A(n14442), .ZN(n15803) );
  INV_X1 U12114 ( .A(n15809), .ZN(n14444) );
  NAND2_X1 U12115 ( .A1(n13424), .A2(n14260), .ZN(n15801) );
  OR2_X1 U12116 ( .A1(n13487), .A2(n13423), .ZN(n13424) );
  NAND2_X1 U12117 ( .A1(n14442), .A2(n14123), .ZN(n14086) );
  INV_X1 U12118 ( .A(n14086), .ZN(n14118) );
  BUF_X1 U12119 ( .A(n19884), .Z(n20709) );
  BUF_X1 U12120 ( .A(n19883), .Z(n19875) );
  NOR2_X1 U12121 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13578), .ZN(n19884) );
  XNOR2_X1 U12122 ( .A(n13791), .B(n13790), .ZN(n14450) );
  OAI21_X1 U12123 ( .B1(n14521), .B2(n11609), .A(n14705), .ZN(n15810) );
  CLKBUF_X1 U12124 ( .A(n14053), .Z(n14054) );
  CLKBUF_X1 U12125 ( .A(n14051), .Z(n14052) );
  AND2_X1 U12126 ( .A1(n14069), .A2(n14085), .ZN(n15847) );
  XNOR2_X1 U12127 ( .A(n9776), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14454) );
  OAI21_X1 U12128 ( .B1(n14455), .B2(n9775), .A(n9675), .ZN(n9776) );
  OAI21_X1 U12129 ( .B1(n14685), .B2(n19970), .A(n14658), .ZN(n14713) );
  NAND2_X1 U12130 ( .A1(n9969), .A2(n11595), .ZN(n14034) );
  NAND2_X1 U12131 ( .A1(n13833), .A2(n11549), .ZN(n15865) );
  OR2_X1 U12132 ( .A1(n20001), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19985) );
  OR2_X1 U12133 ( .A1(n14661), .A2(n19968), .ZN(n19986) );
  INV_X1 U12134 ( .A(n19979), .ZN(n19995) );
  NAND2_X1 U12135 ( .A1(n12723), .A2(n12719), .ZN(n19992) );
  NAND2_X1 U12136 ( .A1(n11684), .A2(n9667), .ZN(n9772) );
  INV_X1 U12137 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20690) );
  INV_X1 U12138 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20681) );
  INV_X1 U12139 ( .A(n9617), .ZN(n20674) );
  CLKBUF_X1 U12140 ( .A(n13554), .Z(n20678) );
  NOR2_X1 U12141 ( .A1(n20214), .A2(n20525), .ZN(n20664) );
  NOR2_X1 U12142 ( .A1(n11701), .A2(n20674), .ZN(n20665) );
  NOR2_X1 U12143 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15945) );
  OAI211_X1 U12144 ( .C1(n20050), .C2(n20780), .A(n20350), .B(n20017), .ZN(
        n20053) );
  INV_X1 U12145 ( .A(n20084), .ZN(n20075) );
  NOR2_X1 U12146 ( .A1(n20446), .A2(n20261), .ZN(n20283) );
  OAI22_X1 U12147 ( .A1(n20354), .A2(n20353), .B1(n20352), .B2(n20472), .ZN(
        n20371) );
  OAI211_X1 U12148 ( .C1(n20509), .C2(n20479), .A(n20478), .B(n20477), .ZN(
        n20513) );
  INV_X1 U12149 ( .A(n20215), .ZN(n20523) );
  AND2_X1 U12150 ( .A1(n20029), .A2(n20049), .ZN(n20540) );
  AND2_X1 U12151 ( .A1(n11340), .A2(n20049), .ZN(n20546) );
  AND2_X1 U12152 ( .A1(n20040), .A2(n20049), .ZN(n20558) );
  AND2_X1 U12153 ( .A1(n20044), .A2(n20049), .ZN(n20564) );
  AND2_X1 U12154 ( .A1(n11310), .A2(n20049), .ZN(n20571) );
  OR2_X1 U12155 ( .A1(n20582), .A2(n20702), .ZN(n19763) );
  AND2_X1 U12156 ( .A1(n15598), .A2(n15597), .ZN(n15610) );
  NAND2_X1 U12157 ( .A1(n13792), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20582) );
  INV_X1 U12158 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20780) );
  INV_X1 U12159 ( .A(n16159), .ZN(n19732) );
  INV_X1 U12160 ( .A(n14199), .ZN(n14983) );
  INV_X1 U12161 ( .A(n9819), .ZN(n15968) );
  NAND2_X1 U12162 ( .A1(n9807), .A2(n9809), .ZN(n15982) );
  AND2_X1 U12163 ( .A1(n12410), .A2(n12547), .ZN(n15977) );
  NOR2_X1 U12164 ( .A1(n14798), .A2(n16031), .ZN(n14797) );
  NAND2_X1 U12165 ( .A1(n9812), .A2(n9811), .ZN(n13209) );
  NAND2_X1 U12166 ( .A1(n10466), .A2(n9813), .ZN(n9811) );
  INV_X1 U12167 ( .A(n15042), .ZN(n9813) );
  AND2_X1 U12168 ( .A1(n9815), .A2(n13945), .ZN(n13210) );
  NOR2_X1 U12169 ( .A1(n12308), .A2(n12307), .ZN(n12282) );
  NAND2_X1 U12170 ( .A1(n18643), .A2(n11169), .ZN(n18852) );
  INV_X1 U12171 ( .A(n18870), .ZN(n18840) );
  NOR2_X1 U12172 ( .A1(n13945), .A2(n18877), .ZN(n18857) );
  INV_X1 U12173 ( .A(n18836), .ZN(n18863) );
  OR2_X1 U12174 ( .A1(n11061), .A2(n11060), .ZN(n18883) );
  OR2_X1 U12175 ( .A1(n11047), .A2(n11046), .ZN(n18884) );
  OR2_X1 U12176 ( .A1(n11029), .A2(n11028), .ZN(n18890) );
  OR2_X1 U12177 ( .A1(n11015), .A2(n11014), .ZN(n18891) );
  INV_X1 U12178 ( .A(n10000), .ZN(n9999) );
  NAND2_X1 U12179 ( .A1(n9998), .A2(n10000), .ZN(n9997) );
  INV_X1 U12180 ( .A(n18899), .ZN(n18893) );
  NAND2_X1 U12181 ( .A1(n13020), .A2(n10071), .ZN(n10006) );
  INV_X1 U12182 ( .A(n10007), .ZN(n14866) );
  NAND2_X1 U12183 ( .A1(n18926), .A2(n9736), .ZN(n16017) );
  INV_X1 U12184 ( .A(n14918), .ZN(n18909) );
  AND2_X1 U12185 ( .A1(n13180), .A2(n19025), .ZN(n18908) );
  NAND2_X1 U12186 ( .A1(n13362), .A2(n13361), .ZN(n13386) );
  AND2_X1 U12187 ( .A1(n13164), .A2(n13460), .ZN(n18926) );
  OR2_X1 U12188 ( .A1(n13456), .A2(n13163), .ZN(n13164) );
  INV_X1 U12189 ( .A(n18912), .ZN(n16018) );
  INV_X1 U12190 ( .A(n16024), .ZN(n18930) );
  NOR2_X1 U12191 ( .A1(n13345), .A2(n13344), .ZN(n19287) );
  INV_X1 U12192 ( .A(n18926), .ZN(n18921) );
  AND2_X1 U12193 ( .A1(n18926), .A2(n19071), .ZN(n18912) );
  OAI21_X1 U12194 ( .B1(n13319), .B2(n13318), .A(n13317), .ZN(n13320) );
  INV_X1 U12195 ( .A(n16001), .ZN(n12833) );
  NAND2_X1 U12196 ( .A1(n9797), .A2(n9795), .ZN(n15076) );
  INV_X1 U12197 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20750) );
  AND2_X1 U12198 ( .A1(n15281), .A2(n15280), .ZN(n18695) );
  INV_X1 U12199 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16095) );
  INV_X1 U12200 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15113) );
  INV_X1 U12201 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20762) );
  BUF_X2 U12202 ( .A(n12875), .Z(n13950) );
  INV_X1 U12203 ( .A(n16113), .ZN(n18980) );
  INV_X1 U12204 ( .A(n16117), .ZN(n18977) );
  NOR2_X1 U12205 ( .A1(n9856), .A2(n12848), .ZN(n9855) );
  NOR2_X1 U12206 ( .A1(n12847), .A2(n12846), .ZN(n12848) );
  INV_X1 U12207 ( .A(n12832), .ZN(n9856) );
  NAND2_X1 U12208 ( .A1(n9606), .A2(n9721), .ZN(n12553) );
  NAND2_X1 U12209 ( .A1(n9612), .A2(n15048), .ZN(n10057) );
  AND2_X1 U12210 ( .A1(n10063), .A2(n10058), .ZN(n15385) );
  INV_X1 U12211 ( .A(n14175), .ZN(n9836) );
  NAND2_X1 U12212 ( .A1(n9878), .A2(n9886), .ZN(n13889) );
  OR2_X1 U12213 ( .A1(n12850), .A2(n12849), .ZN(n18996) );
  OR2_X1 U12214 ( .A1(n19000), .A2(n19002), .ZN(n15452) );
  INV_X1 U12215 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19729) );
  INV_X1 U12216 ( .A(n19287), .ZN(n19724) );
  OR2_X1 U12217 ( .A1(n19549), .A2(n14021), .ZN(n19721) );
  INV_X1 U12218 ( .A(n19715), .ZN(n19712) );
  AND2_X1 U12219 ( .A1(n9921), .A2(n9922), .ZN(n13733) );
  INV_X1 U12220 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15625) );
  XNOR2_X1 U12221 ( .A(n13375), .B(n13374), .ZN(n19715) );
  INV_X1 U12222 ( .A(n13392), .ZN(n13393) );
  INV_X1 U12223 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19044) );
  INV_X1 U12224 ( .A(n19236), .ZN(n19254) );
  NOR2_X2 U12225 ( .A1(n19503), .A2(n19232), .ZN(n19283) );
  OAI21_X1 U12226 ( .B1(n19265), .B2(n19691), .A(n19264), .ZN(n19284) );
  OAI21_X1 U12227 ( .B1(n19310), .B2(n19291), .A(n19554), .ZN(n19312) );
  NOR2_X1 U12228 ( .A1(n19452), .A2(n19327), .ZN(n19350) );
  OAI21_X1 U12229 ( .B1(n19383), .B2(n19348), .A(n19347), .ZN(n19370) );
  NOR2_X2 U12230 ( .A1(n19504), .A2(n19384), .ZN(n19404) );
  OR2_X1 U12231 ( .A1(n19447), .A2(n19442), .ZN(n19495) );
  INV_X1 U12232 ( .A(n19563), .ZN(n19510) );
  INV_X1 U12233 ( .A(n19569), .ZN(n19518) );
  INV_X1 U12234 ( .A(n19575), .ZN(n19522) );
  INV_X1 U12235 ( .A(n19581), .ZN(n19526) );
  INV_X1 U12236 ( .A(n19587), .ZN(n19530) );
  INV_X1 U12237 ( .A(n19593), .ZN(n19534) );
  OAI21_X1 U12238 ( .B1(n19514), .B2(n19513), .A(n19512), .ZN(n19544) );
  INV_X1 U12239 ( .A(n19610), .ZN(n19543) );
  NOR2_X2 U12240 ( .A1(n19452), .A2(n19451), .ZN(n19542) );
  NOR2_X2 U12241 ( .A1(n19504), .A2(n19503), .ZN(n19605) );
  AND2_X1 U12242 ( .A1(n19555), .A2(n19551), .ZN(n19603) );
  INV_X1 U12243 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19751) );
  AND3_X1 U12244 ( .A1(n19622), .A2(n19675), .A3(n19628), .ZN(n19752) );
  INV_X1 U12245 ( .A(n9758), .ZN(n16313) );
  NAND2_X1 U12246 ( .A1(n18617), .A2(n18451), .ZN(n16314) );
  INV_X1 U12247 ( .A(n9735), .ZN(n16360) );
  AND2_X1 U12248 ( .A1(n9735), .A2(n9734), .ZN(n16359) );
  OR2_X1 U12249 ( .A1(n16370), .A2(n9733), .ZN(n9735) );
  NOR2_X1 U12250 ( .A1(n16391), .A2(n9733), .ZN(n16381) );
  NOR2_X1 U12251 ( .A1(n16392), .A2(n17310), .ZN(n16391) );
  NOR2_X1 U12252 ( .A1(n16412), .A2(n9733), .ZN(n16404) );
  NOR2_X1 U12253 ( .A1(n16404), .A2(n17321), .ZN(n16403) );
  NOR2_X1 U12254 ( .A1(n16422), .A2(n17353), .ZN(n16421) );
  NOR2_X1 U12255 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16494), .ZN(n16477) );
  NOR2_X1 U12256 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16564), .ZN(n16542) );
  NOR2_X1 U12257 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16588), .ZN(n16569) );
  NOR2_X1 U12258 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16612), .ZN(n16597) );
  INV_X1 U12259 ( .A(n9591), .ZN(n16659) );
  INV_X1 U12260 ( .A(n16674), .ZN(n16662) );
  INV_X1 U12261 ( .A(n16631), .ZN(n16673) );
  NOR2_X2 U12262 ( .A1(n18634), .A2(n10424), .ZN(n16676) );
  NOR2_X1 U12263 ( .A1(n16518), .A2(n16884), .ZN(n16869) );
  NAND2_X1 U12264 ( .A1(n16985), .A2(n15549), .ZN(n16884) );
  INV_X1 U12265 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16976) );
  INV_X1 U12266 ( .A(n16998), .ZN(n16994) );
  NAND2_X1 U12267 ( .A1(n17017), .A2(n9652), .ZN(n17008) );
  INV_X1 U12268 ( .A(n17022), .ZN(n17017) );
  NAND2_X1 U12269 ( .A1(n17017), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17016) );
  NOR2_X1 U12270 ( .A1(n17066), .A2(n9911), .ZN(n17027) );
  NAND2_X1 U12271 ( .A1(n9912), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n9911) );
  INV_X1 U12272 ( .A(n17031), .ZN(n9912) );
  NOR2_X1 U12273 ( .A1(n10286), .A2(n9909), .ZN(n9908) );
  INV_X1 U12274 ( .A(n17059), .ZN(n17055) );
  NAND2_X1 U12275 ( .A1(n17070), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17066) );
  NAND2_X1 U12276 ( .A1(n17096), .A2(n9913), .ZN(n17075) );
  AND2_X1 U12277 ( .A1(n16988), .A2(n9720), .ZN(n9913) );
  NOR2_X1 U12278 ( .A1(n17180), .A2(n17098), .ZN(n17096) );
  NOR2_X1 U12279 ( .A1(n17999), .A2(n17130), .ZN(n17097) );
  INV_X1 U12280 ( .A(n17097), .ZN(n17123) );
  INV_X1 U12281 ( .A(n17133), .ZN(n17128) );
  INV_X1 U12282 ( .A(n10371), .ZN(n17131) );
  AND2_X1 U12283 ( .A1(n18418), .A2(n16987), .ZN(n17132) );
  INV_X1 U12284 ( .A(n16987), .ZN(n17130) );
  CLKBUF_X1 U12286 ( .A(n17246), .Z(n17239) );
  INV_X1 U12287 ( .A(n17249), .ZN(n17240) );
  OR2_X1 U12288 ( .A1(n18453), .A2(n17200), .ZN(n17249) );
  NOR2_X1 U12289 ( .A1(n17239), .A2(n17971), .ZN(n17247) );
  AND2_X1 U12290 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17524) );
  INV_X1 U12291 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17526) );
  INV_X1 U12292 ( .A(n17470), .ZN(n17533) );
  INV_X1 U12293 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20781) );
  AND2_X1 U12294 ( .A1(n17582), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17567) );
  NAND2_X1 U12295 ( .A1(n18254), .A2(n18303), .ZN(n17991) );
  NOR2_X1 U12296 ( .A1(n18619), .A2(n16314), .ZN(n17611) );
  OAI21_X1 U12297 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18616), .A(n16314), 
        .ZN(n17622) );
  INV_X1 U12298 ( .A(n17611), .ZN(n17626) );
  NAND2_X1 U12299 ( .A1(n17362), .A2(n10221), .ZN(n17309) );
  INV_X1 U12300 ( .A(n17862), .ZN(n17807) );
  NAND2_X1 U12301 ( .A1(n9986), .A2(n9987), .ZN(n17553) );
  NAND2_X1 U12302 ( .A1(n17564), .A2(n9988), .ZN(n9986) );
  NAND2_X1 U12303 ( .A1(n17564), .A2(n17565), .ZN(n17563) );
  AOI21_X2 U12304 ( .B1(n14131), .B2(n12517), .A(n18459), .ZN(n17934) );
  CLKBUF_X1 U12305 ( .A(n17835), .Z(n17950) );
  INV_X1 U12306 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20778) );
  INV_X1 U12307 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18584) );
  AOI211_X2 U12308 ( .C1(n18617), .C2(n18439), .A(n17967), .B(n14132), .ZN(
        n18599) );
  INV_X1 U12309 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18566) );
  INV_X1 U12310 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18488) );
  NAND2_X1 U12311 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18488), .ZN(n18629) );
  AND2_X2 U12312 ( .A1(n13205), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20007)
         );
  CLKBUF_X1 U12313 ( .A(n16296), .Z(n16298) );
  INV_X1 U12314 ( .A(n14584), .ZN(n14330) );
  AOI21_X1 U12315 ( .B1(n12153), .B2(n19934), .A(n12152), .ZN(n12154) );
  NAND2_X1 U12316 ( .A1(n14584), .A2(n19979), .ZN(n9789) );
  NOR2_X1 U12317 ( .A1(n9816), .A2(n14770), .ZN(n14771) );
  INV_X1 U12318 ( .A(n13191), .ZN(n13192) );
  OAI21_X1 U12319 ( .B1(n14199), .B2(n18888), .A(n13190), .ZN(n13191) );
  NOR2_X1 U12320 ( .A1(n9868), .A2(n14982), .ZN(n9867) );
  AOI21_X1 U12321 ( .B1(n16043), .B2(n16112), .A(n16042), .ZN(n16044) );
  AOI21_X1 U12322 ( .B1(n14203), .B2(n18993), .A(n10073), .ZN(n14204) );
  AOI211_X1 U12323 ( .C1(n15139), .C2(n16152), .A(n15138), .B(n15137), .ZN(
        n15140) );
  INV_X1 U12324 ( .A(n9840), .ZN(n15163) );
  NAND2_X1 U12325 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15299) );
  AOI21_X1 U12326 ( .B1(n17264), .B2(n17263), .A(n17262), .ZN(n17265) );
  NAND2_X1 U12327 ( .A1(n9752), .A2(n9671), .ZN(P3_U2803) );
  NAND2_X1 U12328 ( .A1(n9754), .A2(n9753), .ZN(n9752) );
  NOR2_X1 U12329 ( .A1(n9751), .A2(n9749), .ZN(n9748) );
  AND2_X2 U12330 ( .A1(n11193), .A2(n13475), .ZN(n11272) );
  INV_X2 U12331 ( .A(n10235), .ZN(n16933) );
  AND2_X1 U12332 ( .A1(n13342), .A2(n12808), .ZN(n10869) );
  OR3_X1 U12333 ( .A1(n10465), .A2(n9821), .A3(n9820), .ZN(n9635) );
  NOR2_X1 U12334 ( .A1(n13940), .A2(n9645), .ZN(n13523) );
  NAND2_X1 U12335 ( .A1(n12604), .A2(n12623), .ZN(n9768) );
  INV_X1 U12336 ( .A(n12536), .ZN(n9894) );
  XNOR2_X1 U12337 ( .A(n12163), .B(n12165), .ZN(n12857) );
  AND2_X1 U12338 ( .A1(n14823), .A2(n15052), .ZN(n9636) );
  NAND2_X1 U12339 ( .A1(n15271), .A2(n9706), .ZN(n14807) );
  NAND2_X1 U12340 ( .A1(n12373), .A2(n9689), .ZN(n9637) );
  NOR2_X1 U12341 ( .A1(n15058), .A2(n9845), .ZN(n15029) );
  NAND2_X1 U12342 ( .A1(n14364), .A2(n14365), .ZN(n14362) );
  NAND2_X1 U12343 ( .A1(n12202), .A2(n12203), .ZN(n12256) );
  OR2_X1 U12344 ( .A1(n13864), .A2(n11747), .ZN(n9638) );
  NOR2_X1 U12345 ( .A1(n10463), .A2(n18736), .ZN(n10451) );
  OAI21_X1 U12346 ( .B1(n9894), .B2(n12539), .A(n9902), .ZN(n9901) );
  AND2_X1 U12347 ( .A1(n9992), .A2(n17428), .ZN(n9640) );
  AND2_X1 U12348 ( .A1(n12886), .A2(n10072), .ZN(n9641) );
  INV_X1 U12349 ( .A(n11596), .ZN(n9970) );
  AND2_X1 U12350 ( .A1(n13745), .A2(n13746), .ZN(n9642) );
  AND2_X1 U12351 ( .A1(n12312), .A2(n9695), .ZN(n9643) );
  AND2_X1 U12352 ( .A1(n9809), .A2(n13945), .ZN(n9644) );
  INV_X1 U12353 ( .A(n9885), .ZN(n9884) );
  NAND2_X1 U12354 ( .A1(n13955), .A2(n16155), .ZN(n9885) );
  OR2_X1 U12355 ( .A1(n9717), .A2(n13939), .ZN(n9645) );
  AND2_X1 U12356 ( .A1(n12470), .A2(n9839), .ZN(n9646) );
  AND2_X1 U12357 ( .A1(n10021), .A2(n18878), .ZN(n9647) );
  NOR3_X1 U12358 ( .A1(n10980), .A2(n13387), .A3(n9928), .ZN(n13388) );
  NAND2_X1 U12359 ( .A1(n10446), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10444) );
  NOR3_X1 U12360 ( .A1(n10465), .A2(n9821), .A3(n15039), .ZN(n10447) );
  NOR2_X1 U12361 ( .A1(n10463), .A2(n9824), .ZN(n10450) );
  NOR2_X1 U12362 ( .A1(n10465), .A2(n16037), .ZN(n10448) );
  NAND2_X1 U12363 ( .A1(n9935), .A2(n9693), .ZN(n14970) );
  AND2_X1 U12364 ( .A1(n13590), .A2(n10021), .ZN(n9648) );
  NAND2_X1 U12365 ( .A1(n9698), .A2(n9831), .ZN(n12820) );
  AND2_X1 U12366 ( .A1(n10035), .A2(n14062), .ZN(n9649) );
  OR2_X1 U12367 ( .A1(n12850), .A2(n12793), .ZN(n16137) );
  INV_X1 U12368 ( .A(n16137), .ZN(n19008) );
  AND2_X1 U12369 ( .A1(n12562), .A2(n16108), .ZN(n9650) );
  AND2_X1 U12370 ( .A1(n13523), .A2(n13531), .ZN(n13530) );
  AND2_X2 U12371 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13475) );
  AND2_X1 U12372 ( .A1(n12840), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9651) );
  AND2_X1 U12373 ( .A1(n9910), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9652) );
  INV_X1 U12374 ( .A(n9768), .ZN(n12680) );
  INV_X1 U12375 ( .A(n16804), .ZN(n16941) );
  NAND2_X1 U12376 ( .A1(n12478), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15037) );
  INV_X1 U12377 ( .A(n11445), .ZN(n10027) );
  INV_X2 U12378 ( .A(n10661), .ZN(n10675) );
  NOR2_X1 U12379 ( .A1(n14053), .A2(n10033), .ZN(n14119) );
  NOR2_X1 U12380 ( .A1(n10064), .A2(n10066), .ZN(n15057) );
  NOR2_X1 U12381 ( .A1(n14312), .A2(n14315), .ZN(n14314) );
  NAND2_X1 U12382 ( .A1(n12479), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12552) );
  AND2_X1 U12383 ( .A1(n14364), .A2(n10039), .ZN(n14344) );
  AND2_X1 U12384 ( .A1(n14364), .A2(n10041), .ZN(n14350) );
  INV_X1 U12385 ( .A(n11317), .ZN(n12713) );
  NAND2_X1 U12386 ( .A1(n12373), .A2(n9949), .ZN(n9653) );
  OR2_X1 U12387 ( .A1(n14705), .A2(n15911), .ZN(n9654) );
  AND4_X1 U12388 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(
        n9655) );
  NAND2_X1 U12389 ( .A1(n14848), .A2(n9864), .ZN(n12480) );
  NAND2_X1 U12390 ( .A1(n10032), .A2(n11863), .ZN(n14107) );
  AND4_X1 U12391 ( .A1(n10187), .A2(n10186), .A3(n10185), .A4(n10184), .ZN(
        n9656) );
  NAND2_X1 U12392 ( .A1(n9967), .A2(n9968), .ZN(n14534) );
  NAND2_X1 U12393 ( .A1(n12199), .A2(n12182), .ZN(n19022) );
  INV_X1 U12394 ( .A(n19022), .ZN(n19033) );
  INV_X1 U12395 ( .A(n11444), .ZN(n10028) );
  NAND2_X1 U12396 ( .A1(n9898), .A2(n9899), .ZN(n14990) );
  NAND2_X1 U12397 ( .A1(n10063), .A2(n12323), .ZN(n15406) );
  NOR2_X1 U12398 ( .A1(n16380), .A2(n9733), .ZN(n9658) );
  NAND2_X1 U12399 ( .A1(n12869), .A2(n12860), .ZN(n13391) );
  NAND2_X1 U12400 ( .A1(n10057), .A2(n15047), .ZN(n15043) );
  AND4_X1 U12401 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n9659) );
  INV_X1 U12402 ( .A(n13645), .ZN(n10577) );
  AND4_X1 U12403 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n9660) );
  NAND2_X1 U12404 ( .A1(n9969), .A2(n9599), .ZN(n14568) );
  AND4_X1 U12405 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n9661) );
  NOR2_X1 U12406 ( .A1(n15316), .A2(n15289), .ZN(n15291) );
  INV_X1 U12407 ( .A(n15291), .ZN(n9742) );
  NOR3_X1 U12408 ( .A1(n12543), .A2(n12280), .A3(n14201), .ZN(n9662) );
  NOR2_X1 U12409 ( .A1(n13104), .A2(n10008), .ZN(n14842) );
  NOR2_X1 U12410 ( .A1(n10660), .A2(n12810), .ZN(n9663) );
  NOR2_X1 U12411 ( .A1(n16351), .A2(n16352), .ZN(n9664) );
  AND2_X1 U12412 ( .A1(n12179), .A2(n19007), .ZN(n12233) );
  NOR2_X1 U12413 ( .A1(n17138), .A2(n17999), .ZN(n9665) );
  XNOR2_X1 U12414 ( .A(n14764), .B(n12554), .ZN(n14199) );
  OR2_X1 U12415 ( .A1(n12851), .A2(n18996), .ZN(n9666) );
  AND2_X1 U12417 ( .A1(n9773), .A2(n11444), .ZN(n9667) );
  OR2_X1 U12418 ( .A1(n12851), .A2(n18980), .ZN(n9668) );
  NAND2_X1 U12419 ( .A1(n12162), .A2(n12166), .ZN(n18871) );
  AND2_X1 U12420 ( .A1(n11408), .A2(n9771), .ZN(n9670) );
  AND2_X1 U12421 ( .A1(n17274), .A2(n9748), .ZN(n9671) );
  NOR2_X1 U12422 ( .A1(n15161), .A2(n9841), .ZN(n9672) );
  NAND2_X1 U12423 ( .A1(n12202), .A2(n13653), .ZN(n19174) );
  AND2_X1 U12424 ( .A1(n14930), .A2(n14791), .ZN(n14789) );
  AND2_X1 U12425 ( .A1(n14539), .A2(n15911), .ZN(n9673) );
  AND2_X1 U12426 ( .A1(n10027), .A2(n11444), .ZN(n9674) );
  NOR3_X1 U12427 ( .A1(n15060), .A2(n9860), .A3(n9858), .ZN(n9857) );
  INV_X1 U12428 ( .A(n10206), .ZN(n9983) );
  AND2_X1 U12429 ( .A1(n19055), .A2(n19071), .ZN(n9676) );
  OR2_X1 U12430 ( .A1(n9662), .A2(n9904), .ZN(n9677) );
  INV_X1 U12431 ( .A(n17428), .ZN(n17531) );
  OR2_X1 U12432 ( .A1(n10360), .A2(n17971), .ZN(n9678) );
  AND2_X1 U12433 ( .A1(n12680), .A2(n9764), .ZN(n9679) );
  AND2_X1 U12434 ( .A1(n12276), .A2(n12281), .ZN(n9680) );
  OR2_X1 U12435 ( .A1(n10437), .A2(n10436), .ZN(n9681) );
  AND2_X1 U12436 ( .A1(n9848), .A2(n9847), .ZN(n9682) );
  NOR2_X1 U12437 ( .A1(n14582), .A2(n14583), .ZN(n9683) );
  AND2_X1 U12438 ( .A1(n12424), .A2(n15176), .ZN(n12538) );
  INV_X1 U12439 ( .A(n12538), .ZN(n9903) );
  OR2_X1 U12440 ( .A1(n16349), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n9684) );
  INV_X1 U12441 ( .A(n10846), .ZN(n12804) );
  NAND2_X1 U12442 ( .A1(n13381), .A2(n13382), .ZN(n13383) );
  NAND2_X1 U12443 ( .A1(n9960), .A2(n12411), .ZN(n12314) );
  NAND2_X1 U12444 ( .A1(n12313), .A2(n12312), .ZN(n14169) );
  NOR2_X1 U12445 ( .A1(n16119), .A2(n9937), .ZN(n14969) );
  NOR2_X1 U12446 ( .A1(n14878), .A2(n14880), .ZN(n14879) );
  NOR2_X1 U12447 ( .A1(n13902), .A2(n9869), .ZN(n13821) );
  NOR2_X1 U12448 ( .A1(n16119), .A2(n16118), .ZN(n13810) );
  NAND2_X1 U12449 ( .A1(n13987), .A2(n9783), .ZN(n14073) );
  AND2_X1 U12450 ( .A1(n17567), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10413) );
  NOR2_X1 U12451 ( .A1(n10457), .A2(n20762), .ZN(n10454) );
  NOR2_X1 U12452 ( .A1(n10460), .A2(n16095), .ZN(n10453) );
  NOR2_X1 U12453 ( .A1(n10462), .A2(n16079), .ZN(n10452) );
  NOR2_X1 U12454 ( .A1(n10464), .A2(n20750), .ZN(n10449) );
  INV_X1 U12455 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11184) );
  AND2_X1 U12456 ( .A1(n10037), .A2(n10038), .ZN(n9685) );
  AND2_X1 U12457 ( .A1(n17017), .A2(n9910), .ZN(n9686) );
  NAND2_X2 U12458 ( .A1(n17403), .A2(n17428), .ZN(n17362) );
  INV_X1 U12459 ( .A(n9756), .ZN(n14126) );
  NAND2_X1 U12460 ( .A1(n9758), .A2(n9757), .ZN(n9756) );
  NAND2_X1 U12461 ( .A1(n10037), .A2(n9649), .ZN(n14061) );
  INV_X1 U12462 ( .A(n10612), .ZN(n12795) );
  OAI22_X1 U12463 ( .A1(n13935), .A2(n13936), .B1(n18833), .B2(n13938), .ZN(
        n15430) );
  OR3_X1 U12464 ( .A1(n14705), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9687) );
  XNOR2_X1 U12465 ( .A(n12446), .B(n12445), .ZN(n13932) );
  NAND2_X1 U12466 ( .A1(n15121), .A2(n12470), .ZN(n15107) );
  AND2_X1 U12467 ( .A1(n13781), .A2(n12879), .ZN(n13382) );
  OR2_X1 U12468 ( .A1(n10885), .A2(n10884), .ZN(n11146) );
  OR2_X1 U12469 ( .A1(n16382), .A2(n17310), .ZN(n9688) );
  NOR2_X1 U12470 ( .A1(n17379), .A2(n17380), .ZN(n10407) );
  AND2_X1 U12471 ( .A1(n13821), .A2(n13927), .ZN(n13926) );
  NOR2_X1 U12472 ( .A1(n10456), .A2(n20802), .ZN(n10455) );
  NOR2_X1 U12473 ( .A1(n15060), .A2(n15061), .ZN(n14816) );
  AND2_X1 U12474 ( .A1(n12365), .A2(n9952), .ZN(n9689) );
  OR2_X1 U12475 ( .A1(n10463), .A2(n9825), .ZN(n9690) );
  AND2_X1 U12476 ( .A1(n10454), .A2(n9822), .ZN(n9691) );
  AND2_X1 U12477 ( .A1(n9822), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9692) );
  OR2_X1 U12478 ( .A1(n10926), .A2(n10925), .ZN(n12229) );
  NOR2_X1 U12479 ( .A1(n9937), .A2(n9936), .ZN(n9693) );
  INV_X1 U12480 ( .A(n13864), .ZN(n10037) );
  INV_X1 U12481 ( .A(n11488), .ZN(n20158) );
  NAND2_X1 U12482 ( .A1(n11486), .A2(n11485), .ZN(n11488) );
  INV_X1 U12483 ( .A(n14878), .ZN(n10014) );
  AND3_X1 U12484 ( .A1(n13211), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n12548), .ZN(n9694) );
  AND2_X1 U12485 ( .A1(n10088), .A2(n12320), .ZN(n9695) );
  INV_X1 U12486 ( .A(n14053), .ZN(n10032) );
  INV_X1 U12487 ( .A(n9932), .ZN(n15634) );
  NAND2_X1 U12488 ( .A1(n15271), .A2(n9933), .ZN(n9932) );
  INV_X1 U12489 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20702) );
  OR2_X1 U12490 ( .A1(n12307), .A2(n9946), .ZN(n9696) );
  INV_X1 U12491 ( .A(n10036), .ZN(n10035) );
  NAND2_X1 U12492 ( .A1(n10038), .A2(n13985), .ZN(n10036) );
  AND2_X1 U12493 ( .A1(n9884), .A2(n12548), .ZN(n9697) );
  INV_X1 U12494 ( .A(n9859), .ZN(n14817) );
  NOR2_X1 U12495 ( .A1(n15060), .A2(n9860), .ZN(n9859) );
  AND2_X1 U12496 ( .A1(n10613), .A2(n9833), .ZN(n9698) );
  AND2_X1 U12497 ( .A1(n13216), .A2(n13217), .ZN(n13214) );
  INV_X1 U12498 ( .A(n9880), .ZN(n9879) );
  NAND2_X1 U12499 ( .A1(n13891), .A2(n9881), .ZN(n9880) );
  AND2_X1 U12500 ( .A1(n14345), .A2(n10039), .ZN(n9699) );
  AND2_X1 U12501 ( .A1(n12680), .A2(n9765), .ZN(n9700) );
  NOR2_X1 U12502 ( .A1(n14797), .A2(n10466), .ZN(n9701) );
  AND2_X1 U12503 ( .A1(n10007), .A2(n10006), .ZN(n9702) );
  OR2_X1 U12504 ( .A1(n10465), .A2(n9821), .ZN(n9703) );
  AND2_X1 U12505 ( .A1(n20700), .A2(n20771), .ZN(n14157) );
  NAND2_X1 U12506 ( .A1(n9921), .A2(n9919), .ZN(n13732) );
  NAND2_X1 U12507 ( .A1(n13590), .A2(n9641), .ZN(n13816) );
  AND2_X1 U12508 ( .A1(n13590), .A2(n12886), .ZN(n9704) );
  INV_X1 U12509 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U12510 ( .A1(n13530), .A2(n9848), .ZN(n13540) );
  NOR2_X1 U12511 ( .A1(n9635), .A2(n16029), .ZN(n10446) );
  OR2_X1 U12512 ( .A1(n10443), .A2(n12489), .ZN(n9705) );
  AND2_X2 U12513 ( .A1(n10823), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12953) );
  INV_X1 U12514 ( .A(n13925), .ZN(n10022) );
  AND2_X1 U12515 ( .A1(n9933), .A2(n14819), .ZN(n9706) );
  NOR2_X1 U12516 ( .A1(n9852), .A2(n9850), .ZN(n13544) );
  AND2_X1 U12517 ( .A1(n13590), .A2(n9647), .ZN(n13991) );
  AOI21_X1 U12518 ( .B1(n13429), .B2(n10889), .A(n10888), .ZN(n10893) );
  AND2_X1 U12519 ( .A1(n13530), .A2(n9682), .ZN(n13591) );
  AND2_X1 U12520 ( .A1(n9925), .A2(n9924), .ZN(n9707) );
  INV_X1 U12521 ( .A(n10980), .ZN(n13362) );
  OAI21_X1 U12522 ( .B1(n10443), .B2(n9805), .A(n9803), .ZN(n12562) );
  AND2_X1 U12523 ( .A1(n9779), .A2(n9778), .ZN(n9708) );
  AND2_X1 U12524 ( .A1(n14366), .A2(n14359), .ZN(n9709) );
  INV_X1 U12525 ( .A(n13530), .ZN(n9852) );
  OR2_X1 U12526 ( .A1(n13940), .A2(n13939), .ZN(n9846) );
  OR2_X1 U12527 ( .A1(n15293), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9710) );
  AND2_X1 U12528 ( .A1(n15019), .A2(n9810), .ZN(n9711) );
  AND2_X1 U12529 ( .A1(n9986), .A2(n9984), .ZN(n9712) );
  AND2_X1 U12530 ( .A1(n9706), .A2(n9931), .ZN(n9713) );
  AND2_X1 U12531 ( .A1(n9640), .A2(n9991), .ZN(n9714) );
  AND2_X1 U12532 ( .A1(n13383), .A2(n12880), .ZN(n9715) );
  INV_X1 U12533 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n9764) );
  AND2_X1 U12534 ( .A1(n9844), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9716) );
  INV_X1 U12535 ( .A(n12984), .ZN(n13615) );
  INV_X1 U12536 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13879) );
  NAND2_X1 U12537 ( .A1(n13500), .A2(n13499), .ZN(n13744) );
  INV_X1 U12538 ( .A(n13744), .ZN(n9777) );
  AND2_X1 U12539 ( .A1(n10609), .A2(n10608), .ZN(n9717) );
  AND2_X1 U12540 ( .A1(n12680), .A2(n20798), .ZN(n9718) );
  INV_X1 U12541 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n9726) );
  INV_X1 U12542 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9765) );
  OR2_X1 U12543 ( .A1(n15950), .A2(n20380), .ZN(n20006) );
  INV_X1 U12544 ( .A(n20006), .ZN(n19934) );
  INV_X1 U12545 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n9950) );
  INV_X1 U12546 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9727) );
  INV_X1 U12547 ( .A(n17452), .ZN(n16532) );
  INV_X1 U12548 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n9839) );
  OR2_X1 U12549 ( .A1(n11613), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9719) );
  AND2_X1 U12550 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n9720) );
  AND2_X1 U12551 ( .A1(n10070), .A2(n10069), .ZN(n9721) );
  INV_X1 U12552 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9767) );
  INV_X1 U12553 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n9786) );
  INV_X1 U12554 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9823) );
  INV_X1 U12555 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9723) );
  INV_X1 U12556 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9770) );
  INV_X1 U12557 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n9959) );
  AOI22_X2 U12558 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20048), .B1(DATAI_21_), 
        .B2(n20008), .ZN(n20504) );
  AOI22_X2 U12559 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20048), .B1(DATAI_16_), 
        .B2(n20008), .ZN(n20484) );
  AOI22_X2 U12560 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20048), .B1(DATAI_18_), 
        .B2(n20008), .ZN(n20492) );
  AOI22_X2 U12561 ( .A1(DATAI_22_), .A2(n20008), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20048), .ZN(n20508) );
  NOR3_X4 U12562 ( .A1(n18249), .A2(n18133), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18222) );
  NAND3_X1 U12563 ( .A1(n16347), .A2(n16348), .A3(n9684), .ZN(P3_U2642) );
  INV_X1 U12564 ( .A(n9728), .ZN(n10420) );
  CLKBUF_X1 U12565 ( .A(n16603), .Z(n9733) );
  NAND2_X2 U12566 ( .A1(n9736), .A2(n13342), .ZN(n10846) );
  NAND4_X1 U12567 ( .A1(n9736), .A2(n12747), .A3(n13165), .A4(n12816), .ZN(
        n10628) );
  NAND2_X1 U12568 ( .A1(n12226), .A2(n13231), .ZN(n9744) );
  AND2_X2 U12569 ( .A1(n9743), .A2(n12211), .ZN(n12287) );
  NAND4_X1 U12570 ( .A1(n12207), .A2(n12206), .A3(n12208), .A4(n12209), .ZN(
        n9743) );
  NAND2_X2 U12571 ( .A1(n9744), .A2(n12228), .ZN(n12286) );
  NAND2_X1 U12572 ( .A1(n15083), .A2(n15343), .ZN(n9745) );
  NAND2_X1 U12573 ( .A1(n15083), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16104) );
  NAND2_X1 U12574 ( .A1(n15083), .A2(n15085), .ZN(n15263) );
  NOR2_X1 U12575 ( .A1(n15083), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16101) );
  NAND2_X1 U12576 ( .A1(n12464), .A2(n9827), .ZN(n9826) );
  NAND2_X1 U12577 ( .A1(n9747), .A2(n9746), .ZN(n15441) );
  NAND2_X1 U12578 ( .A1(n12459), .A2(n13933), .ZN(n9747) );
  INV_X2 U12579 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18598) );
  OAI22_X2 U12580 ( .A1(n17494), .A2(n17818), .B1(n17820), .B2(n17626), .ZN(
        n17483) );
  NOR2_X2 U12581 ( .A1(n17625), .A2(n17103), .ZN(n17529) );
  NAND2_X2 U12582 ( .A1(n11494), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11495) );
  NAND2_X1 U12583 ( .A1(n12680), .A2(n9767), .ZN(n9766) );
  AOI22_X1 U12584 ( .A1(n12601), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n9768), .B2(P1_EBX_REG_30__SCAN_IN), .ZN(n14278) );
  AOI22_X1 U12585 ( .A1(n12601), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n9768), .B2(P1_EBX_REG_31__SCAN_IN), .ZN(n12600) );
  NAND2_X1 U12586 ( .A1(n12680), .A2(n9770), .ZN(n9769) );
  AOI21_X2 U12587 ( .B1(n14455), .B2(n9634), .A(n12566), .ZN(n12567) );
  OR3_X1 U12588 ( .A1(n12566), .A2(n9634), .A3(n9687), .ZN(n9774) );
  OR2_X1 U12589 ( .A1(n12566), .A2(n9687), .ZN(n9775) );
  AND2_X2 U12590 ( .A1(n15826), .A2(n15825), .ZN(n11608) );
  NOR2_X2 U12591 ( .A1(n13754), .A2(n13755), .ZN(n15934) );
  INV_X1 U12592 ( .A(n9782), .ZN(n14296) );
  NAND2_X1 U12593 ( .A1(n12623), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12611) );
  NAND2_X1 U12594 ( .A1(n12623), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12619) );
  OAI22_X1 U12595 ( .A1(n9633), .A2(n13802), .B1(n12623), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13519) );
  NAND2_X1 U12596 ( .A1(n12623), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n9784) );
  OAI21_X1 U12597 ( .B1(n12601), .B2(P1_EBX_REG_3__SCAN_IN), .A(n12623), .ZN(
        n9788) );
  OAI211_X1 U12598 ( .C1(n14585), .C2(n19996), .A(n9683), .B(n9789), .ZN(
        P1_U3001) );
  XNOR2_X1 U12599 ( .A(n14279), .B(n9790), .ZN(n14584) );
  OR2_X2 U12600 ( .A1(n14361), .A2(n14353), .ZN(n14355) );
  OAI21_X2 U12601 ( .B1(n12463), .B2(n12548), .A(n18809), .ZN(n12311) );
  OAI21_X1 U12602 ( .B1(n10577), .B2(n10627), .A(n12765), .ZN(n10780) );
  INV_X1 U12603 ( .A(n14798), .ZN(n9808) );
  NAND3_X1 U12604 ( .A1(n9636), .A2(n9814), .A3(n9813), .ZN(n9812) );
  NAND2_X1 U12605 ( .A1(n9814), .A2(n14823), .ZN(n14803) );
  INV_X1 U12606 ( .A(n9815), .ZN(n14802) );
  NAND2_X1 U12607 ( .A1(n9827), .A2(n15439), .ZN(n12469) );
  OAI211_X2 U12608 ( .C1(n9827), .C2(n12468), .A(n9826), .B(n12466), .ZN(
        n15122) );
  INV_X1 U12609 ( .A(n9831), .ZN(n9829) );
  NAND3_X1 U12610 ( .A1(n10613), .A2(n19045), .A3(n9833), .ZN(n9830) );
  AND2_X1 U12611 ( .A1(n10837), .A2(n10841), .ZN(n12814) );
  NAND2_X2 U12612 ( .A1(n9676), .A2(n9832), .ZN(n10622) );
  NAND2_X1 U12613 ( .A1(n10837), .A2(n10610), .ZN(n9831) );
  INV_X1 U12614 ( .A(n9996), .ZN(n9833) );
  NAND2_X1 U12615 ( .A1(n9646), .A2(n15121), .ZN(n9837) );
  NAND3_X1 U12616 ( .A1(n9837), .A2(n14174), .A3(n9836), .ZN(n14173) );
  OAI21_X2 U12617 ( .B1(n15121), .B2(n9839), .A(n9838), .ZN(n14174) );
  OR2_X1 U12618 ( .A1(n12479), .A2(n18996), .ZN(n9843) );
  INV_X1 U12619 ( .A(n9846), .ZN(n13522) );
  NAND3_X1 U12620 ( .A1(n9666), .A2(n9854), .A3(n9853), .ZN(P2_U3015) );
  NAND2_X1 U12621 ( .A1(n16001), .A2(n19008), .ZN(n9853) );
  INV_X1 U12622 ( .A(n9857), .ZN(n14859) );
  NAND2_X1 U12623 ( .A1(n14848), .A2(n14847), .ZN(n14850) );
  AOI21_X1 U12624 ( .B1(n14985), .B2(n16113), .A(n9866), .ZN(n14986) );
  OAI21_X1 U12625 ( .B1(n14199), .B2(n19026), .A(n9867), .ZN(n9866) );
  INV_X1 U12626 ( .A(n12808), .ZN(n10578) );
  NOR2_X1 U12627 ( .A1(n12875), .A2(n12172), .ZN(n12179) );
  NAND2_X1 U12628 ( .A1(n15376), .A2(n12343), .ZN(n9872) );
  NAND2_X1 U12629 ( .A1(n9872), .A2(n9873), .ZN(n12393) );
  OAI21_X1 U12630 ( .B1(n13894), .B2(n12548), .A(n9884), .ZN(n13890) );
  NAND2_X1 U12631 ( .A1(n13894), .A2(n9877), .ZN(n9876) );
  NAND2_X1 U12632 ( .A1(n12537), .A2(n12536), .ZN(n9898) );
  NAND2_X1 U12633 ( .A1(n9895), .A2(n9887), .ZN(n12551) );
  AOI21_X2 U12634 ( .B1(n9901), .B2(n9890), .A(n9677), .ZN(n9889) );
  NAND2_X1 U12635 ( .A1(n9897), .A2(n14988), .ZN(n9896) );
  NAND2_X1 U12636 ( .A1(n15628), .A2(n18617), .ZN(n9915) );
  NAND2_X1 U12637 ( .A1(n14128), .A2(n14127), .ZN(n9918) );
  OR3_X1 U12638 ( .A1(n10893), .A2(n13603), .A3(n10890), .ZN(n9921) );
  INV_X1 U12639 ( .A(n10893), .ZN(n9922) );
  NAND2_X2 U12640 ( .A1(n10560), .A2(n10559), .ZN(n10841) );
  NAND3_X1 U12641 ( .A1(n10560), .A2(n10559), .A3(n19700), .ZN(n10847) );
  AND2_X2 U12642 ( .A1(n10612), .A2(n12808), .ZN(n9996) );
  NAND2_X1 U12643 ( .A1(n12795), .A2(n12808), .ZN(n10837) );
  NOR2_X2 U12644 ( .A1(n12534), .A2(n12427), .ZN(n12537) );
  OR2_X2 U12645 ( .A1(n9940), .A2(n15011), .ZN(n12534) );
  NOR2_X4 U12646 ( .A1(n12368), .A2(n9942), .ZN(n12360) );
  NAND3_X1 U12647 ( .A1(n9945), .A2(n9680), .A3(n11148), .ZN(n9944) );
  NOR2_X2 U12648 ( .A1(n9944), .A2(n9943), .ZN(n12319) );
  NAND2_X1 U12649 ( .A1(n12373), .A2(n12365), .ZN(n12364) );
  NOR2_X2 U12650 ( .A1(n14482), .A2(n12736), .ZN(n12566) );
  OAI21_X2 U12651 ( .B1(n13769), .B2(n9964), .A(n9961), .ZN(n19929) );
  NAND2_X1 U12652 ( .A1(n11495), .A2(n9963), .ZN(n9962) );
  INV_X1 U12653 ( .A(n11495), .ZN(n9964) );
  NAND2_X1 U12654 ( .A1(n13767), .A2(n11495), .ZN(n19931) );
  NAND2_X1 U12655 ( .A1(n13769), .A2(n13768), .ZN(n13767) );
  XNOR2_X1 U12656 ( .A(n11494), .B(n12614), .ZN(n13769) );
  NAND2_X1 U12657 ( .A1(n14010), .A2(n9599), .ZN(n9967) );
  NAND2_X2 U12658 ( .A1(n9972), .A2(n11606), .ZN(n15826) );
  AND2_X1 U12659 ( .A1(n9973), .A2(n11388), .ZN(n11353) );
  NAND2_X1 U12660 ( .A1(n11339), .A2(n11338), .ZN(n9973) );
  NAND2_X1 U12661 ( .A1(n11608), .A2(n9977), .ZN(n9976) );
  NAND2_X1 U12662 ( .A1(n17564), .A2(n9982), .ZN(n9981) );
  INV_X1 U12663 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9990) );
  NAND3_X1 U12664 ( .A1(n9640), .A2(n9991), .A3(n17847), .ZN(n17502) );
  INV_X1 U12665 ( .A(n17536), .ZN(n9991) );
  NOR2_X2 U12666 ( .A1(n17279), .A2(n10226), .ZN(n10227) );
  NOR2_X2 U12667 ( .A1(n16663), .A2(n10103), .ZN(n10143) );
  INV_X1 U12668 ( .A(n13382), .ZN(n9998) );
  OAI211_X1 U12669 ( .C1(n13381), .C2(n9999), .A(n9997), .B(n13779), .ZN(
        n13521) );
  NOR2_X1 U12670 ( .A1(n14878), .A2(n10019), .ZN(n14872) );
  AND2_X2 U12671 ( .A1(n13476), .A2(n13475), .ZN(n11283) );
  AND2_X2 U12672 ( .A1(n13476), .A2(n11195), .ZN(n11271) );
  AND2_X2 U12673 ( .A1(n11194), .A2(n13476), .ZN(n11766) );
  AND2_X2 U12674 ( .A1(n11191), .A2(n13476), .ZN(n11392) );
  AND2_X2 U12675 ( .A1(n11185), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13476) );
  NAND2_X1 U12676 ( .A1(n11684), .A2(n10026), .ZN(n10025) );
  INV_X1 U12677 ( .A(n14053), .ZN(n10029) );
  NAND2_X1 U12678 ( .A1(n10029), .A2(n10030), .ZN(n14120) );
  NOR2_X2 U12679 ( .A1(n13864), .A2(n10036), .ZN(n13982) );
  AND2_X2 U12680 ( .A1(n14364), .A2(n9699), .ZN(n14337) );
  NAND2_X1 U12681 ( .A1(n14303), .A2(n10045), .ZN(n14272) );
  NAND2_X1 U12682 ( .A1(n10048), .A2(n10547), .ZN(n10047) );
  NAND4_X1 U12683 ( .A1(n10497), .A2(n10498), .A3(n10496), .A4(n10495), .ZN(
        n10048) );
  NAND2_X1 U12684 ( .A1(n10050), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10049) );
  NAND4_X1 U12685 ( .A1(n10501), .A2(n10502), .A3(n10499), .A4(n10500), .ZN(
        n10050) );
  NAND2_X1 U12686 ( .A1(n15049), .A2(n10052), .ZN(n10051) );
  XNOR2_X2 U12687 ( .A(n12157), .B(n12156), .ZN(n12875) );
  NAND2_X1 U12688 ( .A1(n10063), .A2(n10059), .ZN(n15376) );
  NAND2_X1 U12689 ( .A1(n15082), .A2(n10065), .ZN(n15058) );
  INV_X1 U12690 ( .A(n15058), .ZN(n12478) );
  NAND2_X1 U12691 ( .A1(n15082), .A2(n12477), .ZN(n15244) );
  NAND3_X2 U12692 ( .A1(n12286), .A2(n12287), .A3(n12229), .ZN(n12279) );
  NOR2_X1 U12693 ( .A1(n15001), .A2(n10068), .ZN(n14992) );
  AND2_X1 U12694 ( .A1(n20010), .A2(n11681), .ZN(n20469) );
  NAND2_X1 U12695 ( .A1(n15098), .A2(n15099), .ZN(n15097) );
  AOI21_X1 U12696 ( .B1(n14985), .B2(n16152), .A(n14206), .ZN(n14207) );
  NAND2_X1 U12697 ( .A1(n14239), .A2(n20044), .ZN(n13408) );
  NAND4_X1 U12698 ( .A1(n14251), .A2(n13425), .A3(n14239), .A4(n13557), .ZN(
        n12701) );
  XNOR2_X1 U12699 ( .A(n11455), .B(n11453), .ZN(n11673) );
  NAND2_X1 U12700 ( .A1(n15068), .A2(n15067), .ZN(n15069) );
  OR2_X1 U12701 ( .A1(n12791), .A2(n16147), .ZN(n12852) );
  NAND4_X2 U12702 ( .A1(n11258), .A2(n11257), .A3(n11256), .A4(n11255), .ZN(
        n11325) );
  OAI21_X2 U12703 ( .B1(n13829), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11368), 
        .ZN(n11369) );
  INV_X1 U12704 ( .A(n11352), .ZN(n20120) );
  INV_X1 U12705 ( .A(n19737), .ZN(n13646) );
  NAND2_X1 U12706 ( .A1(n14272), .A2(n12145), .ZN(n14208) );
  XNOR2_X1 U12707 ( .A(n13020), .B(n10071), .ZN(n14868) );
  INV_X1 U12708 ( .A(n11673), .ZN(n11675) );
  INV_X1 U12709 ( .A(n12462), .ZN(n12461) );
  NOR2_X1 U12710 ( .A1(n9613), .A2(n12467), .ZN(n12464) );
  OAI22_X1 U12711 ( .A1(n10681), .A2(n12156), .B1(n10680), .B2(n10679), .ZN(
        n13940) );
  INV_X1 U12712 ( .A(n12862), .ZN(n13375) );
  OAI21_X1 U12713 ( .B1(n18853), .B2(n12874), .A(n12861), .ZN(n12862) );
  OR2_X1 U12714 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  NAND2_X1 U12715 ( .A1(n12859), .A2(n12858), .ZN(n12869) );
  AOI22_X1 U12716 ( .A1(n13141), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10815), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U12717 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12205), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12206) );
  OAI21_X1 U12718 ( .B1(n9626), .B2(n12874), .A(n12856), .ZN(n12859) );
  AND2_X1 U12719 ( .A1(n9626), .A2(n12191), .ZN(n12183) );
  AND2_X1 U12720 ( .A1(n9626), .A2(n18853), .ZN(n12182) );
  XOR2_X1 U12721 ( .A(n13036), .B(n13039), .Z(n10071) );
  NAND2_X1 U12722 ( .A1(n14919), .A2(n13065), .ZN(n13081) );
  AND2_X1 U12723 ( .A1(n13813), .A2(n13817), .ZN(n10072) );
  NOR2_X1 U12724 ( .A1(n14202), .A2(n14201), .ZN(n10073) );
  OR3_X1 U12725 ( .A1(n15131), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15130), .ZN(n10074) );
  NOR2_X1 U12726 ( .A1(n18429), .A2(n10103), .ZN(n16697) );
  AND4_X1 U12727 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n10075) );
  AND2_X1 U12728 ( .A1(n14437), .A2(n14166), .ZN(n10076) );
  AND2_X1 U12729 ( .A1(n17437), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10077) );
  OR3_X1 U12730 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17340), .ZN(n10078) );
  AND2_X1 U12731 ( .A1(n10869), .A2(n12548), .ZN(n10079) );
  NOR2_X1 U12732 ( .A1(n12563), .A2(n9650), .ZN(n10080) );
  OR2_X1 U12733 ( .A1(n16603), .A2(n10415), .ZN(n10081) );
  AND2_X1 U12734 ( .A1(n13081), .A2(n10090), .ZN(n10082) );
  INV_X1 U12735 ( .A(n20636), .ZN(n20715) );
  OR2_X1 U12736 ( .A1(n14918), .A2(n14397), .ZN(n10083) );
  NOR2_X1 U12737 ( .A1(n20010), .A2(n11681), .ZN(n10084) );
  AND4_X1 U12738 ( .A1(n12242), .A2(n12241), .A3(n12240), .A4(n12239), .ZN(
        n10085) );
  INV_X1 U12739 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11864) );
  AND2_X1 U12740 ( .A1(n12746), .A2(n12745), .ZN(n10086) );
  INV_X1 U12741 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13792) );
  INV_X1 U12742 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11729) );
  INV_X2 U12743 ( .A(n16982), .ZN(n16969) );
  AND4_X1 U12744 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10087) );
  INV_X1 U12745 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15947) );
  INV_X1 U12746 ( .A(n15321), .ZN(n15066) );
  INV_X1 U12747 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15715) );
  INV_X1 U12748 ( .A(n12112), .ZN(n11685) );
  INV_X1 U12749 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20802) );
  INV_X1 U12750 ( .A(n14157), .ZN(n12120) );
  INV_X1 U12751 ( .A(n15110), .ZN(n12320) );
  NOR2_X1 U12752 ( .A1(n17475), .A2(n17364), .ZN(n17605) );
  OR2_X1 U12753 ( .A1(n12321), .A2(n14181), .ZN(n10088) );
  INV_X1 U12754 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15561) );
  INV_X1 U12755 ( .A(n19026), .ZN(n18985) );
  AND4_X1 U12756 ( .A1(n12237), .A2(n12236), .A3(n12235), .A4(n12234), .ZN(
        n10089) );
  AND2_X1 U12757 ( .A1(n13080), .A2(n13099), .ZN(n10090) );
  AND2_X2 U12758 ( .A1(n11195), .A2(n13479), .ZN(n11502) );
  INV_X1 U12759 ( .A(n12229), .ZN(n12445) );
  OR2_X1 U12760 ( .A1(n15232), .A2(n15231), .ZN(n10091) );
  INV_X1 U12761 ( .A(n12518), .ZN(n10214) );
  AND2_X1 U12762 ( .A1(n11179), .A2(n11178), .ZN(n10092) );
  AND2_X2 U12763 ( .A1(n18969), .A2(n13322), .ZN(n18967) );
  OR2_X1 U12764 ( .A1(n16481), .A2(n16463), .ZN(n10093) );
  AND2_X1 U12765 ( .A1(n12538), .A2(n12425), .ZN(n10095) );
  INV_X1 U12766 ( .A(n14286), .ZN(n14304) );
  AND4_X1 U12767 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(
        n10097) );
  INV_X1 U12768 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12187) );
  OR2_X1 U12769 ( .A1(n11367), .A2(n11366), .ZN(n11447) );
  NAND2_X1 U12770 ( .A1(n12174), .A2(n12173), .ZN(n12175) );
  AOI22_X1 U12771 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U12772 ( .A1(n11630), .A2(n11629), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20681), .ZN(n11626) );
  INV_X1 U12773 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11186) );
  OR2_X1 U12774 ( .A1(n11455), .A2(n11454), .ZN(n11456) );
  OR2_X1 U12775 ( .A1(n11559), .A2(n11558), .ZN(n11579) );
  OR2_X1 U12776 ( .A1(n11509), .A2(n11508), .ZN(n11541) );
  AOI22_X1 U12777 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11232) );
  AND2_X1 U12778 ( .A1(n10789), .A2(n10788), .ZN(n10791) );
  OAI21_X1 U12779 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18584), .A(
        n10248), .ZN(n10249) );
  NOR3_X1 U12780 ( .A1(n20012), .A2(n11308), .A3(n11325), .ZN(n11259) );
  NOR2_X1 U12781 ( .A1(n11626), .A2(n11627), .ZN(n11625) );
  INV_X1 U12782 ( .A(n14109), .ZN(n11863) );
  AND2_X1 U12783 ( .A1(n14083), .A2(n14067), .ZN(n11827) );
  INV_X1 U12784 ( .A(n13915), .ZN(n11764) );
  INV_X1 U12785 ( .A(n13584), .ZN(n11719) );
  INV_X1 U12786 ( .A(n11564), .ZN(n11562) );
  INV_X1 U12787 ( .A(n12367), .ZN(n11154) );
  INV_X1 U12788 ( .A(n10610), .ZN(n10623) );
  INV_X1 U12789 ( .A(n13334), .ZN(n10839) );
  OR2_X1 U12790 ( .A1(n12280), .A2(n18740), .ZN(n12389) );
  OR2_X1 U12791 ( .A1(n10910), .A2(n10909), .ZN(n12227) );
  NAND2_X1 U12792 ( .A1(n11474), .A2(n11473), .ZN(n11634) );
  AND2_X1 U12793 ( .A1(n12116), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12117) );
  INV_X1 U12794 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11808) );
  AND3_X1 U12795 ( .A1(n14535), .A2(n14537), .A3(n11605), .ZN(n11606) );
  NOR2_X1 U12796 ( .A1(n11150), .A2(n11143), .ZN(n12758) );
  INV_X1 U12797 ( .A(n11153), .ZN(n12276) );
  OR2_X1 U12798 ( .A1(n13064), .A2(n13063), .ZN(n13065) );
  NAND2_X1 U12799 ( .A1(n10642), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10644) );
  OR2_X1 U12800 ( .A1(n14777), .A2(n12280), .ZN(n12427) );
  AND3_X1 U12801 ( .A1(n11122), .A2(n11121), .A3(n11120), .ZN(n15633) );
  OR2_X1 U12802 ( .A1(n18760), .A2(n12336), .ZN(n15377) );
  NAND2_X1 U12803 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10184) );
  NAND2_X1 U12804 ( .A1(n17531), .A2(n17762), .ZN(n10216) );
  AND2_X1 U12805 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10205), .ZN(
        n10206) );
  OAI22_X1 U12806 ( .A1(n18584), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18442), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10255) );
  NOR2_X1 U12807 ( .A1(n11652), .A2(n11623), .ZN(n11655) );
  AND2_X1 U12808 ( .A1(n12689), .A2(n12688), .ZN(n14611) );
  AND2_X1 U12809 ( .A1(n12662), .A2(n12661), .ZN(n14380) );
  NAND2_X1 U12810 ( .A1(n14137), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13791) );
  NAND2_X1 U12811 ( .A1(n12117), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13788) );
  NOR2_X1 U12812 ( .A1(n11823), .A2(n11808), .ZN(n11829) );
  NAND2_X1 U12813 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11694) );
  NOR2_X2 U12814 ( .A1(n20044), .A2(n20700), .ZN(n11856) );
  AND2_X1 U12815 ( .A1(n15833), .A2(n11601), .ZN(n14540) );
  AND2_X1 U12816 ( .A1(n14661), .A2(n19985), .ZN(n14736) );
  NAND2_X1 U12817 ( .A1(n10028), .A2(n11445), .ZN(n11408) );
  NAND2_X1 U12818 ( .A1(n12562), .A2(n19751), .ZN(n10440) );
  NAND2_X1 U12819 ( .A1(n13945), .A2(n14822), .ZN(n14823) );
  AND2_X1 U12820 ( .A1(n12333), .A2(n12332), .ZN(n12335) );
  NOR2_X1 U12821 ( .A1(n16017), .A2(n18918), .ZN(n13177) );
  OR2_X1 U12822 ( .A1(n12898), .A2(n12897), .ZN(n18878) );
  NOR2_X1 U12823 ( .A1(n15972), .A2(n12280), .ZN(n12536) );
  INV_X1 U12824 ( .A(n15013), .ZN(n15014) );
  OR2_X1 U12825 ( .A1(n11116), .A2(n11115), .ZN(n14971) );
  INV_X1 U12826 ( .A(n15378), .ZN(n12334) );
  NAND2_X1 U12827 ( .A1(n16334), .A2(n16691), .ZN(n10433) );
  BUF_X1 U12828 ( .A(n10280), .Z(n15524) );
  NOR2_X1 U12829 ( .A1(n17108), .A2(n10204), .ZN(n10207) );
  INV_X1 U12830 ( .A(n17409), .ZN(n10222) );
  OAI211_X1 U12831 ( .C1(n10256), .C2(n10255), .A(n10257), .B(n10254), .ZN(
        n10359) );
  NOR2_X1 U12832 ( .A1(n12070), .A2(n15662), .ZN(n12071) );
  INV_X1 U12833 ( .A(n12026), .ZN(n12027) );
  NAND2_X1 U12834 ( .A1(n11847), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11865) );
  INV_X1 U12835 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13921) );
  INV_X1 U12836 ( .A(n19790), .ZN(n19793) );
  NAND2_X1 U12837 ( .A1(n11472), .A2(n11471), .ZN(n20159) );
  NAND2_X1 U12838 ( .A1(n13796), .A2(n13800), .ZN(n15685) );
  AND2_X1 U12839 ( .A1(n12676), .A2(n12675), .ZN(n14359) );
  OR2_X1 U12840 ( .A1(n13422), .A2(n12601), .ZN(n13411) );
  NOR2_X1 U12841 ( .A1(n11967), .A2(n15715), .ZN(n11968) );
  NOR2_X1 U12842 ( .A1(n11765), .A2(n13921), .ZN(n11782) );
  NAND2_X1 U12843 ( .A1(n20040), .A2(n20025), .ZN(n11623) );
  AND2_X1 U12844 ( .A1(n14631), .A2(n12731), .ZN(n14610) );
  AND2_X1 U12845 ( .A1(n14700), .A2(n11604), .ZN(n14537) );
  OR2_X1 U12846 ( .A1(n14539), .A2(n14711), .ZN(n14700) );
  AND2_X1 U12847 ( .A1(n12646), .A2(n12645), .ZN(n15780) );
  INV_X1 U12848 ( .A(n14736), .ZN(n19970) );
  AND2_X1 U12849 ( .A1(n12723), .A2(n12716), .ZN(n19991) );
  INV_X1 U12850 ( .A(n20377), .ZN(n20519) );
  NAND2_X1 U12851 ( .A1(n20700), .A2(n20780), .ZN(n20377) );
  AND2_X1 U12852 ( .A1(n10800), .A2(n12438), .ZN(n13633) );
  INV_X1 U12853 ( .A(n13214), .ZN(n13215) );
  OR2_X1 U12854 ( .A1(n12883), .A2(n13548), .ZN(n13538) );
  AND4_X1 U12855 ( .A1(n10931), .A2(n10930), .A3(n10929), .A4(n10928), .ZN(
        n13775) );
  AND2_X1 U12856 ( .A1(n10753), .A2(n10752), .ZN(n14787) );
  INV_X1 U12857 ( .A(n12164), .ZN(n12165) );
  INV_X1 U12858 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12846) );
  AND2_X1 U12859 ( .A1(n13974), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15110) );
  INV_X1 U12860 ( .A(n18839), .ZN(n18772) );
  INV_X1 U12861 ( .A(n13185), .ZN(n13660) );
  INV_X1 U12862 ( .A(n19451), .ZN(n19446) );
  INV_X1 U12863 ( .A(n12253), .ZN(n19319) );
  OR2_X1 U12864 ( .A1(n19177), .A2(n19712), .ZN(n19384) );
  INV_X1 U12865 ( .A(n19696), .ZN(n19503) );
  OR3_X1 U12866 ( .A1(n12233), .A2(n19600), .A3(n19549), .ZN(n19555) );
  NOR2_X1 U12867 ( .A1(n17975), .A2(n10348), .ZN(n12505) );
  OAI211_X1 U12868 ( .C1(n10435), .C2(n10434), .A(n10433), .B(n10432), .ZN(
        n10436) );
  INV_X1 U12869 ( .A(n16650), .ZN(n16571) );
  INV_X1 U12870 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16632) );
  NAND2_X1 U12871 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16802), .ZN(n16773) );
  AOI221_X1 U12872 ( .B1(n15460), .B2(n15459), .C1(n15458), .C2(n15459), .A(
        n18459), .ZN(n15627) );
  AND2_X1 U12873 ( .A1(n17328), .A2(n17259), .ZN(n17261) );
  NOR2_X1 U12874 ( .A1(n17649), .A2(n17290), .ZN(n17638) );
  AND2_X1 U12875 ( .A1(n17430), .A2(n10402), .ZN(n17670) );
  INV_X1 U12876 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17477) );
  NAND2_X1 U12877 ( .A1(n10400), .A2(n17522), .ZN(n17493) );
  INV_X1 U12878 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12521) );
  NOR2_X1 U12879 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17531), .ZN(
        n17393) );
  NOR2_X1 U12880 ( .A1(n12518), .A2(n17818), .ZN(n17691) );
  OR2_X1 U12881 ( .A1(n18593), .A2(n18468), .ZN(n17966) );
  NOR2_X1 U12882 ( .A1(n12509), .A2(n12508), .ZN(n14131) );
  INV_X1 U12883 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18423) );
  NAND2_X1 U12884 ( .A1(n11664), .A2(n11663), .ZN(n14252) );
  NAND2_X1 U12885 ( .A1(n12071), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12115) );
  NAND2_X1 U12886 ( .A1(n11935), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11967) );
  AND2_X1 U12887 ( .A1(n15659), .A2(n13793), .ZN(n19802) );
  INV_X1 U12888 ( .A(n15685), .ZN(n19831) );
  INV_X1 U12889 ( .A(n14394), .ZN(n19850) );
  INV_X1 U12890 ( .A(n19927), .ZN(n19922) );
  INV_X1 U12891 ( .A(n19888), .ZN(n19925) );
  NAND2_X1 U12892 ( .A1(n11912), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U12893 ( .A1(n11866), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11911) );
  NAND2_X1 U12894 ( .A1(n11783), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11823) );
  OR2_X1 U12895 ( .A1(n11726), .A2(n11729), .ZN(n11748) );
  NAND2_X1 U12896 ( .A1(n11712), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11711) );
  INV_X1 U12897 ( .A(n15823), .ZN(n19939) );
  AND2_X1 U12898 ( .A1(n14538), .A2(n14537), .ZN(n14549) );
  NOR2_X1 U12899 ( .A1(n19961), .A2(n14041), .ZN(n15937) );
  INV_X1 U12900 ( .A(n19996), .ZN(n19957) );
  INV_X1 U12901 ( .A(n19992), .ZN(n19968) );
  AND2_X1 U12902 ( .A1(n12723), .A2(n13506), .ZN(n20001) );
  INV_X1 U12903 ( .A(n15599), .ZN(n14753) );
  OAI22_X1 U12904 ( .A1(n20021), .A2(n20020), .B1(n20352), .B2(n20160), .ZN(
        n20052) );
  OAI21_X1 U12905 ( .B1(n20181), .B2(n20165), .A(n20478), .ZN(n20183) );
  INV_X1 U12906 ( .A(n20203), .ZN(n20210) );
  INV_X1 U12907 ( .A(n20214), .ZN(n20262) );
  INV_X1 U12908 ( .A(n11681), .ZN(n20259) );
  INV_X1 U12909 ( .A(n20282), .ZN(n20313) );
  INV_X1 U12910 ( .A(n20404), .ZN(n20289) );
  AND2_X1 U12911 ( .A1(n20665), .A2(n10084), .ZN(n20370) );
  AND2_X1 U12912 ( .A1(n20665), .A2(n20383), .ZN(n20437) );
  NOR2_X2 U12913 ( .A1(n20443), .A2(n20404), .ZN(n20465) );
  INV_X1 U12914 ( .A(n20480), .ZN(n20512) );
  AND2_X1 U12915 ( .A1(n20025), .A2(n20049), .ZN(n20534) );
  AND2_X1 U12916 ( .A1(n20036), .A2(n20049), .ZN(n20552) );
  NOR2_X2 U12917 ( .A1(n20443), .A2(n20011), .ZN(n20575) );
  NAND2_X1 U12918 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n14252), .ZN(n15599) );
  INV_X1 U12919 ( .A(n20708), .ZN(n15619) );
  INV_X1 U12920 ( .A(n20646), .ZN(n20649) );
  AND2_X1 U12921 ( .A1(n13633), .A2(n13460), .ZN(n13222) );
  OR2_X1 U12922 ( .A1(n18643), .A2(n11172), .ZN(n18774) );
  INV_X1 U12923 ( .A(n18852), .ZN(n18865) );
  INV_X1 U12924 ( .A(n18774), .ZN(n18867) );
  OR2_X1 U12925 ( .A1(n11075), .A2(n11074), .ZN(n13813) );
  AND2_X1 U12926 ( .A1(n13179), .A2(n13178), .ZN(n13182) );
  AND2_X1 U12927 ( .A1(n18926), .A2(n10839), .ZN(n16024) );
  INV_X1 U12928 ( .A(n13269), .ZN(n18970) );
  INV_X2 U12929 ( .A(n13317), .ZN(n18974) );
  OAI21_X1 U12930 ( .B1(n15151), .B2(n18980), .A(n12494), .ZN(n12495) );
  AND2_X1 U12931 ( .A1(n16041), .A2(n16113), .ZN(n16042) );
  AND2_X1 U12932 ( .A1(n13906), .A2(n13905), .ZN(n16084) );
  AND2_X1 U12933 ( .A1(n16117), .A2(n13305), .ZN(n16108) );
  NAND2_X1 U12934 ( .A1(n12161), .A2(n12160), .ZN(n12162) );
  INV_X1 U12935 ( .A(n19017), .ZN(n18822) );
  AND2_X1 U12936 ( .A1(n13823), .A2(n13822), .ZN(n18742) );
  AND2_X1 U12937 ( .A1(n19693), .A2(n11170), .ZN(n18839) );
  INV_X1 U12938 ( .A(n16146), .ZN(n18993) );
  XNOR2_X1 U12939 ( .A(n13391), .B(n13393), .ZN(n19177) );
  OAI21_X1 U12940 ( .B1(n19036), .B2(n19035), .A(n19034), .ZN(n19078) );
  NOR2_X2 U12941 ( .A1(n19327), .A2(n19232), .ZN(n19105) );
  INV_X1 U12942 ( .A(n19327), .ZN(n19321) );
  NOR2_X2 U12943 ( .A1(n19232), .A2(n19384), .ZN(n19166) );
  AND2_X1 U12944 ( .A1(n19258), .A2(n19375), .ZN(n19178) );
  OAI21_X1 U12945 ( .B1(n19209), .B2(n19208), .A(n19207), .ZN(n19225) );
  OAI21_X1 U12946 ( .B1(n19234), .B2(n19416), .A(n19231), .ZN(n19253) );
  NAND2_X1 U12947 ( .A1(n19295), .A2(n19294), .ZN(n19311) );
  NOR2_X2 U12948 ( .A1(n19504), .A2(n19327), .ZN(n19342) );
  OAI21_X1 U12949 ( .B1(n19354), .B2(n19369), .A(n19554), .ZN(n19371) );
  INV_X1 U12950 ( .A(n19384), .ZN(n19375) );
  NOR2_X1 U12951 ( .A1(n19504), .A2(n19451), .ZN(n19439) );
  INV_X1 U12952 ( .A(n19599), .ZN(n19538) );
  AND2_X1 U12953 ( .A1(n19554), .A2(n19030), .ZN(n19553) );
  INV_X1 U12954 ( .A(n19474), .ZN(n19582) );
  INV_X1 U12955 ( .A(n19493), .ZN(n19601) );
  INV_X1 U12956 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19549) );
  INV_X1 U12957 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19634) );
  NAND2_X1 U12958 ( .A1(n17968), .A2(n18619), .ZN(n10349) );
  NAND2_X1 U12959 ( .A1(n12516), .A2(n12507), .ZN(n18405) );
  NOR2_X1 U12960 ( .A1(n18541), .A2(n16377), .ZN(n16362) );
  OR3_X1 U12961 ( .A1(n16676), .A2(n16398), .A3(n18539), .ZN(n16385) );
  NOR2_X1 U12962 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16441), .ZN(n16433) );
  OR2_X1 U12963 ( .A1(n16458), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n16441) );
  NOR2_X1 U12964 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16517), .ZN(n16498) );
  NOR2_X1 U12965 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16537), .ZN(n16521) );
  INV_X1 U12966 ( .A(n18467), .ZN(n16650) );
  NOR2_X2 U12967 ( .A1(n18452), .A2(n10429), .ZN(n16646) );
  INV_X1 U12968 ( .A(n16814), .ZN(n16790) );
  NOR2_X1 U12969 ( .A1(n16495), .A2(n16868), .ZN(n16843) );
  NAND3_X1 U12970 ( .A1(n15627), .A2(n18619), .A3(n17138), .ZN(n16978) );
  NOR2_X1 U12971 ( .A1(n17160), .A2(n17054), .ZN(n17048) );
  INV_X1 U12972 ( .A(n17968), .ZN(n17138) );
  NAND2_X1 U12973 ( .A1(n18617), .A2(n18403), .ZN(n17200) );
  INV_X1 U12974 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20869) );
  NAND3_X1 U12975 ( .A1(n10181), .A2(n10180), .A3(n10179), .ZN(n17103) );
  NOR2_X2 U12976 ( .A1(n18577), .A2(n17551), .ZN(n17475) );
  INV_X1 U12977 ( .A(n18043), .ZN(n18254) );
  NOR2_X1 U12978 ( .A1(n17940), .A2(n17934), .ZN(n17896) );
  NOR2_X1 U12979 ( .A1(n17801), .A2(n17951), .ZN(n17947) );
  NOR2_X1 U12980 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18566), .ZN(
        n18593) );
  INV_X1 U12981 ( .A(n18102), .ZN(n18104) );
  INV_X1 U12982 ( .A(n18132), .ZN(n18125) );
  INV_X1 U12983 ( .A(n18150), .ZN(n18153) );
  INV_X1 U12984 ( .A(n18367), .ZN(n18314) );
  INV_X1 U12985 ( .A(n18380), .ZN(n18390) );
  INV_X1 U12986 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18622) );
  INV_X1 U12987 ( .A(U212), .ZN(n16260) );
  NAND2_X1 U12988 ( .A1(n14252), .A2(n13238), .ZN(n13695) );
  INV_X1 U12989 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20771) );
  INV_X1 U12990 ( .A(n19838), .ZN(n19813) );
  INV_X1 U12991 ( .A(n19833), .ZN(n15773) );
  INV_X1 U12992 ( .A(n19802), .ZN(n15779) );
  OR2_X1 U12993 ( .A1(n12149), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19964) );
  NAND2_X1 U12994 ( .A1(n19854), .A2(n11310), .ZN(n14394) );
  NAND2_X1 U12995 ( .A1(n19854), .A2(n14166), .ZN(n14383) );
  OR2_X1 U12996 ( .A1(n14123), .A2(n20005), .ZN(n15809) );
  INV_X1 U12997 ( .A(n15847), .ZN(n15778) );
  INV_X1 U12998 ( .A(n15801), .ZN(n14437) );
  NAND2_X1 U12999 ( .A1(n19855), .A2(n13399), .ZN(n13692) );
  INV_X1 U13000 ( .A(n19855), .ZN(n19886) );
  OR2_X1 U13001 ( .A1(n19920), .A2(n20025), .ZN(n19888) );
  OR3_X1 U13002 ( .A1(n13695), .A2(n12599), .A3(n15619), .ZN(n19927) );
  OR2_X1 U13003 ( .A1(n19935), .A2(n12146), .ZN(n15823) );
  INV_X1 U13004 ( .A(n15849), .ZN(n19942) );
  OR2_X1 U13005 ( .A1(n12598), .A2(n12597), .ZN(n19996) );
  INV_X1 U13006 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20446) );
  NAND2_X1 U13007 ( .A1(n20118), .A2(n20289), .ZN(n20084) );
  NAND2_X1 U13008 ( .A1(n20118), .A2(n10084), .ZN(n20117) );
  NAND2_X1 U13009 ( .A1(n20118), .A2(n20469), .ZN(n20152) );
  NAND2_X1 U13010 ( .A1(n20118), .A2(n20383), .ZN(n20186) );
  NAND2_X1 U13011 ( .A1(n20262), .A2(n20289), .ZN(n20203) );
  NAND2_X1 U13012 ( .A1(n20262), .A2(n10084), .ZN(n20253) );
  NAND2_X1 U13013 ( .A1(n20664), .A2(n11681), .ZN(n20288) );
  NAND2_X1 U13014 ( .A1(n20665), .A2(n20289), .ZN(n20343) );
  NAND2_X1 U13015 ( .A1(n20665), .A2(n20469), .ZN(n20403) );
  AOI22_X1 U13016 ( .A1(n20412), .A2(n20409), .B1(n20408), .B2(n20414), .ZN(
        n20442) );
  NAND2_X1 U13017 ( .A1(n20470), .A2(n10084), .ZN(n20480) );
  NAND2_X1 U13018 ( .A1(n20470), .A2(n20469), .ZN(n20579) );
  INV_X2 U13019 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20700) );
  INV_X1 U13020 ( .A(n20663), .ZN(n20659) );
  INV_X1 U13021 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20598) );
  INV_X1 U13022 ( .A(n20715), .ZN(n20712) );
  INV_X1 U13023 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19622) );
  OR3_X1 U13024 ( .A1(n12784), .A2(n19028), .A3(n16167), .ZN(n13230) );
  AND2_X1 U13025 ( .A1(n11180), .A2(n10092), .ZN(n11181) );
  NAND2_X1 U13026 ( .A1(n18643), .A2(n10802), .ZN(n18870) );
  OR2_X1 U13027 ( .A1(n18867), .A2(n19700), .ZN(n18832) );
  INV_X1 U13028 ( .A(n18827), .ZN(n18877) );
  INV_X1 U13029 ( .A(n16084), .ZN(n18889) );
  INV_X2 U13030 ( .A(n18903), .ZN(n18888) );
  AND2_X2 U13031 ( .A1(n13187), .A2(n13460), .ZN(n18903) );
  OR2_X1 U13032 ( .A1(n13181), .A2(n13272), .ZN(n14918) );
  NOR2_X1 U13033 ( .A1(n16024), .A2(n18912), .ZN(n18936) );
  NAND2_X1 U13034 ( .A1(n13335), .A2(n13334), .ZN(n18928) );
  OR2_X1 U13035 ( .A1(n18969), .A2(n13321), .ZN(n20720) );
  NAND2_X1 U13036 ( .A1(n13320), .A2(n19752), .ZN(n18969) );
  OR2_X1 U13037 ( .A1(n13233), .A2(n13231), .ZN(n13317) );
  INV_X1 U13038 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18736) );
  INV_X1 U13039 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16079) );
  INV_X1 U13040 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18794) );
  INV_X1 U13041 ( .A(n16112), .ZN(n18981) );
  INV_X1 U13042 ( .A(n18992), .ZN(n16147) );
  INV_X1 U13043 ( .A(n15562), .ZN(n15559) );
  AOI21_X1 U13044 ( .B1(n19031), .B2(n19035), .A(n19024), .ZN(n19082) );
  NAND2_X1 U13045 ( .A1(n19321), .A2(n19258), .ZN(n19140) );
  AOI21_X1 U13046 ( .B1(n19145), .B2(n19149), .A(n19144), .ZN(n19170) );
  INV_X1 U13047 ( .A(n19178), .ZN(n19201) );
  INV_X1 U13048 ( .A(n19249), .ZN(n19257) );
  NAND2_X1 U13049 ( .A1(n19696), .A2(n19258), .ZN(n19315) );
  INV_X1 U13050 ( .A(n19350), .ZN(n19374) );
  NAND2_X1 U13051 ( .A1(n19376), .A2(n19375), .ZN(n19438) );
  INV_X1 U13052 ( .A(n19439), .ZN(n19500) );
  AOI211_X2 U13053 ( .C1(n19511), .C2(n19513), .A(n19509), .B(n19508), .ZN(
        n19547) );
  NAND2_X1 U13054 ( .A1(n19376), .A2(n19696), .ZN(n19609) );
  NAND2_X1 U13055 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19622), .ZN(n19758) );
  INV_X1 U13056 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16309) );
  INV_X1 U13057 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17463) );
  INV_X1 U13058 ( .A(n10431), .ZN(n16674) );
  NAND2_X1 U13059 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16737), .ZN(n16728) );
  AND2_X1 U13060 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16790), .ZN(n16802) );
  INV_X1 U13061 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16953) );
  INV_X1 U13062 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16964) );
  INV_X1 U13063 ( .A(n16978), .ZN(n16985) );
  INV_X1 U13064 ( .A(n17065), .ZN(n17058) );
  NOR2_X1 U13065 ( .A1(n10113), .A2(n10112), .ZN(n17108) );
  NOR2_X1 U13066 ( .A1(n10124), .A2(n10123), .ZN(n17115) );
  INV_X1 U13067 ( .A(n17132), .ZN(n17125) );
  NAND2_X1 U13068 ( .A1(n17139), .A2(n17138), .ZN(n17165) );
  NAND2_X1 U13069 ( .A1(n17198), .A2(n17137), .ZN(n17196) );
  INV_X1 U13070 ( .A(n17247), .ZN(n17242) );
  AND2_X1 U13071 ( .A1(n10405), .A2(n10404), .ZN(n10406) );
  INV_X1 U13072 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17809) );
  INV_X1 U13073 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17608) );
  INV_X1 U13074 ( .A(n17934), .ZN(n17951) );
  INV_X1 U13075 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17847) );
  INV_X1 U13076 ( .A(n17947), .ZN(n17930) );
  INV_X1 U13077 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18442) );
  INV_X1 U13078 ( .A(n18599), .ZN(n18596) );
  INV_X1 U13079 ( .A(n18617), .ZN(n18459) );
  INV_X1 U13080 ( .A(n17457), .ZN(n18472) );
  NOR2_X1 U13081 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13208), .ZN(n16296)
         );
  INV_X1 U13082 ( .A(n16251), .ZN(n16263) );
  NAND2_X1 U13083 ( .A1(n11182), .A2(n11181), .ZN(P2_U2825) );
  OR4_X1 U13084 ( .A1(n13221), .A2(n13220), .A3(n13219), .A4(n13218), .ZN(
        P2_U2832) );
  OAI21_X1 U13085 ( .B1(n16208), .B2(n17470), .A(n10406), .ZN(P3_U2799) );
  AOI22_X1 U13086 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U13087 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U13088 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9608), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U13089 ( .A1(n16921), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10098) );
  NAND4_X1 U13090 ( .A1(n10101), .A2(n10100), .A3(n10099), .A4(n10098), .ZN(
        n10113) );
  AOI22_X1 U13091 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U13092 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10110) );
  NOR2_X2 U13093 ( .A1(n10104), .A2(n16663), .ZN(n10311) );
  AOI22_X1 U13094 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U13095 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9600), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10108) );
  NAND4_X1 U13096 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10112) );
  AOI22_X1 U13097 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U13098 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U13099 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(n9609), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U13100 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10115) );
  NAND4_X1 U13101 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10124) );
  AOI22_X1 U13102 ( .A1(n16819), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U13103 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10121) );
  AOI22_X1 U13104 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10120) );
  INV_X2 U13105 ( .A(n16705), .ZN(n16754) );
  AOI22_X1 U13106 ( .A1(n16939), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10119) );
  NAND4_X1 U13107 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10123) );
  AOI22_X1 U13108 ( .A1(n16819), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U13109 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U13110 ( .A1(n10150), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10270), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U13111 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10125) );
  NAND4_X1 U13112 ( .A1(n10128), .A2(n10127), .A3(n10126), .A4(n10125), .ZN(
        n10134) );
  AOI22_X1 U13113 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9608), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U13114 ( .A1(n16931), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U13115 ( .A1(n16939), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U13116 ( .A1(n10280), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10129) );
  NAND4_X1 U13117 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .ZN(
        n10133) );
  AOI22_X1 U13118 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10299), .B1(
        n10136), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10142) );
  AOI22_X1 U13119 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10137), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U13120 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9608), .ZN(n10140) );
  AOI22_X1 U13121 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n9609), .B1(
        n10270), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U13122 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10143), .B1(
        n16931), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U13123 ( .A1(n10280), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n16754), .ZN(n10147) );
  AOI22_X1 U13124 ( .A1(n10150), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10311), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U13125 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n10144), .ZN(n10145) );
  AOI22_X1 U13126 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13127 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10159) );
  INV_X1 U13128 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U13129 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10151) );
  OAI21_X1 U13130 ( .B1(n16622), .B2(n16970), .A(n10151), .ZN(n10157) );
  AOI22_X1 U13131 ( .A1(n16819), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9604), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U13132 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9608), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10154) );
  INV_X1 U13133 ( .A(n10094), .ZN(n16931) );
  AOI22_X1 U13134 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U13135 ( .A1(n16754), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10152) );
  NAND4_X1 U13136 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10156) );
  AOI211_X1 U13137 ( .C1(n16932), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n10157), .B(n10156), .ZN(n10158) );
  NAND3_X1 U13138 ( .A1(n10160), .A2(n10159), .A3(n10158), .ZN(n10196) );
  NAND2_X1 U13139 ( .A1(n10197), .A2(n10196), .ZN(n10199) );
  AOI22_X1 U13140 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13141 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U13142 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10161) );
  OAI21_X1 U13143 ( .B1(n16622), .B2(n16964), .A(n10161), .ZN(n10167) );
  AOI22_X1 U13144 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U13145 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U13146 ( .A1(n16819), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U13147 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10162) );
  NAND4_X1 U13148 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10166) );
  AOI211_X1 U13149 ( .C1(n16932), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n10167), .B(n10166), .ZN(n10168) );
  NAND3_X1 U13150 ( .A1(n10170), .A2(n10169), .A3(n10168), .ZN(n10202) );
  NAND2_X1 U13151 ( .A1(n10203), .A2(n10202), .ZN(n10204) );
  AOI22_X1 U13152 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10181) );
  BUF_X2 U13153 ( .A(n16938), .Z(n16919) );
  AOI22_X1 U13154 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13155 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9609), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10172) );
  OAI21_X1 U13156 ( .B1(n16622), .B2(n16953), .A(n10172), .ZN(n10178) );
  AOI22_X1 U13157 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U13158 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13159 ( .A1(n16819), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U13160 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10173) );
  NAND4_X1 U13161 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  AOI211_X1 U13162 ( .C1(n15537), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n10178), .B(n10177), .ZN(n10179) );
  INV_X1 U13163 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18575) );
  AOI22_X1 U13164 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17428), .B1(
        n17531), .B2(n18575), .ZN(n10234) );
  INV_X1 U13165 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17659) );
  INV_X1 U13166 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n20816) );
  AOI22_X1 U13167 ( .A1(n10270), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10182) );
  OAI21_X1 U13168 ( .B1(n10240), .B2(n20816), .A(n10182), .ZN(n10183) );
  INV_X1 U13169 ( .A(n10183), .ZN(n10187) );
  AOI22_X1 U13170 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U13171 ( .A1(n10280), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13172 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10150), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U13173 ( .A1(n16938), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13174 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13175 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10189) );
  NAND2_X1 U13176 ( .A1(n17620), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17619) );
  NOR2_X1 U13177 ( .A1(n17613), .A2(n17619), .ZN(n17612) );
  INV_X1 U13178 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18576) );
  NOR2_X1 U13179 ( .A1(n17131), .A2(n18576), .ZN(n10193) );
  NOR2_X1 U13180 ( .A1(n17612), .A2(n10193), .ZN(n17600) );
  INV_X1 U13181 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17913) );
  XNOR2_X1 U13182 ( .A(n17913), .B(n10194), .ZN(n17599) );
  NOR2_X1 U13183 ( .A1(n17600), .A2(n17599), .ZN(n17598) );
  NOR2_X1 U13184 ( .A1(n17913), .A2(n10194), .ZN(n10195) );
  INV_X1 U13185 ( .A(n10196), .ZN(n17118) );
  XOR2_X1 U13186 ( .A(n17118), .B(n10197), .Z(n17592) );
  NOR2_X1 U13187 ( .A1(n17591), .A2(n17592), .ZN(n10198) );
  NAND2_X1 U13188 ( .A1(n17591), .A2(n17592), .ZN(n17590) );
  XOR2_X1 U13189 ( .A(n17115), .B(n10199), .Z(n10200) );
  XNOR2_X1 U13190 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n10200), .ZN(
        n17580) );
  NOR2_X1 U13191 ( .A1(n17579), .A2(n17580), .ZN(n17578) );
  NOR2_X2 U13192 ( .A1(n17578), .A2(n10201), .ZN(n17564) );
  INV_X1 U13193 ( .A(n10202), .ZN(n17111) );
  XOR2_X1 U13194 ( .A(n17111), .B(n10203), .Z(n17565) );
  XOR2_X1 U13195 ( .A(n17108), .B(n10204), .Z(n10205) );
  XNOR2_X1 U13196 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n10205), .ZN(
        n17552) );
  OAI21_X1 U13197 ( .B1(n10207), .B2(n17103), .A(n17428), .ZN(n10208) );
  NOR2_X1 U13198 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  XNOR2_X1 U13199 ( .A(n10209), .B(n10208), .ZN(n17537) );
  INV_X1 U13200 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17542) );
  NOR2_X1 U13201 ( .A1(n17537), .A2(n17542), .ZN(n17536) );
  INV_X1 U13202 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17859) );
  NOR2_X1 U13203 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17502), .ZN(
        n10211) );
  INV_X1 U13204 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17485) );
  NAND2_X1 U13205 ( .A1(n10211), .A2(n17485), .ZN(n17471) );
  NOR3_X1 U13206 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10212) );
  AND2_X2 U13207 ( .A1(n17818), .A2(n10213), .ZN(n17864) );
  NAND2_X1 U13208 ( .A1(n17531), .A2(n17864), .ZN(n17530) );
  NAND2_X1 U13209 ( .A1(n10213), .A2(n17530), .ZN(n17448) );
  INV_X1 U13210 ( .A(n17448), .ZN(n10215) );
  INV_X1 U13211 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20872) );
  INV_X1 U13212 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17841) );
  NOR2_X1 U13213 ( .A1(n17847), .A2(n17841), .ZN(n17827) );
  NAND2_X1 U13214 ( .A1(n17827), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17798) );
  NOR2_X1 U13215 ( .A1(n17798), .A2(n17809), .ZN(n17780) );
  NAND2_X1 U13216 ( .A1(n17780), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17765) );
  NOR2_X1 U13217 ( .A1(n20872), .A2(n17765), .ZN(n17757) );
  NAND2_X1 U13218 ( .A1(n17757), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12518) );
  INV_X1 U13219 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17762) );
  NAND2_X1 U13220 ( .A1(n10217), .A2(n10216), .ZN(n10218) );
  INV_X1 U13221 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17747) );
  NAND2_X2 U13222 ( .A1(n17404), .A2(n17747), .ZN(n17403) );
  INV_X1 U13223 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20785) );
  NOR2_X1 U13224 ( .A1(n17762), .A2(n17747), .ZN(n17738) );
  INV_X1 U13225 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17351) );
  NAND2_X1 U13226 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17358) );
  NOR2_X1 U13227 ( .A1(n17351), .A2(n17358), .ZN(n17689) );
  NAND2_X1 U13228 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17689), .ZN(
        n17341) );
  INV_X1 U13229 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17700) );
  NOR2_X1 U13230 ( .A1(n17341), .A2(n17700), .ZN(n15563) );
  NAND2_X1 U13231 ( .A1(n17738), .A2(n15563), .ZN(n17300) );
  NOR2_X1 U13232 ( .A1(n20785), .A2(n17300), .ZN(n10402) );
  INV_X1 U13233 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17730) );
  NAND2_X1 U13234 ( .A1(n17393), .A2(n17730), .ZN(n10219) );
  NOR2_X1 U13235 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n10219), .ZN(
        n17350) );
  NAND2_X1 U13236 ( .A1(n17350), .A2(n17351), .ZN(n17340) );
  NAND2_X1 U13237 ( .A1(n17738), .A2(n10222), .ZN(n17349) );
  NAND2_X2 U13238 ( .A1(n17362), .A2(n17349), .ZN(n17394) );
  NAND2_X1 U13239 ( .A1(n15563), .A2(n17394), .ZN(n17318) );
  NOR3_X2 U13240 ( .A1(n17308), .A2(n17318), .A3(n20785), .ZN(n10224) );
  NAND2_X1 U13241 ( .A1(n17428), .A2(n17304), .ZN(n10223) );
  OAI221_X1 U13242 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17428), 
        .C1(n17659), .C2(n10224), .A(n10223), .ZN(n17280) );
  NOR2_X1 U13243 ( .A1(n17280), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17279) );
  NOR2_X1 U13244 ( .A1(n10224), .A2(n17428), .ZN(n17303) );
  NAND2_X1 U13245 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12504) );
  AND2_X1 U13246 ( .A1(n17531), .A2(n12504), .ZN(n10225) );
  AND2_X1 U13247 ( .A1(n10227), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17270) );
  NAND2_X1 U13248 ( .A1(n17531), .A2(n17270), .ZN(n12499) );
  NOR2_X1 U13249 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17428), .ZN(
        n12525) );
  AOI21_X2 U13250 ( .B1(n12499), .B2(n10228), .A(n12525), .ZN(n15573) );
  NAND2_X1 U13251 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15573), .ZN(
        n15572) );
  INV_X1 U13252 ( .A(n10230), .ZN(n10229) );
  NAND2_X1 U13253 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15612), .ZN(
        n15611) );
  NAND2_X1 U13254 ( .A1(n10230), .A2(n15611), .ZN(n10233) );
  INV_X1 U13255 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16177) );
  OAI211_X1 U13256 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16177), .A(
        n10230), .B(n15572), .ZN(n10231) );
  NAND2_X1 U13257 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16177), .ZN(
        n16200) );
  NAND3_X1 U13258 ( .A1(n10234), .A2(n10231), .A3(n16200), .ZN(n10232) );
  OAI21_X1 U13259 ( .B1(n10234), .B2(n10233), .A(n10232), .ZN(n16208) );
  AOI22_X1 U13260 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U13261 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13262 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13263 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10236) );
  NAND4_X1 U13264 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10246) );
  AOI22_X1 U13265 ( .A1(n16939), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U13266 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15537), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13267 ( .A1(n16921), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n16940), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U13268 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10241) );
  NAND4_X1 U13269 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10245) );
  INV_X1 U13270 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18577) );
  NAND2_X1 U13271 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18577), .ZN(n17621) );
  AOI22_X1 U13272 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18423), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18592), .ZN(n10354) );
  NAND2_X1 U13273 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10249), .ZN(
        n10251) );
  OAI22_X1 U13274 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10249), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20778), .ZN(n10253) );
  AOI21_X1 U13275 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n10251), .A(
        n10253), .ZN(n10250) );
  NOR2_X1 U13276 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20778), .ZN(
        n10252) );
  AOI22_X1 U13277 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n10253), .B1(
        n10252), .B2(n10251), .ZN(n10257) );
  NAND2_X1 U13278 ( .A1(n10256), .A2(n10255), .ZN(n10254) );
  AOI21_X1 U13279 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n18598), .A(
        n10355), .ZN(n10353) );
  NAND3_X1 U13280 ( .A1(n10354), .A2(n10257), .A3(n10353), .ZN(n10258) );
  NAND3_X1 U13281 ( .A1(n10356), .A2(n10359), .A3(n10258), .ZN(n15458) );
  AOI22_X1 U13282 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U13283 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U13284 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9609), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13285 ( .A1(n16921), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10259) );
  NAND4_X1 U13286 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10268) );
  AOI22_X1 U13287 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13288 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U13289 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16940), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U13290 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10263) );
  NAND4_X1 U13291 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(n10263), .ZN(
        n10267) );
  NAND2_X1 U13292 ( .A1(n17971), .A2(n17138), .ZN(n10333) );
  NAND2_X1 U13293 ( .A1(n10349), .A2(n10333), .ZN(n18633) );
  AOI22_X1 U13294 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U13295 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13296 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10269) );
  OAI21_X1 U13297 ( .B1(n10235), .B2(n16976), .A(n10269), .ZN(n10276) );
  AOI22_X1 U13298 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U13299 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U13300 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16940), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13301 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10271) );
  NAND4_X1 U13302 ( .A1(n10274), .A2(n10273), .A3(n10272), .A4(n10271), .ZN(
        n10275) );
  AOI211_X1 U13303 ( .C1(n16932), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n10276), .B(n10275), .ZN(n10277) );
  NAND3_X1 U13304 ( .A1(n10279), .A2(n10278), .A3(n10277), .ZN(n10345) );
  AOI22_X1 U13305 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13306 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13307 ( .A1(n10311), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10281) );
  OAI21_X1 U13308 ( .B1(n10235), .B2(n16953), .A(n10281), .ZN(n10286) );
  AOI22_X1 U13309 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10150), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U13310 ( .A1(n16940), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13311 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13312 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13313 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13314 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16940), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13315 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10289) );
  OAI21_X1 U13316 ( .B1(n10235), .B2(n16970), .A(n10289), .ZN(n10295) );
  AOI22_X1 U13317 ( .A1(n16921), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13318 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13319 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U13320 ( .A1(n10188), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10290) );
  NAND4_X1 U13321 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n10294) );
  AOI211_X1 U13322 ( .C1(n16903), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n10295), .B(n10294), .ZN(n10296) );
  NAND3_X1 U13323 ( .A1(n10298), .A2(n10297), .A3(n10296), .ZN(n10344) );
  INV_X1 U13324 ( .A(n10347), .ZN(n10331) );
  AOI22_X1 U13325 ( .A1(n16940), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13326 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9600), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13327 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U13328 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10300) );
  NAND4_X1 U13329 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n10309) );
  AOI22_X1 U13330 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13331 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13332 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13333 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16920), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10304) );
  NAND4_X1 U13334 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10308) );
  AOI22_X1 U13335 ( .A1(n16921), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13336 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15537), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10319) );
  INV_X1 U13337 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16959) );
  AOI22_X1 U13338 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10310) );
  OAI21_X1 U13339 ( .B1(n10235), .B2(n16959), .A(n10310), .ZN(n10317) );
  AOI22_X1 U13340 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U13341 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13342 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16919), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U13343 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n9609), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10312) );
  NAND4_X1 U13344 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10316) );
  AOI211_X1 U13345 ( .C1(n16939), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n10317), .B(n10316), .ZN(n10318) );
  NAND3_X1 U13346 ( .A1(n10320), .A2(n10319), .A3(n10318), .ZN(n10332) );
  NOR2_X1 U13347 ( .A1(n17983), .A2(n10332), .ZN(n10351) );
  AOI22_X1 U13348 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16919), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13349 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13350 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10321) );
  OAI21_X1 U13351 ( .B1(n10235), .B2(n16964), .A(n10321), .ZN(n10327) );
  AOI22_X1 U13352 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10188), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13353 ( .A1(n10150), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13354 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13355 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10322) );
  NAND4_X1 U13356 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10326) );
  NAND3_X1 U13357 ( .A1(n10331), .A2(n10351), .A3(n16992), .ZN(n15460) );
  NAND4_X1 U13358 ( .A1(n17979), .A2(n17983), .A3(n10338), .A4(n9665), .ZN(
        n10348) );
  NAND2_X1 U13359 ( .A1(n17975), .A2(n16992), .ZN(n12513) );
  NAND2_X1 U13360 ( .A1(n17993), .A2(n16992), .ZN(n10334) );
  AOI21_X1 U13361 ( .B1(n17032), .B2(n10334), .A(n10333), .ZN(n12509) );
  AOI21_X1 U13362 ( .B1(n10346), .B2(n12513), .A(n12509), .ZN(n10343) );
  INV_X1 U13363 ( .A(n9665), .ZN(n10342) );
  INV_X1 U13364 ( .A(n10338), .ZN(n10336) );
  AOI21_X1 U13365 ( .B1(n17975), .B2(n17968), .A(n18418), .ZN(n10335) );
  AOI21_X1 U13366 ( .B1(n10336), .B2(n10346), .A(n10335), .ZN(n10341) );
  NOR2_X1 U13367 ( .A1(n17999), .A2(n10338), .ZN(n10339) );
  NAND2_X1 U13368 ( .A1(n10349), .A2(n17975), .ZN(n10362) );
  INV_X1 U13369 ( .A(n10362), .ZN(n10337) );
  OAI22_X1 U13370 ( .A1(n17983), .A2(n10339), .B1(n10338), .B2(n10337), .ZN(
        n10340) );
  INV_X1 U13371 ( .A(n10353), .ZN(n10358) );
  XNOR2_X1 U13372 ( .A(n10355), .B(n10354), .ZN(n10357) );
  OAI21_X1 U13373 ( .B1(n10359), .B2(n10358), .A(n18403), .ZN(n12510) );
  NAND2_X1 U13374 ( .A1(n17975), .A2(n18619), .ZN(n12511) );
  NOR2_X1 U13375 ( .A1(n17993), .A2(n12511), .ZN(n12516) );
  NOR2_X1 U13376 ( .A1(n17993), .A2(n16992), .ZN(n15456) );
  OAI21_X1 U13377 ( .B1(n17983), .B2(n18418), .A(n10360), .ZN(n10361) );
  NOR2_X2 U13378 ( .A1(n17971), .A2(n16314), .ZN(n17614) );
  NAND2_X1 U13379 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17581) );
  NOR2_X1 U13380 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18632) );
  INV_X1 U13381 ( .A(n18632), .ZN(n18580) );
  NAND2_X1 U13382 ( .A1(n18631), .A2(n18566), .ZN(n16307) );
  NAND2_X1 U13383 ( .A1(n18580), .A2(n16307), .ZN(n17957) );
  INV_X1 U13384 ( .A(n17957), .ZN(n18616) );
  NAND2_X1 U13385 ( .A1(n10413), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17452) );
  INV_X1 U13386 ( .A(n17458), .ZN(n10363) );
  NAND2_X1 U13387 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17414) );
  NAND2_X1 U13388 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17380) );
  INV_X1 U13389 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17336) );
  NOR2_X1 U13390 ( .A1(n20869), .A2(n17336), .ZN(n17335) );
  NAND2_X1 U13391 ( .A1(n17335), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10408) );
  NAND3_X1 U13392 ( .A1(n17295), .A2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17282) );
  INV_X1 U13393 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17281) );
  NOR2_X2 U13394 ( .A1(n17282), .A2(n17281), .ZN(n17253) );
  INV_X1 U13395 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17617) );
  INV_X1 U13396 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16182) );
  NAND2_X1 U13397 ( .A1(n10422), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10364) );
  XOR2_X2 U13398 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n10364), .Z(
        n16603) );
  INV_X1 U13399 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18549) );
  NAND3_X1 U13400 ( .A1(n18632), .A2(n18622), .A3(n18631), .ZN(n17835) );
  NOR2_X1 U13401 ( .A1(n18549), .A2(n17835), .ZN(n16202) );
  OR2_X1 U13402 ( .A1(n17254), .A2(n9727), .ZN(n16183) );
  NOR2_X1 U13403 ( .A1(n16182), .A2(n16183), .ZN(n10365) );
  NOR2_X1 U13404 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18631), .ZN(n17457) );
  NAND2_X1 U13405 ( .A1(n17457), .A2(n17622), .ZN(n17333) );
  NOR2_X1 U13406 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18625) );
  AOI21_X1 U13407 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18625), .ZN(n18468) );
  NOR3_X2 U13408 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n16309), .ZN(n18303) );
  OAI21_X1 U13409 ( .B1(n17333), .B2(n17617), .A(n17991), .ZN(n17294) );
  NAND2_X1 U13410 ( .A1(n10365), .A2(n17294), .ZN(n16174) );
  INV_X1 U13411 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10368) );
  XOR2_X1 U13412 ( .A(n10368), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n10369) );
  NOR2_X1 U13413 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17333), .ZN(
        n16194) );
  INV_X1 U13414 ( .A(n10365), .ZN(n10366) );
  AOI22_X1 U13415 ( .A1(n18344), .A2(n10366), .B1(n17457), .B2(n10423), .ZN(
        n10367) );
  NAND2_X1 U13416 ( .A1(n10367), .A2(n17622), .ZN(n16185) );
  NOR2_X1 U13417 ( .A1(n16194), .A2(n16185), .ZN(n16172) );
  OAI22_X1 U13418 ( .A1(n16174), .A2(n10369), .B1(n16172), .B2(n10368), .ZN(
        n10370) );
  AOI211_X1 U13419 ( .C1(n17475), .C2(n10414), .A(n16202), .B(n10370), .ZN(
        n10405) );
  INV_X1 U13420 ( .A(n17103), .ZN(n12526) );
  INV_X1 U13421 ( .A(n17620), .ZN(n15631) );
  NOR2_X1 U13422 ( .A1(n15631), .A2(n10371), .ZN(n10382) );
  INV_X1 U13423 ( .A(n17124), .ZN(n10372) );
  NOR2_X1 U13424 ( .A1(n10382), .A2(n10372), .ZN(n10380) );
  NOR2_X1 U13425 ( .A1(n10380), .A2(n17118), .ZN(n10379) );
  INV_X1 U13426 ( .A(n17115), .ZN(n10373) );
  NAND2_X1 U13427 ( .A1(n10379), .A2(n10373), .ZN(n10377) );
  NOR2_X1 U13428 ( .A1(n17111), .A2(n10377), .ZN(n10376) );
  INV_X1 U13429 ( .A(n17108), .ZN(n10374) );
  NAND2_X1 U13430 ( .A1(n10376), .A2(n10374), .ZN(n10375) );
  NOR2_X1 U13431 ( .A1(n12526), .A2(n10375), .ZN(n10399) );
  XNOR2_X1 U13432 ( .A(n10375), .B(n17103), .ZN(n17541) );
  XNOR2_X1 U13433 ( .A(n10376), .B(n17108), .ZN(n10392) );
  XOR2_X1 U13434 ( .A(n10377), .B(n17111), .Z(n10378) );
  NAND2_X1 U13435 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n10378), .ZN(
        n10391) );
  XNOR2_X1 U13436 ( .A(n9990), .B(n10378), .ZN(n17562) );
  XNOR2_X1 U13437 ( .A(n10379), .B(n17115), .ZN(n10389) );
  XOR2_X1 U13438 ( .A(n17118), .B(n10380), .Z(n10381) );
  NAND2_X1 U13439 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n10381), .ZN(
        n10387) );
  INV_X1 U13440 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17905) );
  XNOR2_X1 U13441 ( .A(n17905), .B(n10381), .ZN(n17588) );
  XNOR2_X1 U13442 ( .A(n17124), .B(n10382), .ZN(n10385) );
  OR2_X1 U13443 ( .A1(n17913), .A2(n10385), .ZN(n10386) );
  AOI21_X1 U13444 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17131), .A(
        n17620), .ZN(n10384) );
  INV_X1 U13445 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18595) );
  NOR2_X1 U13446 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17131), .ZN(
        n10383) );
  AOI221_X1 U13447 ( .B1(n17620), .B2(n17131), .C1(n10384), .C2(n18595), .A(
        n10383), .ZN(n17603) );
  XNOR2_X1 U13448 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10385), .ZN(
        n17602) );
  NAND2_X1 U13449 ( .A1(n17603), .A2(n17602), .ZN(n17601) );
  NAND2_X1 U13450 ( .A1(n10386), .A2(n17601), .ZN(n17587) );
  NAND2_X1 U13451 ( .A1(n17588), .A2(n17587), .ZN(n17586) );
  NAND2_X1 U13452 ( .A1(n10387), .A2(n17586), .ZN(n10388) );
  NAND2_X1 U13453 ( .A1(n10389), .A2(n10388), .ZN(n10390) );
  XOR2_X1 U13454 ( .A(n10389), .B(n10388), .Z(n17574) );
  NAND2_X1 U13455 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17574), .ZN(
        n17573) );
  NAND2_X1 U13456 ( .A1(n10390), .A2(n17573), .ZN(n17561) );
  NAND2_X1 U13457 ( .A1(n17562), .A2(n17561), .ZN(n17560) );
  NAND2_X1 U13458 ( .A1(n10391), .A2(n17560), .ZN(n10393) );
  NAND2_X1 U13459 ( .A1(n10392), .A2(n10393), .ZN(n10394) );
  XOR2_X1 U13460 ( .A(n10393), .B(n10392), .Z(n17550) );
  NAND2_X1 U13461 ( .A1(n17550), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17549) );
  NAND2_X1 U13462 ( .A1(n10394), .A2(n17549), .ZN(n17540) );
  NAND2_X1 U13463 ( .A1(n10399), .A2(n10395), .ZN(n10400) );
  INV_X1 U13464 ( .A(n10395), .ZN(n10398) );
  NAND2_X1 U13465 ( .A1(n17541), .A2(n17540), .ZN(n10397) );
  NAND2_X1 U13466 ( .A1(n10399), .A2(n10398), .ZN(n10396) );
  OAI211_X1 U13467 ( .C1(n10399), .C2(n10398), .A(n10397), .B(n10396), .ZN(
        n17523) );
  NAND2_X1 U13468 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17523), .ZN(
        n17522) );
  NAND2_X1 U13469 ( .A1(n10214), .A2(n17493), .ZN(n17771) );
  INV_X1 U13470 ( .A(n17771), .ZN(n17430) );
  NAND2_X1 U13471 ( .A1(n17670), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17302) );
  INV_X1 U13472 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17627) );
  NOR2_X1 U13473 ( .A1(n17627), .A2(n12521), .ZN(n15566) );
  NAND2_X1 U13474 ( .A1(n17628), .A2(n15566), .ZN(n16187) );
  NAND3_X1 U13475 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n18575), .ZN(n16199) );
  AND2_X1 U13476 ( .A1(n15566), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16178) );
  NAND2_X1 U13477 ( .A1(n17628), .A2(n16178), .ZN(n16169) );
  OAI21_X1 U13478 ( .B1(n16177), .B2(n16169), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10401) );
  OAI21_X1 U13479 ( .B1(n16187), .B2(n16199), .A(n10401), .ZN(n16204) );
  INV_X1 U13480 ( .A(n17614), .ZN(n17625) );
  INV_X1 U13481 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17649) );
  INV_X1 U13482 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17676) );
  NAND2_X1 U13483 ( .A1(n10402), .A2(n17691), .ZN(n17315) );
  NOR2_X1 U13484 ( .A1(n17676), .A2(n17315), .ZN(n17291) );
  NAND2_X1 U13485 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17291), .ZN(
        n17290) );
  NAND2_X1 U13486 ( .A1(n15566), .A2(n17638), .ZN(n16189) );
  NAND2_X1 U13487 ( .A1(n16178), .A2(n17638), .ZN(n16170) );
  OAI21_X1 U13488 ( .B1(n16177), .B2(n16170), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10403) );
  OAI21_X1 U13489 ( .B1(n16199), .B2(n16189), .A(n10403), .ZN(n16205) );
  AOI22_X1 U13490 ( .A1(n9632), .A2(n16204), .B1(n17529), .B2(n16205), .ZN(
        n10404) );
  XOR2_X1 U13491 ( .A(n10422), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16330) );
  OAI21_X1 U13492 ( .B1(n10420), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n10423), .ZN(n17267) );
  INV_X1 U13493 ( .A(n17267), .ZN(n16352) );
  INV_X1 U13494 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17296) );
  INV_X1 U13495 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17366) );
  NAND2_X1 U13496 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10407), .ZN(
        n17330) );
  INV_X1 U13497 ( .A(n10417), .ZN(n10416) );
  NOR2_X1 U13498 ( .A1(n10408), .A2(n10416), .ZN(n10418) );
  INV_X1 U13499 ( .A(n10418), .ZN(n10410) );
  NOR2_X1 U13500 ( .A1(n17296), .A2(n10410), .ZN(n10419) );
  NAND2_X1 U13501 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n10419), .ZN(
        n17251) );
  INV_X1 U13502 ( .A(n17251), .ZN(n10409) );
  NAND2_X1 U13503 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n10409), .ZN(
        n10421) );
  OAI21_X1 U13504 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n10409), .A(
        n10421), .ZN(n17283) );
  INV_X1 U13505 ( .A(n17283), .ZN(n16371) );
  AOI21_X1 U13506 ( .B1(n17296), .B2(n10410), .A(n10419), .ZN(n17310) );
  NAND2_X1 U13507 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n10417), .ZN(
        n10412) );
  NAND2_X1 U13508 ( .A1(n17335), .A2(n10417), .ZN(n17293) );
  INV_X1 U13509 ( .A(n17293), .ZN(n10411) );
  AOI21_X1 U13510 ( .B1(n17336), .B2(n10412), .A(n10411), .ZN(n17334) );
  INV_X1 U13511 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17425) );
  INV_X1 U13512 ( .A(n17437), .ZN(n17460) );
  INV_X1 U13513 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17555) );
  NAND2_X1 U13514 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10413), .ZN(
        n16604) );
  NOR2_X1 U13515 ( .A1(n17555), .A2(n16604), .ZN(n16592) );
  NAND2_X1 U13516 ( .A1(n17454), .A2(n16592), .ZN(n17456) );
  NOR2_X1 U13517 ( .A1(n17460), .A2(n17456), .ZN(n16509) );
  NAND2_X1 U13518 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16509), .ZN(
        n17411) );
  NOR2_X1 U13519 ( .A1(n17425), .A2(n17411), .ZN(n16487) );
  INV_X1 U13520 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16675) );
  NAND2_X1 U13521 ( .A1(n16487), .A2(n16675), .ZN(n16481) );
  NAND3_X1 U13522 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17398), .A3(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16463) );
  INV_X1 U13523 ( .A(n17380), .ZN(n10415) );
  AOI21_X1 U13524 ( .B1(n17366), .B2(n17330), .A(n10417), .ZN(n17371) );
  NOR2_X1 U13525 ( .A1(n16430), .A2(n16603), .ZN(n16422) );
  AOI22_X1 U13526 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n10417), .B1(
        n10416), .B2(n20869), .ZN(n17353) );
  INV_X1 U13527 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17324) );
  AOI21_X1 U13528 ( .B1(n17324), .B2(n17293), .A(n10418), .ZN(n17321) );
  NOR2_X1 U13529 ( .A1(n16403), .A2(n16603), .ZN(n16392) );
  OAI21_X1 U13530 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n10419), .A(
        n17251), .ZN(n17297) );
  INV_X1 U13531 ( .A(n17297), .ZN(n16382) );
  AOI21_X1 U13532 ( .B1(n9726), .B2(n10421), .A(n10420), .ZN(n17276) );
  NOR2_X1 U13533 ( .A1(n9664), .A2(n9733), .ZN(n16342) );
  AOI21_X1 U13534 ( .B1(n10423), .B2(n16182), .A(n10422), .ZN(n16343) );
  NOR2_X1 U13535 ( .A1(n16341), .A2(n16603), .ZN(n16329) );
  NAND4_X1 U13536 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18631), .A3(n18622), 
        .A4(n16309), .ZN(n18467) );
  NOR4_X1 U13537 ( .A1(n16330), .A2(n16329), .A3(n16603), .A4(n18467), .ZN(
        n10438) );
  INV_X2 U13538 ( .A(n18629), .ZN(n18610) );
  NAND2_X2 U13539 ( .A1(n18610), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18552) );
  INV_X1 U13540 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18483) );
  INV_X1 U13541 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18490) );
  NAND2_X1 U13542 ( .A1(n18483), .A2(n18490), .ZN(n18474) );
  NAND3_X1 U13543 ( .A1(n18488), .A2(n18552), .A3(n18474), .ZN(n18478) );
  INV_X1 U13544 ( .A(n18478), .ZN(n18618) );
  NAND2_X1 U13545 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18613) );
  OAI211_X1 U13546 ( .C1(n18619), .C2(n18618), .A(n18613), .B(n16309), .ZN(
        n18452) );
  NAND3_X1 U13547 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n10425) );
  INV_X1 U13548 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18541) );
  NAND2_X1 U13549 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18631), .ZN(n18462) );
  OAI211_X1 U13550 ( .C1(n17621), .C2(n18462), .A(n16571), .B(n17835), .ZN(
        n10424) );
  INV_X1 U13551 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18535) );
  INV_X1 U13552 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18530) );
  INV_X1 U13553 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18526) );
  INV_X1 U13554 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18524) );
  INV_X1 U13555 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18513) );
  INV_X1 U13556 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18505) );
  INV_X1 U13557 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18500) );
  INV_X1 U13558 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18496) );
  NAND3_X1 U13559 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16629) );
  NOR2_X1 U13560 ( .A1(n18496), .A2(n16629), .ZN(n16611) );
  NAND2_X1 U13561 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16611), .ZN(n16602) );
  NOR2_X1 U13562 ( .A1(n18500), .A2(n16602), .ZN(n16580) );
  NAND2_X1 U13563 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16580), .ZN(n16579) );
  NOR2_X1 U13564 ( .A1(n18505), .A2(n16579), .ZN(n16568) );
  NAND4_X1 U13565 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16568), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16508) );
  NOR2_X1 U13566 ( .A1(n18513), .A2(n16508), .ZN(n16501) );
  NAND3_X1 U13567 ( .A1(n16501), .A2(P3_REIP_REG_14__SCAN_IN), .A3(
        P3_REIP_REG_13__SCAN_IN), .ZN(n16446) );
  NAND3_X1 U13568 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16448) );
  NOR4_X1 U13569 ( .A1(n18526), .A2(n18524), .A3(n16446), .A4(n16448), .ZN(
        n16436) );
  NAND2_X1 U13570 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16436), .ZN(n16420) );
  NOR2_X1 U13571 ( .A1(n18530), .A2(n16420), .ZN(n16411) );
  NAND2_X1 U13572 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16411), .ZN(n16402) );
  NOR2_X1 U13573 ( .A1(n18535), .A2(n16402), .ZN(n16397) );
  NAND2_X1 U13574 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16397), .ZN(n10426) );
  AND2_X1 U13575 ( .A1(n10426), .A2(n16646), .ZN(n16398) );
  INV_X1 U13576 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18539) );
  NOR2_X1 U13577 ( .A1(n16646), .A2(n16676), .ZN(n16479) );
  INV_X1 U13578 ( .A(n16479), .ZN(n16679) );
  OAI21_X1 U13579 ( .B1(n18541), .B2(n16385), .A(n16679), .ZN(n16378) );
  INV_X1 U13580 ( .A(n16378), .ZN(n16363) );
  AOI21_X1 U13581 ( .B1(n16646), .B2(n10425), .A(n16363), .ZN(n16338) );
  NOR2_X1 U13582 ( .A1(n16666), .A2(n10426), .ZN(n16384) );
  NAND2_X1 U13583 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16384), .ZN(n16377) );
  NAND4_X1 U13584 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16362), .ZN(n10435) );
  NOR2_X1 U13585 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n10435), .ZN(n16333) );
  INV_X1 U13586 ( .A(n16333), .ZN(n10427) );
  AOI21_X1 U13587 ( .B1(n16338), .B2(n10427), .A(n18549), .ZN(n10437) );
  NAND2_X1 U13588 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18549), .ZN(n10434) );
  NAND2_X1 U13589 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18619), .ZN(n10428) );
  AOI211_X4 U13590 ( .C1(n16309), .C2(n18613), .A(n10429), .B(n10428), .ZN(
        n16631) );
  INV_X1 U13591 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16462) );
  NOR3_X1 U13592 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16644) );
  NAND2_X1 U13593 ( .A1(n16644), .A2(n16632), .ZN(n16630) );
  NOR2_X1 U13594 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16630), .ZN(n16616) );
  INV_X1 U13595 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16896) );
  NAND2_X1 U13596 ( .A1(n16616), .A2(n16896), .ZN(n16612) );
  INV_X1 U13597 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16589) );
  NAND2_X1 U13598 ( .A1(n16597), .A2(n16589), .ZN(n16588) );
  INV_X1 U13599 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16567) );
  NAND2_X1 U13600 ( .A1(n16569), .A2(n16567), .ZN(n16564) );
  INV_X1 U13601 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16538) );
  NAND2_X1 U13602 ( .A1(n16542), .A2(n16538), .ZN(n16537) );
  INV_X1 U13603 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16518) );
  NAND2_X1 U13604 ( .A1(n16521), .A2(n16518), .ZN(n16517) );
  INV_X1 U13605 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16495) );
  NAND2_X1 U13606 ( .A1(n16498), .A2(n16495), .ZN(n16494) );
  INV_X1 U13607 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16475) );
  NAND2_X1 U13608 ( .A1(n16477), .A2(n16475), .ZN(n16472) );
  INV_X1 U13609 ( .A(n16472), .ZN(n16459) );
  NAND2_X1 U13610 ( .A1(n16462), .A2(n16459), .ZN(n16458) );
  INV_X1 U13611 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16774) );
  NAND2_X1 U13612 ( .A1(n16433), .A2(n16774), .ZN(n16427) );
  NOR2_X1 U13613 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16427), .ZN(n16414) );
  INV_X1 U13614 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16682) );
  NAND2_X1 U13615 ( .A1(n16414), .A2(n16682), .ZN(n16407) );
  NOR2_X1 U13616 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16407), .ZN(n16379) );
  INV_X1 U13617 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16388) );
  NAND2_X1 U13618 ( .A1(n16379), .A2(n16388), .ZN(n16369) );
  NOR2_X1 U13619 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16369), .ZN(n16368) );
  INV_X1 U13620 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16684) );
  NAND2_X1 U13621 ( .A1(n16368), .A2(n16684), .ZN(n16364) );
  NOR2_X1 U13622 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16364), .ZN(n16350) );
  INV_X1 U13623 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16721) );
  NAND2_X1 U13624 ( .A1(n16350), .A2(n16721), .ZN(n16331) );
  NOR2_X1 U13625 ( .A1(n16673), .A2(n16331), .ZN(n16334) );
  INV_X1 U13626 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16691) );
  INV_X1 U13627 ( .A(n18452), .ZN(n10430) );
  AOI211_X1 U13628 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18619), .A(n10430), .B(
        n10429), .ZN(n10431) );
  AOI22_X1 U13629 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n9591), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16662), .ZN(n10432) );
  OR2_X1 U13630 ( .A1(n10438), .A2(n9681), .ZN(P3_U2640) );
  INV_X1 U13631 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16037) );
  INV_X1 U13632 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15039) );
  INV_X1 U13633 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16029) );
  INV_X1 U13634 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15000) );
  INV_X1 U13635 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12489) );
  INV_X1 U13636 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10442) );
  XNOR2_X1 U13637 ( .A(n10441), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14984) );
  INV_X1 U13638 ( .A(n14984), .ZN(n10468) );
  NAND2_X1 U13639 ( .A1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10439) );
  NAND2_X2 U13640 ( .A1(n10440), .A2(n10439), .ZN(n13945) );
  AOI21_X1 U13641 ( .B1(n10442), .B2(n9705), .A(n10441), .ZN(n14993) );
  INV_X1 U13642 ( .A(n10443), .ZN(n10445) );
  OAI21_X1 U13643 ( .B1(n10445), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n9705), .ZN(n12491) );
  INV_X1 U13644 ( .A(n12491), .ZN(n15970) );
  AOI21_X1 U13645 ( .B1(n15000), .B2(n10444), .A(n10445), .ZN(n15004) );
  OAI21_X1 U13646 ( .B1(n10446), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n10444), .ZN(n15019) );
  INV_X1 U13647 ( .A(n15019), .ZN(n15983) );
  AOI21_X1 U13648 ( .B1(n16029), .B2(n9635), .A(n10446), .ZN(n16031) );
  OAI21_X1 U13649 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n10447), .A(
        n9635), .ZN(n15031) );
  INV_X1 U13650 ( .A(n15031), .ZN(n15994) );
  AOI21_X1 U13651 ( .B1(n15039), .B2(n9703), .A(n10447), .ZN(n15042) );
  OAI21_X1 U13652 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10448), .A(
        n9703), .ZN(n15052) );
  INV_X1 U13653 ( .A(n15052), .ZN(n14804) );
  AOI21_X1 U13654 ( .B1(n16037), .B2(n10465), .A(n10448), .ZN(n16040) );
  INV_X1 U13655 ( .A(n16040), .ZN(n14826) );
  AOI21_X1 U13656 ( .B1(n20750), .B2(n10464), .A(n10449), .ZN(n18679) );
  AOI21_X1 U13657 ( .B1(n18703), .B2(n9690), .A(n10450), .ZN(n18702) );
  AOI21_X1 U13658 ( .B1(n18736), .B2(n10463), .A(n10451), .ZN(n18729) );
  AOI21_X1 U13659 ( .B1(n16079), .B2(n10462), .A(n10452), .ZN(n18755) );
  AOI21_X1 U13660 ( .B1(n16095), .B2(n10460), .A(n10453), .ZN(n18764) );
  AOI21_X1 U13661 ( .B1(n18794), .B2(n10459), .A(n10461), .ZN(n18787) );
  AOI21_X1 U13662 ( .B1(n15113), .B2(n10458), .A(n9691), .ZN(n15114) );
  AOI21_X1 U13663 ( .B1(n20762), .B2(n10457), .A(n10454), .ZN(n18825) );
  AOI21_X1 U13664 ( .B1(n20802), .B2(n10456), .A(n10455), .ZN(n13948) );
  OAI22_X1 U13665 ( .A1(n19751), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n14020) );
  INV_X1 U13666 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18856) );
  OAI22_X1 U13667 ( .A1(n19751), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n18856), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14019) );
  AND2_X1 U13668 ( .A1(n14020), .A2(n14019), .ZN(n13966) );
  OAI21_X1 U13669 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n10456), .ZN(n13968) );
  NAND2_X1 U13670 ( .A1(n13966), .A2(n13968), .ZN(n13946) );
  NOR2_X1 U13671 ( .A1(n13948), .A2(n13946), .ZN(n18841) );
  OAI21_X1 U13672 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10455), .A(
        n10457), .ZN(n18988) );
  NAND2_X1 U13673 ( .A1(n18841), .A2(n18988), .ZN(n18823) );
  NOR2_X1 U13674 ( .A1(n18825), .A2(n18823), .ZN(n18811) );
  OAI21_X1 U13675 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10454), .A(
        n10458), .ZN(n18812) );
  NAND2_X1 U13676 ( .A1(n18811), .A2(n18812), .ZN(n13972) );
  NOR2_X1 U13677 ( .A1(n15114), .A2(n13972), .ZN(n18795) );
  OAI21_X1 U13678 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n9691), .A(
        n10459), .ZN(n18796) );
  NAND2_X1 U13679 ( .A1(n18795), .A2(n18796), .ZN(n18785) );
  NOR2_X1 U13680 ( .A1(n18787), .A2(n18785), .ZN(n18776) );
  OAI21_X1 U13681 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10461), .A(
        n10460), .ZN(n18777) );
  NAND2_X1 U13682 ( .A1(n18776), .A2(n18777), .ZN(n18762) );
  NOR2_X1 U13683 ( .A1(n18764), .A2(n18762), .ZN(n13899) );
  OAI21_X1 U13684 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10453), .A(
        n10462), .ZN(n16087) );
  NAND2_X1 U13685 ( .A1(n13899), .A2(n16087), .ZN(n18747) );
  NOR2_X1 U13686 ( .A1(n18755), .A2(n18747), .ZN(n18737) );
  OAI21_X1 U13687 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10452), .A(
        n10463), .ZN(n18738) );
  NAND2_X1 U13688 ( .A1(n18737), .A2(n18738), .ZN(n18727) );
  NOR2_X1 U13689 ( .A1(n18729), .A2(n18727), .ZN(n18714) );
  OAI21_X1 U13690 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10451), .A(
        n9690), .ZN(n18715) );
  NAND2_X1 U13691 ( .A1(n18714), .A2(n18715), .ZN(n18700) );
  NOR2_X1 U13692 ( .A1(n18702), .A2(n18700), .ZN(n18689) );
  OAI21_X1 U13693 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n10450), .A(
        n10464), .ZN(n18690) );
  NAND2_X1 U13694 ( .A1(n18689), .A2(n18690), .ZN(n18677) );
  NOR2_X1 U13695 ( .A1(n18679), .A2(n18677), .ZN(n18664) );
  OAI21_X1 U13696 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10449), .A(
        n10465), .ZN(n15059) );
  NAND2_X1 U13697 ( .A1(n18664), .A2(n15059), .ZN(n14822) );
  NOR2_X1 U13698 ( .A1(n10466), .A2(n13209), .ZN(n15993) );
  NOR2_X1 U13699 ( .A1(n15994), .A2(n15993), .ZN(n15992) );
  NOR2_X1 U13700 ( .A1(n10466), .A2(n15992), .ZN(n14798) );
  NOR2_X1 U13701 ( .A1(n15004), .A2(n14782), .ZN(n14781) );
  NOR2_X1 U13702 ( .A1(n10466), .A2(n14781), .ZN(n15969) );
  NOR2_X1 U13703 ( .A1(n10466), .A2(n14770), .ZN(n10469) );
  NOR2_X1 U13704 ( .A1(n10468), .A2(n10469), .ZN(n15960) );
  INV_X1 U13705 ( .A(n15960), .ZN(n10471) );
  INV_X1 U13706 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19692) );
  NAND3_X1 U13707 ( .A1(n19549), .A2(n19751), .A3(n19692), .ZN(n10467) );
  NOR2_X2 U13708 ( .A1(n14021), .A2(n10467), .ZN(n18827) );
  AOI21_X1 U13709 ( .B1(n10469), .B2(n10468), .A(n18877), .ZN(n10470) );
  NAND2_X1 U13710 ( .A1(n10471), .A2(n10470), .ZN(n11182) );
  INV_X1 U13711 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n13908) );
  AND2_X4 U13712 ( .A1(n13619), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13146) );
  INV_X2 U13713 ( .A(n13027), .ZN(n10823) );
  AOI22_X1 U13714 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10477) );
  AND2_X2 U13715 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13716 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10476) );
  AND2_X2 U13717 ( .A1(n10473), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10821) );
  AND2_X4 U13718 ( .A1(n10821), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13149) );
  AOI22_X1 U13719 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10475) );
  AND2_X4 U13720 ( .A1(n13619), .A2(n10814), .ZN(n10812) );
  AOI22_X1 U13721 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10474) );
  NAND4_X1 U13722 ( .A1(n10477), .A2(n10476), .A3(n10475), .A4(n10474), .ZN(
        n10584) );
  NAND2_X1 U13723 ( .A1(n10584), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10483) );
  AOI22_X1 U13724 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13725 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13726 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13727 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10478) );
  NAND4_X1 U13728 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10591) );
  NAND2_X1 U13729 ( .A1(n10591), .A2(n10547), .ZN(n10482) );
  NAND2_X2 U13730 ( .A1(n10483), .A2(n10482), .ZN(n10611) );
  INV_X1 U13731 ( .A(n10611), .ZN(n10494) );
  AOI22_X1 U13732 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13733 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13734 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13735 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U13736 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10587) );
  NAND2_X1 U13737 ( .A1(n10587), .A2(n10547), .ZN(n10493) );
  AOI22_X1 U13738 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13739 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10490) );
  NAND4_X1 U13740 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10580) );
  NAND2_X1 U13741 ( .A1(n10580), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10492) );
  NOR2_X2 U13742 ( .A1(n10494), .A2(n12785), .ZN(n10575) );
  AOI22_X1 U13743 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13744 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13745 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13746 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13747 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13748 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U13749 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13750 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13751 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13752 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U13753 ( .A1(n10812), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13754 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10503) );
  NAND4_X1 U13755 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10579) );
  NAND2_X1 U13756 ( .A1(n10579), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10512) );
  AOI22_X1 U13757 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13758 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13759 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13760 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10507) );
  NAND4_X1 U13761 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10586) );
  NAND2_X1 U13762 ( .A1(n10586), .A2(n10547), .ZN(n10511) );
  NAND2_X2 U13763 ( .A1(n10512), .A2(n10511), .ZN(n10610) );
  AND2_X2 U13764 ( .A1(n10575), .A2(n10513), .ZN(n10616) );
  AOI22_X1 U13765 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13766 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13767 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13768 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10815), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10514) );
  NAND4_X1 U13769 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10590) );
  NAND2_X1 U13770 ( .A1(n10590), .A2(n10547), .ZN(n10523) );
  AOI22_X1 U13771 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13772 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13773 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10519) );
  NAND4_X1 U13774 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10583) );
  NAND2_X1 U13775 ( .A1(n10583), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10522) );
  NAND2_X2 U13776 ( .A1(n10523), .A2(n10522), .ZN(n10612) );
  AOI22_X1 U13777 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13778 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13779 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13780 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10524) );
  NAND4_X1 U13781 ( .A1(n10527), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(
        n10528) );
  NAND2_X1 U13782 ( .A1(n10528), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10535) );
  AOI22_X1 U13783 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13784 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13785 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13786 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10529) );
  NAND4_X1 U13787 ( .A1(n10532), .A2(n10531), .A3(n10530), .A4(n10529), .ZN(
        n10533) );
  NOR2_X1 U13788 ( .A1(n13165), .A2(n12808), .ZN(n10536) );
  NAND2_X2 U13789 ( .A1(n10616), .A2(n10536), .ZN(n10627) );
  NAND2_X1 U13790 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10540) );
  NAND2_X1 U13791 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10539) );
  NAND2_X1 U13792 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10538) );
  NAND2_X1 U13793 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10537) );
  NAND4_X1 U13794 ( .A1(n10540), .A2(n10539), .A3(n10538), .A4(n10537), .ZN(
        n10546) );
  NAND2_X1 U13795 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10544) );
  NAND2_X1 U13796 ( .A1(n10812), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10543) );
  NAND2_X1 U13797 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10542) );
  OR2_X1 U13798 ( .A1(n13027), .A2(n19044), .ZN(n10541) );
  NAND4_X1 U13799 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10545) );
  NOR2_X1 U13800 ( .A1(n10546), .A2(n10545), .ZN(n10589) );
  NAND2_X1 U13801 ( .A1(n10589), .A2(n10547), .ZN(n10560) );
  NAND2_X1 U13802 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10551) );
  NAND2_X1 U13803 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10550) );
  NAND2_X1 U13804 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10549) );
  NAND2_X1 U13805 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10548) );
  NAND4_X1 U13806 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n10558) );
  NAND2_X1 U13807 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10556) );
  NAND2_X1 U13808 ( .A1(n10812), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10555) );
  NAND2_X1 U13809 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10554) );
  OR2_X1 U13810 ( .A1(n13027), .A2(n12187), .ZN(n10553) );
  NAND4_X1 U13811 ( .A1(n10556), .A2(n10555), .A3(n10554), .A4(n10553), .ZN(
        n10557) );
  NOR2_X1 U13812 ( .A1(n10558), .A2(n10557), .ZN(n10582) );
  NAND2_X1 U13813 ( .A1(n10582), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10559) );
  AOI22_X1 U13814 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13815 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13816 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13817 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10561) );
  NAND4_X1 U13818 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n10570) );
  AOI22_X1 U13819 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13820 ( .A1(n10552), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13821 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13822 ( .A1(n10815), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10565) );
  NAND4_X1 U13823 ( .A1(n10568), .A2(n10567), .A3(n10566), .A4(n10565), .ZN(
        n10569) );
  MUX2_X2 U13824 ( .A(n10570), .B(n10569), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13645) );
  AND2_X1 U13825 ( .A1(n13162), .A2(n10637), .ZN(n10661) );
  NAND2_X1 U13826 ( .A1(n10774), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10572) );
  NAND2_X1 U13827 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10571) );
  OAI211_X1 U13828 ( .C1(n13908), .C2(n9622), .A(n10572), .B(n10571), .ZN(
        n10573) );
  INV_X1 U13829 ( .A(n10573), .ZN(n10603) );
  INV_X1 U13830 ( .A(n10614), .ZN(n10574) );
  AND2_X1 U13831 ( .A1(n10841), .A2(n13645), .ZN(n19734) );
  NAND2_X1 U13832 ( .A1(n12774), .A2(n19734), .ZN(n13671) );
  INV_X1 U13833 ( .A(n10579), .ZN(n10581) );
  NAND4_X1 U13834 ( .A1(n10582), .A2(n10581), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(n10580), .ZN(n10597) );
  INV_X1 U13835 ( .A(n10583), .ZN(n10585) );
  NAND2_X1 U13836 ( .A1(n10585), .A2(n10584), .ZN(n10596) );
  INV_X1 U13837 ( .A(n10586), .ZN(n10588) );
  NAND4_X1 U13838 ( .A1(n10589), .A2(n10588), .A3(n10547), .A4(n10587), .ZN(
        n10594) );
  INV_X1 U13839 ( .A(n10590), .ZN(n10592) );
  NAND2_X1 U13840 ( .A1(n10592), .A2(n10591), .ZN(n10593) );
  OAI21_X1 U13841 ( .B1(n10597), .B2(n10596), .A(n10595), .ZN(n10598) );
  NAND3_X1 U13842 ( .A1(n10600), .A2(n13671), .A3(n13437), .ZN(n10601) );
  INV_X1 U13844 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15364) );
  OR2_X1 U13845 ( .A1(n10689), .A2(n15364), .ZN(n10602) );
  INV_X1 U13846 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U13847 ( .A1(n10774), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10605) );
  NAND2_X1 U13848 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10604) );
  OAI211_X1 U13849 ( .C1(n9622), .C2(n10606), .A(n10605), .B(n10604), .ZN(
        n10607) );
  INV_X1 U13850 ( .A(n10607), .ZN(n10609) );
  INV_X1 U13851 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12460) );
  OR2_X1 U13852 ( .A1(n10689), .A2(n12460), .ZN(n10608) );
  MUX2_X1 U13853 ( .A(n10612), .B(n10611), .S(n12785), .Z(n10613) );
  NOR2_X1 U13854 ( .A1(n13645), .A2(n19751), .ZN(n19744) );
  NAND2_X1 U13855 ( .A1(n10615), .A2(n19744), .ZN(n10619) );
  AND2_X1 U13856 ( .A1(n19045), .A2(n10806), .ZN(n10617) );
  NAND2_X1 U13857 ( .A1(n19737), .A2(n10617), .ZN(n12799) );
  NAND3_X1 U13858 ( .A1(n12799), .A2(n12743), .A3(n10627), .ZN(n10618) );
  AND2_X2 U13859 ( .A1(n10619), .A2(n10618), .ZN(n10648) );
  NAND2_X1 U13860 ( .A1(n10837), .A2(n12785), .ZN(n12767) );
  AND2_X1 U13861 ( .A1(n12767), .A2(n13188), .ZN(n10621) );
  NAND2_X1 U13862 ( .A1(n10620), .A2(n10837), .ZN(n12772) );
  NAND2_X1 U13863 ( .A1(n12772), .A2(n19055), .ZN(n12769) );
  NAND2_X1 U13864 ( .A1(n12811), .A2(n10610), .ZN(n10625) );
  NAND2_X1 U13865 ( .A1(n10651), .A2(n10637), .ZN(n10626) );
  NAND2_X1 U13866 ( .A1(n9614), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10631) );
  INV_X1 U13867 ( .A(n10780), .ZN(n10629) );
  NAND2_X2 U13868 ( .A1(n10629), .A2(n10628), .ZN(n13656) );
  AOI22_X1 U13869 ( .A1(n13656), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13672), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10630) );
  NAND2_X1 U13870 ( .A1(n10631), .A2(n10630), .ZN(n10656) );
  AND2_X1 U13871 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10632) );
  INV_X1 U13872 ( .A(n9621), .ZN(n10633) );
  NAND2_X1 U13873 ( .A1(n10633), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10634) );
  NAND2_X1 U13874 ( .A1(n10635), .A2(n10634), .ZN(n10636) );
  AOI21_X2 U13875 ( .B1(n9615), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10636), .ZN(n10655) );
  XNOR2_X1 U13876 ( .A(n10656), .B(n10655), .ZN(n12167) );
  INV_X1 U13877 ( .A(n10637), .ZN(n10638) );
  NOR2_X1 U13878 ( .A1(n10638), .A2(n12768), .ZN(n10639) );
  AOI22_X1 U13879 ( .A1(n12792), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13672), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U13880 ( .A1(n10641), .A2(n10640), .ZN(n12158) );
  NAND2_X1 U13881 ( .A1(n10661), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10646) );
  INV_X1 U13882 ( .A(n13672), .ZN(n10645) );
  INV_X1 U13883 ( .A(n9621), .ZN(n10642) );
  NAND2_X1 U13884 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10643) );
  NAND2_X1 U13885 ( .A1(n9616), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10653) );
  INV_X1 U13886 ( .A(n10649), .ZN(n10650) );
  NAND3_X1 U13887 ( .A1(n10651), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10650), 
        .ZN(n10652) );
  NAND2_X1 U13888 ( .A1(n12167), .A2(n12166), .ZN(n10659) );
  INV_X1 U13889 ( .A(n10655), .ZN(n10657) );
  NAND2_X1 U13890 ( .A1(n10659), .A2(n10658), .ZN(n12163) );
  INV_X1 U13891 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12810) );
  INV_X1 U13892 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13394) );
  INV_X1 U13893 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n14224) );
  NAND2_X1 U13894 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10662) );
  NOR2_X1 U13895 ( .A1(n9663), .A2(n10664), .ZN(n10667) );
  NAND2_X1 U13896 ( .A1(n9614), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10666) );
  AOI21_X1 U13897 ( .B1(n19751), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U13898 ( .A1(n10666), .A2(n10665), .ZN(n10668) );
  XNOR2_X1 U13899 ( .A(n10667), .B(n10668), .ZN(n12164) );
  NAND2_X1 U13900 ( .A1(n12163), .A2(n12164), .ZN(n10671) );
  INV_X1 U13901 ( .A(n10667), .ZN(n10669) );
  OR2_X1 U13902 ( .A1(n10669), .A2(n10668), .ZN(n10670) );
  NAND2_X2 U13903 ( .A1(n10671), .A2(n10670), .ZN(n12157) );
  INV_X1 U13904 ( .A(n12157), .ZN(n10681) );
  NAND2_X1 U13905 ( .A1(n9614), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10674) );
  NAND2_X1 U13906 ( .A1(n13672), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10673) );
  INV_X1 U13907 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10678) );
  INV_X1 U13908 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16155) );
  AOI22_X1 U13909 ( .A1(n12555), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10676) );
  INV_X1 U13910 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13938) );
  AOI22_X1 U13911 ( .A1(n12555), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10683) );
  NAND2_X1 U13912 ( .A1(n10774), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10682) );
  OAI211_X1 U13913 ( .C1(n10689), .C2(n13938), .A(n10683), .B(n10682), .ZN(
        n10684) );
  INV_X1 U13914 ( .A(n10684), .ZN(n13939) );
  INV_X1 U13915 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13534) );
  AOI22_X1 U13916 ( .A1(n12555), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10686) );
  INV_X1 U13917 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12828) );
  OR2_X1 U13918 ( .A1(n10689), .A2(n12828), .ZN(n10685) );
  OAI211_X1 U13919 ( .C1(n13534), .C2(n10675), .A(n10686), .B(n10685), .ZN(
        n13531) );
  AOI22_X1 U13920 ( .A1(n12555), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10688) );
  NAND2_X1 U13921 ( .A1(n10774), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10687) );
  OAI211_X1 U13922 ( .C1(n10689), .C2(n9839), .A(n10688), .B(n10687), .ZN(
        n13597) );
  INV_X1 U13923 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14181) );
  AOI22_X1 U13924 ( .A1(n12555), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10691) );
  NAND2_X1 U13925 ( .A1(n10774), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10690) );
  OAI211_X1 U13926 ( .C1(n10689), .C2(n14181), .A(n10691), .B(n10690), .ZN(
        n13545) );
  INV_X1 U13927 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U13928 ( .A1(n12555), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10693) );
  INV_X1 U13929 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15412) );
  OR2_X1 U13930 ( .A1(n10689), .A2(n15412), .ZN(n10692) );
  OAI211_X1 U13931 ( .C1(n12324), .C2(n10675), .A(n10693), .B(n10692), .ZN(
        n13539) );
  INV_X1 U13932 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11030) );
  NAND2_X1 U13933 ( .A1(n10774), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10695) );
  NAND2_X1 U13934 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10694) );
  OAI211_X1 U13935 ( .C1(n9622), .C2(n11030), .A(n10695), .B(n10694), .ZN(
        n10696) );
  INV_X1 U13936 ( .A(n10696), .ZN(n10698) );
  INV_X1 U13937 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15393) );
  OR2_X1 U13938 ( .A1(n10689), .A2(n15393), .ZN(n10697) );
  INV_X1 U13939 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13940 ( .A1(n12555), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10700) );
  INV_X1 U13941 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15367) );
  OR2_X1 U13942 ( .A1(n10689), .A2(n15367), .ZN(n10699) );
  OAI211_X1 U13943 ( .C1(n10701), .C2(n10675), .A(n10700), .B(n10699), .ZN(
        n13592) );
  INV_X1 U13944 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U13945 ( .A1(n12555), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10703) );
  NAND2_X1 U13946 ( .A1(n10774), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10702) );
  OAI211_X1 U13947 ( .C1(n10689), .C2(n12384), .A(n10703), .B(n10702), .ZN(
        n13763) );
  INV_X1 U13948 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13949 ( .A1(n10774), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U13950 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10704) );
  OAI211_X1 U13951 ( .C1(n9622), .C2(n11095), .A(n10705), .B(n10704), .ZN(
        n10706) );
  INV_X1 U13952 ( .A(n10706), .ZN(n10708) );
  INV_X1 U13953 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16069) );
  OR2_X1 U13954 ( .A1(n10689), .A2(n16069), .ZN(n10707) );
  INV_X1 U13955 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n10711) );
  NAND2_X1 U13956 ( .A1(n10774), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10710) );
  NAND2_X1 U13957 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10709) );
  OAI211_X1 U13958 ( .C1(n9622), .C2(n10711), .A(n10710), .B(n10709), .ZN(
        n10712) );
  INV_X1 U13959 ( .A(n10712), .ZN(n10714) );
  INV_X1 U13960 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15315) );
  OR2_X1 U13961 ( .A1(n10689), .A2(n15315), .ZN(n10713) );
  NAND2_X1 U13962 ( .A1(n10714), .A2(n10713), .ZN(n13927) );
  INV_X1 U13963 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U13964 ( .A1(n10774), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10716) );
  NAND2_X1 U13965 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10715) );
  OAI211_X1 U13966 ( .C1(n11111), .C2(n9622), .A(n10716), .B(n10715), .ZN(
        n10717) );
  INV_X1 U13967 ( .A(n10717), .ZN(n10719) );
  INV_X1 U13968 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15289) );
  OR2_X1 U13969 ( .A1(n10689), .A2(n15289), .ZN(n10718) );
  NAND2_X1 U13970 ( .A1(n10719), .A2(n10718), .ZN(n15101) );
  INV_X1 U13971 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19656) );
  NAND2_X1 U13972 ( .A1(n10774), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10721) );
  NAND2_X1 U13973 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10720) );
  OAI211_X1 U13974 ( .C1(n19656), .C2(n9622), .A(n10721), .B(n10720), .ZN(
        n10722) );
  INV_X1 U13975 ( .A(n10722), .ZN(n10724) );
  INV_X1 U13976 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n20868) );
  OR2_X1 U13977 ( .A1(n10689), .A2(n20868), .ZN(n10723) );
  INV_X1 U13978 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n10807) );
  NAND2_X1 U13979 ( .A1(n10774), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10726) );
  NAND2_X1 U13980 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10725) );
  OAI211_X1 U13981 ( .C1(n10807), .C2(n9622), .A(n10726), .B(n10725), .ZN(
        n10727) );
  INV_X1 U13982 ( .A(n10727), .ZN(n10729) );
  INV_X1 U13983 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15275) );
  OR2_X1 U13984 ( .A1(n10689), .A2(n15275), .ZN(n10728) );
  INV_X1 U13985 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11158) );
  AOI22_X1 U13986 ( .A1(n12555), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10731) );
  INV_X1 U13987 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15259) );
  OR2_X1 U13988 ( .A1(n10689), .A2(n15259), .ZN(n10730) );
  OAI211_X1 U13989 ( .C1(n11158), .C2(n10675), .A(n10731), .B(n10730), .ZN(
        n14877) );
  INV_X1 U13990 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U13991 ( .A1(n10774), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10733) );
  NAND2_X1 U13992 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10732) );
  OAI211_X1 U13993 ( .C1(n9622), .C2(n11119), .A(n10733), .B(n10732), .ZN(
        n10734) );
  INV_X1 U13994 ( .A(n10734), .ZN(n10736) );
  INV_X1 U13995 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15636) );
  OR2_X1 U13996 ( .A1(n10689), .A2(n15636), .ZN(n10735) );
  AOI22_X1 U13997 ( .A1(n12555), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10738) );
  INV_X1 U13998 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15227) );
  OR2_X1 U13999 ( .A1(n10689), .A2(n15227), .ZN(n10737) );
  OAI211_X1 U14000 ( .C1(n10675), .C2(n9950), .A(n10738), .B(n10737), .ZN(
        n14818) );
  INV_X1 U14001 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15218) );
  AOI22_X1 U14002 ( .A1(n12555), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10740) );
  NAND2_X1 U14003 ( .A1(n10774), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10739) );
  OAI211_X1 U14004 ( .C1(n10689), .C2(n15218), .A(n10740), .B(n10739), .ZN(
        n14811) );
  INV_X1 U14005 ( .A(n14811), .ZN(n10741) );
  INV_X1 U14006 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11161) );
  AOI22_X1 U14007 ( .A1(n12555), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10743) );
  INV_X1 U14008 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15205) );
  OR2_X1 U14009 ( .A1(n10689), .A2(n15205), .ZN(n10742) );
  OAI211_X1 U14010 ( .C1(n11161), .C2(n10675), .A(n10743), .B(n10742), .ZN(
        n13213) );
  INV_X1 U14011 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n11127) );
  NAND2_X1 U14012 ( .A1(n10774), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10745) );
  NAND2_X1 U14013 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10744) );
  OAI211_X1 U14014 ( .C1(n9622), .C2(n11127), .A(n10745), .B(n10744), .ZN(
        n10746) );
  INV_X1 U14015 ( .A(n10746), .ZN(n10748) );
  INV_X1 U14016 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15195) );
  OR2_X1 U14017 ( .A1(n10689), .A2(n15195), .ZN(n10747) );
  NAND2_X1 U14018 ( .A1(n10748), .A2(n10747), .ZN(n14858) );
  INV_X1 U14019 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n14792) );
  NAND2_X1 U14020 ( .A1(n10774), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U14021 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10749) );
  OAI211_X1 U14022 ( .C1(n9622), .C2(n14792), .A(n10750), .B(n10749), .ZN(
        n10751) );
  INV_X1 U14023 ( .A(n10751), .ZN(n10753) );
  INV_X1 U14024 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15187) );
  OR2_X1 U14025 ( .A1(n10689), .A2(n15187), .ZN(n10752) );
  INV_X1 U14026 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11163) );
  INV_X1 U14027 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15166) );
  OR2_X1 U14028 ( .A1(n10689), .A2(n15166), .ZN(n10757) );
  INV_X1 U14029 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15016) );
  INV_X1 U14030 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n14021) );
  INV_X1 U14031 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10754) );
  OAI22_X1 U14032 ( .A1(n9622), .A2(n15016), .B1(n14021), .B2(n10754), .ZN(
        n10755) );
  INV_X1 U14033 ( .A(n10755), .ZN(n10756) );
  OAI211_X1 U14034 ( .C1(n10675), .C2(n11163), .A(n10757), .B(n10756), .ZN(
        n14847) );
  INV_X1 U14035 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19670) );
  NAND2_X1 U14036 ( .A1(n10774), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U14037 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10758) );
  OAI211_X1 U14038 ( .C1(n9622), .C2(n19670), .A(n10759), .B(n10758), .ZN(
        n10761) );
  INV_X1 U14039 ( .A(n10761), .ZN(n10763) );
  INV_X1 U14040 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n20763) );
  OR2_X1 U14041 ( .A1(n10689), .A2(n20763), .ZN(n10762) );
  AND2_X1 U14042 ( .A1(n10763), .A2(n10762), .ZN(n14775) );
  INV_X1 U14043 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19671) );
  NAND2_X1 U14044 ( .A1(n10774), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10765) );
  NAND2_X1 U14045 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10764) );
  OAI211_X1 U14046 ( .C1(n9622), .C2(n19671), .A(n10765), .B(n10764), .ZN(
        n10766) );
  INV_X1 U14047 ( .A(n10766), .ZN(n10768) );
  INV_X1 U14048 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12539) );
  OR2_X1 U14049 ( .A1(n10689), .A2(n12539), .ZN(n10767) );
  AND2_X1 U14050 ( .A1(n10768), .A2(n10767), .ZN(n12481) );
  INV_X1 U14051 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19673) );
  NAND2_X1 U14052 ( .A1(n10774), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U14053 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10769) );
  OAI211_X1 U14054 ( .C1(n9622), .C2(n19673), .A(n10770), .B(n10769), .ZN(
        n10771) );
  INV_X1 U14055 ( .A(n10771), .ZN(n10773) );
  INV_X1 U14056 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15128) );
  OR2_X1 U14057 ( .A1(n10689), .A2(n15128), .ZN(n10772) );
  NAND2_X1 U14058 ( .A1(n10773), .A2(n10772), .ZN(n14761) );
  NAND2_X1 U14059 ( .A1(n14762), .A2(n14761), .ZN(n14764) );
  INV_X1 U14060 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19676) );
  NAND2_X1 U14061 ( .A1(n10774), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U14062 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10775) );
  OAI211_X1 U14063 ( .C1(n9622), .C2(n19676), .A(n10776), .B(n10775), .ZN(
        n10777) );
  INV_X1 U14064 ( .A(n10777), .ZN(n10779) );
  INV_X1 U14065 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14201) );
  OR2_X1 U14066 ( .A1(n10689), .A2(n14201), .ZN(n10778) );
  AND2_X1 U14067 ( .A1(n10779), .A2(n10778), .ZN(n12554) );
  MUX2_X1 U14068 ( .A(n19719), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12746) );
  NAND2_X1 U14069 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19729), .ZN(
        n12297) );
  NOR2_X1 U14070 ( .A1(n12746), .A2(n10781), .ZN(n12436) );
  INV_X1 U14071 ( .A(n12436), .ZN(n10782) );
  NAND2_X1 U14072 ( .A1(n12746), .A2(n10781), .ZN(n10784) );
  NAND2_X1 U14073 ( .A1(n10782), .A2(n10784), .ZN(n12751) );
  NAND2_X1 U14074 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19719), .ZN(
        n10783) );
  NAND2_X1 U14075 ( .A1(n10784), .A2(n10783), .ZN(n10792) );
  NAND2_X1 U14076 ( .A1(n19710), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10787) );
  NAND2_X1 U14077 ( .A1(n10785), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10786) );
  NAND2_X1 U14078 ( .A1(n10792), .A2(n10793), .ZN(n10796) );
  NAND2_X1 U14079 ( .A1(n10796), .A2(n10787), .ZN(n10789) );
  XNOR2_X1 U14080 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10788) );
  AOI21_X1 U14081 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19704), .A(
        n10791), .ZN(n10799) );
  AND3_X1 U14082 ( .A1(n15561), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10799), .ZN(n11150) );
  NOR2_X1 U14083 ( .A1(n10789), .A2(n10788), .ZN(n10790) );
  OR2_X1 U14084 ( .A1(n10791), .A2(n10790), .ZN(n11143) );
  INV_X1 U14085 ( .A(n10792), .ZN(n10795) );
  INV_X1 U14086 ( .A(n10793), .ZN(n10794) );
  NAND2_X1 U14087 ( .A1(n10795), .A2(n10794), .ZN(n10797) );
  AND2_X1 U14088 ( .A1(n10797), .A2(n10796), .ZN(n12748) );
  NAND2_X1 U14089 ( .A1(n12758), .A2(n12748), .ZN(n12440) );
  NOR2_X1 U14090 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15625), .ZN(
        n10798) );
  INV_X1 U14091 ( .A(n12762), .ZN(n12438) );
  NAND2_X1 U14092 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14021), .ZN(n19612) );
  INV_X1 U14093 ( .A(n19612), .ZN(n10801) );
  NAND2_X1 U14094 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10801), .ZN(n16167) );
  NAND2_X1 U14095 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19747) );
  INV_X1 U14096 ( .A(n19747), .ZN(n19618) );
  NOR2_X1 U14097 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19618), .ZN(n10804) );
  INV_X1 U14098 ( .A(n10804), .ZN(n11175) );
  NOR2_X1 U14099 ( .A1(n19731), .A2(n11175), .ZN(n10802) );
  NAND2_X1 U14100 ( .A1(n13222), .A2(n13645), .ZN(n10803) );
  NAND2_X2 U14101 ( .A1(n19761), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19675) );
  INV_X1 U14102 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20756) );
  NAND2_X1 U14103 ( .A1(n20756), .A2(n19634), .ZN(n19628) );
  NAND2_X1 U14104 ( .A1(n19752), .A2(n10804), .ZN(n13673) );
  INV_X1 U14105 ( .A(n13673), .ZN(n10805) );
  AOI222_X1 U14106 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n12804), .B1(n10838), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .C1(n12803), .C2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n11141) );
  OR2_X1 U14107 ( .A1(n10846), .A2(n10807), .ZN(n10811) );
  OR2_X1 U14108 ( .A1(n10847), .A2(n15275), .ZN(n10810) );
  INV_X1 U14109 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n10808) );
  OR2_X1 U14110 ( .A1(n11140), .A2(n10808), .ZN(n10809) );
  INV_X1 U14111 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19517) );
  AND2_X2 U14112 ( .A1(n13146), .A2(n10547), .ZN(n13002) );
  AOI22_X1 U14113 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10819) );
  AND2_X2 U14114 ( .A1(n10812), .A2(n10547), .ZN(n10870) );
  AND2_X2 U14115 ( .A1(n10812), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10920) );
  AOI22_X1 U14116 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U14117 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10817) );
  INV_X1 U14118 ( .A(n10815), .ZN(n12984) );
  AND2_X2 U14119 ( .A1(n10815), .A2(n10547), .ZN(n13439) );
  AOI22_X1 U14120 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10816) );
  NAND4_X1 U14121 ( .A1(n10819), .A2(n10818), .A3(n10817), .A4(n10816), .ZN(
        n10833) );
  AND2_X2 U14122 ( .A1(n10820), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13007) );
  AND2_X2 U14123 ( .A1(n9602), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12969) );
  AOI22_X1 U14124 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10831) );
  AND2_X2 U14125 ( .A1(n13443), .A2(n10822), .ZN(n13008) );
  AOI22_X1 U14126 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10825) );
  NAND2_X1 U14127 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10824) );
  AND2_X1 U14128 ( .A1(n10825), .A2(n10824), .ZN(n10830) );
  AND2_X2 U14129 ( .A1(n10826), .A2(n13443), .ZN(n13012) );
  AND2_X2 U14130 ( .A1(n13443), .A2(n10827), .ZN(n13011) );
  AOI22_X1 U14131 ( .A1(n13012), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10829) );
  NAND2_X1 U14132 ( .A1(n13446), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12978) );
  NAND2_X1 U14133 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10828) );
  NAND4_X1 U14134 ( .A1(n10831), .A2(n10830), .A3(n10829), .A4(n10828), .ZN(
        n10832) );
  NAND2_X1 U14135 ( .A1(n10869), .A2(n12449), .ZN(n10836) );
  OAI22_X1 U14136 ( .A1(n13188), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19729), 
        .B2(n19700), .ZN(n10834) );
  INV_X1 U14137 ( .A(n10834), .ZN(n10835) );
  NAND2_X1 U14138 ( .A1(n10839), .A2(n10838), .ZN(n10886) );
  INV_X1 U14139 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18657) );
  INV_X1 U14140 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13370) );
  OAI21_X1 U14141 ( .B1(n10841), .B2(n13370), .A(n19700), .ZN(n10844) );
  INV_X1 U14142 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n10842) );
  NOR2_X1 U14143 ( .A1(n13188), .A2(n10842), .ZN(n10843) );
  NOR2_X1 U14144 ( .A1(n10844), .A2(n10843), .ZN(n10845) );
  OAI21_X1 U14145 ( .B1(n10846), .B2(n18657), .A(n10845), .ZN(n13336) );
  INV_X1 U14146 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19636) );
  NOR2_X1 U14147 ( .A1(n10846), .A2(n19636), .ZN(n10849) );
  INV_X1 U14148 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15446) );
  INV_X1 U14149 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18966) );
  OAI22_X1 U14150 ( .A1(n15446), .A2(n10847), .B1(n11140), .B2(n18966), .ZN(
        n10848) );
  OR2_X1 U14151 ( .A1(n10849), .A2(n10848), .ZN(n10868) );
  INV_X1 U14152 ( .A(n10868), .ZN(n10850) );
  AOI22_X1 U14153 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U14154 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13013), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U14155 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U14156 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10852) );
  NAND4_X1 U14157 ( .A1(n10855), .A2(n10854), .A3(n10853), .A4(n10852), .ZN(
        n10862) );
  AOI22_X1 U14158 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U14159 ( .A1(n13012), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U14160 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U14161 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10857) );
  NAND4_X1 U14162 ( .A1(n10860), .A2(n10859), .A3(n10858), .A4(n10857), .ZN(
        n10861) );
  NOR2_X1 U14163 ( .A1(n10862), .A2(n10861), .ZN(n12448) );
  INV_X1 U14164 ( .A(n10869), .ZN(n10863) );
  OR2_X1 U14165 ( .A1(n12448), .A2(n10863), .ZN(n10867) );
  AND2_X1 U14166 ( .A1(n13188), .A2(n19700), .ZN(n10865) );
  NOR2_X1 U14167 ( .A1(n19719), .A2(n19700), .ZN(n10864) );
  AOI21_X1 U14168 ( .B1(n13334), .B2(n10865), .A(n10864), .ZN(n10866) );
  AND2_X1 U14169 ( .A1(n10867), .A2(n10866), .ZN(n13430) );
  NAND2_X1 U14170 ( .A1(n13431), .A2(n13430), .ZN(n13429) );
  OR2_X1 U14171 ( .A1(n13339), .A2(n10868), .ZN(n10889) );
  AOI22_X1 U14172 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13002), .B1(
        n9618), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U14173 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U14174 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U14175 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10871) );
  NAND4_X1 U14176 ( .A1(n10874), .A2(n10873), .A3(n10872), .A4(n10871), .ZN(
        n10885) );
  AOI22_X1 U14177 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U14178 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10882) );
  INV_X1 U14179 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10878) );
  NAND2_X1 U14180 ( .A1(n13012), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10877) );
  NAND2_X1 U14181 ( .A1(n13011), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10876) );
  OAI211_X1 U14182 ( .C1(n12978), .C2(n10878), .A(n10877), .B(n10876), .ZN(
        n10879) );
  INV_X1 U14183 ( .A(n10879), .ZN(n10881) );
  NAND2_X1 U14184 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10880) );
  NAND4_X1 U14185 ( .A1(n10883), .A2(n10882), .A3(n10881), .A4(n10880), .ZN(
        n10884) );
  NAND2_X1 U14186 ( .A1(n10869), .A2(n11146), .ZN(n10887) );
  OAI211_X1 U14187 ( .C1(n19700), .C2(n19710), .A(n10887), .B(n10886), .ZN(
        n10888) );
  AND3_X1 U14188 ( .A1(n13429), .A2(n10889), .A3(n10888), .ZN(n10890) );
  NOR2_X1 U14189 ( .A1(n10846), .A2(n14224), .ZN(n10892) );
  INV_X1 U14190 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18964) );
  OAI22_X1 U14191 ( .A1(n12810), .A2(n10847), .B1(n11140), .B2(n18964), .ZN(
        n10891) );
  OR2_X1 U14192 ( .A1(n10892), .A2(n10891), .ZN(n13603) );
  INV_X1 U14193 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10913) );
  INV_X1 U14194 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n10894) );
  OR2_X1 U14195 ( .A1(n11140), .A2(n10894), .ZN(n10896) );
  NAND2_X1 U14196 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10895) );
  OAI211_X1 U14197 ( .C1(n10847), .C2(n16155), .A(n10896), .B(n10895), .ZN(
        n10897) );
  INV_X1 U14198 ( .A(n10897), .ZN(n10912) );
  AOI22_X1 U14199 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10851), .B1(
        n13007), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U14200 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10875), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U14201 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10898) );
  AND2_X1 U14202 ( .A1(n10899), .A2(n10898), .ZN(n10902) );
  AOI22_X1 U14203 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13012), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10901) );
  NAND2_X1 U14204 ( .A1(n10856), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10900) );
  NAND4_X1 U14205 ( .A1(n10903), .A2(n10902), .A3(n10901), .A4(n10900), .ZN(
        n10910) );
  AOI22_X1 U14206 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U14207 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n9619), .B1(
        n10904), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U14208 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13013), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U14209 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n13439), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10905) );
  NAND4_X1 U14210 ( .A1(n10908), .A2(n10907), .A3(n10906), .A4(n10905), .ZN(
        n10909) );
  NAND2_X1 U14211 ( .A1(n10869), .A2(n12227), .ZN(n10911) );
  OAI211_X1 U14212 ( .C1(n10846), .C2(n10913), .A(n10912), .B(n10911), .ZN(
        n13734) );
  AOI22_X1 U14213 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10851), .B1(
        n13007), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U14214 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10915) );
  NAND2_X1 U14215 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10914) );
  AND2_X1 U14216 ( .A1(n10915), .A2(n10914), .ZN(n10918) );
  AOI22_X1 U14217 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10917) );
  NAND2_X1 U14218 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10916) );
  NAND4_X1 U14219 ( .A1(n10919), .A2(n10918), .A3(n10917), .A4(n10916), .ZN(
        n10926) );
  AOI22_X1 U14220 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10920), .B1(
        n10904), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U14221 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13002), .B1(
        n9619), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U14222 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U14223 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13439), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10921) );
  NAND4_X1 U14224 ( .A1(n10924), .A2(n10923), .A3(n10922), .A4(n10921), .ZN(
        n10925) );
  NAND2_X1 U14225 ( .A1(n10869), .A2(n12229), .ZN(n10931) );
  INV_X1 U14226 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10927) );
  OR2_X1 U14227 ( .A1(n10846), .A2(n10927), .ZN(n10930) );
  OR2_X1 U14228 ( .A1(n10847), .A2(n13938), .ZN(n10929) );
  INV_X1 U14229 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n13783) );
  OR2_X1 U14230 ( .A1(n11140), .A2(n13783), .ZN(n10928) );
  AOI22_X1 U14231 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10851), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U14232 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10933) );
  NAND2_X1 U14233 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10932) );
  AND2_X1 U14234 ( .A1(n10933), .A2(n10932), .ZN(n10936) );
  AOI22_X1 U14235 ( .A1(n13012), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10935) );
  NAND2_X1 U14236 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10934) );
  NAND4_X1 U14237 ( .A1(n10937), .A2(n10936), .A3(n10935), .A4(n10934), .ZN(
        n10943) );
  AOI22_X1 U14238 ( .A1(n9619), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10870), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14239 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14240 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U14241 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10938) );
  NAND4_X1 U14242 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n10942) );
  NAND2_X1 U14243 ( .A1(n12244), .A2(n12403), .ZN(n11152) );
  INV_X1 U14244 ( .A(n11152), .ZN(n10944) );
  AOI22_X1 U14245 ( .A1(n12804), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n13342), 
        .B2(n10944), .ZN(n10946) );
  AOI22_X1 U14246 ( .A1(n10838), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n12803), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U14247 ( .A1(n10946), .A2(n10945), .ZN(n15432) );
  NAND2_X1 U14248 ( .A1(n15433), .A2(n15432), .ZN(n15431) );
  AOI22_X1 U14249 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13002), .B1(
        n10904), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U14250 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U14251 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U14252 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10947) );
  NAND4_X1 U14253 ( .A1(n10950), .A2(n10949), .A3(n10948), .A4(n10947), .ZN(
        n10958) );
  AOI22_X1 U14254 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U14255 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10952) );
  NAND2_X1 U14256 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10951) );
  AND2_X1 U14257 ( .A1(n10952), .A2(n10951), .ZN(n10955) );
  AOI22_X1 U14258 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10954) );
  NAND2_X1 U14259 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10953) );
  NAND4_X1 U14260 ( .A1(n10956), .A2(n10955), .A3(n10954), .A4(n10953), .ZN(
        n10957) );
  INV_X1 U14261 ( .A(n12269), .ZN(n10959) );
  NAND2_X1 U14262 ( .A1(n10869), .A2(n10959), .ZN(n10960) );
  INV_X1 U14263 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19641) );
  NOR2_X1 U14264 ( .A1(n10846), .A2(n19641), .ZN(n10962) );
  INV_X1 U14265 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18958) );
  OAI22_X1 U14266 ( .A1(n10847), .A2(n12828), .B1(n11140), .B2(n18958), .ZN(
        n10961) );
  NAND2_X1 U14267 ( .A1(n9619), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10967) );
  NAND2_X1 U14268 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10966) );
  NAND2_X1 U14269 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10965) );
  NAND2_X1 U14270 ( .A1(n10856), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10964) );
  NAND2_X1 U14271 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10971) );
  NAND2_X1 U14272 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10970) );
  NAND2_X1 U14273 ( .A1(n10920), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10969) );
  NAND2_X1 U14274 ( .A1(n13439), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10968) );
  AOI22_X1 U14275 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U14276 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U14277 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U14278 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10973) );
  NAND2_X1 U14279 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10972) );
  AND4_X2 U14280 ( .A1(n10979), .A2(n10978), .A3(n10977), .A4(n10976), .ZN(
        n12280) );
  AOI21_X1 U14281 ( .B1(n13360), .B2(n13359), .A(n10079), .ZN(n10980) );
  INV_X1 U14282 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19643) );
  NOR2_X1 U14283 ( .A1(n10846), .A2(n19643), .ZN(n10982) );
  INV_X1 U14284 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18956) );
  OAI22_X1 U14285 ( .A1(n9839), .A2(n10847), .B1(n11140), .B2(n18956), .ZN(
        n10981) );
  NAND2_X1 U14286 ( .A1(n10920), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10986) );
  NAND2_X1 U14287 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10985) );
  NAND2_X1 U14288 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10984) );
  NAND2_X1 U14289 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10983) );
  AND4_X1 U14290 ( .A1(n10986), .A2(n10985), .A3(n10984), .A4(n10983), .ZN(
        n10997) );
  NAND2_X1 U14291 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10990) );
  NAND2_X1 U14292 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10989) );
  NAND2_X1 U14293 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10988) );
  NAND2_X1 U14294 ( .A1(n13439), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10987) );
  AND4_X1 U14295 ( .A1(n10990), .A2(n10989), .A3(n10988), .A4(n10987), .ZN(
        n10996) );
  AOI22_X1 U14296 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U14297 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14298 ( .A1(n13012), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10993) );
  NAND2_X1 U14299 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10992) );
  NAND2_X1 U14300 ( .A1(n10856), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10991) );
  NAND4_X1 U14301 ( .A1(n10997), .A2(n10996), .A3(n10995), .A4(n10075), .ZN(
        n13550) );
  NAND2_X1 U14302 ( .A1(n10869), .A2(n13550), .ZN(n11003) );
  INV_X1 U14303 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10998) );
  OR2_X1 U14304 ( .A1(n10846), .A2(n10998), .ZN(n11002) );
  OR2_X1 U14305 ( .A1(n10847), .A2(n14181), .ZN(n11001) );
  INV_X1 U14306 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n10999) );
  OR2_X1 U14307 ( .A1(n11140), .A2(n10999), .ZN(n11000) );
  AOI22_X1 U14308 ( .A1(n12804), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n12803), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U14309 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11007) );
  AOI22_X1 U14310 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U14311 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U14312 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11004) );
  NAND4_X1 U14313 ( .A1(n11007), .A2(n11006), .A3(n11005), .A4(n11004), .ZN(
        n11015) );
  AOI22_X1 U14314 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14315 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U14316 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11008) );
  AND2_X1 U14317 ( .A1(n11009), .A2(n11008), .ZN(n11012) );
  AOI22_X1 U14318 ( .A1(n13012), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U14319 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11010) );
  NAND4_X1 U14320 ( .A1(n11013), .A2(n11012), .A3(n11011), .A4(n11010), .ZN(
        n11014) );
  AOI22_X1 U14321 ( .A1(n10869), .A2(n18891), .B1(n10838), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11016) );
  NAND2_X1 U14322 ( .A1(n11017), .A2(n11016), .ZN(n13416) );
  AOI22_X1 U14323 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10851), .B1(
        n13007), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U14324 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11019) );
  NAND2_X1 U14325 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11018) );
  AND2_X1 U14326 ( .A1(n11019), .A2(n11018), .ZN(n11022) );
  AOI22_X1 U14327 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11021) );
  NAND2_X1 U14328 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11020) );
  NAND4_X1 U14329 ( .A1(n11023), .A2(n11022), .A3(n11021), .A4(n11020), .ZN(
        n11029) );
  AOI22_X1 U14330 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13002), .B1(
        n9619), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14331 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U14332 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U14333 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n13439), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11024) );
  NAND4_X1 U14334 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n11028) );
  NAND2_X1 U14335 ( .A1(n10869), .A2(n18890), .ZN(n11035) );
  OR2_X1 U14336 ( .A1(n10846), .A2(n11030), .ZN(n11034) );
  OR2_X1 U14337 ( .A1(n10847), .A2(n15393), .ZN(n11033) );
  INV_X1 U14338 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n11031) );
  OR2_X1 U14339 ( .A1(n11140), .A2(n11031), .ZN(n11032) );
  AOI22_X1 U14340 ( .A1(n12804), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n12803), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U14341 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13002), .B1(
        n10904), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U14342 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U14343 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U14344 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11036) );
  NAND4_X1 U14345 ( .A1(n11039), .A2(n11038), .A3(n11037), .A4(n11036), .ZN(
        n11047) );
  AOI22_X1 U14346 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U14347 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11041) );
  NAND2_X1 U14348 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11040) );
  AND2_X1 U14349 ( .A1(n11041), .A2(n11040), .ZN(n11044) );
  AOI22_X1 U14350 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U14351 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11042) );
  NAND4_X1 U14352 ( .A1(n11045), .A2(n11044), .A3(n11043), .A4(n11042), .ZN(
        n11046) );
  AOI22_X1 U14353 ( .A1(n10869), .A2(n18884), .B1(n10838), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11048) );
  NAND2_X1 U14354 ( .A1(n11049), .A2(n11048), .ZN(n13536) );
  NAND2_X1 U14355 ( .A1(n13537), .A2(n13536), .ZN(n13535) );
  AOI22_X1 U14356 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10851), .B1(
        n13007), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14357 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10875), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11051) );
  NAND2_X1 U14358 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11050) );
  AND2_X1 U14359 ( .A1(n11051), .A2(n11050), .ZN(n11054) );
  AOI22_X1 U14360 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13012), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U14361 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11052) );
  NAND4_X1 U14362 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11061) );
  AOI22_X1 U14363 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13002), .B1(
        n9619), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14364 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10870), .B1(
        n10904), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14365 ( .A1(n10920), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14366 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13439), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11056) );
  NAND4_X1 U14367 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n11060) );
  AOI22_X1 U14368 ( .A1(n10838), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12803), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n11062) );
  OAI21_X1 U14369 ( .B1(n10846), .B2(n13908), .A(n11062), .ZN(n11063) );
  AOI21_X1 U14370 ( .B1(n10869), .B2(n18883), .A(n11063), .ZN(n13677) );
  AOI22_X1 U14371 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14372 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14373 ( .A1(n9619), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14374 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11064) );
  NAND4_X1 U14375 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n11075) );
  AOI22_X1 U14376 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U14377 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11069) );
  NAND2_X1 U14378 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11068) );
  AND2_X1 U14379 ( .A1(n11069), .A2(n11068), .ZN(n11072) );
  AOI22_X1 U14380 ( .A1(n13012), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11071) );
  NAND2_X1 U14381 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11070) );
  NAND4_X1 U14382 ( .A1(n11073), .A2(n11072), .A3(n11071), .A4(n11070), .ZN(
        n11074) );
  AOI22_X1 U14383 ( .A1(n12804), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n10869), 
        .B2(n13813), .ZN(n11077) );
  AOI22_X1 U14384 ( .A1(n10838), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n12803), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U14385 ( .A1(n11077), .A2(n11076), .ZN(n13730) );
  NAND2_X1 U14386 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11081) );
  NAND2_X1 U14387 ( .A1(n9619), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11080) );
  NAND2_X1 U14388 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11079) );
  NAND2_X1 U14389 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11078) );
  AND4_X1 U14390 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n11093) );
  NAND2_X1 U14391 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11085) );
  NAND2_X1 U14392 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11084) );
  NAND2_X1 U14393 ( .A1(n10920), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11083) );
  NAND2_X1 U14394 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11082) );
  AND4_X1 U14395 ( .A1(n11085), .A2(n11084), .A3(n11083), .A4(n11082), .ZN(
        n11092) );
  AOI22_X1 U14396 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U14397 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10875), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14398 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13012), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11088) );
  NAND2_X1 U14399 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11087) );
  NAND2_X1 U14400 ( .A1(n10856), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11086) );
  AND4_X1 U14401 ( .A1(n11089), .A2(n11088), .A3(n11087), .A4(n11086), .ZN(
        n11090) );
  NAND4_X1 U14402 ( .A1(n11093), .A2(n11092), .A3(n11091), .A4(n11090), .ZN(
        n13817) );
  AOI22_X1 U14403 ( .A1(n10838), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n12803), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11094) );
  OAI21_X1 U14404 ( .B1(n10846), .B2(n11095), .A(n11094), .ZN(n11096) );
  AOI21_X1 U14405 ( .B1(n10869), .B2(n13817), .A(n11096), .ZN(n16118) );
  AOI22_X1 U14406 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13002), .B1(
        n10904), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U14407 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14408 ( .A1(n9619), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14409 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11097) );
  NAND4_X1 U14410 ( .A1(n11100), .A2(n11099), .A3(n11098), .A4(n11097), .ZN(
        n11108) );
  AOI22_X1 U14411 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14412 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U14413 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11101) );
  AND2_X1 U14414 ( .A1(n11102), .A2(n11101), .ZN(n11105) );
  AOI22_X1 U14415 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11104) );
  NAND2_X1 U14416 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11103) );
  NAND4_X1 U14417 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n11107) );
  NOR2_X1 U14418 ( .A1(n11108), .A2(n11107), .ZN(n13925) );
  AOI22_X1 U14419 ( .A1(n12804), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n10869), 
        .B2(n10022), .ZN(n11110) );
  AOI22_X1 U14420 ( .A1(n10838), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12803), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11109) );
  NAND2_X1 U14421 ( .A1(n11110), .A2(n11109), .ZN(n13811) );
  NOR2_X1 U14422 ( .A1(n10846), .A2(n11111), .ZN(n11114) );
  INV_X1 U14423 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n11112) );
  OAI22_X1 U14424 ( .A1(n10847), .A2(n15289), .B1(n11140), .B2(n11112), .ZN(
        n11113) );
  NOR2_X1 U14425 ( .A1(n11114), .A2(n11113), .ZN(n15304) );
  NOR2_X1 U14426 ( .A1(n10846), .A2(n19656), .ZN(n11116) );
  INV_X1 U14427 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14972) );
  OAI22_X1 U14428 ( .A1(n10847), .A2(n20868), .B1(n11140), .B2(n14972), .ZN(
        n11115) );
  INV_X1 U14429 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20834) );
  NOR2_X1 U14430 ( .A1(n10846), .A2(n20834), .ZN(n11118) );
  INV_X1 U14431 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14960) );
  OAI22_X1 U14432 ( .A1(n10847), .A2(n15259), .B1(n11140), .B2(n14960), .ZN(
        n11117) );
  OR2_X1 U14433 ( .A1(n10846), .A2(n11119), .ZN(n11122) );
  OR2_X1 U14434 ( .A1(n10847), .A2(n15636), .ZN(n11121) );
  INV_X1 U14435 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n20719) );
  OR2_X1 U14436 ( .A1(n11140), .A2(n20719), .ZN(n11120) );
  INV_X1 U14437 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19661) );
  NOR2_X1 U14438 ( .A1(n10846), .A2(n19661), .ZN(n11124) );
  INV_X1 U14439 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n20852) );
  OAI22_X1 U14440 ( .A1(n10847), .A2(n15227), .B1(n11140), .B2(n20852), .ZN(
        n11123) );
  OR2_X1 U14441 ( .A1(n11124), .A2(n11123), .ZN(n14819) );
  AOI222_X1 U14442 ( .A1(n12804), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n10838), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C1(n12803), .C2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n14808) );
  INV_X1 U14443 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n11126) );
  INV_X1 U14444 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n11125) );
  OAI222_X1 U14445 ( .A1(n11126), .A2(n11140), .B1(n11125), .B2(n10846), .C1(
        n10847), .C2(n15205), .ZN(n13217) );
  NOR2_X1 U14446 ( .A1(n10846), .A2(n11127), .ZN(n11130) );
  INV_X1 U14447 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n11128) );
  OAI22_X1 U14448 ( .A1(n15195), .A2(n10847), .B1(n11140), .B2(n11128), .ZN(
        n11129) );
  OR2_X1 U14449 ( .A1(n11130), .A2(n11129), .ZN(n14932) );
  NOR2_X1 U14450 ( .A1(n10846), .A2(n14792), .ZN(n11132) );
  INV_X1 U14451 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14922) );
  OAI22_X1 U14452 ( .A1(n15187), .A2(n10847), .B1(n11140), .B2(n14922), .ZN(
        n11131) );
  OR2_X1 U14453 ( .A1(n11132), .A2(n11131), .ZN(n14791) );
  NOR2_X1 U14454 ( .A1(n10846), .A2(n15016), .ZN(n11135) );
  INV_X1 U14455 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n11133) );
  OAI22_X1 U14456 ( .A1(n15166), .A2(n10847), .B1(n11140), .B2(n11133), .ZN(
        n11134) );
  OR2_X1 U14457 ( .A1(n11135), .A2(n11134), .ZN(n14909) );
  NOR2_X1 U14458 ( .A1(n10846), .A2(n19670), .ZN(n11137) );
  INV_X1 U14459 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14902) );
  OAI22_X1 U14460 ( .A1(n20763), .A2(n10847), .B1(n11140), .B2(n14902), .ZN(
        n11136) );
  OR2_X1 U14461 ( .A1(n11137), .A2(n11136), .ZN(n14776) );
  NOR2_X1 U14462 ( .A1(n10846), .A2(n19671), .ZN(n11139) );
  INV_X1 U14463 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n20796) );
  OAI22_X1 U14464 ( .A1(n12539), .A2(n10847), .B1(n11140), .B2(n20796), .ZN(
        n11138) );
  NOR2_X1 U14465 ( .A1(n11139), .A2(n11138), .ZN(n14892) );
  INV_X1 U14466 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14885) );
  OAI222_X1 U14467 ( .A1(n19673), .A2(n10846), .B1(n10847), .B2(n15128), .C1(
        n11140), .C2(n14885), .ZN(n14766) );
  AOI21_X1 U14468 ( .B1(n11141), .B2(n14765), .A(n12806), .ZN(n14203) );
  AOI22_X1 U14469 ( .A1(n14983), .A2(n18840), .B1(n18863), .B2(n14203), .ZN(
        n11180) );
  INV_X1 U14470 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13376) );
  INV_X1 U14471 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13372) );
  NAND2_X1 U14472 ( .A1(n13376), .A2(n13372), .ZN(n11142) );
  MUX2_X1 U14473 ( .A(n12448), .B(n11142), .S(n19061), .Z(n12296) );
  OR2_X1 U14474 ( .A1(n19731), .A2(n19061), .ZN(n12302) );
  AND2_X1 U14475 ( .A1(n19731), .A2(n12808), .ZN(n12298) );
  NAND2_X1 U14476 ( .A1(n12298), .A2(n11143), .ZN(n11145) );
  NAND2_X1 U14477 ( .A1(n19061), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11144) );
  OAI211_X1 U14478 ( .C1(n12302), .C2(n12227), .A(n11145), .B(n11144), .ZN(
        n12291) );
  INV_X1 U14479 ( .A(n11146), .ZN(n12210) );
  INV_X1 U14480 ( .A(n12748), .ZN(n11147) );
  INV_X1 U14481 ( .A(n12293), .ZN(n11148) );
  OAI22_X1 U14482 ( .A1(n12302), .A2(n12445), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n12403), .ZN(n11151) );
  OAI21_X1 U14483 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n12808), .A(n11152), .ZN(
        n12281) );
  MUX2_X1 U14484 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12269), .S(n12808), .Z(
        n11153) );
  INV_X1 U14485 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13602) );
  MUX2_X1 U14486 ( .A(n13602), .B(n12548), .S(n12403), .Z(n12317) );
  NAND2_X1 U14487 ( .A1(n12319), .A2(n12317), .ZN(n12315) );
  NAND2_X1 U14488 ( .A1(n12330), .A2(n10701), .ZN(n12340) );
  NAND2_X1 U14489 ( .A1(n19061), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12339) );
  NAND2_X1 U14490 ( .A1(n19061), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12367) );
  INV_X1 U14491 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13826) );
  INV_X1 U14492 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n18724) );
  NAND2_X1 U14493 ( .A1(n13826), .A2(n18724), .ZN(n11155) );
  NAND2_X1 U14494 ( .A1(n19061), .A2(n11155), .ZN(n11156) );
  OAI21_X1 U14495 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(P2_EBX_REG_16__SCAN_IN), 
        .A(n19061), .ZN(n11157) );
  AND2_X2 U14496 ( .A1(n12360), .A2(n11157), .ZN(n12373) );
  NAND2_X1 U14497 ( .A1(n19061), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12365) );
  NOR2_X1 U14498 ( .A1(n12403), .A2(n11158), .ZN(n12362) );
  INV_X1 U14499 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U14500 ( .A1(n9653), .A2(n12411), .ZN(n11160) );
  NAND2_X1 U14501 ( .A1(n19061), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12394) );
  NAND2_X1 U14502 ( .A1(n11160), .A2(n12394), .ZN(n12400) );
  NOR2_X1 U14503 ( .A1(n12808), .A2(n11161), .ZN(n12399) );
  INV_X1 U14504 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11162) );
  NAND2_X1 U14505 ( .A1(n12415), .A2(n11163), .ZN(n12418) );
  INV_X1 U14506 ( .A(n12547), .ZN(n11165) );
  NAND2_X1 U14507 ( .A1(n19061), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11164) );
  INV_X1 U14508 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11166) );
  NOR2_X1 U14509 ( .A1(n12808), .A2(n11166), .ZN(n12429) );
  OR2_X2 U14510 ( .A1(n12430), .A2(n12429), .ZN(n12432) );
  INV_X2 U14511 ( .A(n12432), .ZN(n12541) );
  NAND2_X1 U14512 ( .A1(n19061), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12540) );
  NAND2_X1 U14513 ( .A1(n12541), .A2(n12540), .ZN(n12545) );
  NAND2_X1 U14514 ( .A1(n19061), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11167) );
  XNOR2_X1 U14515 ( .A(n12545), .B(n11167), .ZN(n12542) );
  INV_X1 U14516 ( .A(n12542), .ZN(n12543) );
  NAND2_X1 U14517 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n11175), .ZN(n11168) );
  NOR2_X1 U14518 ( .A1(n19731), .A2(n11168), .ZN(n11169) );
  NOR2_X1 U14519 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19693) );
  NOR2_X1 U14520 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11170) );
  NAND2_X1 U14521 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19549), .ZN(n19083) );
  NOR2_X1 U14522 ( .A1(n19612), .A2(n19083), .ZN(n16157) );
  INV_X1 U14523 ( .A(n16157), .ZN(n11171) );
  NAND3_X1 U14524 ( .A1(n18877), .A2(n18772), .A3(n11171), .ZN(n11172) );
  INV_X2 U14525 ( .A(n18832), .ZN(n18874) );
  AOI22_X1 U14526 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n18867), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18874), .ZN(n11173) );
  OAI21_X1 U14527 ( .B1(n12543), .B2(n18852), .A(n11173), .ZN(n11174) );
  INV_X1 U14528 ( .A(n11174), .ZN(n11179) );
  AND2_X1 U14529 ( .A1(n18974), .A2(n13673), .ZN(n15959) );
  INV_X1 U14530 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12557) );
  NAND2_X1 U14531 ( .A1(n12557), .A2(n11175), .ZN(n11176) );
  NOR2_X1 U14532 ( .A1(n13233), .A2(n11176), .ZN(n11177) );
  OR2_X2 U14533 ( .A1(n15959), .A2(n11177), .ZN(n18866) );
  NAND2_X1 U14534 ( .A1(n18866), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11178) );
  INV_X1 U14535 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14536 ( .A1(n11502), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11503), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11190) );
  AND2_X2 U14537 ( .A1(n11194), .A2(n11192), .ZN(n11523) );
  AOI22_X1 U14538 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11523), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14539 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11264), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14540 ( .A1(n11272), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11361), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11187) );
  AND2_X2 U14541 ( .A1(n11195), .A2(n11193), .ZN(n11250) );
  AOI22_X1 U14542 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14139), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11199) );
  AND2_X2 U14543 ( .A1(n11195), .A2(n11192), .ZN(n11360) );
  AND2_X2 U14544 ( .A1(n13479), .A2(n11194), .ZN(n11391) );
  AOI22_X1 U14545 ( .A1(n11360), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9630), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14546 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11197) );
  AND2_X4 U14547 ( .A1(n13479), .A2(n13475), .ZN(n11496) );
  AOI22_X1 U14548 ( .A1(n11271), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14549 ( .A1(n11502), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11503), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14550 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11523), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14551 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11264), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14552 ( .A1(n11272), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14553 ( .A1(n11271), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14554 ( .A1(n11360), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9630), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14555 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11206) );
  AOI22_X1 U14556 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14139), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11205) );
  INV_X1 U14557 ( .A(n11320), .ZN(n11383) );
  NAND2_X1 U14558 ( .A1(n11360), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11212) );
  NAND2_X1 U14559 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11211) );
  NAND2_X1 U14560 ( .A1(n11271), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11210) );
  NAND2_X1 U14561 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11209) );
  NAND2_X1 U14562 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11216) );
  NAND2_X1 U14563 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11215) );
  NAND2_X1 U14564 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11214) );
  NAND2_X1 U14565 ( .A1(n14139), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11213) );
  NAND2_X1 U14566 ( .A1(n11502), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11220) );
  NAND2_X1 U14567 ( .A1(n11503), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11219) );
  NAND2_X1 U14568 ( .A1(n11361), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11218) );
  NAND2_X1 U14569 ( .A1(n11272), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11217) );
  NAND2_X1 U14570 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11224) );
  NAND2_X1 U14571 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14572 ( .A1(n11523), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11222) );
  NAND2_X1 U14573 ( .A1(n11264), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11221) );
  AOI22_X1 U14574 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11523), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14575 ( .A1(n11502), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14576 ( .A1(n11503), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14577 ( .A1(n11271), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14578 ( .A1(n11272), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9623), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11233) );
  NAND2_X1 U14579 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11241) );
  NAND2_X1 U14580 ( .A1(n11503), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11240) );
  NAND2_X1 U14581 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11239) );
  NAND2_X1 U14582 ( .A1(n11523), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11238) );
  NAND2_X1 U14583 ( .A1(n11502), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11245) );
  NAND2_X1 U14584 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11244) );
  NAND2_X1 U14585 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11243) );
  NAND2_X1 U14586 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11242) );
  NAND2_X1 U14587 ( .A1(n11360), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11249) );
  NAND2_X1 U14588 ( .A1(n9630), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11248) );
  NAND2_X1 U14589 ( .A1(n11272), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11247) );
  NAND2_X1 U14590 ( .A1(n11264), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11246) );
  NAND2_X1 U14591 ( .A1(n11271), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11254) );
  NAND2_X1 U14592 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11253) );
  NAND2_X1 U14593 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11252) );
  NAND2_X1 U14594 ( .A1(n14139), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11251) );
  AND2_X2 U14595 ( .A1(n11383), .A2(n11259), .ZN(n14240) );
  AOI22_X1 U14596 ( .A1(n11360), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9630), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U14597 ( .A1(n11271), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U14598 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14599 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14139), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14600 ( .A1(n11502), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11503), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14601 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11523), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U14602 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14603 ( .A1(n11272), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11361), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14604 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11503), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11276) );
  AOI22_X1 U14605 ( .A1(n11271), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11250), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U14606 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14607 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11272), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11273) );
  NAND4_X1 U14608 ( .A1(n11276), .A2(n11275), .A3(n11274), .A4(n11273), .ZN(
        n11282) );
  AOI22_X1 U14609 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11523), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14610 ( .A1(n11502), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11264), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U14611 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14139), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11278) );
  AOI22_X1 U14612 ( .A1(n11360), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11277) );
  NAND4_X1 U14613 ( .A1(n11280), .A2(n11279), .A3(n11278), .A4(n11277), .ZN(
        n11281) );
  NAND2_X2 U14614 ( .A1(n14240), .A2(n13489), .ZN(n12700) );
  INV_X1 U14615 ( .A(n12700), .ZN(n11304) );
  NAND2_X1 U14616 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11287) );
  NAND2_X1 U14617 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11286) );
  NAND2_X1 U14618 ( .A1(n11523), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11285) );
  NAND2_X1 U14619 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11284) );
  NAND2_X1 U14620 ( .A1(n11360), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11291) );
  NAND2_X1 U14621 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11290) );
  NAND2_X1 U14622 ( .A1(n11271), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11289) );
  NAND2_X1 U14623 ( .A1(n11496), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11288) );
  AND4_X2 U14624 ( .A1(n11291), .A2(n11290), .A3(n11289), .A4(n11288), .ZN(
        n11302) );
  NAND2_X1 U14625 ( .A1(n11502), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11295) );
  NAND2_X1 U14626 ( .A1(n11503), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11294) );
  NAND2_X1 U14627 ( .A1(n11361), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11293) );
  NAND2_X1 U14628 ( .A1(n11272), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11292) );
  NAND2_X1 U14629 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11299) );
  NAND2_X1 U14630 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11298) );
  NAND2_X1 U14631 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11297) );
  NAND2_X1 U14632 ( .A1(n14139), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11296) );
  NAND4_X4 U14633 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n20025) );
  NAND2_X1 U14634 ( .A1(n11304), .A2(n20025), .ZN(n12591) );
  INV_X1 U14635 ( .A(n12591), .ZN(n11307) );
  XNOR2_X1 U14636 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12574) );
  OAI21_X1 U14637 ( .B1(n12700), .B2(n12574), .A(n12701), .ZN(n11306) );
  NOR2_X1 U14638 ( .A1(n11307), .A2(n11306), .ZN(n11318) );
  INV_X2 U14639 ( .A(n11308), .ZN(n11682) );
  INV_X1 U14640 ( .A(n11340), .ZN(n11316) );
  NAND2_X2 U14641 ( .A1(n11309), .A2(n20040), .ZN(n11321) );
  AOI21_X2 U14642 ( .B1(n11321), .B2(n20029), .A(n14166), .ZN(n11315) );
  NAND2_X1 U14643 ( .A1(n12580), .A2(n20040), .ZN(n11312) );
  OAI21_X1 U14644 ( .B1(n11312), .B2(n11682), .A(n11311), .ZN(n11313) );
  INV_X1 U14645 ( .A(n11313), .ZN(n11314) );
  NAND2_X1 U14646 ( .A1(n11318), .A2(n12592), .ZN(n11319) );
  OAI21_X1 U14647 ( .B1(n11317), .B2(n13557), .A(n20012), .ZN(n11330) );
  NAND2_X2 U14648 ( .A1(n11340), .A2(n20025), .ZN(n12623) );
  NAND2_X1 U14649 ( .A1(n20012), .A2(n20025), .ZN(n14257) );
  NAND2_X1 U14650 ( .A1(n12709), .A2(n14257), .ZN(n11323) );
  OR2_X1 U14651 ( .A1(n20012), .A2(n20025), .ZN(n14258) );
  INV_X1 U14652 ( .A(n20012), .ZN(n13399) );
  NAND2_X1 U14653 ( .A1(n13399), .A2(n20029), .ZN(n11322) );
  OAI211_X1 U14654 ( .C1(n14258), .C2(n13409), .A(n13467), .B(n11322), .ZN(
        n11347) );
  NOR2_X1 U14655 ( .A1(n11323), .A2(n11347), .ZN(n11329) );
  NAND2_X1 U14656 ( .A1(n12584), .A2(n13409), .ZN(n11324) );
  INV_X1 U14657 ( .A(n12704), .ZN(n11326) );
  NAND2_X1 U14658 ( .A1(n12586), .A2(n14742), .ZN(n11328) );
  NAND3_X1 U14659 ( .A1(n11330), .A2(n11329), .A3(n11328), .ZN(n12718) );
  NAND2_X1 U14660 ( .A1(n12718), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U14661 ( .A1(n11419), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11334) );
  NAND2_X1 U14662 ( .A1(n15945), .A2(n20702), .ZN(n12149) );
  NAND2_X1 U14663 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11421) );
  OAI21_X1 U14664 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11421), .ZN(n20348) );
  NAND2_X1 U14665 ( .A1(n20582), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11416) );
  OAI21_X1 U14666 ( .B1(n12149), .B2(n20348), .A(n11416), .ZN(n11332) );
  INV_X1 U14667 ( .A(n11332), .ZN(n11333) );
  NAND2_X1 U14668 ( .A1(n11334), .A2(n11333), .ZN(n11336) );
  NAND2_X1 U14669 ( .A1(n11419), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11339) );
  INV_X1 U14670 ( .A(n20582), .ZN(n11337) );
  MUX2_X1 U14671 ( .A(n11337), .B(n12149), .S(n20446), .Z(n11338) );
  NAND3_X1 U14672 ( .A1(n12586), .A2(n20025), .A3(n14742), .ZN(n11351) );
  INV_X1 U14673 ( .A(n14251), .ZN(n13421) );
  NAND3_X1 U14674 ( .A1(n13421), .A2(n11341), .A3(n11340), .ZN(n11342) );
  NAND2_X1 U14675 ( .A1(n11317), .A2(n11342), .ZN(n11350) );
  INV_X1 U14676 ( .A(n14258), .ZN(n20701) );
  INV_X1 U14677 ( .A(n11343), .ZN(n11344) );
  NAND2_X1 U14678 ( .A1(n20701), .A2(n11344), .ZN(n11346) );
  NAND2_X1 U14679 ( .A1(n15945), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19766) );
  INV_X1 U14680 ( .A(n19766), .ZN(n11345) );
  NAND2_X1 U14681 ( .A1(n13557), .A2(n11682), .ZN(n12714) );
  NAND4_X1 U14682 ( .A1(n11346), .A2(n11345), .A3(n12714), .A4(n14257), .ZN(
        n11348) );
  NOR2_X1 U14683 ( .A1(n11348), .A2(n11347), .ZN(n11349) );
  NAND3_X1 U14684 ( .A1(n11351), .A2(n11350), .A3(n11349), .ZN(n11388) );
  INV_X1 U14685 ( .A(n11353), .ZN(n11354) );
  INV_X1 U14686 ( .A(n11473), .ZN(n11449) );
  AOI22_X1 U14687 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14688 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11355), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14689 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14690 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11523), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11356) );
  NAND4_X1 U14691 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11367) );
  AOI22_X1 U14692 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14693 ( .A1(n12058), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14694 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14695 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11362) );
  NAND4_X1 U14696 ( .A1(n11365), .A2(n11364), .A3(n11363), .A4(n11362), .ZN(
        n11366) );
  NAND2_X1 U14697 ( .A1(n11449), .A2(n11447), .ZN(n11368) );
  INV_X1 U14698 ( .A(n11369), .ZN(n11674) );
  NAND2_X1 U14699 ( .A1(n11674), .A2(n20025), .ZN(n11387) );
  AOI22_X1 U14700 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12131), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14702 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14703 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14704 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11372) );
  NAND4_X1 U14705 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n11382) );
  AOI22_X1 U14706 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14707 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11523), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14708 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14709 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11377) );
  NAND4_X1 U14710 ( .A1(n11380), .A2(n11379), .A3(n11378), .A4(n11377), .ZN(
        n11381) );
  NAND2_X1 U14711 ( .A1(n11447), .A2(n11409), .ZN(n11492) );
  OAI21_X1 U14712 ( .B1(n11447), .B2(n11409), .A(n11492), .ZN(n11384) );
  OAI211_X1 U14713 ( .C1(n11384), .C2(n14258), .A(n11383), .B(n20040), .ZN(
        n11385) );
  INV_X1 U14714 ( .A(n11385), .ZN(n11386) );
  INV_X1 U14715 ( .A(n11388), .ZN(n11389) );
  INV_X1 U14716 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11404) );
  AOI21_X1 U14717 ( .B1(n20012), .B2(n11409), .A(n20702), .ZN(n11403) );
  AOI22_X1 U14718 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9631), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14719 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14720 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14721 ( .A1(n11250), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11393) );
  NAND4_X1 U14722 ( .A1(n11396), .A2(n11395), .A3(n11394), .A4(n11393), .ZN(
        n11402) );
  AOI22_X1 U14723 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14724 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11523), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14725 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14726 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11397) );
  NAND4_X1 U14727 ( .A1(n11400), .A2(n11399), .A3(n11398), .A4(n11397), .ZN(
        n11401) );
  NAND2_X1 U14728 ( .A1(n13409), .A2(n11581), .ZN(n11446) );
  OAI211_X1 U14729 ( .C1(n11652), .C2(n11404), .A(n11403), .B(n11446), .ZN(
        n11445) );
  INV_X1 U14730 ( .A(n11581), .ZN(n11592) );
  NAND2_X1 U14731 ( .A1(n11592), .A2(n13409), .ZN(n11405) );
  MUX2_X1 U14732 ( .A(n11446), .B(n11405), .S(n11409), .Z(n11406) );
  INV_X1 U14733 ( .A(n11406), .ZN(n11407) );
  NAND2_X1 U14734 ( .A1(n11407), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U14735 ( .A1(n20012), .A2(n11340), .ZN(n11461) );
  OAI21_X1 U14736 ( .B1(n14258), .B2(n11409), .A(n11461), .ZN(n11410) );
  INV_X1 U14737 ( .A(n11410), .ZN(n11411) );
  OAI21_X1 U14738 ( .B1(n11681), .B2(n11623), .A(n11411), .ZN(n13349) );
  NAND2_X1 U14739 ( .A1(n13349), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11412) );
  NAND2_X1 U14740 ( .A1(n19941), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19940) );
  INV_X1 U14741 ( .A(n11412), .ZN(n11414) );
  NAND2_X1 U14742 ( .A1(n11414), .A2(n11413), .ZN(n11415) );
  INV_X1 U14743 ( .A(n11335), .ZN(n11418) );
  NAND2_X1 U14744 ( .A1(n11416), .A2(n11186), .ZN(n11417) );
  NAND2_X1 U14745 ( .A1(n11418), .A2(n11417), .ZN(n11427) );
  NAND2_X1 U14746 ( .A1(n11429), .A2(n11427), .ZN(n11425) );
  NAND2_X1 U14747 ( .A1(n9610), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11424) );
  INV_X1 U14748 ( .A(n11421), .ZN(n11420) );
  NAND2_X1 U14749 ( .A1(n11420), .A2(n20681), .ZN(n20375) );
  NAND2_X1 U14750 ( .A1(n11421), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11422) );
  NAND2_X1 U14751 ( .A1(n20375), .A2(n11422), .ZN(n20019) );
  INV_X1 U14752 ( .A(n12149), .ZN(n11470) );
  AOI22_X1 U14753 ( .A1(n20019), .A2(n11470), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20582), .ZN(n11423) );
  INV_X1 U14754 ( .A(n11426), .ZN(n11428) );
  NAND3_X1 U14755 ( .A1(n11429), .A2(n11428), .A3(n11427), .ZN(n11430) );
  NAND2_X1 U14756 ( .A1(n11468), .A2(n11430), .ZN(n13554) );
  AOI22_X1 U14757 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14758 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14759 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14760 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11431) );
  NAND4_X1 U14761 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(
        n11440) );
  AOI22_X1 U14762 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14763 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14764 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14765 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11435) );
  NAND4_X1 U14766 ( .A1(n11438), .A2(n11437), .A3(n11436), .A4(n11435), .ZN(
        n11439) );
  OAI22_X2 U14767 ( .A1(n13554), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11491), 
        .B2(n11473), .ZN(n11443) );
  INV_X1 U14768 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U14769 ( .A1(n20012), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11474) );
  OAI22_X1 U14770 ( .A1(n11652), .A2(n11441), .B1(n11474), .B2(n11491), .ZN(
        n11442) );
  XNOR2_X1 U14771 ( .A(n11443), .B(n11442), .ZN(n11459) );
  INV_X1 U14772 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11452) );
  INV_X1 U14773 ( .A(n11447), .ZN(n11448) );
  OR2_X1 U14774 ( .A1(n11448), .A2(n11474), .ZN(n11451) );
  NAND2_X1 U14775 ( .A1(n11449), .A2(n11592), .ZN(n11450) );
  OAI211_X1 U14776 ( .C1(n11652), .C2(n11452), .A(n11451), .B(n11450), .ZN(
        n11454) );
  INV_X1 U14777 ( .A(n11454), .ZN(n11453) );
  NAND2_X1 U14778 ( .A1(n11673), .A2(n11674), .ZN(n11457) );
  NAND2_X1 U14779 ( .A1(n11457), .A2(n11456), .ZN(n11458) );
  OR2_X2 U14780 ( .A1(n11459), .A2(n11458), .ZN(n11489) );
  NAND2_X1 U14781 ( .A1(n11459), .A2(n11458), .ZN(n11460) );
  NAND2_X1 U14782 ( .A1(n11489), .A2(n11460), .ZN(n20009) );
  OR2_X1 U14783 ( .A1(n20009), .A2(n11623), .ZN(n11465) );
  XNOR2_X1 U14784 ( .A(n11492), .B(n11491), .ZN(n11463) );
  INV_X1 U14785 ( .A(n11461), .ZN(n11462) );
  AOI21_X1 U14786 ( .B1(n11463), .B2(n20701), .A(n11462), .ZN(n11464) );
  NAND2_X1 U14787 ( .A1(n11466), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11467) );
  INV_X1 U14788 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12614) );
  INV_X1 U14789 ( .A(n11489), .ZN(n11487) );
  NAND2_X1 U14790 ( .A1(n9610), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11472) );
  NOR3_X1 U14791 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20681), .A3(
        n20690), .ZN(n20266) );
  INV_X1 U14792 ( .A(n20266), .ZN(n20261) );
  NAND3_X1 U14793 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20473) );
  INV_X1 U14794 ( .A(n20473), .ZN(n20529) );
  NAND2_X1 U14795 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20529), .ZN(
        n20518) );
  OAI21_X1 U14796 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20283), .A(
        n20518), .ZN(n20290) );
  INV_X1 U14797 ( .A(n20290), .ZN(n11469) );
  AOI22_X1 U14798 ( .A1(n11470), .A2(n11469), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20582), .ZN(n11471) );
  AOI22_X1 U14799 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14800 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14801 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14802 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11475) );
  NAND4_X1 U14803 ( .A1(n11478), .A2(n11477), .A3(n11476), .A4(n11475), .ZN(
        n11484) );
  AOI22_X1 U14804 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14805 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14806 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14807 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U14808 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11483) );
  AOI22_X1 U14809 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11656), .B1(
        n11634), .B2(n11542), .ZN(n11485) );
  NAND2_X1 U14810 ( .A1(n11489), .A2(n20158), .ZN(n11490) );
  NAND2_X1 U14811 ( .A1(n11492), .A2(n11491), .ZN(n11544) );
  XNOR2_X1 U14812 ( .A(n11544), .B(n11542), .ZN(n11493) );
  OAI22_X1 U14813 ( .A1(n11701), .A2(n11623), .B1(n14258), .B2(n11493), .ZN(
        n13768) );
  NAND2_X1 U14814 ( .A1(n11656), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11511) );
  AOI22_X1 U14815 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14816 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14817 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11370), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14818 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11988), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11498) );
  NAND4_X1 U14819 ( .A1(n11501), .A2(n11500), .A3(n11499), .A4(n11498), .ZN(
        n11509) );
  AOI22_X1 U14820 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14821 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12130), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14822 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n14144), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14823 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11504) );
  NAND4_X1 U14824 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n11508) );
  NAND2_X1 U14825 ( .A1(n11634), .A2(n11541), .ZN(n11510) );
  NAND2_X1 U14826 ( .A1(n11511), .A2(n11510), .ZN(n11534) );
  INV_X1 U14827 ( .A(n11623), .ZN(n11577) );
  NAND2_X1 U14828 ( .A1(n11716), .A2(n11577), .ZN(n11515) );
  NAND2_X1 U14829 ( .A1(n11544), .A2(n11542), .ZN(n11512) );
  XNOR2_X1 U14830 ( .A(n11512), .B(n11541), .ZN(n11513) );
  NAND2_X1 U14831 ( .A1(n11513), .A2(n20701), .ZN(n11514) );
  NAND2_X1 U14832 ( .A1(n11515), .A2(n11514), .ZN(n11517) );
  INV_X1 U14833 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11516) );
  XNOR2_X1 U14834 ( .A(n11517), .B(n11516), .ZN(n19930) );
  NAND2_X1 U14835 ( .A1(n11517), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11518) );
  INV_X1 U14836 ( .A(n11538), .ZN(n11533) );
  NAND2_X1 U14837 ( .A1(n11656), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11531) );
  AOI22_X1 U14838 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14839 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14840 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14841 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11519) );
  NAND4_X1 U14842 ( .A1(n11522), .A2(n11521), .A3(n11520), .A4(n11519), .ZN(
        n11529) );
  AOI22_X1 U14843 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14844 ( .A1(n12058), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14845 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14846 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11524) );
  NAND4_X1 U14847 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n11528) );
  NAND2_X1 U14848 ( .A1(n11634), .A2(n11566), .ZN(n11530) );
  NAND2_X1 U14849 ( .A1(n11531), .A2(n11530), .ZN(n11535) );
  INV_X1 U14850 ( .A(n11534), .ZN(n11537) );
  INV_X1 U14851 ( .A(n11535), .ZN(n11536) );
  OAI21_X1 U14852 ( .B1(n11538), .B2(n11537), .A(n11536), .ZN(n11539) );
  INV_X1 U14853 ( .A(n11706), .ZN(n11540) );
  OR2_X1 U14854 ( .A1(n11540), .A2(n11623), .ZN(n11547) );
  AND2_X1 U14855 ( .A1(n11542), .A2(n11541), .ZN(n11543) );
  NAND2_X1 U14856 ( .A1(n11544), .A2(n11543), .ZN(n11568) );
  XNOR2_X1 U14857 ( .A(n11568), .B(n11566), .ZN(n11545) );
  NAND2_X1 U14858 ( .A1(n11545), .A2(n20701), .ZN(n11546) );
  NAND2_X1 U14859 ( .A1(n11547), .A2(n11546), .ZN(n11548) );
  INV_X1 U14860 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20804) );
  XNOR2_X1 U14861 ( .A(n11548), .B(n20804), .ZN(n13834) );
  NAND2_X1 U14862 ( .A1(n11548), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11549) );
  INV_X1 U14863 ( .A(n11565), .ZN(n11563) );
  NAND2_X1 U14864 ( .A1(n11656), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11561) );
  AOI22_X1 U14865 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14866 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14867 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14868 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11550) );
  NAND4_X1 U14869 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11559) );
  AOI22_X1 U14870 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14871 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14872 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14873 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11554) );
  NAND4_X1 U14874 ( .A1(n11557), .A2(n11556), .A3(n11555), .A4(n11554), .ZN(
        n11558) );
  NAND2_X1 U14875 ( .A1(n11634), .A2(n11579), .ZN(n11560) );
  NAND2_X1 U14876 ( .A1(n11565), .A2(n11564), .ZN(n11724) );
  NAND3_X1 U14877 ( .A1(n11591), .A2(n11724), .A3(n11577), .ZN(n11571) );
  INV_X1 U14878 ( .A(n11566), .ZN(n11567) );
  OR2_X1 U14879 ( .A1(n11568), .A2(n11567), .ZN(n11578) );
  XNOR2_X1 U14880 ( .A(n11578), .B(n11579), .ZN(n11569) );
  NAND2_X1 U14881 ( .A1(n11569), .A2(n20701), .ZN(n11570) );
  NAND2_X1 U14882 ( .A1(n11571), .A2(n11570), .ZN(n11572) );
  XNOR2_X1 U14883 ( .A(n11572), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15864) );
  OR2_X1 U14884 ( .A1(n11572), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11573) );
  INV_X1 U14885 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11575) );
  NAND2_X1 U14886 ( .A1(n11634), .A2(n11581), .ZN(n11574) );
  OAI21_X1 U14887 ( .B1(n11575), .B2(n11652), .A(n11574), .ZN(n11576) );
  NAND2_X1 U14888 ( .A1(n11725), .A2(n11577), .ZN(n11584) );
  INV_X1 U14889 ( .A(n11578), .ZN(n11580) );
  NAND2_X1 U14890 ( .A1(n11580), .A2(n11579), .ZN(n11593) );
  XNOR2_X1 U14891 ( .A(n11593), .B(n11581), .ZN(n11582) );
  NAND2_X1 U14892 ( .A1(n11582), .A2(n20701), .ZN(n11583) );
  NAND2_X1 U14893 ( .A1(n11584), .A2(n11583), .ZN(n11586) );
  INV_X1 U14894 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11585) );
  XNOR2_X1 U14895 ( .A(n11586), .B(n11585), .ZN(n15861) );
  NAND2_X1 U14896 ( .A1(n15860), .A2(n15861), .ZN(n11588) );
  OR2_X1 U14897 ( .A1(n11586), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11587) );
  NOR2_X1 U14898 ( .A1(n11589), .A2(n11623), .ZN(n11590) );
  OR3_X1 U14899 ( .A1(n11593), .A2(n11592), .A3(n14258), .ZN(n11594) );
  NAND2_X1 U14900 ( .A1(n14539), .A2(n11594), .ZN(n14011) );
  NOR2_X1 U14901 ( .A1(n14011), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11596) );
  NAND2_X1 U14902 ( .A1(n14011), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11595) );
  INV_X1 U14903 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15911) );
  INV_X1 U14904 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14711) );
  NAND2_X1 U14905 ( .A1(n14539), .A2(n14711), .ZN(n11597) );
  NAND2_X1 U14906 ( .A1(n14700), .A2(n11597), .ZN(n14561) );
  INV_X1 U14907 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20856) );
  NAND2_X1 U14908 ( .A1(n14705), .A2(n20856), .ZN(n14560) );
  NAND2_X1 U14909 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11598) );
  NAND2_X1 U14910 ( .A1(n14539), .A2(n11598), .ZN(n14555) );
  NAND2_X1 U14911 ( .A1(n14560), .A2(n14555), .ZN(n11599) );
  OR2_X1 U14912 ( .A1(n14539), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14541) );
  NAND2_X1 U14913 ( .A1(n14539), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U14914 ( .A1(n14541), .A2(n11600), .ZN(n15833) );
  INV_X1 U14915 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15895) );
  NAND2_X1 U14916 ( .A1(n14539), .A2(n15895), .ZN(n11601) );
  INV_X1 U14917 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14704) );
  NAND2_X1 U14918 ( .A1(n14539), .A2(n14704), .ZN(n14536) );
  NAND2_X1 U14919 ( .A1(n14705), .A2(n14682), .ZN(n11602) );
  NAND4_X1 U14920 ( .A1(n14702), .A2(n14540), .A3(n14536), .A4(n11602), .ZN(
        n11607) );
  OR2_X1 U14921 ( .A1(n14539), .A2(n20856), .ZN(n14559) );
  NOR2_X1 U14922 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11603) );
  OR2_X1 U14923 ( .A1(n14539), .A2(n11603), .ZN(n14557) );
  OR2_X1 U14924 ( .A1(n14539), .A2(n14704), .ZN(n11604) );
  NAND2_X1 U14925 ( .A1(n15895), .A2(n9765), .ZN(n15834) );
  OAI21_X1 U14926 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15834), .A(
        n9634), .ZN(n11605) );
  XNOR2_X1 U14927 ( .A(n14705), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15825) );
  NAND2_X1 U14928 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11609) );
  INV_X1 U14929 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12720) );
  NAND2_X1 U14930 ( .A1(n14663), .A2(n12720), .ZN(n11610) );
  NOR2_X2 U14931 ( .A1(n15826), .A2(n11610), .ZN(n14651) );
  INV_X1 U14932 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14668) );
  INV_X1 U14933 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11611) );
  NAND2_X1 U14934 ( .A1(n9669), .A2(n11611), .ZN(n11612) );
  NAND2_X1 U14935 ( .A1(n11612), .A2(n9634), .ZN(n15811) );
  INV_X1 U14936 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14621) );
  INV_X1 U14937 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U14938 ( .A1(n14621), .A2(n14512), .ZN(n11613) );
  INV_X1 U14939 ( .A(n11618), .ZN(n11615) );
  INV_X1 U14940 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11616) );
  NAND2_X1 U14941 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12734) );
  NOR2_X1 U14942 ( .A1(n12734), .A2(n14621), .ZN(n12729) );
  NAND2_X1 U14943 ( .A1(n11618), .A2(n12729), .ZN(n14482) );
  NAND2_X1 U14944 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12736) );
  XNOR2_X1 U14945 ( .A(n9634), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11619) );
  XNOR2_X1 U14946 ( .A(n12567), .B(n11619), .ZN(n14594) );
  XNOR2_X1 U14947 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11633) );
  NAND2_X1 U14948 ( .A1(n20446), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11636) );
  NAND2_X1 U14949 ( .A1(n11633), .A2(n11632), .ZN(n11621) );
  NAND2_X1 U14950 ( .A1(n20690), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11620) );
  XNOR2_X1 U14951 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11629) );
  INV_X1 U14952 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20004) );
  NOR2_X1 U14953 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20004), .ZN(
        n11622) );
  NAND2_X1 U14954 ( .A1(n12573), .A2(n11655), .ZN(n11664) );
  NAND2_X1 U14955 ( .A1(n12573), .A2(n11634), .ZN(n11662) );
  NAND3_X1 U14956 ( .A1(n15947), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n11624), .ZN(n12571) );
  INV_X1 U14957 ( .A(n11655), .ZN(n11659) );
  AOI21_X1 U14958 ( .B1(n11627), .B2(n11626), .A(n11625), .ZN(n11628) );
  INV_X1 U14959 ( .A(n11628), .ZN(n12568) );
  XNOR2_X1 U14960 ( .A(n11630), .B(n11629), .ZN(n12569) );
  INV_X1 U14961 ( .A(n11634), .ZN(n11651) );
  OR2_X1 U14962 ( .A1(n20040), .A2(n20012), .ZN(n11631) );
  NAND2_X1 U14963 ( .A1(n11631), .A2(n12599), .ZN(n11650) );
  XNOR2_X1 U14964 ( .A(n11633), .B(n11632), .ZN(n12570) );
  AOI22_X1 U14965 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14239), .B1(n11634), 
        .B2(n20025), .ZN(n11645) );
  INV_X1 U14966 ( .A(n11645), .ZN(n11635) );
  NOR2_X1 U14967 ( .A1(n12570), .A2(n11635), .ZN(n11641) );
  OAI21_X1 U14968 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20446), .A(
        n11636), .ZN(n11637) );
  NOR2_X1 U14969 ( .A1(n11651), .A2(n11637), .ZN(n11640) );
  INV_X1 U14970 ( .A(n11637), .ZN(n11638) );
  OAI211_X1 U14971 ( .C1(n20012), .C2(n11321), .A(n11638), .B(n11650), .ZN(
        n11639) );
  OAI21_X1 U14972 ( .B1(n11655), .B2(n11640), .A(n11639), .ZN(n11642) );
  AND2_X1 U14973 ( .A1(n11641), .A2(n11642), .ZN(n11649) );
  INV_X1 U14974 ( .A(n12570), .ZN(n11644) );
  NOR2_X1 U14975 ( .A1(n11645), .A2(n11642), .ZN(n11643) );
  AOI211_X1 U14976 ( .C1(n11645), .C2(n20025), .A(n11644), .B(n11643), .ZN(
        n11648) );
  OAI21_X1 U14977 ( .B1(n11651), .B2(n12569), .A(n11650), .ZN(n11646) );
  AOI21_X1 U14978 ( .B1(n11656), .B2(n12569), .A(n11646), .ZN(n11647) );
  OAI33_X1 U14979 ( .A1(n12569), .A2(n11651), .A3(n11650), .B1(n11649), .B2(
        n11648), .B3(n11647), .ZN(n11654) );
  NAND2_X1 U14980 ( .A1(n11652), .A2(n12568), .ZN(n11653) );
  AOI22_X1 U14981 ( .A1(n11655), .A2(n12568), .B1(n11654), .B2(n11653), .ZN(
        n11658) );
  NOR2_X1 U14982 ( .A1(n11656), .A2(n12571), .ZN(n11657) );
  OAI22_X1 U14983 ( .A1(n12571), .A2(n11659), .B1(n11658), .B2(n11657), .ZN(
        n11660) );
  AOI21_X1 U14984 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20702), .A(
        n11660), .ZN(n11661) );
  NAND2_X1 U14985 ( .A1(n11662), .A2(n11661), .ZN(n11663) );
  NOR2_X1 U14986 ( .A1(n12704), .A2(n11320), .ZN(n11666) );
  NAND2_X1 U14987 ( .A1(n14742), .A2(n20012), .ZN(n11665) );
  NAND2_X1 U14988 ( .A1(n11666), .A2(n11665), .ZN(n13417) );
  NOR2_X1 U14989 ( .A1(n13417), .A2(n11321), .ZN(n11667) );
  OR2_X2 U14990 ( .A1(n14594), .A2(n19943), .ZN(n12155) );
  INV_X1 U14991 ( .A(n11856), .ZN(n11811) );
  NAND2_X1 U14992 ( .A1(n13425), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11709) );
  XNOR2_X1 U14993 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13513) );
  AOI21_X1 U14994 ( .B1(n14157), .B2(n13513), .A(n14163), .ZN(n11669) );
  NAND2_X1 U14995 ( .A1(n14164), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11668) );
  OAI211_X1 U14996 ( .C1(n11709), .C2(n11185), .A(n11669), .B(n11668), .ZN(
        n11670) );
  INV_X1 U14997 ( .A(n11670), .ZN(n11671) );
  NAND2_X1 U14998 ( .A1(n14163), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11692) );
  NAND2_X1 U14999 ( .A1(n11672), .A2(n11692), .ZN(n13501) );
  INV_X1 U15000 ( .A(n13501), .ZN(n11691) );
  XNOR2_X2 U15001 ( .A(n11675), .B(n11369), .ZN(n20010) );
  NAND2_X1 U15002 ( .A1(n20010), .A2(n11856), .ZN(n11680) );
  AOI22_X1 U15003 ( .A1(n14164), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20700), .ZN(n11678) );
  INV_X1 U15004 ( .A(n11709), .ZN(n11676) );
  NAND2_X1 U15005 ( .A1(n11676), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11677) );
  AND2_X1 U15006 ( .A1(n11678), .A2(n11677), .ZN(n11679) );
  NAND2_X1 U15007 ( .A1(n11681), .A2(n11682), .ZN(n11683) );
  NAND2_X1 U15008 ( .A1(n11683), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13352) );
  NAND2_X1 U15009 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20700), .ZN(
        n11687) );
  NAND2_X1 U15010 ( .A1(n11685), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11686) );
  OAI211_X1 U15011 ( .C1(n11709), .C2(n11183), .A(n11687), .B(n11686), .ZN(
        n11688) );
  AOI21_X1 U15012 ( .B1(n11684), .B2(n11856), .A(n11688), .ZN(n13353) );
  OR2_X1 U15013 ( .A1(n13352), .A2(n13353), .ZN(n13350) );
  NAND2_X1 U15014 ( .A1(n13353), .A2(n14157), .ZN(n11689) );
  NAND2_X1 U15015 ( .A1(n13350), .A2(n11689), .ZN(n13414) );
  NAND2_X1 U15016 ( .A1(n11691), .A2(n11690), .ZN(n13503) );
  INV_X1 U15017 ( .A(n11694), .ZN(n11693) );
  INV_X1 U15018 ( .A(n11712), .ZN(n11696) );
  INV_X1 U15019 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13856) );
  NAND2_X1 U15020 ( .A1(n13856), .A2(n11694), .ZN(n11695) );
  NAND2_X1 U15021 ( .A1(n11696), .A2(n11695), .ZN(n13855) );
  AOI22_X1 U15022 ( .A1(n13855), .A2(n14157), .B1(n14163), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11698) );
  NAND2_X1 U15023 ( .A1(n14164), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11697) );
  OAI211_X1 U15024 ( .C1(n11709), .C2(n11184), .A(n11698), .B(n11697), .ZN(
        n11699) );
  INV_X1 U15025 ( .A(n11699), .ZN(n11700) );
  NAND2_X1 U15026 ( .A1(n13587), .A2(n13586), .ZN(n13584) );
  INV_X1 U15027 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11704) );
  AND2_X1 U15028 ( .A1(n11711), .A2(n19812), .ZN(n11702) );
  OR2_X1 U15029 ( .A1(n11702), .A2(n11720), .ZN(n19819) );
  AOI22_X1 U15030 ( .A1(n19819), .A2(n14157), .B1(n14163), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11703) );
  OAI21_X1 U15031 ( .B1(n12112), .B2(n11704), .A(n11703), .ZN(n11705) );
  INV_X1 U15032 ( .A(n13751), .ZN(n11718) );
  NAND2_X1 U15033 ( .A1(n20700), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11708) );
  NAND2_X1 U15034 ( .A1(n14164), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11707) );
  OAI211_X1 U15035 ( .C1(n11709), .C2(n15947), .A(n11708), .B(n11707), .ZN(
        n11710) );
  NAND2_X1 U15036 ( .A1(n11710), .A2(n12120), .ZN(n11714) );
  OAI21_X1 U15037 ( .B1(n11712), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11711), .ZN(n19938) );
  NAND2_X1 U15038 ( .A1(n19938), .A2(n14157), .ZN(n11713) );
  NAND2_X1 U15039 ( .A1(n11714), .A2(n11713), .ZN(n11715) );
  INV_X1 U15040 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13847) );
  OR2_X1 U15041 ( .A1(n11720), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U15042 ( .A1(n11726), .A2(n11721), .ZN(n19805) );
  AOI22_X1 U15043 ( .A1(n19805), .A2(n14157), .B1(n14163), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11722) );
  OAI21_X1 U15044 ( .B1(n12112), .B2(n13847), .A(n11722), .ZN(n11723) );
  NOR2_X2 U15045 ( .A1(n13750), .A2(n13844), .ZN(n13863) );
  NAND2_X1 U15046 ( .A1(n11725), .A2(n11856), .ZN(n11732) );
  INV_X1 U15047 ( .A(n14163), .ZN(n11893) );
  NAND2_X1 U15048 ( .A1(n11726), .A2(n11729), .ZN(n11727) );
  NAND2_X1 U15049 ( .A1(n11748), .A2(n11727), .ZN(n19797) );
  NAND2_X1 U15050 ( .A1(n19797), .A2(n14157), .ZN(n11728) );
  OAI21_X1 U15051 ( .B1(n11729), .B2(n11893), .A(n11728), .ZN(n11730) );
  AOI21_X1 U15052 ( .B1(n14164), .B2(P1_EAX_REG_7__SCAN_IN), .A(n11730), .ZN(
        n11731) );
  NAND2_X1 U15053 ( .A1(n11732), .A2(n11731), .ZN(n13862) );
  NAND2_X1 U15054 ( .A1(n13863), .A2(n13862), .ZN(n13864) );
  AOI22_X1 U15055 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U15056 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U15057 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U15058 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11733) );
  NAND4_X1 U15059 ( .A1(n11736), .A2(n11735), .A3(n11734), .A4(n11733), .ZN(
        n11742) );
  AOI22_X1 U15060 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U15061 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U15062 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U15063 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11737) );
  NAND4_X1 U15064 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n11741) );
  OAI21_X1 U15065 ( .B1(n11742), .B2(n11741), .A(n11856), .ZN(n11746) );
  NAND2_X1 U15066 ( .A1(n14164), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11745) );
  XNOR2_X1 U15067 ( .A(n11748), .B(n13879), .ZN(n14013) );
  NAND2_X1 U15068 ( .A1(n14013), .A2(n14157), .ZN(n11744) );
  NAND2_X1 U15069 ( .A1(n14163), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11743) );
  NAND4_X1 U15070 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n13870) );
  INV_X1 U15071 ( .A(n13870), .ZN(n11747) );
  XNOR2_X1 U15072 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11765), .ZN(
        n14035) );
  INV_X1 U15073 ( .A(n14035), .ZN(n11763) );
  AOI22_X1 U15074 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U15075 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U15076 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U15077 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11749) );
  NAND4_X1 U15078 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n11758) );
  AOI22_X1 U15079 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U15080 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U15081 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U15082 ( .A1(n12058), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11753) );
  NAND4_X1 U15083 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n11753), .ZN(
        n11757) );
  OAI21_X1 U15084 ( .B1(n11758), .B2(n11757), .A(n11856), .ZN(n11761) );
  NAND2_X1 U15085 ( .A1(n14164), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U15086 ( .A1(n14163), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11759) );
  NAND3_X1 U15087 ( .A1(n11761), .A2(n11760), .A3(n11759), .ZN(n11762) );
  AOI21_X1 U15088 ( .B1(n11763), .B2(n14157), .A(n11762), .ZN(n13915) );
  XNOR2_X1 U15089 ( .A(n11782), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14574) );
  NAND2_X1 U15090 ( .A1(n14574), .A2(n14157), .ZN(n11781) );
  AOI22_X1 U15091 ( .A1(n11766), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U15092 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U15093 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U15094 ( .A1(n12058), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11767) );
  NAND4_X1 U15095 ( .A1(n11770), .A2(n11769), .A3(n11768), .A4(n11767), .ZN(
        n11776) );
  AOI22_X1 U15096 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U15097 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U15098 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U15099 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11771) );
  NAND4_X1 U15100 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n11775) );
  OAI21_X1 U15101 ( .B1(n11776), .B2(n11775), .A(n11856), .ZN(n11779) );
  NAND2_X1 U15102 ( .A1(n11685), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11778) );
  NAND2_X1 U15103 ( .A1(n14163), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11777) );
  AND3_X1 U15104 ( .A1(n11779), .A2(n11778), .A3(n11777), .ZN(n11780) );
  NAND2_X1 U15105 ( .A1(n11781), .A2(n11780), .ZN(n13985) );
  NAND2_X1 U15106 ( .A1(n11685), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11785) );
  OAI21_X1 U15107 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11783), .A(
        n11823), .ZN(n15859) );
  AOI22_X1 U15108 ( .A1(n14157), .A2(n15859), .B1(n14163), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11784) );
  NAND2_X1 U15109 ( .A1(n11785), .A2(n11784), .ZN(n14062) );
  AOI22_X1 U15110 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U15111 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U15112 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U15113 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11786) );
  NAND4_X1 U15114 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11795) );
  AOI22_X1 U15115 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U15116 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U15117 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U15118 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11790) );
  NAND4_X1 U15119 ( .A1(n11793), .A2(n11792), .A3(n11791), .A4(n11790), .ZN(
        n11794) );
  OR2_X1 U15120 ( .A1(n11795), .A2(n11794), .ZN(n11796) );
  NAND2_X1 U15121 ( .A1(n13982), .A2(n14078), .ZN(n11797) );
  NAND2_X1 U15122 ( .A1(n14061), .A2(n11797), .ZN(n11828) );
  AOI22_X1 U15123 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11355), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U15124 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U15125 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U15126 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11798) );
  NAND4_X1 U15127 ( .A1(n11801), .A2(n11800), .A3(n11799), .A4(n11798), .ZN(
        n11807) );
  AOI22_X1 U15128 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11988), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U15129 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U15130 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U15131 ( .A1(n14145), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11802) );
  NAND4_X1 U15132 ( .A1(n11805), .A2(n11804), .A3(n11803), .A4(n11802), .ZN(
        n11806) );
  NOR2_X1 U15133 ( .A1(n11807), .A2(n11806), .ZN(n11812) );
  XNOR2_X1 U15134 ( .A(n11829), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14564) );
  NAND2_X1 U15135 ( .A1(n14564), .A2(n14157), .ZN(n11810) );
  AOI22_X1 U15136 ( .A1(n11685), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n14163), 
        .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11809) );
  OAI211_X1 U15137 ( .C1(n11812), .C2(n11811), .A(n11810), .B(n11809), .ZN(
        n14083) );
  INV_X1 U15138 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U15139 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n14144), .B1(
        n12130), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U15140 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12131), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U15141 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11988), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U15142 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11813) );
  NAND4_X1 U15143 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n11822) );
  AOI22_X1 U15144 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U15145 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11370), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U15146 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U15147 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11371), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11817) );
  NAND4_X1 U15148 ( .A1(n11820), .A2(n11819), .A3(n11818), .A4(n11817), .ZN(
        n11821) );
  OAI21_X1 U15149 ( .B1(n11822), .B2(n11821), .A(n11856), .ZN(n11826) );
  XNOR2_X1 U15150 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11823), .ZN(
        n15848) );
  OAI22_X1 U15151 ( .A1(n15848), .A2(n12120), .B1(n11893), .B2(n11808), .ZN(
        n11824) );
  INV_X1 U15152 ( .A(n11824), .ZN(n11825) );
  OAI211_X1 U15153 ( .C1(n12112), .C2(n14081), .A(n11826), .B(n11825), .ZN(
        n14067) );
  NAND2_X1 U15154 ( .A1(n11828), .A2(n11827), .ZN(n14051) );
  INV_X1 U15155 ( .A(n14051), .ZN(n11846) );
  XOR2_X1 U15156 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11847), .Z(
        n15842) );
  INV_X1 U15157 ( .A(n15842), .ZN(n11844) );
  AOI22_X1 U15158 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U15159 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U15160 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U15161 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11830) );
  NAND4_X1 U15162 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n11839) );
  AOI22_X1 U15163 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U15164 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U15165 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U15166 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11834) );
  NAND4_X1 U15167 ( .A1(n11837), .A2(n11836), .A3(n11835), .A4(n11834), .ZN(
        n11838) );
  OAI21_X1 U15168 ( .B1(n11839), .B2(n11838), .A(n11856), .ZN(n11842) );
  NAND2_X1 U15169 ( .A1(n11685), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11841) );
  NAND2_X1 U15170 ( .A1(n14163), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11840) );
  NAND3_X1 U15171 ( .A1(n11842), .A2(n11841), .A3(n11840), .ZN(n11843) );
  AOI21_X1 U15172 ( .B1(n11844), .B2(n14157), .A(n11843), .ZN(n14055) );
  NAND2_X1 U15173 ( .A1(n11846), .A2(n11845), .ZN(n14053) );
  XNOR2_X1 U15174 ( .A(n11865), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15756) );
  INV_X1 U15175 ( .A(n15756), .ZN(n14551) );
  AOI22_X1 U15176 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12131), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U15177 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U15178 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U15179 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11848) );
  NAND4_X1 U15180 ( .A1(n11851), .A2(n11850), .A3(n11849), .A4(n11848), .ZN(
        n11858) );
  AOI22_X1 U15181 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U15182 ( .A1(n14145), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U15183 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U15184 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11852) );
  NAND4_X1 U15185 ( .A1(n11855), .A2(n11854), .A3(n11853), .A4(n11852), .ZN(
        n11857) );
  OAI21_X1 U15186 ( .B1(n11858), .B2(n11857), .A(n11856), .ZN(n11861) );
  NAND2_X1 U15187 ( .A1(n14164), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U15188 ( .A1(n14163), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11859) );
  NAND3_X1 U15189 ( .A1(n11861), .A2(n11860), .A3(n11859), .ZN(n11862) );
  AOI21_X1 U15190 ( .B1(n14551), .B2(n14157), .A(n11862), .ZN(n14109) );
  OR2_X1 U15191 ( .A1(n11866), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11867) );
  NAND2_X1 U15192 ( .A1(n11867), .A2(n11911), .ZN(n15841) );
  AOI22_X1 U15193 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U15194 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U15195 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U15196 ( .A1(n14145), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11868) );
  NAND4_X1 U15197 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11877) );
  AOI22_X1 U15198 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U15199 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U15200 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U15201 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U15202 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11876) );
  NOR2_X1 U15203 ( .A1(n11877), .A2(n11876), .ZN(n11880) );
  OAI21_X1 U15204 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20771), .A(
        n20700), .ZN(n11879) );
  NAND2_X1 U15205 ( .A1(n14164), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n11878) );
  OAI211_X1 U15206 ( .C1(n14160), .C2(n11880), .A(n11879), .B(n11878), .ZN(
        n11881) );
  OAI21_X1 U15207 ( .B1(n15841), .B2(n12120), .A(n11881), .ZN(n14386) );
  AOI22_X1 U15208 ( .A1(n14145), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U15209 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11370), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U15210 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U15211 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11882) );
  NAND4_X1 U15212 ( .A1(n11885), .A2(n11884), .A3(n11883), .A4(n11882), .ZN(
        n11891) );
  AOI22_X1 U15213 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12131), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U15214 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U15215 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U15216 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11886) );
  NAND4_X1 U15217 ( .A1(n11889), .A2(n11888), .A3(n11887), .A4(n11886), .ZN(
        n11890) );
  NOR2_X1 U15218 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  OR2_X1 U15219 ( .A1(n14160), .A2(n11892), .ZN(n11896) );
  XNOR2_X1 U15220 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11911), .ZN(
        n15733) );
  INV_X1 U15221 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14543) );
  OAI22_X1 U15222 ( .A1(n15733), .A2(n12120), .B1(n11893), .B2(n14543), .ZN(
        n11894) );
  AOI21_X1 U15223 ( .B1(n14164), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11894), .ZN(
        n11895) );
  NAND2_X1 U15224 ( .A1(n11896), .A2(n11895), .ZN(n14121) );
  INV_X1 U15225 ( .A(n14120), .ZN(n11916) );
  AOI22_X1 U15226 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U15227 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U15228 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U15229 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11897) );
  NAND4_X1 U15230 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11897), .ZN(
        n11906) );
  AOI22_X1 U15231 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U15232 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U15233 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U15234 ( .A1(n14145), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11901) );
  NAND4_X1 U15235 ( .A1(n11904), .A2(n11903), .A3(n11902), .A4(n11901), .ZN(
        n11905) );
  NOR2_X1 U15236 ( .A1(n11906), .A2(n11905), .ZN(n11910) );
  NAND2_X1 U15237 ( .A1(n20700), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11907) );
  NAND2_X1 U15238 ( .A1(n12120), .A2(n11907), .ZN(n11908) );
  AOI21_X1 U15239 ( .B1(n14164), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11908), .ZN(
        n11909) );
  OAI21_X1 U15240 ( .B1(n14160), .B2(n11910), .A(n11909), .ZN(n11914) );
  OAI21_X1 U15241 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11912), .A(
        n11934), .ZN(n15831) );
  OR2_X1 U15242 ( .A1(n12120), .A2(n15831), .ZN(n11913) );
  NAND2_X1 U15243 ( .A1(n11914), .A2(n11913), .ZN(n14377) );
  NAND2_X1 U15244 ( .A1(n11916), .A2(n11915), .ZN(n14312) );
  AOI22_X1 U15245 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U15246 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15247 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U15248 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11917) );
  NAND4_X1 U15249 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(
        n11926) );
  AOI22_X1 U15250 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11370), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15251 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U15252 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U15253 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11921) );
  NAND4_X1 U15254 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11925) );
  NOR2_X1 U15255 ( .A1(n11926), .A2(n11925), .ZN(n11930) );
  NAND2_X1 U15256 ( .A1(n20700), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11927) );
  NAND2_X1 U15257 ( .A1(n12120), .A2(n11927), .ZN(n11928) );
  AOI21_X1 U15258 ( .B1(n14164), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11928), .ZN(
        n11929) );
  OAI21_X1 U15259 ( .B1(n14160), .B2(n11930), .A(n11929), .ZN(n11932) );
  XNOR2_X1 U15260 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n11934), .ZN(
        n14529) );
  NAND2_X1 U15261 ( .A1(n14157), .A2(n14529), .ZN(n11931) );
  NAND2_X1 U15262 ( .A1(n11932), .A2(n11931), .ZN(n14315) );
  INV_X1 U15263 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11933) );
  OR2_X1 U15264 ( .A1(n11935), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11936) );
  NAND2_X1 U15265 ( .A1(n11936), .A2(n11967), .ZN(n15817) );
  AOI22_X1 U15266 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11355), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15267 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12131), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15268 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11988), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15269 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11937) );
  NAND4_X1 U15270 ( .A1(n11940), .A2(n11939), .A3(n11938), .A4(n11937), .ZN(
        n11946) );
  AOI22_X1 U15271 ( .A1(n14145), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U15272 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12130), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U15273 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n14144), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U15274 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11370), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11941) );
  NAND4_X1 U15275 ( .A1(n11944), .A2(n11943), .A3(n11942), .A4(n11941), .ZN(
        n11945) );
  NOR2_X1 U15276 ( .A1(n11946), .A2(n11945), .ZN(n11949) );
  OAI21_X1 U15277 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20771), .A(
        n20700), .ZN(n11948) );
  NAND2_X1 U15278 ( .A1(n14164), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n11947) );
  OAI211_X1 U15279 ( .C1(n14160), .C2(n11949), .A(n11948), .B(n11947), .ZN(
        n11950) );
  OAI21_X1 U15280 ( .B1(n15817), .B2(n12120), .A(n11950), .ZN(n11951) );
  INV_X1 U15281 ( .A(n11951), .ZN(n15720) );
  AOI22_X1 U15282 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15283 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15284 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U15285 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11952) );
  NAND4_X1 U15286 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n11961) );
  AOI22_X1 U15287 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15288 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U15289 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15290 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U15291 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11960) );
  NOR2_X1 U15292 ( .A1(n11961), .A2(n11960), .ZN(n11964) );
  AOI21_X1 U15293 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15715), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11962) );
  AOI21_X1 U15294 ( .B1(n14164), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11962), .ZN(
        n11963) );
  OAI21_X1 U15295 ( .B1(n14160), .B2(n11964), .A(n11963), .ZN(n11966) );
  XNOR2_X1 U15296 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n11967), .ZN(
        n15712) );
  NAND2_X1 U15297 ( .A1(n14157), .A2(n15712), .ZN(n11965) );
  OR2_X1 U15298 ( .A1(n11968), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11969) );
  NAND2_X1 U15299 ( .A1(n11969), .A2(n12026), .ZN(n15816) );
  AOI22_X1 U15300 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12131), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U15301 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15302 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15303 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11970) );
  NAND4_X1 U15304 ( .A1(n11973), .A2(n11972), .A3(n11971), .A4(n11970), .ZN(
        n11979) );
  AOI22_X1 U15305 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12130), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15306 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15307 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15308 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11974) );
  NAND4_X1 U15309 ( .A1(n11977), .A2(n11976), .A3(n11975), .A4(n11974), .ZN(
        n11978) );
  NOR2_X1 U15310 ( .A1(n11979), .A2(n11978), .ZN(n11982) );
  OAI21_X1 U15311 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20771), .A(
        n20700), .ZN(n11981) );
  NAND2_X1 U15312 ( .A1(n14164), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n11980) );
  OAI211_X1 U15313 ( .C1(n14160), .C2(n11982), .A(n11981), .B(n11980), .ZN(
        n11983) );
  OAI21_X1 U15314 ( .B1(n15816), .B2(n12120), .A(n11983), .ZN(n14363) );
  AOI22_X1 U15315 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U15316 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15317 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U15318 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11984) );
  NAND4_X1 U15319 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n11984), .ZN(
        n11994) );
  AOI22_X1 U15320 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15321 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15322 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15323 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11989) );
  NAND4_X1 U15324 ( .A1(n11992), .A2(n11991), .A3(n11990), .A4(n11989), .ZN(
        n11993) );
  NOR2_X1 U15325 ( .A1(n11994), .A2(n11993), .ZN(n12010) );
  AOI22_X1 U15326 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15327 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15328 ( .A1(n11371), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15329 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11995) );
  NAND4_X1 U15330 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        n12004) );
  AOI22_X1 U15331 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15332 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11988), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15333 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15334 ( .A1(n14145), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14138), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11999) );
  NAND4_X1 U15335 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n12003) );
  NOR2_X1 U15336 ( .A1(n12004), .A2(n12003), .ZN(n12011) );
  XNOR2_X1 U15337 ( .A(n12010), .B(n12011), .ZN(n12007) );
  INV_X1 U15338 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15695) );
  OAI21_X1 U15339 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15695), .A(n12120), 
        .ZN(n12005) );
  AOI21_X1 U15340 ( .B1(n14164), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12005), .ZN(
        n12006) );
  OAI21_X1 U15341 ( .B1(n14160), .B2(n12007), .A(n12006), .ZN(n12009) );
  XNOR2_X1 U15342 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12026), .ZN(
        n15692) );
  NAND2_X1 U15343 ( .A1(n14157), .A2(n15692), .ZN(n12008) );
  NAND2_X1 U15344 ( .A1(n12009), .A2(n12008), .ZN(n14352) );
  NOR2_X1 U15345 ( .A1(n12011), .A2(n12010), .ZN(n12033) );
  AOI22_X1 U15346 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15347 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15348 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15349 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U15350 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12021) );
  INV_X1 U15351 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n20849) );
  AOI22_X1 U15352 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15353 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15354 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15355 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U15356 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12020) );
  OR2_X1 U15357 ( .A1(n12021), .A2(n12020), .ZN(n12032) );
  INV_X1 U15358 ( .A(n12032), .ZN(n12022) );
  XNOR2_X1 U15359 ( .A(n12033), .B(n12022), .ZN(n12023) );
  NAND2_X1 U15360 ( .A1(n12023), .A2(n12140), .ZN(n12031) );
  NAND2_X1 U15361 ( .A1(n20700), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12024) );
  NAND2_X1 U15362 ( .A1(n12120), .A2(n12024), .ZN(n12025) );
  AOI21_X1 U15363 ( .B1(n14164), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12025), .ZN(
        n12030) );
  OAI21_X1 U15364 ( .B1(n12028), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n12070), .ZN(n15683) );
  NOR2_X1 U15365 ( .A1(n15683), .A2(n12120), .ZN(n12029) );
  AOI21_X1 U15366 ( .B1(n12031), .B2(n12030), .A(n12029), .ZN(n14345) );
  NAND2_X1 U15367 ( .A1(n12033), .A2(n12032), .ZN(n12050) );
  AOI22_X1 U15368 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15369 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15370 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U15371 ( .A1(n11371), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12034) );
  NAND4_X1 U15372 ( .A1(n12037), .A2(n12036), .A3(n12035), .A4(n12034), .ZN(
        n12044) );
  AOI22_X1 U15373 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15374 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11988), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15375 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15376 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12039) );
  NAND4_X1 U15377 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12043) );
  NOR2_X1 U15378 ( .A1(n12044), .A2(n12043), .ZN(n12051) );
  XOR2_X1 U15379 ( .A(n12050), .B(n12051), .Z(n12045) );
  NAND2_X1 U15380 ( .A1(n12045), .A2(n12140), .ZN(n12049) );
  INV_X1 U15381 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15662) );
  OAI21_X1 U15382 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15662), .A(n12120), 
        .ZN(n12046) );
  AOI21_X1 U15383 ( .B1(n11685), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12046), .ZN(
        n12048) );
  XNOR2_X1 U15384 ( .A(n12070), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15666) );
  AOI21_X1 U15385 ( .B1(n12049), .B2(n12048), .A(n12047), .ZN(n14338) );
  NOR2_X1 U15386 ( .A1(n12051), .A2(n12050), .ZN(n12078) );
  AOI22_X1 U15387 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9631), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15388 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15389 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15390 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12053) );
  NAND4_X1 U15391 ( .A1(n12056), .A2(n12055), .A3(n12054), .A4(n12053), .ZN(
        n12064) );
  AOI22_X1 U15392 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15393 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15394 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15395 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12059) );
  NAND4_X1 U15396 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12063) );
  OR2_X1 U15397 ( .A1(n12064), .A2(n12063), .ZN(n12077) );
  INV_X1 U15398 ( .A(n12077), .ZN(n12065) );
  XNOR2_X1 U15399 ( .A(n12078), .B(n12065), .ZN(n12069) );
  INV_X1 U15400 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12067) );
  NAND2_X1 U15401 ( .A1(n20700), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12066) );
  OAI211_X1 U15402 ( .C1(n12112), .C2(n12067), .A(n12120), .B(n12066), .ZN(
        n12068) );
  AOI21_X1 U15403 ( .B1(n12069), .B2(n12140), .A(n12068), .ZN(n12076) );
  INV_X1 U15404 ( .A(n12071), .ZN(n12073) );
  INV_X1 U15405 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12072) );
  NAND2_X1 U15406 ( .A1(n12073), .A2(n12072), .ZN(n12074) );
  NAND2_X1 U15407 ( .A1(n12115), .A2(n12074), .ZN(n15657) );
  NOR2_X1 U15408 ( .A1(n15657), .A2(n12120), .ZN(n12075) );
  NAND2_X1 U15409 ( .A1(n12078), .A2(n12077), .ZN(n12097) );
  AOI22_X1 U15410 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n14146), .B1(
        n12131), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15411 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11370), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15412 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11355), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15413 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12080) );
  NAND4_X1 U15414 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(
        n12089) );
  AOI22_X1 U15415 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12130), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15416 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11371), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15417 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15418 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11497), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12084) );
  NAND4_X1 U15419 ( .A1(n12087), .A2(n12086), .A3(n12085), .A4(n12084), .ZN(
        n12088) );
  NOR2_X1 U15420 ( .A1(n12089), .A2(n12088), .ZN(n12098) );
  XOR2_X1 U15421 ( .A(n12097), .B(n12098), .Z(n12090) );
  NAND2_X1 U15422 ( .A1(n12090), .A2(n12140), .ZN(n12093) );
  INV_X1 U15423 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14486) );
  AOI21_X1 U15424 ( .B1(n14486), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12091) );
  AOI21_X1 U15425 ( .B1(n11685), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12091), .ZN(
        n12092) );
  NAND2_X1 U15426 ( .A1(n12093), .A2(n12092), .ZN(n12095) );
  XNOR2_X1 U15427 ( .A(n12115), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14484) );
  NAND2_X1 U15428 ( .A1(n14484), .A2(n14157), .ZN(n12094) );
  NAND2_X1 U15429 ( .A1(n12095), .A2(n12094), .ZN(n14305) );
  NOR2_X1 U15430 ( .A1(n12098), .A2(n12097), .ZN(n12125) );
  AOI22_X1 U15431 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9631), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15432 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11496), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15433 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15434 ( .A1(n11988), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U15435 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12108) );
  AOI22_X1 U15436 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15437 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15438 ( .A1(n14144), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15439 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12103) );
  NAND4_X1 U15440 ( .A1(n12106), .A2(n12105), .A3(n12104), .A4(n12103), .ZN(
        n12107) );
  OR2_X1 U15441 ( .A1(n12108), .A2(n12107), .ZN(n12124) );
  INV_X1 U15442 ( .A(n12124), .ZN(n12109) );
  XNOR2_X1 U15443 ( .A(n12125), .B(n12109), .ZN(n12114) );
  INV_X1 U15444 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12111) );
  NAND2_X1 U15445 ( .A1(n20700), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12110) );
  OAI211_X1 U15446 ( .C1(n12112), .C2(n12111), .A(n12120), .B(n12110), .ZN(
        n12113) );
  AOI21_X1 U15447 ( .B1(n12114), .B2(n12140), .A(n12113), .ZN(n12122) );
  INV_X1 U15448 ( .A(n12115), .ZN(n12116) );
  INV_X1 U15449 ( .A(n12117), .ZN(n12118) );
  INV_X1 U15450 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14292) );
  NAND2_X1 U15451 ( .A1(n12118), .A2(n14292), .ZN(n12119) );
  NAND2_X1 U15452 ( .A1(n13788), .A2(n12119), .ZN(n14477) );
  NOR2_X1 U15453 ( .A1(n14477), .A2(n12120), .ZN(n12121) );
  XNOR2_X1 U15454 ( .A(n13788), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14215) );
  NAND2_X1 U15455 ( .A1(n12125), .A2(n12124), .ZN(n14153) );
  AOI22_X1 U15456 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15457 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11988), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15458 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15459 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12126) );
  NAND4_X1 U15460 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12137) );
  AOI22_X1 U15461 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15462 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9631), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15463 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15464 ( .A1(n11371), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U15465 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12136) );
  NOR2_X1 U15466 ( .A1(n12137), .A2(n12136), .ZN(n14154) );
  XOR2_X1 U15467 ( .A(n14153), .B(n14154), .Z(n12141) );
  INV_X1 U15468 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14218) );
  NAND2_X1 U15469 ( .A1(n14164), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12138) );
  OAI211_X1 U15470 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n14218), .A(n12138), 
        .B(n12120), .ZN(n12139) );
  AOI21_X1 U15471 ( .B1(n12141), .B2(n12140), .A(n12139), .ZN(n12142) );
  AOI21_X1 U15472 ( .B1(n14157), .B2(n14215), .A(n12142), .ZN(n12144) );
  NAND2_X1 U15473 ( .A1(n20702), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15950) );
  NAND2_X1 U15474 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20519), .ZN(n20380) );
  NAND2_X1 U15475 ( .A1(n12149), .A2(n20377), .ZN(n20707) );
  AND2_X1 U15476 ( .A1(n20707), .A2(n20702), .ZN(n12146) );
  NAND2_X1 U15477 ( .A1(n20702), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15601) );
  NAND2_X1 U15478 ( .A1(n20771), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12147) );
  AND2_X1 U15479 ( .A1(n15601), .A2(n12147), .ZN(n13354) );
  INV_X1 U15480 ( .A(n13354), .ZN(n12148) );
  INV_X2 U15481 ( .A(n19964), .ZN(n19977) );
  NAND2_X1 U15482 ( .A1(n19977), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14589) );
  OAI21_X1 U15483 ( .B1(n15823), .B2(n14218), .A(n14589), .ZN(n12150) );
  AOI21_X1 U15484 ( .B1(n15849), .B2(n14215), .A(n12150), .ZN(n12151) );
  INV_X1 U15485 ( .A(n12151), .ZN(n12152) );
  NAND2_X1 U15486 ( .A1(n12155), .A2(n12154), .ZN(P1_U2970) );
  INV_X1 U15487 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12170) );
  INV_X1 U15488 ( .A(n12158), .ZN(n12161) );
  INV_X1 U15489 ( .A(n12159), .ZN(n12160) );
  XNOR2_X2 U15490 ( .A(n12166), .B(n12171), .ZN(n18853) );
  INV_X1 U15491 ( .A(n18853), .ZN(n12203) );
  AND2_X2 U15492 ( .A1(n12200), .A2(n12168), .ZN(n12231) );
  INV_X1 U15493 ( .A(n12231), .ZN(n19352) );
  INV_X1 U15494 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12169) );
  OAI22_X1 U15495 ( .A1(n12170), .A2(n19114), .B1(n19352), .B2(n12169), .ZN(
        n12176) );
  NOR2_X1 U15496 ( .A1(n18871), .A2(n12171), .ZN(n12191) );
  INV_X1 U15497 ( .A(n12191), .ZN(n12172) );
  NOR2_X1 U15498 ( .A1(n12176), .A2(n12175), .ZN(n12209) );
  INV_X1 U15499 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12181) );
  INV_X1 U15500 ( .A(n18871), .ZN(n12177) );
  AND2_X1 U15501 ( .A1(n12177), .A2(n12171), .ZN(n12189) );
  INV_X1 U15502 ( .A(n12189), .ZN(n12178) );
  INV_X1 U15503 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12180) );
  OAI22_X1 U15504 ( .A1(n12181), .A2(n19319), .B1(n19382), .B2(n12180), .ZN(
        n12198) );
  AND2_X2 U15505 ( .A1(n13950), .A2(n12183), .ZN(n19141) );
  AOI21_X1 U15506 ( .B1(n19141), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n12750), .ZN(n12186) );
  INV_X1 U15507 ( .A(n9626), .ZN(n19007) );
  AND2_X1 U15508 ( .A1(n19007), .A2(n12189), .ZN(n12184) );
  AND2_X2 U15509 ( .A1(n12184), .A2(n13950), .ZN(n19206) );
  NAND2_X1 U15510 ( .A1(n19206), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12185) );
  OAI211_X1 U15511 ( .C1(n12212), .C2(n12187), .A(n12186), .B(n12185), .ZN(
        n12197) );
  NAND2_X1 U15512 ( .A1(n12188), .A2(n19007), .ZN(n12220) );
  INV_X1 U15513 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12195) );
  AND2_X1 U15514 ( .A1(n9626), .A2(n12189), .ZN(n12190) );
  NAND2_X1 U15515 ( .A1(n19084), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12194) );
  AND2_X2 U15516 ( .A1(n12192), .A2(n13950), .ZN(n12238) );
  NAND2_X1 U15517 ( .A1(n12238), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12193) );
  OAI211_X1 U15518 ( .C1(n12220), .C2(n12195), .A(n12194), .B(n12193), .ZN(
        n12196) );
  INV_X1 U15519 ( .A(n12203), .ZN(n13653) );
  NOR2_X2 U15520 ( .A1(n12204), .A2(n12203), .ZN(n12249) );
  NAND2_X1 U15521 ( .A1(n12750), .A2(n12449), .ZN(n13303) );
  OR2_X1 U15522 ( .A1(n12448), .A2(n13303), .ZN(n12453) );
  NAND2_X1 U15523 ( .A1(n12453), .A2(n12210), .ZN(n12211) );
  AOI22_X1 U15524 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n12253), .B1(
        n12233), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15525 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19033), .B1(
        n12231), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12215) );
  INV_X1 U15526 ( .A(n12212), .ZN(n12232) );
  AOI22_X1 U15527 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19110), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U15528 ( .A1(n12248), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12213) );
  AOI22_X1 U15529 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19084), .B1(
        n19141), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12219) );
  NAND2_X1 U15530 ( .A1(n12249), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12218) );
  AOI22_X1 U15531 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19206), .B1(
        n12238), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12217) );
  NAND3_X1 U15532 ( .A1(n12219), .A2(n12218), .A3(n12217), .ZN(n12223) );
  INV_X1 U15533 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n20825) );
  INV_X1 U15534 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12221) );
  OAI22_X1 U15535 ( .A1(n20825), .A2(n12220), .B1(n19382), .B2(n12221), .ZN(
        n12222) );
  NOR2_X1 U15536 ( .A1(n12223), .A2(n12222), .ZN(n12225) );
  AOI22_X1 U15537 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12205), .B1(
        n12201), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12224) );
  NAND3_X1 U15538 ( .A1(n9661), .A2(n12225), .A3(n12224), .ZN(n12226) );
  NAND2_X1 U15539 ( .A1(n12750), .A2(n12227), .ZN(n12228) );
  INV_X1 U15540 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12949) );
  INV_X1 U15541 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12951) );
  OAI22_X1 U15542 ( .A1(n12949), .A2(n12256), .B1(n19174), .B2(n12951), .ZN(
        n12230) );
  INV_X1 U15543 ( .A(n12230), .ZN(n12243) );
  AOI22_X1 U15544 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19033), .B1(
        n12231), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15545 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19110), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15546 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n12253), .B1(
        n12233), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12235) );
  NAND2_X1 U15547 ( .A1(n12248), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12234) );
  INV_X1 U15548 ( .A(n12220), .ZN(n12261) );
  AOI22_X1 U15549 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n12261), .B1(
        n19379), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15550 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19084), .B1(
        n19141), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12241) );
  NAND2_X1 U15551 ( .A1(n12249), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12240) );
  AOI22_X1 U15552 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19206), .B1(
        n12238), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12239) );
  NAND3_X1 U15553 ( .A1(n12243), .A2(n10089), .A3(n10085), .ZN(n12247) );
  INV_X1 U15554 ( .A(n12244), .ZN(n12245) );
  NAND2_X1 U15555 ( .A1(n12245), .A2(n12750), .ZN(n12246) );
  INV_X1 U15556 ( .A(n12274), .ZN(n12273) );
  INV_X1 U15557 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12970) );
  INV_X1 U15558 ( .A(n12248), .ZN(n12252) );
  INV_X1 U15559 ( .A(n12249), .ZN(n12250) );
  INV_X1 U15560 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12251) );
  OAI22_X1 U15561 ( .A1(n12970), .A2(n12252), .B1(n12250), .B2(n12251), .ZN(
        n12268) );
  AOI22_X1 U15562 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19110), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15563 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12253), .B1(
        n12233), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12259) );
  INV_X1 U15564 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19070) );
  INV_X1 U15565 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12254) );
  OAI22_X1 U15566 ( .A1(n19070), .A2(n19022), .B1(n19352), .B2(n12254), .ZN(
        n12255) );
  INV_X1 U15567 ( .A(n12255), .ZN(n12258) );
  NAND2_X1 U15568 ( .A1(n12205), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12257) );
  NAND4_X1 U15569 ( .A1(n12260), .A2(n12259), .A3(n12258), .A4(n12257), .ZN(
        n12267) );
  AOI22_X1 U15570 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12261), .B1(
        n19379), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15571 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19206), .B1(
        n12238), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12264) );
  NAND2_X1 U15572 ( .A1(n12201), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12263) );
  AOI22_X1 U15573 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19084), .B1(
        n19141), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12262) );
  NAND4_X1 U15574 ( .A1(n12265), .A2(n12264), .A3(n12263), .A4(n12262), .ZN(
        n12266) );
  NAND2_X1 U15575 ( .A1(n12269), .A2(n12750), .ZN(n12270) );
  NAND2_X2 U15576 ( .A1(n12273), .A2(n12272), .ZN(n12471) );
  NAND2_X1 U15577 ( .A1(n12274), .A2(n12465), .ZN(n12275) );
  NOR2_X1 U15578 ( .A1(n12284), .A2(n12276), .ZN(n12277) );
  OR2_X1 U15579 ( .A1(n12319), .A2(n12277), .ZN(n18809) );
  XNOR2_X2 U15580 ( .A(n12279), .B(n12278), .ZN(n12462) );
  NAND2_X1 U15581 ( .A1(n12462), .A2(n12280), .ZN(n12285) );
  NOR2_X1 U15582 ( .A1(n12282), .A2(n12281), .ZN(n12283) );
  OR2_X1 U15583 ( .A1(n12284), .A2(n12283), .ZN(n18820) );
  NAND2_X2 U15584 ( .A1(n12285), .A2(n18820), .ZN(n12309) );
  INV_X1 U15585 ( .A(n12286), .ZN(n12289) );
  INV_X1 U15586 ( .A(n12287), .ZN(n12288) );
  OAI21_X1 U15587 ( .B1(n12293), .B2(n12296), .A(n12291), .ZN(n12292) );
  NAND2_X1 U15588 ( .A1(n12308), .A2(n12292), .ZN(n13955) );
  XNOR2_X1 U15589 ( .A(n12293), .B(n12296), .ZN(n12305) );
  XNOR2_X1 U15590 ( .A(n12305), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14232) );
  AND2_X1 U15591 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12294) );
  NAND2_X1 U15592 ( .A1(n19061), .A2(n12294), .ZN(n12295) );
  NAND2_X1 U15593 ( .A1(n12296), .A2(n12295), .ZN(n18851) );
  INV_X1 U15594 ( .A(n12449), .ZN(n12301) );
  OAI21_X1 U15595 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19729), .A(
        n12297), .ZN(n12749) );
  INV_X1 U15596 ( .A(n12749), .ZN(n12745) );
  NAND2_X1 U15597 ( .A1(n12298), .A2(n12745), .ZN(n12300) );
  NAND2_X1 U15598 ( .A1(n19061), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12299) );
  OAI211_X1 U15599 ( .C1(n12302), .C2(n12301), .A(n12300), .B(n12299), .ZN(
        n18864) );
  NAND2_X1 U15600 ( .A1(n18864), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13308) );
  OAI21_X1 U15601 ( .B1(n18851), .B2(n15446), .A(n13308), .ZN(n12304) );
  NAND2_X1 U15602 ( .A1(n18851), .A2(n15446), .ZN(n12303) );
  AND2_X1 U15603 ( .A1(n12304), .A2(n12303), .ZN(n14233) );
  NAND2_X1 U15604 ( .A1(n14232), .A2(n14233), .ZN(n18991) );
  INV_X1 U15605 ( .A(n12305), .ZN(n13964) );
  NAND2_X1 U15606 ( .A1(n13964), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12306) );
  AND2_X1 U15607 ( .A1(n18991), .A2(n12306), .ZN(n13891) );
  XNOR2_X1 U15608 ( .A(n12308), .B(n12307), .ZN(n18833) );
  XNOR2_X1 U15609 ( .A(n18833), .B(n13938), .ZN(n13936) );
  NAND2_X1 U15610 ( .A1(n12309), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12310) );
  NAND2_X1 U15611 ( .A1(n12311), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12312) );
  AND3_X1 U15612 ( .A1(n12315), .A2(n19061), .A3(P2_EBX_REG_8__SCAN_IN), .ZN(
        n12316) );
  NOR2_X1 U15613 ( .A1(n12314), .A2(n12316), .ZN(n18798) );
  NAND2_X1 U15614 ( .A1(n18798), .A2(n12548), .ZN(n12321) );
  INV_X1 U15615 ( .A(n12317), .ZN(n12318) );
  XNOR2_X1 U15616 ( .A(n12319), .B(n12318), .ZN(n13974) );
  NAND2_X1 U15617 ( .A1(n12321), .A2(n14181), .ZN(n14170) );
  INV_X1 U15618 ( .A(n13974), .ZN(n12322) );
  NAND2_X1 U15619 ( .A1(n12322), .A2(n9839), .ZN(n15111) );
  AND2_X1 U15620 ( .A1(n14170), .A2(n15111), .ZN(n12323) );
  NOR2_X1 U15621 ( .A1(n12403), .A2(n12324), .ZN(n12325) );
  XNOR2_X1 U15622 ( .A(n12314), .B(n12325), .ZN(n18782) );
  AOI21_X1 U15623 ( .B1(n18782), .B2(n12548), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15405) );
  NAND2_X1 U15624 ( .A1(n19061), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12327) );
  MUX2_X1 U15625 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n12327), .S(n12326), .Z(
        n12328) );
  AND2_X1 U15626 ( .A1(n12328), .A2(n12411), .ZN(n18771) );
  NAND2_X1 U15627 ( .A1(n18771), .A2(n12548), .ZN(n12338) );
  NAND2_X1 U15628 ( .A1(n12338), .A2(n15393), .ZN(n15387) );
  NAND2_X1 U15629 ( .A1(n19061), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12329) );
  OR2_X1 U15630 ( .A1(n12330), .A2(n12329), .ZN(n12333) );
  INV_X1 U15631 ( .A(n12331), .ZN(n12332) );
  AOI21_X1 U15632 ( .B1(n12335), .B2(n12548), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15378) );
  INV_X1 U15633 ( .A(n12335), .ZN(n18760) );
  OR2_X1 U15634 ( .A1(n12280), .A2(n15367), .ZN(n12336) );
  NOR2_X1 U15635 ( .A1(n12280), .A2(n15412), .ZN(n12337) );
  NAND2_X1 U15636 ( .A1(n18782), .A2(n12337), .ZN(n15384) );
  OR2_X1 U15637 ( .A1(n15393), .A2(n12338), .ZN(n15386) );
  AND2_X1 U15638 ( .A1(n15384), .A2(n15386), .ZN(n15375) );
  NAND2_X1 U15639 ( .A1(n15377), .A2(n15375), .ZN(n15351) );
  INV_X1 U15640 ( .A(n12339), .ZN(n12341) );
  NAND2_X1 U15641 ( .A1(n12341), .A2(n12340), .ZN(n12342) );
  AND2_X1 U15642 ( .A1(n12368), .A2(n12342), .ZN(n13911) );
  AND2_X1 U15643 ( .A1(n13911), .A2(n12548), .ZN(n12366) );
  AND2_X1 U15644 ( .A1(n12366), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15355) );
  NOR2_X1 U15645 ( .A1(n15351), .A2(n15355), .ZN(n12343) );
  INV_X1 U15646 ( .A(n12360), .ZN(n12345) );
  NAND2_X1 U15647 ( .A1(n12346), .A2(n13826), .ZN(n12349) );
  NAND3_X1 U15648 ( .A1(n12349), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n19061), 
        .ZN(n12344) );
  NAND2_X1 U15649 ( .A1(n12345), .A2(n12344), .ZN(n18725) );
  NOR2_X1 U15650 ( .A1(n12280), .A2(n18725), .ZN(n12390) );
  NOR2_X1 U15651 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n12390), .ZN(
        n15319) );
  INV_X1 U15652 ( .A(n15319), .ZN(n12372) );
  INV_X1 U15653 ( .A(n12346), .ZN(n12347) );
  NAND2_X1 U15654 ( .A1(n12347), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12348) );
  MUX2_X1 U15655 ( .A(n12348), .B(n12347), .S(n12403), .Z(n12350) );
  NAND2_X1 U15656 ( .A1(n12350), .A2(n12349), .ZN(n18740) );
  NAND2_X1 U15657 ( .A1(n16069), .A2(n12389), .ZN(n15320) );
  NAND2_X1 U15658 ( .A1(n12354), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12351) );
  OAI21_X1 U15659 ( .B1(n12351), .B2(n12808), .A(n12411), .ZN(n12352) );
  INV_X1 U15660 ( .A(n12352), .ZN(n12353) );
  OAI21_X1 U15661 ( .B1(n12354), .B2(P2_EBX_REG_21__SCAN_IN), .A(n12353), .ZN(
        n14815) );
  OR2_X1 U15662 ( .A1(n14815), .A2(n12280), .ZN(n12355) );
  NAND2_X1 U15663 ( .A1(n19061), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12356) );
  XNOR2_X1 U15664 ( .A(n9637), .B(n12356), .ZN(n18668) );
  NAND2_X1 U15665 ( .A1(n18668), .A2(n12548), .ZN(n12357) );
  NAND2_X1 U15666 ( .A1(n12357), .A2(n15636), .ZN(n15077) );
  INV_X1 U15667 ( .A(n15077), .ZN(n15075) );
  NAND2_X1 U15668 ( .A1(n19061), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12359) );
  INV_X1 U15669 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12358) );
  NAND2_X1 U15670 ( .A1(n12360), .A2(n12358), .ZN(n12374) );
  OAI211_X1 U15671 ( .C1(n12360), .C2(n12359), .A(n12411), .B(n12374), .ZN(
        n18718) );
  OR2_X1 U15672 ( .A1(n18718), .A2(n12280), .ZN(n12361) );
  XNOR2_X1 U15673 ( .A(n12361), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15099) );
  NAND2_X1 U15674 ( .A1(n12364), .A2(n12362), .ZN(n12363) );
  NAND2_X1 U15675 ( .A1(n9637), .A2(n12363), .ZN(n18680) );
  NOR2_X1 U15676 ( .A1(n18680), .A2(n12280), .ZN(n12381) );
  NOR2_X1 U15677 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n12381), .ZN(
        n15246) );
  OAI21_X1 U15678 ( .B1(n12373), .B2(n12365), .A(n12364), .ZN(n18693) );
  NOR2_X1 U15679 ( .A1(n18693), .A2(n12280), .ZN(n12382) );
  NOR2_X1 U15680 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n12382), .ZN(
        n15265) );
  NOR2_X1 U15681 ( .A1(n15246), .A2(n15265), .ZN(n15072) );
  NOR2_X1 U15682 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n12366), .ZN(
        n15336) );
  INV_X1 U15683 ( .A(n15336), .ZN(n15354) );
  XNOR2_X1 U15684 ( .A(n12368), .B(n12367), .ZN(n18748) );
  NAND2_X1 U15685 ( .A1(n18748), .A2(n12548), .ZN(n12385) );
  NAND2_X1 U15686 ( .A1(n12384), .A2(n12385), .ZN(n15338) );
  NAND2_X1 U15687 ( .A1(n15354), .A2(n15338), .ZN(n15322) );
  INV_X1 U15688 ( .A(n15322), .ZN(n12369) );
  NAND3_X1 U15689 ( .A1(n15099), .A2(n15072), .A3(n12369), .ZN(n12370) );
  NOR3_X1 U15690 ( .A1(n15231), .A2(n15075), .A3(n12370), .ZN(n12371) );
  NAND3_X1 U15691 ( .A1(n12372), .A2(n15320), .A3(n12371), .ZN(n12377) );
  INV_X1 U15692 ( .A(n12373), .ZN(n12376) );
  NAND3_X1 U15693 ( .A1(n12374), .A2(n19061), .A3(P2_EBX_REG_17__SCAN_IN), 
        .ZN(n12375) );
  NAND2_X1 U15694 ( .A1(n12376), .A2(n12375), .ZN(n18704) );
  NOR2_X1 U15695 ( .A1(n12280), .A2(n18704), .ZN(n12379) );
  NOR2_X1 U15696 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n12379), .ZN(
        n15089) );
  NOR2_X1 U15697 ( .A1(n12377), .A2(n15089), .ZN(n12378) );
  AND2_X1 U15698 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n12379), .ZN(
        n15088) );
  OR2_X1 U15699 ( .A1(n12280), .A2(n15289), .ZN(n12380) );
  NOR2_X1 U15700 ( .A1(n18718), .A2(n12380), .ZN(n15087) );
  NOR2_X1 U15701 ( .A1(n15088), .A2(n15087), .ZN(n15071) );
  NAND2_X1 U15702 ( .A1(n12381), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15247) );
  NAND2_X1 U15703 ( .A1(n12382), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15267) );
  NAND2_X1 U15704 ( .A1(n15247), .A2(n15267), .ZN(n15073) );
  INV_X1 U15705 ( .A(n15073), .ZN(n12388) );
  OR2_X1 U15706 ( .A1(n12280), .A2(n15227), .ZN(n12383) );
  NOR2_X1 U15707 ( .A1(n14815), .A2(n12383), .ZN(n15232) );
  NOR2_X1 U15708 ( .A1(n12385), .A2(n12384), .ZN(n15321) );
  NOR2_X1 U15709 ( .A1(n15232), .A2(n15321), .ZN(n12387) );
  NOR2_X1 U15710 ( .A1(n12280), .A2(n15636), .ZN(n12386) );
  NAND2_X1 U15711 ( .A1(n18668), .A2(n12386), .ZN(n15230) );
  NAND4_X1 U15712 ( .A1(n15071), .A2(n12388), .A3(n12387), .A4(n15230), .ZN(
        n12391) );
  NOR2_X1 U15713 ( .A1(n16069), .A2(n12389), .ZN(n15323) );
  AND2_X1 U15714 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n12390), .ZN(
        n15318) );
  NOR2_X1 U15715 ( .A1(n12391), .A2(n15065), .ZN(n12392) );
  INV_X1 U15716 ( .A(n12394), .ZN(n12395) );
  NAND2_X1 U15717 ( .A1(n12395), .A2(n9653), .ZN(n12396) );
  NAND2_X1 U15718 ( .A1(n12400), .A2(n12396), .ZN(n14814) );
  OR2_X1 U15719 ( .A1(n14814), .A2(n12280), .ZN(n12397) );
  NAND2_X1 U15720 ( .A1(n12397), .A2(n15218), .ZN(n15048) );
  OR2_X1 U15721 ( .A1(n12280), .A2(n15218), .ZN(n12398) );
  NAND2_X1 U15722 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  NAND2_X1 U15723 ( .A1(n13211), .A2(n12548), .ZN(n12402) );
  XNOR2_X1 U15724 ( .A(n12402), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15044) );
  INV_X1 U15725 ( .A(n12413), .ZN(n12408) );
  INV_X1 U15726 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14865) );
  NOR2_X1 U15727 ( .A1(n12403), .A2(n14865), .ZN(n12405) );
  INV_X1 U15728 ( .A(n12411), .ZN(n12404) );
  AOI21_X1 U15729 ( .B1(n12406), .B2(n12405), .A(n12404), .ZN(n12407) );
  NAND2_X1 U15730 ( .A1(n12408), .A2(n12407), .ZN(n15996) );
  NOR2_X1 U15731 ( .A1(n15008), .A2(n15195), .ZN(n12417) );
  NAND2_X1 U15732 ( .A1(n19061), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12409) );
  OR2_X1 U15733 ( .A1(n12415), .A2(n12409), .ZN(n12410) );
  INV_X1 U15734 ( .A(n15008), .ZN(n15023) );
  NAND2_X1 U15735 ( .A1(n19061), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12412) );
  OAI21_X1 U15736 ( .B1(n12413), .B2(n12412), .A(n12411), .ZN(n12414) );
  OR2_X1 U15737 ( .A1(n12415), .A2(n12414), .ZN(n14793) );
  OAI21_X1 U15738 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15023), .A(
        n15177), .ZN(n12416) );
  NAND3_X1 U15739 ( .A1(n19061), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n12418), 
        .ZN(n12419) );
  NAND2_X1 U15740 ( .A1(n12430), .A2(n12419), .ZN(n14777) );
  INV_X1 U15741 ( .A(n12537), .ZN(n12426) );
  INV_X1 U15742 ( .A(n12420), .ZN(n12421) );
  NAND2_X1 U15743 ( .A1(n12421), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12424) );
  INV_X1 U15744 ( .A(n14793), .ZN(n12423) );
  NOR2_X1 U15745 ( .A1(n12280), .A2(n15187), .ZN(n12422) );
  NAND2_X1 U15746 ( .A1(n12423), .A2(n12422), .ZN(n15176) );
  NAND2_X1 U15747 ( .A1(n12534), .A2(n12427), .ZN(n12425) );
  AOI21_X1 U15748 ( .B1(n12534), .B2(n12538), .A(n12427), .ZN(n12428) );
  NAND2_X1 U15749 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  NAND2_X1 U15750 ( .A1(n12432), .A2(n12431), .ZN(n15972) );
  XOR2_X1 U15751 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n12536), .Z(
        n12433) );
  OAI21_X1 U15752 ( .B1(n12749), .B2(n12436), .A(n12435), .ZN(n12437) );
  NAND2_X1 U15753 ( .A1(n12758), .A2(n12437), .ZN(n12439) );
  NAND2_X1 U15754 ( .A1(n12439), .A2(n12438), .ZN(n19735) );
  INV_X1 U15755 ( .A(n19734), .ZN(n19750) );
  OAI21_X1 U15756 ( .B1(n12749), .B2(n12440), .A(n13633), .ZN(n12441) );
  INV_X1 U15757 ( .A(n12441), .ZN(n12443) );
  INV_X1 U15758 ( .A(n13446), .ZN(n12442) );
  NAND2_X1 U15759 ( .A1(n12442), .A2(n15561), .ZN(n15556) );
  INV_X1 U15760 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13642) );
  OAI21_X1 U15761 ( .B1(n10904), .B2(n15556), .A(n13642), .ZN(n19720) );
  MUX2_X1 U15762 ( .A(n12443), .B(n19720), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n16159) );
  OAI22_X1 U15763 ( .A1(n19735), .A2(n19750), .B1(n12750), .B2(n19732), .ZN(
        n12444) );
  NAND2_X1 U15764 ( .A1(n12444), .A2(n13646), .ZN(n12784) );
  NOR2_X2 U15765 ( .A1(n13230), .A2(n12750), .ZN(n16112) );
  NAND2_X1 U15766 ( .A1(n15142), .A2(n16112), .ZN(n12497) );
  INV_X1 U15767 ( .A(n13932), .ZN(n12447) );
  NAND2_X1 U15768 ( .A1(n13932), .A2(n13938), .ZN(n12459) );
  NAND2_X1 U15769 ( .A1(n13303), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13302) );
  INV_X1 U15770 ( .A(n13302), .ZN(n12450) );
  XNOR2_X1 U15771 ( .A(n12449), .B(n12448), .ZN(n12451) );
  NAND2_X1 U15772 ( .A1(n12450), .A2(n12451), .ZN(n12452) );
  XNOR2_X1 U15773 ( .A(n12451), .B(n13302), .ZN(n13311) );
  NAND2_X1 U15774 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13311), .ZN(
        n13310) );
  NAND2_X1 U15775 ( .A1(n12452), .A2(n13310), .ZN(n12455) );
  XNOR2_X1 U15776 ( .A(n12810), .B(n12455), .ZN(n14228) );
  INV_X1 U15777 ( .A(n12453), .ZN(n12454) );
  XNOR2_X1 U15778 ( .A(n11146), .B(n12454), .ZN(n14227) );
  NAND2_X1 U15779 ( .A1(n14228), .A2(n14227), .ZN(n14226) );
  NAND2_X1 U15780 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12455), .ZN(
        n12456) );
  NAND2_X1 U15781 ( .A1(n14226), .A2(n12456), .ZN(n12457) );
  XNOR2_X1 U15782 ( .A(n12457), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13893) );
  NAND2_X1 U15783 ( .A1(n12457), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12458) );
  INV_X1 U15784 ( .A(n9613), .ZN(n12468) );
  NAND2_X1 U15785 ( .A1(n12467), .A2(n12465), .ZN(n12466) );
  NAND2_X1 U15786 ( .A1(n15122), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15121) );
  INV_X1 U15787 ( .A(n12467), .ZN(n15439) );
  NAND2_X1 U15788 ( .A1(n12469), .A2(n12468), .ZN(n12470) );
  XNOR2_X1 U15789 ( .A(n12474), .B(n14181), .ZN(n14175) );
  NAND2_X1 U15790 ( .A1(n12471), .A2(n12280), .ZN(n12473) );
  NAND2_X1 U15791 ( .A1(n12474), .A2(n12473), .ZN(n15108) );
  INV_X1 U15792 ( .A(n12474), .ZN(n12475) );
  NAND2_X1 U15793 ( .A1(n12475), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12476) );
  NAND2_X2 U15794 ( .A1(n14173), .A2(n12476), .ZN(n15082) );
  AND2_X1 U15795 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16120) );
  AND2_X1 U15796 ( .A1(n16120), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15314) );
  AND3_X1 U15797 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15343) );
  NAND2_X1 U15798 ( .A1(n15314), .A2(n15343), .ZN(n15288) );
  NAND3_X1 U15799 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15253) );
  NOR2_X1 U15800 ( .A1(n15288), .A2(n15253), .ZN(n15085) );
  NAND2_X1 U15801 ( .A1(n15085), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12839) );
  INV_X1 U15802 ( .A(n12839), .ZN(n12477) );
  AND2_X1 U15803 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12840) );
  OAI21_X1 U15804 ( .B1(n12479), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12552), .ZN(n15151) );
  NOR2_X2 U15805 ( .A1(n13230), .A2(n13231), .ZN(n16113) );
  AND2_X1 U15806 ( .A1(n12480), .A2(n12481), .ZN(n12482) );
  OR2_X1 U15807 ( .A1(n14762), .A2(n12482), .ZN(n15966) );
  INV_X1 U15808 ( .A(n15966), .ZN(n15148) );
  NAND2_X1 U15809 ( .A1(n19690), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19714) );
  NAND2_X1 U15810 ( .A1(n12762), .A2(n12743), .ZN(n12484) );
  NAND2_X1 U15811 ( .A1(n19751), .A2(n15561), .ZN(n12483) );
  NAND2_X1 U15812 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19751), .ZN(n13461) );
  INV_X1 U15813 ( .A(n13461), .ZN(n12485) );
  OAI21_X1 U15814 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n19751), .ZN(n16162) );
  INV_X1 U15815 ( .A(n16162), .ZN(n19746) );
  NAND2_X1 U15816 ( .A1(n19746), .A2(n19721), .ZN(n12486) );
  OR2_X2 U15817 ( .A1(n19714), .A2(n19509), .ZN(n19026) );
  OR2_X1 U15818 ( .A1(n19690), .A2(n19693), .ZN(n19694) );
  NAND2_X1 U15819 ( .A1(n19694), .A2(n19751), .ZN(n12488) );
  INV_X1 U15820 ( .A(n18839), .ZN(n19017) );
  NAND2_X1 U15821 ( .A1(n18822), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15143) );
  OAI21_X1 U15822 ( .B1(n16117), .B2(n12489), .A(n15143), .ZN(n12493) );
  NAND2_X1 U15823 ( .A1(n19751), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12874) );
  NAND2_X1 U15824 ( .A1(n19692), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12490) );
  NAND2_X1 U15825 ( .A1(n12874), .A2(n12490), .ZN(n13305) );
  NOR2_X1 U15826 ( .A1(n12491), .A2(n18989), .ZN(n12492) );
  AOI211_X1 U15827 ( .C1(n15148), .C2(n18985), .A(n12493), .B(n12492), .ZN(
        n12494) );
  INV_X1 U15828 ( .A(n12495), .ZN(n12496) );
  NAND2_X1 U15829 ( .A1(n12497), .A2(n12496), .ZN(P2_U2986) );
  INV_X1 U15830 ( .A(n16189), .ZN(n15568) );
  NOR2_X1 U15831 ( .A1(n18405), .A2(n17103), .ZN(n17819) );
  INV_X1 U15832 ( .A(n17819), .ZN(n17690) );
  NOR2_X1 U15833 ( .A1(n17271), .A2(n17269), .ZN(n12524) );
  AOI21_X1 U15834 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17428), .A(
        n12525), .ZN(n17258) );
  NOR2_X1 U15835 ( .A1(n12524), .A2(n17258), .ZN(n17257) );
  NOR2_X1 U15836 ( .A1(n18405), .A2(n12526), .ZN(n12498) );
  NAND2_X1 U15837 ( .A1(n12499), .A2(n12498), .ZN(n12501) );
  INV_X1 U15838 ( .A(n17801), .ZN(n18399) );
  NAND2_X1 U15839 ( .A1(n16187), .A2(n18399), .ZN(n12500) );
  INV_X1 U15840 ( .A(n12502), .ZN(n12503) );
  OAI21_X1 U15841 ( .B1(n15568), .B2(n17690), .A(n12503), .ZN(n12523) );
  INV_X1 U15842 ( .A(n9629), .ZN(n17952) );
  NOR2_X1 U15843 ( .A1(n18438), .A2(n17952), .ZN(n17828) );
  NOR2_X1 U15844 ( .A1(n20785), .A2(n17676), .ZN(n17658) );
  INV_X1 U15845 ( .A(n17658), .ZN(n17656) );
  NOR2_X1 U15846 ( .A1(n12504), .A2(n17656), .ZN(n17268) );
  INV_X1 U15847 ( .A(n17268), .ZN(n17634) );
  INV_X1 U15848 ( .A(n17738), .ZN(n17338) );
  NAND3_X1 U15849 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17849) );
  NAND2_X1 U15850 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17857) );
  NOR3_X1 U15851 ( .A1(n17859), .A2(n17849), .A3(n17857), .ZN(n17735) );
  NAND2_X1 U15852 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17894) );
  INV_X1 U15853 ( .A(n17894), .ZN(n17851) );
  NAND2_X1 U15854 ( .A1(n17735), .A2(n17851), .ZN(n17821) );
  NOR2_X1 U15855 ( .A1(n12518), .A2(n17821), .ZN(n17694) );
  INV_X1 U15856 ( .A(n17694), .ZN(n17737) );
  NOR2_X1 U15857 ( .A1(n17338), .A2(n17737), .ZN(n12527) );
  NAND2_X1 U15858 ( .A1(n15563), .A2(n12527), .ZN(n17629) );
  NAND2_X1 U15859 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17694), .ZN(
        n17755) );
  NOR4_X1 U15860 ( .A1(n17300), .A2(n17627), .A3(n17634), .A4(n17755), .ZN(
        n12519) );
  AOI21_X1 U15861 ( .B1(n12507), .B2(n12506), .A(n12505), .ZN(n12508) );
  INV_X1 U15862 ( .A(n12510), .ZN(n18404) );
  INV_X1 U15863 ( .A(n15458), .ZN(n18400) );
  OAI21_X1 U15864 ( .B1(n17975), .B2(n18619), .A(n12511), .ZN(n12512) );
  OAI21_X1 U15865 ( .B1(n18618), .B2(n12512), .A(n18613), .ZN(n16310) );
  NOR2_X1 U15866 ( .A1(n16311), .A2(n16310), .ZN(n12514) );
  MUX2_X1 U15867 ( .A(n18400), .B(n12514), .S(n12513), .Z(n12515) );
  AOI21_X1 U15868 ( .B1(n18404), .B2(n12516), .A(n12515), .ZN(n12517) );
  OAI21_X1 U15869 ( .B1(n18595), .B2(n18576), .A(n17913), .ZN(n17893) );
  NAND2_X1 U15870 ( .A1(n17735), .A2(n17893), .ZN(n17754) );
  NOR3_X1 U15871 ( .A1(n12518), .A2(n17338), .A3(n17754), .ZN(n17692) );
  INV_X1 U15872 ( .A(n18438), .ZN(n17919) );
  AOI21_X1 U15873 ( .B1(n15563), .B2(n17692), .A(n17919), .ZN(n17673) );
  AOI21_X1 U15874 ( .B1(n18438), .B2(n17634), .A(n17673), .ZN(n17637) );
  OAI211_X1 U15875 ( .C1(n18427), .C2(n12519), .A(n17934), .B(n17637), .ZN(
        n12520) );
  AOI221_X1 U15876 ( .B1(n17634), .B2(n17952), .C1(n17629), .C2(n17952), .A(
        n12520), .ZN(n15614) );
  OAI21_X1 U15877 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17828), .A(
        n15614), .ZN(n15571) );
  NOR2_X1 U15878 ( .A1(n17940), .A2(n12521), .ZN(n12522) );
  OAI21_X1 U15879 ( .B1(n12523), .B2(n15571), .A(n12522), .ZN(n12533) );
  NOR2_X1 U15880 ( .A1(n18405), .A2(n17951), .ZN(n17949) );
  NAND3_X1 U15881 ( .A1(n12525), .A2(n17949), .A3(n12524), .ZN(n12532) );
  NOR3_X2 U15882 ( .A1(n18405), .A2(n17951), .A3(n12526), .ZN(n17862) );
  NAND3_X1 U15883 ( .A1(n17271), .A2(n17862), .A3(n17258), .ZN(n12531) );
  INV_X1 U15884 ( .A(n17835), .ZN(n17877) );
  NAND2_X1 U15885 ( .A1(n10214), .A2(n17738), .ZN(n12528) );
  AOI22_X1 U15886 ( .A1(n17493), .A2(n18399), .B1(n17495), .B2(n17819), .ZN(
        n17736) );
  OAI21_X1 U15887 ( .B1(n18427), .B2(n18595), .A(n9629), .ZN(n17917) );
  AOI22_X1 U15888 ( .A1(n18438), .A2(n17692), .B1(n12527), .B2(n17917), .ZN(
        n15565) );
  OAI21_X1 U15889 ( .B1(n12528), .B2(n17736), .A(n15565), .ZN(n12529) );
  INV_X1 U15890 ( .A(n12529), .ZN(n17708) );
  NOR2_X1 U15891 ( .A1(n17708), .A2(n17341), .ZN(n17703) );
  NAND2_X1 U15892 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17703), .ZN(
        n17684) );
  NOR2_X1 U15893 ( .A1(n17951), .A2(n17684), .ZN(n17680) );
  NOR3_X1 U15894 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17627), .A3(
        n17634), .ZN(n17259) );
  AOI22_X1 U15895 ( .A1(n17877), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17680), 
        .B2(n17259), .ZN(n12530) );
  NAND4_X1 U15896 ( .A1(n12533), .A2(n12532), .A3(n12531), .A4(n12530), .ZN(
        P3_U2834) );
  INV_X1 U15897 ( .A(n12534), .ZN(n12535) );
  XNOR2_X1 U15898 ( .A(n12541), .B(n12540), .ZN(n12544) );
  OAI21_X1 U15899 ( .B1(n12544), .B2(n12280), .A(n15128), .ZN(n14988) );
  AOI21_X1 U15900 ( .B1(n12542), .B2(n12548), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14194) );
  INV_X1 U15901 ( .A(n12544), .ZN(n14767) );
  NAND3_X1 U15902 ( .A1(n14767), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12548), .ZN(n14989) );
  NOR2_X1 U15903 ( .A1(n12545), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12546) );
  MUX2_X1 U15904 ( .A(n12547), .B(n12546), .S(n19061), .Z(n15958) );
  NAND2_X1 U15905 ( .A1(n15958), .A2(n12548), .ZN(n12549) );
  XNOR2_X1 U15906 ( .A(n12549), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12550) );
  XNOR2_X1 U15907 ( .A(n12551), .B(n12550), .ZN(n12791) );
  OR2_X1 U15908 ( .A1(n12791), .A2(n18981), .ZN(n12564) );
  XNOR2_X1 U15909 ( .A(n12553), .B(n12846), .ZN(n12851) );
  NOR2_X1 U15910 ( .A1(n14764), .A2(n12554), .ZN(n12560) );
  AOI22_X1 U15911 ( .A1(n12555), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12556) );
  OAI21_X1 U15912 ( .B1(n10675), .B2(n12557), .A(n12556), .ZN(n12558) );
  AOI21_X1 U15913 ( .B1(n9616), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12558), .ZN(n12559) );
  XNOR2_X1 U15914 ( .A(n12560), .B(n12559), .ZN(n16001) );
  NAND2_X1 U15915 ( .A1(n18822), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U15916 ( .A1(n18977), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12561) );
  OAI211_X1 U15917 ( .C1(n12833), .C2(n19026), .A(n12807), .B(n12561), .ZN(
        n12563) );
  NAND3_X1 U15918 ( .A1(n12564), .A2(n9668), .A3(n10080), .ZN(P2_U2983) );
  AND2_X1 U15919 ( .A1(n14539), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12565) );
  INV_X1 U15920 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14462) );
  NOR3_X1 U15921 ( .A1(n12570), .A2(n12569), .A3(n12568), .ZN(n12572) );
  OAI21_X1 U15922 ( .B1(n12573), .B2(n12572), .A(n12571), .ZN(n14245) );
  INV_X1 U15923 ( .A(n12574), .ZN(n12575) );
  NAND2_X1 U15924 ( .A1(n12575), .A2(n20598), .ZN(n15620) );
  NAND2_X1 U15925 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20708) );
  AOI21_X1 U15926 ( .B1(n20025), .B2(n15620), .A(n15619), .ZN(n12576) );
  NAND2_X1 U15927 ( .A1(n14245), .A2(n12576), .ZN(n12582) );
  INV_X1 U15928 ( .A(n15620), .ZN(n13397) );
  OAI21_X1 U15929 ( .B1(n20025), .B2(n13397), .A(n20708), .ZN(n13795) );
  INV_X1 U15930 ( .A(n13795), .ZN(n12577) );
  NAND2_X1 U15931 ( .A1(n12577), .A2(n13489), .ZN(n12578) );
  INV_X1 U15932 ( .A(n13425), .ZN(n13428) );
  NAND3_X1 U15933 ( .A1(n12578), .A2(n13399), .A3(n13428), .ZN(n12579) );
  NAND2_X1 U15934 ( .A1(n14252), .A2(n12579), .ZN(n12581) );
  MUX2_X1 U15935 ( .A(n12582), .B(n12581), .S(n12580), .Z(n12589) );
  AND2_X1 U15936 ( .A1(n12583), .A2(n20012), .ZN(n14246) );
  INV_X1 U15937 ( .A(n14246), .ZN(n12587) );
  NAND2_X1 U15938 ( .A1(n12584), .A2(n20025), .ZN(n12717) );
  AND2_X1 U15939 ( .A1(n12717), .A2(n13399), .ZN(n12585) );
  AND2_X1 U15940 ( .A1(n12586), .A2(n12585), .ZN(n12710) );
  AOI21_X1 U15941 ( .B1(n12587), .B2(n13417), .A(n12710), .ZN(n13491) );
  OR3_X1 U15942 ( .A1(n14252), .A2(n12599), .A3(n14742), .ZN(n12588) );
  NAND3_X1 U15943 ( .A1(n12589), .A2(n13491), .A3(n12588), .ZN(n12590) );
  INV_X1 U15944 ( .A(n12723), .ZN(n12598) );
  NOR2_X1 U15945 ( .A1(n12593), .A2(n14251), .ZN(n12594) );
  OR2_X1 U15946 ( .A1(n13417), .A2(n12594), .ZN(n14242) );
  INV_X1 U15947 ( .A(n12701), .ZN(n12595) );
  NAND2_X1 U15948 ( .A1(n12595), .A2(n20036), .ZN(n12596) );
  AND4_X1 U15949 ( .A1(n12591), .A2(n12592), .A3(n14242), .A4(n12596), .ZN(
        n12597) );
  OR2_X2 U15950 ( .A1(n12599), .A2(n20012), .ZN(n12601) );
  XNOR2_X1 U15951 ( .A(n12600), .B(n14278), .ZN(n12699) );
  INV_X1 U15952 ( .A(n12623), .ZN(n14276) );
  OR2_X1 U15953 ( .A1(n12600), .A2(n14276), .ZN(n12698) );
  INV_X1 U15954 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19987) );
  NAND2_X1 U15955 ( .A1(n12680), .A2(n19987), .ZN(n12602) );
  NAND2_X1 U15956 ( .A1(n12603), .A2(n12602), .ZN(n12606) );
  INV_X1 U15957 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13802) );
  XNOR2_X1 U15958 ( .A(n12606), .B(n13519), .ZN(n13407) );
  NAND2_X1 U15959 ( .A1(n13407), .A2(n12605), .ZN(n12608) );
  INV_X1 U15960 ( .A(n12606), .ZN(n12607) );
  MUX2_X1 U15961 ( .A(n12686), .B(n14276), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12609) );
  NOR2_X1 U15962 ( .A1(n12609), .A2(n9679), .ZN(n13499) );
  INV_X1 U15963 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n12610) );
  NAND2_X1 U15964 ( .A1(n12686), .A2(n12610), .ZN(n12613) );
  OAI211_X1 U15965 ( .C1(n12601), .C2(P1_EBX_REG_4__SCAN_IN), .A(n9633), .B(
        n12611), .ZN(n12612) );
  AND2_X1 U15966 ( .A1(n12613), .A2(n12612), .ZN(n13745) );
  INV_X1 U15967 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13854) );
  NAND2_X1 U15968 ( .A1(n12696), .A2(n13854), .ZN(n12617) );
  NAND2_X1 U15969 ( .A1(n9633), .A2(n12614), .ZN(n12615) );
  NAND2_X1 U15970 ( .A1(n12617), .A2(n12616), .ZN(n13746) );
  INV_X1 U15971 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n12618) );
  NAND2_X1 U15972 ( .A1(n12696), .A2(n12618), .ZN(n12622) );
  NAND2_X1 U15973 ( .A1(n9633), .A2(n12619), .ZN(n12620) );
  OAI21_X1 U15974 ( .B1(n12601), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12620), .ZN(
        n12621) );
  AND2_X1 U15975 ( .A1(n12622), .A2(n12621), .ZN(n13755) );
  INV_X1 U15976 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19853) );
  NAND2_X1 U15977 ( .A1(n12686), .A2(n19853), .ZN(n12626) );
  NAND2_X1 U15978 ( .A1(n12693), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12624) );
  OAI211_X1 U15979 ( .C1(n12601), .C2(P1_EBX_REG_6__SCAN_IN), .A(n9633), .B(
        n12624), .ZN(n12625) );
  AND2_X1 U15980 ( .A1(n12626), .A2(n12625), .ZN(n15933) );
  INV_X1 U15981 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13880) );
  NAND2_X1 U15982 ( .A1(n12686), .A2(n13880), .ZN(n12629) );
  NAND2_X1 U15983 ( .A1(n12693), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12627) );
  OAI211_X1 U15984 ( .C1(n12601), .C2(P1_EBX_REG_8__SCAN_IN), .A(n9633), .B(
        n12627), .ZN(n12628) );
  AND2_X1 U15985 ( .A1(n12629), .A2(n12628), .ZN(n13871) );
  INV_X1 U15986 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U15987 ( .A1(n12696), .A2(n13868), .ZN(n12633) );
  NAND2_X1 U15988 ( .A1(n12693), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12630) );
  NAND2_X1 U15989 ( .A1(n9633), .A2(n12630), .ZN(n12631) );
  OAI21_X1 U15990 ( .B1(n12601), .B2(P1_EBX_REG_7__SCAN_IN), .A(n12631), .ZN(
        n12632) );
  NAND2_X1 U15991 ( .A1(n12633), .A2(n12632), .ZN(n13872) );
  NAND2_X1 U15992 ( .A1(n13871), .A2(n13872), .ZN(n12634) );
  INV_X1 U15993 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U15994 ( .A1(n12696), .A2(n12635), .ZN(n12639) );
  NAND2_X1 U15995 ( .A1(n12693), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12636) );
  NAND2_X1 U15996 ( .A1(n9633), .A2(n12636), .ZN(n12637) );
  OAI21_X1 U15997 ( .B1(n12601), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12637), .ZN(
        n12638) );
  NOR2_X2 U15998 ( .A1(n13917), .A2(n13916), .ZN(n13987) );
  MUX2_X1 U15999 ( .A(n12694), .B(n12693), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12641) );
  INV_X1 U16000 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15917) );
  NAND2_X1 U16001 ( .A1(n15917), .A2(n12680), .ZN(n12640) );
  NAND2_X1 U16002 ( .A1(n12641), .A2(n12640), .ZN(n13989) );
  INV_X1 U16003 ( .A(n13989), .ZN(n12642) );
  INV_X1 U16004 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15797) );
  NAND2_X1 U16005 ( .A1(n12696), .A2(n15797), .ZN(n12646) );
  INV_X1 U16006 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12643) );
  NAND2_X1 U16007 ( .A1(n9633), .A2(n12643), .ZN(n12644) );
  OAI211_X1 U16008 ( .C1(n12601), .C2(P1_EBX_REG_11__SCAN_IN), .A(n12644), .B(
        n12693), .ZN(n12645) );
  INV_X1 U16009 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15769) );
  NAND2_X1 U16010 ( .A1(n12686), .A2(n15769), .ZN(n12649) );
  NAND2_X1 U16011 ( .A1(n12693), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12647) );
  OAI211_X1 U16012 ( .C1(n12601), .C2(P1_EBX_REG_12__SCAN_IN), .A(n9633), .B(
        n12647), .ZN(n12648) );
  NAND2_X1 U16013 ( .A1(n12649), .A2(n12648), .ZN(n14071) );
  NOR2_X1 U16014 ( .A1(n15780), .A2(n14071), .ZN(n12650) );
  INV_X1 U16015 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14099) );
  NAND2_X1 U16016 ( .A1(n12696), .A2(n14099), .ZN(n12653) );
  NAND2_X1 U16017 ( .A1(n9633), .A2(n14711), .ZN(n12651) );
  OAI211_X1 U16018 ( .C1(n12601), .C2(P1_EBX_REG_13__SCAN_IN), .A(n12651), .B(
        n12693), .ZN(n12652) );
  MUX2_X1 U16019 ( .A(n12694), .B(n12693), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12655) );
  NAND2_X1 U16020 ( .A1(n12680), .A2(n14704), .ZN(n12654) );
  NAND2_X1 U16021 ( .A1(n12655), .A2(n12654), .ZN(n14057) );
  INV_X1 U16022 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14113) );
  NAND2_X1 U16023 ( .A1(n12696), .A2(n14113), .ZN(n12658) );
  NAND2_X1 U16024 ( .A1(n9633), .A2(n15895), .ZN(n12656) );
  OAI211_X1 U16025 ( .C1(n12601), .C2(P1_EBX_REG_15__SCAN_IN), .A(n12656), .B(
        n12693), .ZN(n12657) );
  NAND2_X1 U16026 ( .A1(n12658), .A2(n12657), .ZN(n14110) );
  MUX2_X1 U16027 ( .A(n12686), .B(n14276), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12659) );
  NOR2_X1 U16028 ( .A1(n12659), .A2(n9700), .ZN(n14388) );
  NAND2_X1 U16029 ( .A1(n14389), .A2(n14388), .ZN(n14391) );
  INV_X1 U16030 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15731) );
  NAND2_X1 U16031 ( .A1(n12696), .A2(n15731), .ZN(n12662) );
  NAND2_X1 U16032 ( .A1(n9633), .A2(n14682), .ZN(n12660) );
  OAI211_X1 U16033 ( .C1(n12601), .C2(P1_EBX_REG_17__SCAN_IN), .A(n12660), .B(
        n12693), .ZN(n12661) );
  OR2_X2 U16034 ( .A1(n14391), .A2(n14380), .ZN(n14382) );
  MUX2_X1 U16035 ( .A(n12694), .B(n12693), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12664) );
  NAND2_X1 U16036 ( .A1(n12680), .A2(n12720), .ZN(n12663) );
  NAND2_X1 U16037 ( .A1(n12664), .A2(n12663), .ZN(n14374) );
  OR2_X2 U16038 ( .A1(n14382), .A2(n14374), .ZN(n14376) );
  INV_X1 U16039 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n20863) );
  NAND2_X1 U16040 ( .A1(n12696), .A2(n20863), .ZN(n12667) );
  NAND2_X1 U16041 ( .A1(n9633), .A2(n14663), .ZN(n12665) );
  OAI211_X1 U16042 ( .C1(n12601), .C2(P1_EBX_REG_19__SCAN_IN), .A(n12665), .B(
        n12693), .ZN(n12666) );
  NOR2_X2 U16043 ( .A1(n14376), .A2(n14316), .ZN(n14654) );
  INV_X1 U16044 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n20822) );
  NAND2_X1 U16045 ( .A1(n12686), .A2(n20822), .ZN(n12670) );
  NAND2_X1 U16046 ( .A1(n12693), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12668) );
  OAI211_X1 U16047 ( .C1(n12601), .C2(P1_EBX_REG_20__SCAN_IN), .A(n9633), .B(
        n12668), .ZN(n12669) );
  INV_X1 U16048 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14369) );
  NAND2_X1 U16049 ( .A1(n12696), .A2(n14369), .ZN(n12673) );
  NAND2_X1 U16050 ( .A1(n9633), .A2(n11611), .ZN(n12671) );
  OAI211_X1 U16051 ( .C1(n12601), .C2(P1_EBX_REG_21__SCAN_IN), .A(n12671), .B(
        n12693), .ZN(n12672) );
  NAND2_X1 U16052 ( .A1(n12673), .A2(n12672), .ZN(n14366) );
  MUX2_X1 U16053 ( .A(n12694), .B(n12693), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12676) );
  INV_X1 U16054 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12674) );
  NAND2_X1 U16055 ( .A1(n12680), .A2(n12674), .ZN(n12675) );
  INV_X1 U16056 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14356) );
  NAND2_X1 U16057 ( .A1(n12696), .A2(n14356), .ZN(n12679) );
  INV_X1 U16058 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14638) );
  NAND2_X1 U16059 ( .A1(n9633), .A2(n14638), .ZN(n12677) );
  OAI211_X1 U16060 ( .C1(n12601), .C2(P1_EBX_REG_23__SCAN_IN), .A(n12677), .B(
        n12693), .ZN(n12678) );
  MUX2_X1 U16061 ( .A(n12694), .B(n12693), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12682) );
  NAND2_X1 U16062 ( .A1(n12680), .A2(n14512), .ZN(n12681) );
  NAND2_X1 U16063 ( .A1(n12682), .A2(n12681), .ZN(n14348) );
  INV_X1 U16064 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15661) );
  NAND2_X1 U16065 ( .A1(n12696), .A2(n15661), .ZN(n12685) );
  NAND2_X1 U16066 ( .A1(n9633), .A2(n14621), .ZN(n12683) );
  OAI211_X1 U16067 ( .C1(n12601), .C2(P1_EBX_REG_25__SCAN_IN), .A(n12683), .B(
        n12693), .ZN(n12684) );
  NAND2_X1 U16068 ( .A1(n12685), .A2(n12684), .ZN(n14340) );
  AND2_X2 U16069 ( .A1(n14347), .A2(n14340), .ZN(n14612) );
  INV_X1 U16070 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15792) );
  NAND2_X1 U16071 ( .A1(n12686), .A2(n15792), .ZN(n12689) );
  NAND2_X1 U16072 ( .A1(n12693), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12687) );
  OAI211_X1 U16073 ( .C1(n12601), .C2(P1_EBX_REG_26__SCAN_IN), .A(n9633), .B(
        n12687), .ZN(n12688) );
  INV_X1 U16074 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14334) );
  NAND2_X1 U16075 ( .A1(n12696), .A2(n14334), .ZN(n12692) );
  NAND2_X1 U16076 ( .A1(n9633), .A2(n11616), .ZN(n12690) );
  OAI211_X1 U16077 ( .C1(n12601), .C2(P1_EBX_REG_27__SCAN_IN), .A(n12690), .B(
        n12693), .ZN(n12691) );
  AND2_X1 U16078 ( .A1(n12692), .A2(n12691), .ZN(n14300) );
  MUX2_X1 U16079 ( .A(n12694), .B(n12693), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12695) );
  INV_X1 U16080 ( .A(n12696), .ZN(n12697) );
  OAI22_X1 U16081 ( .A1(n14274), .A2(n14276), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12697), .ZN(n14219) );
  MUX2_X1 U16082 ( .A(n12699), .B(n12698), .S(n14277), .Z(n14329) );
  INV_X1 U16083 ( .A(n14329), .ZN(n12741) );
  OR2_X1 U16084 ( .A1(n12700), .A2(n20025), .ZN(n15604) );
  OAI21_X1 U16085 ( .B1(n12701), .B2(n20036), .A(n15604), .ZN(n12702) );
  INV_X1 U16086 ( .A(n14257), .ZN(n12703) );
  AOI22_X1 U16087 ( .A1(n12703), .A2(n11321), .B1(n13557), .B2(n20025), .ZN(
        n12708) );
  NAND2_X1 U16088 ( .A1(n12704), .A2(n14276), .ZN(n12707) );
  NAND2_X1 U16089 ( .A1(n13425), .A2(n20012), .ZN(n12705) );
  NAND2_X1 U16090 ( .A1(n12705), .A2(n20029), .ZN(n12706) );
  AND4_X1 U16091 ( .A1(n12709), .A2(n12708), .A3(n12707), .A4(n12706), .ZN(
        n12712) );
  INV_X1 U16092 ( .A(n12710), .ZN(n12711) );
  OAI211_X1 U16093 ( .C1(n12713), .C2(n13421), .A(n12712), .B(n12711), .ZN(
        n13470) );
  OAI21_X1 U16094 ( .B1(n13467), .B2(n13399), .A(n12714), .ZN(n12715) );
  OR2_X1 U16095 ( .A1(n13470), .A2(n12715), .ZN(n12716) );
  OR2_X1 U16096 ( .A1(n12718), .A2(n12717), .ZN(n14243) );
  INV_X1 U16097 ( .A(n14243), .ZN(n12719) );
  NAND2_X1 U16098 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13838) );
  NAND2_X1 U16099 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19948) );
  OR2_X1 U16100 ( .A1(n20804), .A2(n19948), .ZN(n14041) );
  NOR2_X1 U16101 ( .A1(n13838), .A2(n14041), .ZN(n14732) );
  INV_X1 U16102 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15941) );
  NAND2_X1 U16103 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15919) );
  NOR2_X1 U16104 ( .A1(n15941), .A2(n15919), .ZN(n14042) );
  NAND3_X1 U16105 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n14042), .ZN(n14735) );
  NOR2_X1 U16106 ( .A1(n12643), .A2(n14735), .ZN(n14729) );
  NAND3_X1 U16107 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14732), .A3(
        n14729), .ZN(n14685) );
  INV_X1 U16108 ( .A(n14685), .ZN(n14717) );
  NAND3_X1 U16109 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15884) );
  NOR4_X1 U16110 ( .A1(n12720), .A2(n14711), .A3(n14704), .A4(n15884), .ZN(
        n14657) );
  NAND2_X1 U16111 ( .A1(n14717), .A2(n14657), .ZN(n14662) );
  AOI21_X1 U16112 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13837) );
  NOR2_X1 U16113 ( .A1(n13837), .A2(n14041), .ZN(n14043) );
  NAND2_X1 U16114 ( .A1(n14729), .A2(n14043), .ZN(n14734) );
  NOR2_X1 U16115 ( .A1(n20856), .A2(n14734), .ZN(n14687) );
  NAND2_X1 U16116 ( .A1(n14657), .A2(n14687), .ZN(n14660) );
  NAND2_X1 U16117 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12721) );
  AOI211_X1 U16118 ( .C1(n14662), .C2(n14661), .A(n14660), .B(n12721), .ZN(
        n12722) );
  OR2_X1 U16119 ( .A1(n12722), .A2(n15922), .ZN(n12726) );
  INV_X1 U16120 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20798) );
  NAND2_X1 U16121 ( .A1(n19991), .A2(n20798), .ZN(n12725) );
  OR2_X1 U16122 ( .A1(n12723), .A2(n19977), .ZN(n12724) );
  NAND2_X1 U16123 ( .A1(n12725), .A2(n12724), .ZN(n19981) );
  INV_X1 U16124 ( .A(n19981), .ZN(n14664) );
  AND2_X1 U16125 ( .A1(n12726), .A2(n14664), .ZN(n14644) );
  NAND2_X1 U16126 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15877) );
  NAND2_X1 U16127 ( .A1(n19986), .A2(n15877), .ZN(n12727) );
  AND2_X1 U16128 ( .A1(n14644), .A2(n12727), .ZN(n14637) );
  OR2_X1 U16129 ( .A1(n19992), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12728) );
  AND2_X1 U16130 ( .A1(n14637), .A2(n12728), .ZN(n14631) );
  OR2_X1 U16131 ( .A1(n19968), .A2(n20001), .ZN(n12730) );
  INV_X1 U16132 ( .A(n12729), .ZN(n14471) );
  AOI22_X1 U16133 ( .A1(n12730), .A2(n14471), .B1(n19991), .B2(n12734), .ZN(
        n12731) );
  NAND2_X1 U16134 ( .A1(n14610), .A2(n15922), .ZN(n12733) );
  NAND2_X1 U16135 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14615) );
  NAND2_X1 U16136 ( .A1(n19986), .A2(n14615), .ZN(n12732) );
  NAND2_X1 U16137 ( .A1(n14610), .A2(n12732), .ZN(n14607) );
  AOI21_X1 U16138 ( .B1(n12736), .B2(n12733), .A(n14607), .ZN(n14586) );
  OAI211_X1 U16139 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15922), .A(
        n14586), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14579) );
  NAND3_X1 U16140 ( .A1(n14579), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12733), .ZN(n12739) );
  NAND2_X1 U16141 ( .A1(n19977), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14449) );
  NAND2_X1 U16142 ( .A1(n19968), .A2(n14687), .ZN(n14658) );
  NAND3_X1 U16143 ( .A1(n14657), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14713), .ZN(n14669) );
  NOR2_X1 U16144 ( .A1(n14668), .A2(n14669), .ZN(n15878) );
  NAND3_X1 U16145 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n15878), .ZN(n14639) );
  NOR2_X1 U16146 ( .A1(n12734), .A2(n14639), .ZN(n14622) );
  INV_X1 U16147 ( .A(n14615), .ZN(n12735) );
  NAND2_X1 U16148 ( .A1(n14622), .A2(n12735), .ZN(n14603) );
  NOR2_X1 U16149 ( .A1(n14603), .A2(n12736), .ZN(n14587) );
  INV_X1 U16150 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12737) );
  NAND4_X1 U16151 ( .A1(n14587), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n12737), .ZN(n12738) );
  NAND3_X1 U16152 ( .A1(n12739), .A2(n14449), .A3(n12738), .ZN(n12740) );
  AOI21_X1 U16153 ( .B1(n12741), .B2(n19979), .A(n12740), .ZN(n12742) );
  OAI21_X1 U16154 ( .B1(n14454), .B2(n19996), .A(n12742), .ZN(P1_U3000) );
  INV_X1 U16155 ( .A(n12743), .ZN(n13321) );
  NAND2_X1 U16156 ( .A1(n13321), .A2(n13231), .ZN(n12744) );
  MUX2_X1 U16157 ( .A(n12744), .B(n19731), .S(n12748), .Z(n12757) );
  NAND2_X1 U16158 ( .A1(n12747), .A2(n12748), .ZN(n12755) );
  NAND2_X1 U16159 ( .A1(n12750), .A2(n12749), .ZN(n12753) );
  INV_X1 U16160 ( .A(n12751), .ZN(n12752) );
  NAND3_X1 U16161 ( .A1(n12753), .A2(n19028), .A3(n12752), .ZN(n12754) );
  OAI211_X1 U16162 ( .C1(n10086), .C2(n19731), .A(n12755), .B(n12754), .ZN(
        n12756) );
  NAND2_X1 U16163 ( .A1(n12757), .A2(n12756), .ZN(n12759) );
  MUX2_X1 U16164 ( .A(n19731), .B(n12759), .S(n12758), .Z(n12760) );
  NAND2_X1 U16165 ( .A1(n12760), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12761) );
  NOR2_X1 U16166 ( .A1(n12762), .A2(n12761), .ZN(n12763) );
  NAND2_X1 U16167 ( .A1(n19752), .A2(n19747), .ZN(n13229) );
  NAND2_X1 U16168 ( .A1(n12767), .A2(n19045), .ZN(n12771) );
  NAND2_X1 U16169 ( .A1(n12769), .A2(n12768), .ZN(n12770) );
  AOI21_X1 U16170 ( .B1(n12766), .B2(n12771), .A(n12770), .ZN(n12781) );
  OR2_X1 U16171 ( .A1(n12772), .A2(n19071), .ZN(n12773) );
  NAND2_X1 U16172 ( .A1(n12773), .A2(n19734), .ZN(n12812) );
  INV_X1 U16173 ( .A(n13229), .ZN(n12775) );
  NAND3_X1 U16174 ( .A1(n12774), .A2(n13633), .A3(n12775), .ZN(n12780) );
  NAND2_X1 U16175 ( .A1(n12776), .A2(n12785), .ZN(n12794) );
  NAND2_X1 U16176 ( .A1(n12794), .A2(n19028), .ZN(n12777) );
  NAND2_X1 U16177 ( .A1(n12777), .A2(n13188), .ZN(n12778) );
  NAND2_X1 U16178 ( .A1(n12778), .A2(n19045), .ZN(n12779) );
  MUX2_X1 U16179 ( .A(n12774), .B(n12819), .S(n12750), .Z(n12782) );
  NAND3_X1 U16180 ( .A1(n12782), .A2(n13633), .A3(n19747), .ZN(n12783) );
  AND3_X1 U16181 ( .A1(n12784), .A2(n13454), .A3(n12783), .ZN(n12787) );
  OAI211_X1 U16182 ( .C1(n13645), .C2(n13631), .A(n13319), .B(n12785), .ZN(
        n12786) );
  OAI211_X1 U16183 ( .C1(n13459), .C2(n19045), .A(n12787), .B(n12786), .ZN(
        n12788) );
  INV_X1 U16184 ( .A(n12850), .ZN(n12790) );
  NOR2_X1 U16185 ( .A1(n19737), .A2(n19731), .ZN(n12789) );
  AOI21_X1 U16186 ( .B1(n13656), .B2(n12750), .A(n12792), .ZN(n12793) );
  OR2_X1 U16187 ( .A1(n12794), .A2(n19071), .ZN(n12798) );
  NAND3_X1 U16188 ( .A1(n13334), .A2(n12795), .A3(n12750), .ZN(n12796) );
  MUX2_X1 U16189 ( .A(n12796), .B(n13334), .S(n10610), .Z(n12797) );
  INV_X1 U16190 ( .A(n12799), .ZN(n12800) );
  NAND2_X1 U16191 ( .A1(n13650), .A2(n12800), .ZN(n13634) );
  NAND2_X1 U16192 ( .A1(n13632), .A2(n13231), .ZN(n12801) );
  AND2_X1 U16193 ( .A1(n13634), .A2(n12801), .ZN(n12802) );
  AOI222_X1 U16194 ( .A1(n12804), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n10838), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n12803), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n12805) );
  XNOR2_X1 U16195 ( .A(n12806), .B(n12805), .ZN(n18904) );
  INV_X1 U16196 ( .A(n12807), .ZN(n12831) );
  AND3_X1 U16197 ( .A1(n19045), .A2(n12750), .A3(n12808), .ZN(n12809) );
  NAND2_X1 U16198 ( .A1(n13650), .A2(n12809), .ZN(n13441) );
  NOR2_X1 U16199 ( .A1(n15446), .A2(n13370), .ZN(n19009) );
  INV_X1 U16200 ( .A(n19009), .ZN(n19001) );
  NOR2_X1 U16201 ( .A1(n12810), .A2(n19001), .ZN(n12834) );
  NOR2_X1 U16202 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19009), .ZN(
        n12836) );
  INV_X1 U16203 ( .A(n12836), .ZN(n12827) );
  NAND2_X1 U16204 ( .A1(n12811), .A2(n13231), .ZN(n13648) );
  NAND2_X1 U16205 ( .A1(n13648), .A2(n12812), .ZN(n12813) );
  NAND2_X1 U16206 ( .A1(n12813), .A2(n10610), .ZN(n12825) );
  MUX2_X1 U16207 ( .A(n13639), .B(n12814), .S(n10622), .Z(n12815) );
  NAND2_X1 U16208 ( .A1(n12815), .A2(n12776), .ZN(n12817) );
  NAND2_X1 U16209 ( .A1(n12817), .A2(n12816), .ZN(n12824) );
  NOR2_X1 U16210 ( .A1(n12776), .A2(n19055), .ZN(n12818) );
  AOI21_X1 U16211 ( .B1(n12766), .B2(n12819), .A(n12818), .ZN(n12823) );
  NAND3_X1 U16212 ( .A1(n12820), .A2(n19028), .A3(n12821), .ZN(n12822) );
  NAND4_X1 U16213 ( .A1(n12825), .A2(n12824), .A3(n12823), .A4(n12822), .ZN(
        n13185) );
  INV_X1 U16214 ( .A(n10622), .ZN(n13186) );
  NOR2_X1 U16215 ( .A1(n13185), .A2(n13186), .ZN(n12826) );
  NOR2_X1 U16216 ( .A1(n12850), .A2(n12826), .ZN(n19002) );
  OAI211_X1 U16217 ( .C1(n19000), .C2(n12834), .A(n12827), .B(n15452), .ZN(
        n16154) );
  NAND2_X1 U16218 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15434) );
  NOR2_X1 U16219 ( .A1(n12828), .A2(n15434), .ZN(n12837) );
  NAND2_X1 U16220 ( .A1(n15435), .A2(n12837), .ZN(n16135) );
  NAND2_X1 U16221 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14179) );
  NAND2_X1 U16222 ( .A1(n15085), .A2(n15413), .ZN(n15276) );
  NOR2_X1 U16223 ( .A1(n15275), .A2(n15276), .ZN(n15643) );
  NOR2_X1 U16224 ( .A1(n15636), .A2(n15259), .ZN(n12838) );
  NAND2_X1 U16225 ( .A1(n15643), .A2(n12838), .ZN(n15237) );
  NOR2_X1 U16226 ( .A1(n15227), .A2(n15237), .ZN(n15219) );
  NAND2_X1 U16227 ( .A1(n12840), .A2(n15219), .ZN(n15194) );
  NOR2_X1 U16228 ( .A1(n15194), .A2(n15195), .ZN(n15181) );
  NAND2_X1 U16229 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12842) );
  INV_X1 U16230 ( .A(n12842), .ZN(n12829) );
  NAND2_X1 U16231 ( .A1(n15181), .A2(n12829), .ZN(n15131) );
  NAND3_X1 U16232 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14197) );
  NOR4_X1 U16233 ( .A1(n15131), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14201), .A4(n14197), .ZN(n12830) );
  AOI211_X1 U16234 ( .C1(n18993), .C2(n18904), .A(n12831), .B(n12830), .ZN(
        n12832) );
  INV_X1 U16235 ( .A(n15452), .ZN(n15293) );
  AND2_X1 U16236 ( .A1(n12850), .A2(n19017), .ZN(n13363) );
  INV_X1 U16237 ( .A(n12834), .ZN(n12835) );
  AND2_X1 U16238 ( .A1(n19002), .A2(n12835), .ZN(n19010) );
  AND2_X1 U16239 ( .A1(n19000), .A2(n12836), .ZN(n18999) );
  NOR4_X1 U16240 ( .A1(n19010), .A2(n13363), .A3(n18999), .A4(n16155), .ZN(
        n16156) );
  NAND2_X1 U16241 ( .A1(n12837), .A2(n16156), .ZN(n14177) );
  NOR2_X1 U16242 ( .A1(n14179), .A2(n14177), .ZN(n15409) );
  INV_X1 U16243 ( .A(n12838), .ZN(n15642) );
  NOR3_X1 U16244 ( .A1(n15227), .A2(n12839), .A3(n15642), .ZN(n15203) );
  NAND3_X1 U16245 ( .A1(n12840), .A2(n15409), .A3(n15203), .ZN(n12841) );
  AOI21_X1 U16246 ( .B1(n14178), .B2(n12841), .A(n15195), .ZN(n15193) );
  OR2_X1 U16247 ( .A1(n15193), .A2(n15410), .ZN(n15188) );
  NAND2_X1 U16248 ( .A1(n14178), .A2(n12842), .ZN(n12843) );
  NAND2_X1 U16249 ( .A1(n15188), .A2(n12843), .ZN(n15162) );
  AND2_X1 U16250 ( .A1(n15452), .A2(n14197), .ZN(n12844) );
  NOR2_X1 U16251 ( .A1(n15162), .A2(n12844), .ZN(n14202) );
  OAI21_X1 U16252 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15293), .A(
        n14202), .ZN(n12845) );
  INV_X1 U16253 ( .A(n12845), .ZN(n12847) );
  NAND2_X1 U16254 ( .A1(n13646), .A2(n19734), .ZN(n12849) );
  NAND2_X1 U16255 ( .A1(n13165), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12853) );
  NAND2_X1 U16256 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19378) );
  NAND2_X1 U16257 ( .A1(n19378), .A2(n19710), .ZN(n12855) );
  NAND2_X1 U16258 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19548) );
  INV_X1 U16259 ( .A(n19548), .ZN(n12854) );
  NAND2_X1 U16260 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12854), .ZN(
        n19020) );
  NAND2_X1 U16261 ( .A1(n12855), .A2(n19020), .ZN(n19175) );
  NOR2_X1 U16262 ( .A1(n19175), .A2(n19416), .ZN(n19409) );
  AOI21_X1 U16263 ( .B1(n12872), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n19409), .ZN(n12856) );
  NOR2_X1 U16264 ( .A1(n13165), .A2(n19751), .ZN(n13340) );
  OAI21_X1 U16265 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19378), .ZN(n19408) );
  OR2_X1 U16266 ( .A1(n19408), .A2(n19416), .ZN(n19348) );
  INV_X1 U16267 ( .A(n19348), .ZN(n19111) );
  AOI21_X1 U16268 ( .B1(n12872), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19111), .ZN(n12861) );
  NOR2_X1 U16269 ( .A1(n19416), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12863) );
  INV_X1 U16270 ( .A(n13099), .ZN(n12865) );
  OR2_X1 U16271 ( .A1(n12865), .A2(n19044), .ZN(n12866) );
  NAND2_X1 U16272 ( .A1(n13375), .A2(n13374), .ZN(n12868) );
  INV_X1 U16273 ( .A(n13345), .ZN(n14006) );
  NAND2_X1 U16274 ( .A1(n14006), .A2(n12866), .ZN(n12867) );
  NAND2_X1 U16275 ( .A1(n19020), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12870) );
  NOR2_X1 U16276 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19548), .ZN(
        n19265) );
  NAND2_X1 U16277 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19265), .ZN(
        n19290) );
  NAND2_X1 U16278 ( .A1(n12870), .A2(n19290), .ZN(n12871) );
  AOI22_X1 U16279 ( .A1(n12872), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19690), .B2(n12871), .ZN(n12873) );
  INV_X1 U16280 ( .A(n12881), .ZN(n12878) );
  INV_X1 U16281 ( .A(n12876), .ZN(n12877) );
  NAND2_X1 U16282 ( .A1(n12878), .A2(n12877), .ZN(n12879) );
  NAND2_X1 U16283 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13165), .ZN(
        n12880) );
  NAND2_X1 U16284 ( .A1(n12881), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12882) );
  AND2_X1 U16285 ( .A1(n13099), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13779) );
  AND2_X1 U16286 ( .A1(n18883), .A2(n18884), .ZN(n12885) );
  NAND2_X1 U16287 ( .A1(n18890), .A2(n18891), .ZN(n12884) );
  INV_X1 U16288 ( .A(n13550), .ZN(n12883) );
  INV_X1 U16289 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19081) );
  NAND2_X1 U16290 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13528) );
  OR2_X1 U16291 ( .A1(n19081), .A2(n13528), .ZN(n13548) );
  NOR2_X1 U16292 ( .A1(n12884), .A2(n13538), .ZN(n13589) );
  AOI22_X1 U16293 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16294 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16295 ( .A1(n9619), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U16296 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12887) );
  NAND4_X1 U16297 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n12887), .ZN(
        n12898) );
  AOI22_X1 U16298 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U16299 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U16300 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12891) );
  AND2_X1 U16301 ( .A1(n12892), .A2(n12891), .ZN(n12895) );
  AOI22_X1 U16302 ( .A1(n13012), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U16303 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12893) );
  NAND4_X1 U16304 ( .A1(n12896), .A2(n12895), .A3(n12894), .A4(n12893), .ZN(
        n12897) );
  AOI22_X1 U16305 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U16306 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U16307 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U16308 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12899) );
  NAND4_X1 U16309 ( .A1(n12902), .A2(n12901), .A3(n12900), .A4(n12899), .ZN(
        n12910) );
  AOI22_X1 U16310 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U16311 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U16312 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12903) );
  AND2_X1 U16313 ( .A1(n12904), .A2(n12903), .ZN(n12907) );
  AOI22_X1 U16314 ( .A1(n13012), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12906) );
  NAND2_X1 U16315 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12905) );
  NAND4_X1 U16316 ( .A1(n12908), .A2(n12907), .A3(n12906), .A4(n12905), .ZN(
        n12909) );
  NAND2_X1 U16317 ( .A1(n13991), .A2(n13993), .ZN(n13992) );
  INV_X1 U16318 ( .A(n13992), .ZN(n12924) );
  AOI22_X1 U16319 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10904), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U16320 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12913) );
  AOI22_X1 U16321 ( .A1(n9619), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12912) );
  AOI22_X1 U16322 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12911) );
  NAND4_X1 U16323 ( .A1(n12914), .A2(n12913), .A3(n12912), .A4(n12911), .ZN(
        n12922) );
  AOI22_X1 U16324 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U16325 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12916) );
  NAND2_X1 U16326 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12915) );
  AND2_X1 U16327 ( .A1(n12916), .A2(n12915), .ZN(n12919) );
  AOI22_X1 U16328 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12918) );
  NAND2_X1 U16329 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12917) );
  NAND4_X1 U16330 ( .A1(n12920), .A2(n12919), .A3(n12918), .A4(n12917), .ZN(
        n12921) );
  NOR2_X1 U16331 ( .A1(n12922), .A2(n12921), .ZN(n16014) );
  INV_X1 U16332 ( .A(n16014), .ZN(n12923) );
  AOI22_X1 U16333 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10904), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U16334 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U16335 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U16336 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12925) );
  NAND4_X1 U16337 ( .A1(n12928), .A2(n12927), .A3(n12926), .A4(n12925), .ZN(
        n12936) );
  AOI22_X1 U16338 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U16339 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12930) );
  NAND2_X1 U16340 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12929) );
  AND2_X1 U16341 ( .A1(n12930), .A2(n12929), .ZN(n12933) );
  AOI22_X1 U16342 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12932) );
  NAND2_X1 U16343 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12931) );
  NAND4_X1 U16344 ( .A1(n12934), .A2(n12933), .A3(n12932), .A4(n12931), .ZN(
        n12935) );
  NOR2_X1 U16345 ( .A1(n12936), .A2(n12935), .ZN(n14880) );
  AOI22_X1 U16346 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10904), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16347 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U16348 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U16349 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12937) );
  NAND4_X1 U16350 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        n12948) );
  AOI22_X1 U16351 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U16352 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12942) );
  NAND2_X1 U16353 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12941) );
  AND2_X1 U16354 ( .A1(n12942), .A2(n12941), .ZN(n12945) );
  AOI22_X1 U16355 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12944) );
  NAND2_X1 U16356 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12943) );
  NAND4_X1 U16357 ( .A1(n12946), .A2(n12945), .A3(n12944), .A4(n12943), .ZN(
        n12947) );
  OR2_X1 U16358 ( .A1(n12948), .A2(n12947), .ZN(n16010) );
  INV_X1 U16359 ( .A(n13012), .ZN(n12952) );
  INV_X1 U16360 ( .A(n13011), .ZN(n12950) );
  OAI22_X1 U16361 ( .A1(n12952), .A2(n12951), .B1(n12950), .B2(n12949), .ZN(
        n12957) );
  INV_X1 U16362 ( .A(n12953), .ZN(n12976) );
  INV_X1 U16363 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U16364 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12954) );
  OAI21_X1 U16365 ( .B1(n12976), .B2(n12955), .A(n12954), .ZN(n12956) );
  AOI211_X1 U16366 ( .C1(n13013), .C2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n12957), .B(n12956), .ZN(n12964) );
  AOI22_X1 U16367 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16368 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12961) );
  AOI22_X1 U16369 ( .A1(n10870), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12960) );
  AOI22_X1 U16370 ( .A1(n9619), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U16371 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12958) );
  AND4_X1 U16372 ( .A1(n12961), .A2(n12960), .A3(n12959), .A4(n12958), .ZN(
        n12962) );
  NAND3_X1 U16373 ( .A1(n12964), .A2(n12963), .A3(n12962), .ZN(n14874) );
  AOI22_X1 U16374 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10904), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U16375 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16376 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12966) );
  AOI22_X1 U16377 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12965) );
  NAND4_X1 U16378 ( .A1(n12968), .A2(n12967), .A3(n12966), .A4(n12965), .ZN(
        n12983) );
  INV_X1 U16379 ( .A(n13007), .ZN(n12973) );
  INV_X1 U16380 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12972) );
  INV_X1 U16381 ( .A(n12969), .ZN(n12971) );
  OAI22_X1 U16382 ( .A1(n12973), .A2(n12972), .B1(n12971), .B2(n12970), .ZN(
        n12982) );
  INV_X1 U16383 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U16384 ( .A1(n10875), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12974) );
  OAI21_X1 U16385 ( .B1(n12976), .B2(n12975), .A(n12974), .ZN(n12981) );
  INV_X1 U16386 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12979) );
  AOI22_X1 U16387 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12977) );
  OAI21_X1 U16388 ( .B1(n12979), .B2(n12978), .A(n12977), .ZN(n12980) );
  AOI22_X1 U16389 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16390 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16391 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U16392 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12989) );
  INV_X1 U16393 ( .A(n13443), .ZN(n12987) );
  INV_X1 U16394 ( .A(n12985), .ZN(n12986) );
  NAND2_X1 U16395 ( .A1(n12987), .A2(n12986), .ZN(n13142) );
  NAND2_X1 U16396 ( .A1(n13141), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12988) );
  AND3_X1 U16397 ( .A1(n12989), .A2(n13142), .A3(n12988), .ZN(n12990) );
  NAND4_X1 U16398 ( .A1(n12993), .A2(n12992), .A3(n12991), .A4(n12990), .ZN(
        n13001) );
  AOI22_X1 U16399 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U16400 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16401 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12997) );
  INV_X1 U16402 ( .A(n13142), .ZN(n13152) );
  NAND2_X1 U16403 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12995) );
  NAND2_X1 U16404 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12994) );
  AND3_X1 U16405 ( .A1(n13152), .A2(n12995), .A3(n12994), .ZN(n12996) );
  NAND4_X1 U16406 ( .A1(n12999), .A2(n12998), .A3(n12997), .A4(n12996), .ZN(
        n13000) );
  AND2_X1 U16407 ( .A1(n13001), .A2(n13000), .ZN(n13037) );
  NAND2_X1 U16408 ( .A1(n13231), .A2(n13037), .ZN(n13036) );
  AOI22_X1 U16409 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10904), .B1(
        n13002), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U16410 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10870), .B1(
        n10920), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U16411 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10856), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16412 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13439), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13003) );
  NAND4_X1 U16413 ( .A1(n13006), .A2(n13005), .A3(n13004), .A4(n13003), .ZN(
        n13019) );
  AOI22_X1 U16414 ( .A1(n13007), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U16415 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10875), .B1(
        n13008), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13010) );
  NAND2_X1 U16416 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13009) );
  AND2_X1 U16417 ( .A1(n13010), .A2(n13009), .ZN(n13016) );
  AOI22_X1 U16418 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13012), .B1(
        n13011), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13015) );
  NAND2_X1 U16419 ( .A1(n13013), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13014) );
  NAND4_X1 U16420 ( .A1(n13017), .A2(n13016), .A3(n13015), .A4(n13014), .ZN(
        n13018) );
  NOR2_X1 U16421 ( .A1(n13019), .A2(n13018), .ZN(n13039) );
  NAND2_X1 U16422 ( .A1(n12750), .A2(n13037), .ZN(n14867) );
  AOI22_X1 U16423 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U16424 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U16425 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13024) );
  NAND2_X1 U16426 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13022) );
  NAND2_X1 U16427 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13021) );
  AND3_X1 U16428 ( .A1(n13022), .A2(n13142), .A3(n13021), .ZN(n13023) );
  NAND4_X1 U16429 ( .A1(n13026), .A2(n13025), .A3(n13024), .A4(n13023), .ZN(
        n13035) );
  AOI22_X1 U16430 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U16431 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U16432 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13031) );
  INV_X1 U16433 ( .A(n13027), .ZN(n13140) );
  NAND2_X1 U16434 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13029) );
  NAND2_X1 U16435 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13028) );
  AND3_X1 U16436 ( .A1(n13152), .A2(n13029), .A3(n13028), .ZN(n13030) );
  NAND4_X1 U16437 ( .A1(n13033), .A2(n13032), .A3(n13031), .A4(n13030), .ZN(
        n13034) );
  NAND2_X1 U16438 ( .A1(n13035), .A2(n13034), .ZN(n13042) );
  OAI21_X1 U16439 ( .B1(n13036), .B2(n13039), .A(n13042), .ZN(n13044) );
  INV_X1 U16440 ( .A(n13037), .ZN(n13038) );
  NOR2_X1 U16441 ( .A1(n13042), .A2(n13038), .ZN(n13041) );
  INV_X1 U16442 ( .A(n13039), .ZN(n13040) );
  NAND2_X1 U16443 ( .A1(n13041), .A2(n13040), .ZN(n13059) );
  INV_X1 U16444 ( .A(n13042), .ZN(n13043) );
  AOI22_X1 U16445 ( .A1(n13044), .A2(n13059), .B1(n13043), .B2(n12750), .ZN(
        n14857) );
  AOI22_X1 U16446 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16447 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U16448 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13048) );
  NAND2_X1 U16449 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13046) );
  NAND2_X1 U16450 ( .A1(n13141), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13045) );
  AND3_X1 U16451 ( .A1(n13046), .A2(n13142), .A3(n13045), .ZN(n13047) );
  NAND4_X1 U16452 ( .A1(n13050), .A2(n13049), .A3(n13048), .A4(n13047), .ZN(
        n13058) );
  AOI22_X1 U16453 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U16454 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16455 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U16456 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13052) );
  NAND2_X1 U16457 ( .A1(n13141), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13051) );
  AND3_X1 U16458 ( .A1(n13152), .A2(n13052), .A3(n13051), .ZN(n13053) );
  NAND4_X1 U16459 ( .A1(n13056), .A2(n13055), .A3(n13054), .A4(n13053), .ZN(
        n13057) );
  AND2_X1 U16460 ( .A1(n13058), .A2(n13057), .ZN(n13061) );
  INV_X1 U16461 ( .A(n13059), .ZN(n13060) );
  NAND2_X1 U16462 ( .A1(n13060), .A2(n13061), .ZN(n13084) );
  OAI211_X1 U16463 ( .C1(n13061), .C2(n13060), .A(n13099), .B(n13084), .ZN(
        n13063) );
  INV_X1 U16464 ( .A(n13061), .ZN(n13062) );
  NOR2_X1 U16465 ( .A1(n13231), .A2(n13062), .ZN(n14920) );
  INV_X1 U16466 ( .A(n14856), .ZN(n13064) );
  AOI22_X1 U16467 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16468 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U16469 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13069) );
  NAND2_X1 U16470 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n13067) );
  NAND2_X1 U16471 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13066) );
  AND3_X1 U16472 ( .A1(n13067), .A2(n13142), .A3(n13066), .ZN(n13068) );
  NAND4_X1 U16473 ( .A1(n13071), .A2(n13070), .A3(n13069), .A4(n13068), .ZN(
        n13079) );
  AOI22_X1 U16474 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U16475 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U16476 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13075) );
  NAND2_X1 U16477 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n13073) );
  NAND2_X1 U16478 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13072) );
  AND3_X1 U16479 ( .A1(n13152), .A2(n13073), .A3(n13072), .ZN(n13074) );
  NAND4_X1 U16480 ( .A1(n13077), .A2(n13076), .A3(n13075), .A4(n13074), .ZN(
        n13078) );
  AND2_X1 U16481 ( .A1(n13079), .A2(n13078), .ZN(n13082) );
  XNOR2_X1 U16482 ( .A(n13084), .B(n13082), .ZN(n13080) );
  NAND2_X1 U16483 ( .A1(n12750), .A2(n13082), .ZN(n14852) );
  INV_X1 U16484 ( .A(n13082), .ZN(n13083) );
  NOR2_X1 U16485 ( .A1(n13084), .A2(n13083), .ZN(n13100) );
  AOI22_X1 U16486 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16487 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U16488 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13088) );
  NAND2_X1 U16489 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n13086) );
  NAND2_X1 U16490 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13085) );
  AND3_X1 U16491 ( .A1(n13086), .A2(n13142), .A3(n13085), .ZN(n13087) );
  NAND4_X1 U16492 ( .A1(n13090), .A2(n13089), .A3(n13088), .A4(n13087), .ZN(
        n13098) );
  AOI22_X1 U16493 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U16494 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16495 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13094) );
  NAND2_X1 U16496 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13092) );
  NAND2_X1 U16497 ( .A1(n13141), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13091) );
  AND3_X1 U16498 ( .A1(n13152), .A2(n13092), .A3(n13091), .ZN(n13093) );
  NAND4_X1 U16499 ( .A1(n13096), .A2(n13095), .A3(n13094), .A4(n13093), .ZN(
        n13097) );
  AND2_X1 U16500 ( .A1(n13098), .A2(n13097), .ZN(n13102) );
  NAND2_X1 U16501 ( .A1(n13100), .A2(n13102), .ZN(n14836) );
  OAI211_X1 U16502 ( .C1(n13100), .C2(n13102), .A(n14836), .B(n13099), .ZN(
        n13101) );
  INV_X1 U16503 ( .A(n13102), .ZN(n13103) );
  NOR2_X1 U16504 ( .A1(n13231), .A2(n13103), .ZN(n14844) );
  NAND2_X1 U16505 ( .A1(n14842), .A2(n14844), .ZN(n14843) );
  INV_X1 U16506 ( .A(n13104), .ZN(n14837) );
  AOI22_X1 U16507 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13110) );
  AOI22_X1 U16508 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U16509 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13108) );
  NAND2_X1 U16510 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n13106) );
  NAND2_X1 U16511 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13105) );
  AND3_X1 U16512 ( .A1(n13106), .A2(n13142), .A3(n13105), .ZN(n13107) );
  NAND4_X1 U16513 ( .A1(n13110), .A2(n13109), .A3(n13108), .A4(n13107), .ZN(
        n13118) );
  AOI22_X1 U16514 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16515 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U16516 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13114) );
  NAND2_X1 U16517 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n13112) );
  NAND2_X1 U16518 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13111) );
  AND3_X1 U16519 ( .A1(n13152), .A2(n13112), .A3(n13111), .ZN(n13113) );
  NAND4_X1 U16520 ( .A1(n13116), .A2(n13115), .A3(n13114), .A4(n13113), .ZN(
        n13117) );
  NAND2_X1 U16521 ( .A1(n13118), .A2(n13117), .ZN(n14839) );
  AOI22_X1 U16522 ( .A1(n10813), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13124) );
  NAND2_X1 U16523 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n13120) );
  NAND2_X1 U16524 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n13119) );
  AND3_X1 U16525 ( .A1(n13120), .A2(n13142), .A3(n13119), .ZN(n13123) );
  AOI22_X1 U16526 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16527 ( .A1(n13615), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13121) );
  NAND4_X1 U16528 ( .A1(n13124), .A2(n13123), .A3(n13122), .A4(n13121), .ZN(
        n13132) );
  AOI22_X1 U16529 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U16530 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10813), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U16531 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13128) );
  NAND2_X1 U16532 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n13126) );
  NAND2_X1 U16533 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n13125) );
  AND3_X1 U16534 ( .A1(n13152), .A2(n13126), .A3(n13125), .ZN(n13127) );
  NAND4_X1 U16535 ( .A1(n13130), .A2(n13129), .A3(n13128), .A4(n13127), .ZN(
        n13131) );
  NAND2_X1 U16536 ( .A1(n13132), .A2(n13131), .ZN(n13134) );
  OR3_X1 U16537 ( .A1(n14836), .A2(n12750), .A3(n14839), .ZN(n13133) );
  NOR2_X1 U16538 ( .A1(n13133), .A2(n13134), .ZN(n13135) );
  AOI21_X1 U16539 ( .B1(n13134), .B2(n13133), .A(n13135), .ZN(n14831) );
  NAND2_X1 U16540 ( .A1(n14832), .A2(n14831), .ZN(n14833) );
  INV_X1 U16541 ( .A(n13135), .ZN(n13136) );
  NAND2_X1 U16542 ( .A1(n14833), .A2(n13136), .ZN(n13159) );
  AOI22_X1 U16543 ( .A1(n10813), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U16544 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13138) );
  NAND2_X1 U16545 ( .A1(n13139), .A2(n13138), .ZN(n13157) );
  AOI22_X1 U16546 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13145) );
  NAND2_X1 U16547 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n13144) );
  NAND2_X1 U16548 ( .A1(n13141), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13143) );
  NAND4_X1 U16549 ( .A1(n13145), .A2(n13144), .A3(n13143), .A4(n13142), .ZN(
        n13156) );
  AOI22_X1 U16550 ( .A1(n10813), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13148) );
  AOI22_X1 U16551 ( .A1(n10812), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13147) );
  NAND2_X1 U16552 ( .A1(n13148), .A2(n13147), .ZN(n13155) );
  AOI22_X1 U16553 ( .A1(n13149), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13153) );
  NAND2_X1 U16554 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13151) );
  NAND2_X1 U16555 ( .A1(n13140), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n13150) );
  NAND4_X1 U16556 ( .A1(n13153), .A2(n13152), .A3(n13151), .A4(n13150), .ZN(
        n13154) );
  OAI22_X1 U16557 ( .A1(n13157), .A2(n13156), .B1(n13155), .B2(n13154), .ZN(
        n13158) );
  XNOR2_X1 U16558 ( .A(n13159), .B(n13158), .ZN(n13189) );
  INV_X1 U16559 ( .A(n13441), .ZN(n13636) );
  NAND2_X1 U16560 ( .A1(n13631), .A2(n13636), .ZN(n13161) );
  AND2_X1 U16561 ( .A1(n12776), .A2(n19747), .ZN(n13227) );
  NAND3_X1 U16562 ( .A1(n13632), .A2(n13633), .A3(n13227), .ZN(n13160) );
  NAND2_X1 U16563 ( .A1(n13161), .A2(n13160), .ZN(n13456) );
  AND2_X1 U16564 ( .A1(n13162), .A2(n12747), .ZN(n13163) );
  NAND2_X1 U16565 ( .A1(n13189), .A2(n16024), .ZN(n13184) );
  AOI22_X1 U16566 ( .A1(n18912), .A2(n14203), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n18921), .ZN(n13179) );
  AND2_X1 U16567 ( .A1(n13335), .A2(n13165), .ZN(n13180) );
  NOR4_X1 U16568 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13169) );
  NOR4_X1 U16569 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13168) );
  NOR4_X1 U16570 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13167) );
  NOR4_X1 U16571 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13166) );
  NAND4_X1 U16572 ( .A1(n13169), .A2(n13168), .A3(n13167), .A4(n13166), .ZN(
        n13174) );
  NOR4_X1 U16573 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13172) );
  NOR4_X1 U16574 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13171) );
  NOR4_X1 U16575 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13170) );
  INV_X1 U16576 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19638) );
  NAND4_X1 U16577 ( .A1(n13172), .A2(n13171), .A3(n13170), .A4(n19638), .ZN(
        n13173) );
  INV_X1 U16578 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n13175) );
  NOR2_X1 U16579 ( .A1(n19027), .A2(n13175), .ZN(n13176) );
  AOI21_X1 U16580 ( .B1(BUF1_REG_14__SCAN_IN), .B2(n19027), .A(n13176), .ZN(
        n18918) );
  AOI21_X1 U16581 ( .B1(n18908), .B2(BUF2_REG_30__SCAN_IN), .A(n13177), .ZN(
        n13178) );
  INV_X1 U16582 ( .A(n13180), .ZN(n13181) );
  INV_X1 U16583 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14397) );
  AND2_X1 U16584 ( .A1(n13182), .A2(n10083), .ZN(n13183) );
  NAND2_X1 U16585 ( .A1(n13184), .A2(n13183), .ZN(P2_U2889) );
  NAND2_X1 U16586 ( .A1(n13660), .A2(n13186), .ZN(n13438) );
  NAND2_X1 U16587 ( .A1(n13455), .A2(n13438), .ZN(n13187) );
  NAND2_X1 U16588 ( .A1(n13189), .A2(n18899), .ZN(n13193) );
  NAND2_X1 U16589 ( .A1(n18888), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13190) );
  NAND2_X1 U16590 ( .A1(n13193), .A2(n13192), .ZN(P2_U2857) );
  NOR2_X1 U16591 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13195) );
  NOR4_X1 U16592 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13194) );
  NAND4_X1 U16593 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13195), .A4(n13194), .ZN(n13208) );
  NOR4_X1 U16594 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13199) );
  NOR4_X1 U16595 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13198) );
  NOR4_X1 U16596 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13197) );
  NOR4_X1 U16597 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13196) );
  AND4_X1 U16598 ( .A1(n13199), .A2(n13198), .A3(n13197), .A4(n13196), .ZN(
        n13204) );
  NOR4_X1 U16599 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13202) );
  NOR4_X1 U16600 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13201) );
  NOR4_X1 U16601 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13200) );
  INV_X1 U16602 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20603) );
  AND4_X1 U16603 ( .A1(n13202), .A2(n13201), .A3(n13200), .A4(n20603), .ZN(
        n13203) );
  NAND2_X1 U16604 ( .A1(n13204), .A2(n13203), .ZN(n13205) );
  INV_X1 U16605 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20713) );
  NOR3_X1 U16606 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20713), .ZN(n13207) );
  NOR4_X1 U16607 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13206) );
  NAND4_X1 U16608 ( .A1(n20007), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n13207), .A4(
        n13206), .ZN(U214) );
  NOR2_X1 U16609 ( .A1(n19025), .A2(n13208), .ZN(n16211) );
  NAND2_X1 U16610 ( .A1(n16211), .A2(U214), .ZN(U212) );
  AOI211_X1 U16611 ( .C1(n15042), .C2(n13210), .A(n13209), .B(n18877), .ZN(
        n13221) );
  INV_X1 U16612 ( .A(n13211), .ZN(n13212) );
  OAI22_X1 U16613 ( .A1(n13212), .A2(n18852), .B1(n15039), .B2(n18832), .ZN(
        n13220) );
  INV_X1 U16614 ( .A(n18866), .ZN(n18837) );
  OAI22_X1 U16615 ( .A1(n18837), .A2(n11161), .B1(n11125), .B2(n18774), .ZN(
        n13219) );
  OAI21_X1 U16616 ( .B1(n13213), .B2(n14809), .A(n14859), .ZN(n15208) );
  OAI21_X1 U16617 ( .B1(n13217), .B2(n13216), .A(n13215), .ZN(n15204) );
  OAI22_X1 U16618 ( .A1(n15208), .A2(n18870), .B1(n15204), .B2(n18836), .ZN(
        n13218) );
  INV_X1 U16619 ( .A(n13222), .ZN(n13223) );
  NOR2_X1 U16620 ( .A1(n12766), .A2(n13223), .ZN(n18873) );
  INV_X1 U16621 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19760) );
  NAND2_X1 U16622 ( .A1(n19690), .A2(n14021), .ZN(n18641) );
  OAI211_X1 U16623 ( .C1(n18873), .C2(n19760), .A(n13233), .B(n18641), .ZN(
        P2_U2814) );
  INV_X1 U16624 ( .A(n12776), .ZN(n13226) );
  INV_X1 U16625 ( .A(n18643), .ZN(n19741) );
  INV_X1 U16626 ( .A(n18641), .ZN(n13224) );
  OAI21_X1 U16627 ( .B1(n13224), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19741), 
        .ZN(n13225) );
  OAI21_X1 U16628 ( .B1(n13226), .B2(n19741), .A(n13225), .ZN(P2_U3612) );
  INV_X1 U16629 ( .A(n13227), .ZN(n13228) );
  NAND4_X1 U16630 ( .A1(n13632), .A2(n13633), .A3(n13229), .A4(n13228), .ZN(
        n13640) );
  AND2_X1 U16631 ( .A1(n13640), .A2(n13460), .ZN(n19739) );
  OAI21_X1 U16632 ( .B1(n13642), .B2(n19739), .A(n13230), .ZN(P2_U2819) );
  INV_X1 U16633 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U16634 ( .A1(n13231), .A2(n19747), .ZN(n13232) );
  NOR2_X2 U16635 ( .A1(n13233), .A2(n13232), .ZN(n18972) );
  INV_X1 U16636 ( .A(n18972), .ZN(n13236) );
  AOI22_X1 U16637 ( .A1(n19027), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19025), .ZN(n13812) );
  INV_X1 U16638 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13235) );
  INV_X1 U16639 ( .A(n13233), .ZN(n13234) );
  OAI21_X1 U16640 ( .B1(n12750), .B2(n19747), .A(n13234), .ZN(n13245) );
  INV_X1 U16641 ( .A(n13245), .ZN(n13269) );
  OAI222_X1 U16642 ( .A1(n13237), .A2(n13317), .B1(n13236), .B2(n13812), .C1(
        n13235), .C2(n13269), .ZN(P2_U2982) );
  NOR2_X1 U16643 ( .A1(n12700), .A2(n19763), .ZN(n13238) );
  NAND2_X1 U16644 ( .A1(n14253), .A2(n14260), .ZN(n13298) );
  NOR2_X1 U16645 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20377), .ZN(n13297) );
  AOI21_X1 U16646 ( .B1(n13298), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13297), 
        .ZN(n13239) );
  NAND2_X1 U16647 ( .A1(n13695), .A2(n13239), .ZN(P1_U2801) );
  AOI22_X1 U16648 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13241) );
  AOI22_X1 U16649 ( .A1(n19027), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n13272), .ZN(n14923) );
  INV_X1 U16650 ( .A(n14923), .ZN(n13240) );
  NAND2_X1 U16651 ( .A1(n18972), .A2(n13240), .ZN(n13252) );
  NAND2_X1 U16652 ( .A1(n13241), .A2(n13252), .ZN(P2_U2961) );
  AOI22_X1 U16653 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16654 ( .A1(n19027), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13272), .ZN(n14939) );
  INV_X1 U16655 ( .A(n14939), .ZN(n19075) );
  NAND2_X1 U16656 ( .A1(n18972), .A2(n19075), .ZN(n13258) );
  NAND2_X1 U16657 ( .A1(n13242), .A2(n13258), .ZN(P2_U2959) );
  AOI22_X1 U16658 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U16659 ( .A1(n19027), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13272), .ZN(n14947) );
  INV_X1 U16660 ( .A(n14947), .ZN(n19067) );
  NAND2_X1 U16661 ( .A1(n18972), .A2(n19067), .ZN(n13256) );
  NAND2_X1 U16662 ( .A1(n13243), .A2(n13256), .ZN(P2_U2958) );
  AOI22_X1 U16663 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16664 ( .A1(n19027), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19025), .ZN(n14973) );
  INV_X1 U16665 ( .A(n14973), .ZN(n19041) );
  NAND2_X1 U16666 ( .A1(n18972), .A2(n19041), .ZN(n13285) );
  NAND2_X1 U16667 ( .A1(n13244), .A2(n13285), .ZN(P2_U2953) );
  AOI22_X1 U16668 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16669 ( .A1(n19027), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13272), .ZN(n14929) );
  INV_X1 U16670 ( .A(n14929), .ZN(n13246) );
  NAND2_X1 U16671 ( .A1(n18972), .A2(n13246), .ZN(n13267) );
  NAND2_X1 U16672 ( .A1(n13247), .A2(n13267), .ZN(P2_U2960) );
  INV_X1 U16673 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16246) );
  NOR2_X1 U16674 ( .A1(n19025), .A2(n16246), .ZN(n13248) );
  AOI21_X1 U16675 ( .B1(n19025), .B2(BUF2_REG_10__SCAN_IN), .A(n13248), .ZN(
        n14913) );
  INV_X1 U16676 ( .A(n14913), .ZN(n18922) );
  NAND2_X1 U16677 ( .A1(n18972), .A2(n18922), .ZN(n13271) );
  NAND2_X1 U16678 ( .A1(n18970), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13249) );
  OAI211_X1 U16679 ( .C1(n13317), .C2(n11133), .A(n13271), .B(n13249), .ZN(
        P2_U2962) );
  AOI22_X1 U16680 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U16681 ( .A1(n19027), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19025), .ZN(n14961) );
  INV_X1 U16682 ( .A(n14961), .ZN(n19051) );
  NAND2_X1 U16683 ( .A1(n18972), .A2(n19051), .ZN(n13295) );
  NAND2_X1 U16684 ( .A1(n13250), .A2(n13295), .ZN(P2_U2955) );
  AOI22_X1 U16685 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13251) );
  INV_X1 U16686 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16254) );
  INV_X1 U16687 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n17982) );
  AOI22_X1 U16688 ( .A1(n19027), .A2(n16254), .B1(n17982), .B2(n19025), .ZN(
        n19057) );
  NAND2_X1 U16689 ( .A1(n18972), .A2(n19057), .ZN(n13274) );
  NAND2_X1 U16690 ( .A1(n13251), .A2(n13274), .ZN(P2_U2971) );
  AOI22_X1 U16691 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U16692 ( .A1(n13253), .A2(n13252), .ZN(P2_U2976) );
  AOI22_X1 U16693 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U16694 ( .A1(n19027), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13272), .ZN(n18927) );
  INV_X1 U16695 ( .A(n18927), .ZN(n19063) );
  NAND2_X1 U16696 ( .A1(n18972), .A2(n19063), .ZN(n13283) );
  NAND2_X1 U16697 ( .A1(n13254), .A2(n13283), .ZN(P2_U2972) );
  AOI22_X1 U16698 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13255) );
  INV_X1 U16699 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16258) );
  INV_X1 U16700 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n17974) );
  AOI22_X1 U16701 ( .A1(n19027), .A2(n16258), .B1(n17974), .B2(n13272), .ZN(
        n19047) );
  NAND2_X1 U16702 ( .A1(n18972), .A2(n19047), .ZN(n13291) );
  NAND2_X1 U16703 ( .A1(n13255), .A2(n13291), .ZN(P2_U2954) );
  AOI22_X1 U16704 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13257) );
  NAND2_X1 U16705 ( .A1(n13257), .A2(n13256), .ZN(P2_U2973) );
  AOI22_X1 U16706 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13259) );
  NAND2_X1 U16707 ( .A1(n13259), .A2(n13258), .ZN(P2_U2974) );
  AOI22_X1 U16708 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n13261) );
  AOI22_X1 U16709 ( .A1(n19027), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13272), .ZN(n14891) );
  INV_X1 U16710 ( .A(n14891), .ZN(n13260) );
  NAND2_X1 U16711 ( .A1(n18972), .A2(n13260), .ZN(n13289) );
  NAND2_X1 U16712 ( .A1(n13261), .A2(n13289), .ZN(P2_U2979) );
  AOI22_X1 U16713 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13266) );
  INV_X1 U16714 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13262) );
  OR2_X1 U16715 ( .A1(n19025), .A2(n13262), .ZN(n13264) );
  NAND2_X1 U16716 ( .A1(n19025), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13263) );
  AND2_X1 U16717 ( .A1(n13264), .A2(n13263), .ZN(n14901) );
  INV_X1 U16718 ( .A(n14901), .ZN(n13265) );
  NAND2_X1 U16719 ( .A1(n18972), .A2(n13265), .ZN(n13287) );
  NAND2_X1 U16720 ( .A1(n13266), .A2(n13287), .ZN(P2_U2978) );
  AOI22_X1 U16721 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13268) );
  NAND2_X1 U16722 ( .A1(n13268), .A2(n13267), .ZN(P2_U2975) );
  NAND2_X1 U16723 ( .A1(n18970), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13270) );
  OAI211_X1 U16724 ( .C1(n13317), .C2(n11031), .A(n13271), .B(n13270), .ZN(
        P2_U2977) );
  AOI22_X1 U16725 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13273) );
  INV_X1 U16726 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16264) );
  INV_X1 U16727 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n17964) );
  AOI22_X1 U16728 ( .A1(n19027), .A2(n16264), .B1(n17964), .B2(n13272), .ZN(
        n19030) );
  NAND2_X1 U16729 ( .A1(n18972), .A2(n19030), .ZN(n13293) );
  NAND2_X1 U16730 ( .A1(n13273), .A2(n13293), .ZN(P2_U2967) );
  AOI22_X1 U16731 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13275) );
  NAND2_X1 U16732 ( .A1(n13275), .A2(n13274), .ZN(P2_U2956) );
  AOI22_X1 U16733 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13280) );
  INV_X1 U16734 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13276) );
  OR2_X1 U16735 ( .A1(n19025), .A2(n13276), .ZN(n13278) );
  NAND2_X1 U16736 ( .A1(n19025), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13277) );
  AND2_X1 U16737 ( .A1(n13278), .A2(n13277), .ZN(n14884) );
  INV_X1 U16738 ( .A(n14884), .ZN(n13279) );
  NAND2_X1 U16739 ( .A1(n18972), .A2(n13279), .ZN(n13281) );
  NAND2_X1 U16740 ( .A1(n13280), .A2(n13281), .ZN(P2_U2980) );
  AOI22_X1 U16741 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13282) );
  NAND2_X1 U16742 ( .A1(n13282), .A2(n13281), .ZN(P2_U2965) );
  AOI22_X1 U16743 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n13245), .B1(n18974), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13284) );
  NAND2_X1 U16744 ( .A1(n13284), .A2(n13283), .ZN(P2_U2957) );
  AOI22_X1 U16745 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13286) );
  NAND2_X1 U16746 ( .A1(n13286), .A2(n13285), .ZN(P2_U2968) );
  AOI22_X1 U16747 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n13288) );
  NAND2_X1 U16748 ( .A1(n13288), .A2(n13287), .ZN(P2_U2963) );
  AOI22_X1 U16749 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n13290) );
  NAND2_X1 U16750 ( .A1(n13290), .A2(n13289), .ZN(P2_U2964) );
  AOI22_X1 U16751 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13292) );
  NAND2_X1 U16752 ( .A1(n13292), .A2(n13291), .ZN(P2_U2969) );
  AOI22_X1 U16753 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13294) );
  NAND2_X1 U16754 ( .A1(n13294), .A2(n13293), .ZN(P2_U2952) );
  AOI22_X1 U16755 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13296) );
  NAND2_X1 U16756 ( .A1(n13296), .A2(n13295), .ZN(P2_U2970) );
  NOR2_X1 U16757 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(n13297), .ZN(n13300)
         );
  OAI21_X1 U16758 ( .B1(n14251), .B2(n14276), .A(n20706), .ZN(n13299) );
  OAI21_X1 U16759 ( .B1(n13300), .B2(n20706), .A(n13299), .ZN(P1_U3487) );
  OAI21_X1 U16760 ( .B1(n18864), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13308), .ZN(n13301) );
  INV_X1 U16761 ( .A(n13301), .ZN(n13365) );
  OAI21_X1 U16762 ( .B1(n13303), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13302), .ZN(n13364) );
  NAND2_X1 U16763 ( .A1(n18822), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13366) );
  OAI21_X1 U16764 ( .B1(n18980), .B2(n13364), .A(n13366), .ZN(n13304) );
  AOI21_X1 U16765 ( .B1(n16112), .B2(n13365), .A(n13304), .ZN(n13307) );
  OAI21_X1 U16766 ( .B1(n18977), .B2(n13305), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13306) );
  OAI211_X1 U16767 ( .C1(n19026), .C2(n18871), .A(n13307), .B(n13306), .ZN(
        P2_U3014) );
  XNOR2_X1 U16768 ( .A(n13308), .B(n15446), .ZN(n13309) );
  XNOR2_X1 U16769 ( .A(n18851), .B(n13309), .ZN(n15447) );
  INV_X1 U16770 ( .A(n15447), .ZN(n13315) );
  MUX2_X1 U16771 ( .A(n16108), .B(n18977), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13314) );
  OAI21_X1 U16772 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13311), .A(
        n13310), .ZN(n15450) );
  NOR2_X1 U16773 ( .A1(n18772), .A2(n19636), .ZN(n15449) );
  INV_X1 U16774 ( .A(n15449), .ZN(n13312) );
  OAI21_X1 U16775 ( .B1(n18980), .B2(n15450), .A(n13312), .ZN(n13313) );
  AOI211_X1 U16776 ( .C1(n13315), .C2(n16112), .A(n13314), .B(n13313), .ZN(
        n13316) );
  OAI21_X1 U16777 ( .B1(n18853), .B2(n19026), .A(n13316), .ZN(P2_U3013) );
  OR2_X1 U16778 ( .A1(n12766), .A2(n16167), .ZN(n13318) );
  NOR2_X1 U16779 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19721), .ZN(n13379) );
  INV_X1 U16780 ( .A(n13379), .ZN(n13322) );
  INV_X1 U16781 ( .A(n13322), .ZN(n20716) );
  AOI22_X1 U16782 ( .A1(n20716), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13323) );
  OAI21_X1 U16783 ( .B1(n11112), .B2(n20720), .A(n13323), .ZN(P2_U2935) );
  AOI22_X1 U16784 ( .A1(n20716), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13324) );
  OAI21_X1 U16785 ( .B1(n14902), .B2(n20720), .A(n13324), .ZN(P2_U2924) );
  AOI22_X1 U16786 ( .A1(n20716), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13325) );
  OAI21_X1 U16787 ( .B1(n14885), .B2(n20720), .A(n13325), .ZN(P2_U2922) );
  AOI22_X1 U16788 ( .A1(n13379), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13326) );
  OAI21_X1 U16789 ( .B1(n20852), .B2(n20720), .A(n13326), .ZN(P2_U2930) );
  INV_X1 U16790 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14946) );
  AOI22_X1 U16791 ( .A1(n13379), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13327) );
  OAI21_X1 U16792 ( .B1(n14946), .B2(n20720), .A(n13327), .ZN(P2_U2929) );
  AOI22_X1 U16793 ( .A1(n13379), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13328) );
  OAI21_X1 U16794 ( .B1(n11126), .B2(n20720), .A(n13328), .ZN(P2_U2928) );
  AOI22_X1 U16795 ( .A1(n13379), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13329) );
  OAI21_X1 U16796 ( .B1(n14972), .B2(n20720), .A(n13329), .ZN(P2_U2934) );
  AOI22_X1 U16797 ( .A1(n13379), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13330) );
  OAI21_X1 U16798 ( .B1(n14922), .B2(n20720), .A(n13330), .ZN(P2_U2926) );
  AOI22_X1 U16799 ( .A1(n13379), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13331) );
  OAI21_X1 U16800 ( .B1(n20796), .B2(n20720), .A(n13331), .ZN(P2_U2923) );
  AOI22_X1 U16801 ( .A1(n13379), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13332) );
  OAI21_X1 U16802 ( .B1(n11128), .B2(n20720), .A(n13332), .ZN(P2_U2927) );
  AOI22_X1 U16803 ( .A1(n13379), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13333) );
  OAI21_X1 U16804 ( .B1(n11133), .B2(n20720), .A(n13333), .ZN(P2_U2925) );
  INV_X1 U16805 ( .A(n19030), .ZN(n13348) );
  NOR2_X1 U16806 ( .A1(n13337), .A2(n13336), .ZN(n13338) );
  NOR2_X1 U16807 ( .A1(n13339), .A2(n13338), .ZN(n18862) );
  AOI22_X1 U16808 ( .A1(n18912), .A2(n18862), .B1(n18921), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13347) );
  INV_X1 U16809 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19039) );
  AND2_X1 U16810 ( .A1(n19700), .A2(n19039), .ZN(n13341) );
  OAI21_X1 U16811 ( .B1(n13342), .B2(n13341), .A(n13340), .ZN(n13343) );
  INV_X1 U16812 ( .A(n13343), .ZN(n13344) );
  NAND2_X1 U16813 ( .A1(n19287), .A2(n18862), .ZN(n13432) );
  OAI211_X1 U16814 ( .C1(n19287), .C2(n18862), .A(n16024), .B(n13432), .ZN(
        n13346) );
  OAI211_X1 U16815 ( .C1(n13348), .C2(n18928), .A(n13347), .B(n13346), .ZN(
        P2_U2919) );
  OAI21_X1 U16816 ( .B1(n13349), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11412), .ZN(n19997) );
  INV_X1 U16817 ( .A(n13350), .ZN(n13351) );
  AOI21_X1 U16818 ( .B1(n13353), .B2(n13352), .A(n13351), .ZN(n13520) );
  NAND2_X1 U16819 ( .A1(n13520), .A2(n19934), .ZN(n13358) );
  NAND2_X1 U16820 ( .A1(n13354), .A2(n15823), .ZN(n13356) );
  NAND2_X1 U16821 ( .A1(n19977), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20002) );
  INV_X1 U16822 ( .A(n20002), .ZN(n13355) );
  AOI21_X1 U16823 ( .B1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13356), .A(
        n13355), .ZN(n13357) );
  OAI211_X1 U16824 ( .C1(n19943), .C2(n19997), .A(n13358), .B(n13357), .ZN(
        P1_U2999) );
  XNOR2_X1 U16825 ( .A(n13360), .B(n13359), .ZN(n18818) );
  OAI222_X1 U16826 ( .A1(n18928), .A2(n14947), .B1(n18818), .B2(n18936), .C1(
        n18958), .C2(n18926), .ZN(P2_U2913) );
  XNOR2_X1 U16827 ( .A(n13362), .B(n13361), .ZN(n16138) );
  OAI222_X1 U16828 ( .A1(n18928), .A2(n14939), .B1(n16138), .B2(n18936), .C1(
        n18956), .C2(n18926), .ZN(P2_U2912) );
  INV_X1 U16829 ( .A(n13363), .ZN(n19004) );
  OAI22_X1 U16830 ( .A1(n19004), .A2(n13370), .B1(n18996), .B2(n13364), .ZN(
        n13369) );
  AOI22_X1 U16831 ( .A1(n18993), .A2(n18862), .B1(n18992), .B2(n13365), .ZN(
        n13367) );
  OAI211_X1 U16832 ( .C1(n16137), .C2(n18871), .A(n13367), .B(n13366), .ZN(
        n13368) );
  AOI211_X1 U16833 ( .C1(n13370), .C2(n15452), .A(n13369), .B(n13368), .ZN(
        n13371) );
  INV_X1 U16834 ( .A(n13371), .ZN(P2_U3046) );
  MUX2_X1 U16835 ( .A(n13372), .B(n18871), .S(n18903), .Z(n13373) );
  OAI21_X1 U16836 ( .B1(n18893), .B2(n19724), .A(n13373), .ZN(P2_U2887) );
  MUX2_X1 U16837 ( .A(n13376), .B(n18853), .S(n18903), .Z(n13377) );
  OAI21_X1 U16838 ( .B1(n19712), .B2(n18893), .A(n13377), .ZN(P2_U2886) );
  AOI22_X1 U16839 ( .A1(n13379), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13378) );
  OAI21_X1 U16840 ( .B1(n10808), .B2(n20720), .A(n13378), .ZN(P2_U2933) );
  AOI22_X1 U16841 ( .A1(n13379), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13380) );
  OAI21_X1 U16842 ( .B1(n14960), .B2(n20720), .A(n13380), .ZN(P2_U2932) );
  NOR2_X1 U16843 ( .A1(n13950), .A2(n18888), .ZN(n13384) );
  AOI21_X1 U16844 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n18888), .A(n13384), .ZN(
        n13385) );
  OAI21_X1 U16845 ( .B1(n19320), .B2(n18893), .A(n13385), .ZN(P2_U2884) );
  NAND2_X1 U16846 ( .A1(n13387), .A2(n13386), .ZN(n13390) );
  INV_X1 U16847 ( .A(n13388), .ZN(n13389) );
  NAND2_X1 U16848 ( .A1(n13390), .A2(n13389), .ZN(n18802) );
  OAI222_X1 U16849 ( .A1(n18928), .A2(n14929), .B1(n18802), .B2(n18936), .C1(
        n10999), .C2(n18926), .ZN(P2_U2911) );
  INV_X1 U16850 ( .A(n19177), .ZN(n19705) );
  MUX2_X1 U16851 ( .A(n13394), .B(n14238), .S(n18903), .Z(n13395) );
  OAI21_X1 U16852 ( .B1(n19705), .B2(n18893), .A(n13395), .ZN(P2_U2885) );
  INV_X1 U16853 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13713) );
  NAND3_X1 U16854 ( .A1(n14252), .A2(n14260), .A3(n13506), .ZN(n13396) );
  OAI21_X1 U16855 ( .B1(n13695), .B2(n20025), .A(n13396), .ZN(n13398) );
  NOR2_X1 U16856 ( .A1(n20700), .A2(n13792), .ZN(n15952) );
  INV_X1 U16857 ( .A(n15952), .ZN(n13578) );
  AOI22_X1 U16858 ( .A1(n20709), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13400) );
  OAI21_X1 U16859 ( .B1(n13713), .B2(n13692), .A(n13400), .ZN(P1_U2909) );
  INV_X1 U16860 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13726) );
  AOI22_X1 U16861 ( .A1(n20709), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13401) );
  OAI21_X1 U16862 ( .B1(n13726), .B2(n13692), .A(n13401), .ZN(P1_U2912) );
  INV_X1 U16863 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U16864 ( .A1(n20709), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13402) );
  OAI21_X1 U16865 ( .B1(n13717), .B2(n13692), .A(n13402), .ZN(P1_U2906) );
  AOI22_X1 U16866 ( .A1(n20709), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13403) );
  OAI21_X1 U16867 ( .B1(n12111), .B2(n13692), .A(n13403), .ZN(P1_U2908) );
  INV_X1 U16868 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13706) );
  AOI22_X1 U16869 ( .A1(n20709), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13404) );
  OAI21_X1 U16870 ( .B1(n13706), .B2(n13692), .A(n13404), .ZN(P1_U2907) );
  INV_X1 U16871 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U16872 ( .A1(n20709), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13405) );
  OAI21_X1 U16873 ( .B1(n13702), .B2(n13692), .A(n13405), .ZN(P1_U2911) );
  AOI22_X1 U16874 ( .A1(n20709), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13406) );
  OAI21_X1 U16875 ( .B1(n12067), .B2(n13692), .A(n13406), .ZN(P1_U2910) );
  XNOR2_X1 U16876 ( .A(n13407), .B(n12601), .ZN(n19976) );
  OR2_X1 U16877 ( .A1(n14252), .A2(n14243), .ZN(n13493) );
  INV_X1 U16878 ( .A(n13408), .ZN(n13410) );
  NAND4_X1 U16879 ( .A1(n13410), .A2(n13409), .A3(n14166), .A4(n13557), .ZN(
        n13422) );
  NAND2_X1 U16880 ( .A1(n13493), .A2(n13411), .ZN(n13412) );
  OAI21_X1 U16881 ( .B1(n13415), .B2(n13414), .A(n13413), .ZN(n19947) );
  OAI222_X1 U16882 ( .A1(n19976), .A2(n14383), .B1(n9786), .B2(n19854), .C1(
        n19947), .C2(n14394), .ZN(P1_U2871) );
  INV_X1 U16883 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18953) );
  OAI21_X1 U16884 ( .B1(n13388), .B2(n13416), .A(n15391), .ZN(n18789) );
  OAI222_X1 U16885 ( .A1(n18928), .A2(n14923), .B1(n18926), .B2(n18953), .C1(
        n18936), .C2(n18789), .ZN(P2_U2910) );
  OR2_X1 U16886 ( .A1(n13417), .A2(n13421), .ZN(n13477) );
  OAI21_X1 U16887 ( .B1(n15619), .B2(n12591), .A(n13477), .ZN(n13418) );
  NAND2_X1 U16888 ( .A1(n14252), .A2(n13418), .ZN(n13420) );
  INV_X1 U16889 ( .A(n12592), .ZN(n15944) );
  NAND3_X1 U16890 ( .A1(n15944), .A2(n14245), .A3(n20708), .ZN(n13419) );
  NAND2_X1 U16891 ( .A1(n13420), .A2(n13419), .ZN(n13487) );
  NOR2_X1 U16892 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  OR3_X2 U16893 ( .A1(n15801), .A2(n13489), .A3(n13425), .ZN(n14435) );
  INV_X1 U16894 ( .A(n20007), .ZN(n20005) );
  NAND2_X1 U16895 ( .A1(n20005), .A2(DATAI_1_), .ZN(n13427) );
  NAND2_X1 U16896 ( .A1(n20007), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13426) );
  AND2_X1 U16897 ( .A1(n13427), .A2(n13426), .ZN(n20026) );
  INV_X1 U16898 ( .A(n13489), .ZN(n13468) );
  INV_X1 U16899 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19882) );
  OAI222_X1 U16900 ( .A1(n14435), .A2(n19947), .B1(n20026), .B2(n14118), .C1(
        n14437), .C2(n19882), .ZN(P1_U2903) );
  OAI21_X1 U16901 ( .B1(n13431), .B2(n13430), .A(n13429), .ZN(n19717) );
  NOR2_X1 U16902 ( .A1(n19715), .A2(n19717), .ZN(n13606) );
  AOI21_X1 U16903 ( .B1(n19715), .B2(n19717), .A(n13606), .ZN(n13433) );
  NAND2_X1 U16904 ( .A1(n13433), .A2(n13432), .ZN(n13608) );
  OAI21_X1 U16905 ( .B1(n13433), .B2(n13432), .A(n13608), .ZN(n13434) );
  NAND2_X1 U16906 ( .A1(n13434), .A2(n16024), .ZN(n13436) );
  AOI22_X1 U16907 ( .A1(n18912), .A2(n19717), .B1(n18921), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13435) );
  OAI211_X1 U16908 ( .C1(n14973), .C2(n18928), .A(n13436), .B(n13435), .ZN(
        P2_U2918) );
  INV_X1 U16909 ( .A(n19320), .ZN(n19697) );
  AND2_X1 U16910 ( .A1(n13631), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16163) );
  OR2_X1 U16911 ( .A1(n13950), .A2(n13660), .ZN(n13453) );
  NAND2_X1 U16912 ( .A1(n13438), .A2(n13437), .ZN(n13627) );
  INV_X1 U16913 ( .A(n13439), .ZN(n13440) );
  OAI21_X1 U16914 ( .B1(n13615), .B2(n10547), .A(n13440), .ZN(n13451) );
  NAND2_X1 U16915 ( .A1(n13634), .A2(n13441), .ZN(n13618) );
  INV_X1 U16916 ( .A(n10827), .ZN(n13442) );
  NAND2_X1 U16917 ( .A1(n13442), .A2(n10785), .ZN(n13616) );
  AOI22_X1 U16918 ( .A1(n13616), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13443), .B2(n13442), .ZN(n13444) );
  NAND2_X1 U16919 ( .A1(n13618), .A2(n13444), .ZN(n13449) );
  AOI21_X1 U16920 ( .B1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13445) );
  NOR2_X1 U16921 ( .A1(n13446), .A2(n13445), .ZN(n13447) );
  NAND2_X1 U16922 ( .A1(n13656), .A2(n13447), .ZN(n13448) );
  NAND2_X1 U16923 ( .A1(n13449), .A2(n13448), .ZN(n13450) );
  AOI21_X1 U16924 ( .B1(n13627), .B2(n13451), .A(n13450), .ZN(n13452) );
  NAND2_X1 U16925 ( .A1(n13453), .A2(n13452), .ZN(n13630) );
  AOI22_X1 U16926 ( .A1(n19697), .A2(n16163), .B1(n19693), .B2(n13630), .ZN(
        n13466) );
  NAND2_X1 U16927 ( .A1(n13455), .A2(n13454), .ZN(n13457) );
  NOR2_X1 U16928 ( .A1(n13457), .A2(n13456), .ZN(n13458) );
  OAI21_X1 U16929 ( .B1(n13459), .B2(n12766), .A(n13458), .ZN(n13654) );
  NAND2_X1 U16930 ( .A1(n13654), .A2(n13460), .ZN(n13464) );
  NOR2_X1 U16931 ( .A1(n19751), .A2(n19721), .ZN(n16158) );
  NAND2_X1 U16932 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(n16158), .ZN(n13462) );
  AND2_X1 U16933 ( .A1(n13462), .A2(n13461), .ZN(n13463) );
  NAND2_X1 U16934 ( .A1(n13464), .A2(n13463), .ZN(n15562) );
  NAND2_X1 U16935 ( .A1(n15559), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13465) );
  OAI21_X1 U16936 ( .B1(n13466), .B2(n15559), .A(n13465), .ZN(P2_U3596) );
  NAND2_X1 U16937 ( .A1(n13468), .A2(n13467), .ZN(n13469) );
  NOR2_X1 U16938 ( .A1(n13470), .A2(n13469), .ZN(n13471) );
  NAND2_X1 U16939 ( .A1(n13471), .A2(n12592), .ZN(n14745) );
  NAND2_X1 U16940 ( .A1(n20666), .A2(n14745), .ZN(n13485) );
  AND2_X1 U16941 ( .A1(n13506), .A2(n11186), .ZN(n14744) );
  INV_X1 U16942 ( .A(n13476), .ZN(n13473) );
  NAND2_X1 U16943 ( .A1(n13479), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13472) );
  NAND2_X1 U16944 ( .A1(n13473), .A2(n13472), .ZN(n13474) );
  AOI22_X1 U16945 ( .A1(n14744), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13506), .B2(n13474), .ZN(n13484) );
  MUX2_X1 U16946 ( .A(n13476), .B(n11184), .S(n13475), .Z(n13478) );
  NAND2_X1 U16947 ( .A1(n14243), .A2(n13477), .ZN(n13561) );
  OAI21_X1 U16948 ( .B1(n13479), .B2(n13478), .A(n13561), .ZN(n13483) );
  INV_X1 U16949 ( .A(n14745), .ZN(n13563) );
  AOI21_X1 U16950 ( .B1(n13475), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13480) );
  NOR2_X1 U16951 ( .A1(n13481), .A2(n13480), .ZN(n13486) );
  NAND3_X1 U16952 ( .A1(n13563), .A2(n13557), .A3(n13486), .ZN(n13482) );
  NAND4_X1 U16953 ( .A1(n13485), .A2(n13484), .A3(n13483), .A4(n13482), .ZN(
        n13564) );
  AOI22_X1 U16954 ( .A1(n13564), .A2(n15945), .B1(n13486), .B2(n14753), .ZN(
        n13498) );
  INV_X1 U16955 ( .A(n13487), .ZN(n13496) );
  NOR2_X1 U16956 ( .A1(n15620), .A2(n15619), .ZN(n13488) );
  AND2_X1 U16957 ( .A1(n14252), .A2(n13488), .ZN(n15600) );
  OAI21_X1 U16958 ( .B1(n13489), .B2(n13506), .A(n15600), .ZN(n13495) );
  OR2_X1 U16959 ( .A1(n14257), .A2(n20029), .ZN(n13490) );
  AND2_X1 U16960 ( .A1(n13491), .A2(n13490), .ZN(n13492) );
  AND2_X1 U16961 ( .A1(n13493), .A2(n13492), .ZN(n13494) );
  NAND3_X1 U16962 ( .A1(n13496), .A2(n13495), .A3(n13494), .ZN(n13566) );
  INV_X1 U16963 ( .A(n13566), .ZN(n15579) );
  NAND2_X1 U16964 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15952), .ZN(n15957) );
  INV_X1 U16965 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19770) );
  OAI22_X1 U16966 ( .A1(n15579), .A2(n19763), .B1(n15957), .B2(n19770), .ZN(
        n15943) );
  AOI21_X1 U16967 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20702), .A(n15943), 
        .ZN(n14749) );
  NAND2_X1 U16968 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14749), .ZN(
        n13497) );
  OAI21_X1 U16969 ( .B1(n13498), .B2(n14749), .A(n13497), .ZN(P1_U3469) );
  OAI21_X1 U16970 ( .B1(n13500), .B2(n13499), .A(n13744), .ZN(n19965) );
  INV_X1 U16971 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13504) );
  NAND2_X1 U16972 ( .A1(n13501), .A2(n13413), .ZN(n13502) );
  AND2_X1 U16973 ( .A1(n13503), .A2(n13502), .ZN(n19844) );
  INV_X1 U16974 ( .A(n19844), .ZN(n13720) );
  OAI222_X1 U16975 ( .A1(n19965), .A2(n14383), .B1(n13504), .B2(n19854), .C1(
        n13720), .C2(n14394), .ZN(P1_U2870) );
  INV_X1 U16976 ( .A(n11684), .ZN(n20121) );
  OAI22_X1 U16977 ( .A1(n20121), .A2(n13563), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14742), .ZN(n15578) );
  OAI22_X1 U16978 ( .A1(n13792), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15599), .ZN(n13505) );
  AOI21_X1 U16979 ( .B1(n15578), .B2(n15945), .A(n13505), .ZN(n13508) );
  INV_X1 U16980 ( .A(n13506), .ZN(n13555) );
  NOR2_X1 U16981 ( .A1(n13555), .A2(n11183), .ZN(n15577) );
  AOI22_X1 U16982 ( .A1(n15577), .A2(n15945), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14749), .ZN(n13507) );
  OAI21_X1 U16983 ( .B1(n13508), .B2(n14749), .A(n13507), .ZN(P1_U3474) );
  NOR2_X1 U16984 ( .A1(n13510), .A2(n13509), .ZN(n19969) );
  INV_X1 U16985 ( .A(n19969), .ZN(n13512) );
  NAND3_X1 U16986 ( .A1(n13512), .A2(n19935), .A3(n13511), .ZN(n13518) );
  INV_X1 U16987 ( .A(n13513), .ZN(n19836) );
  INV_X1 U16988 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13515) );
  INV_X1 U16989 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13514) );
  OAI22_X1 U16990 ( .A1(n15823), .A2(n13515), .B1(n19964), .B2(n13514), .ZN(
        n13516) );
  AOI21_X1 U16991 ( .B1(n19836), .B2(n15849), .A(n13516), .ZN(n13517) );
  OAI211_X1 U16992 ( .C1(n20006), .C2(n13720), .A(n13518), .B(n13517), .ZN(
        P1_U2997) );
  OR2_X1 U16993 ( .A1(n9718), .A2(n13519), .ZN(n19994) );
  INV_X1 U16994 ( .A(n13520), .ZN(n13809) );
  OAI222_X1 U16995 ( .A1(n19994), .A2(n14383), .B1(n13802), .B2(n19854), .C1(
        n13809), .C2(n14394), .ZN(P1_U2872) );
  XOR2_X1 U16996 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n9625), .Z(n13526)
         );
  NAND2_X1 U16997 ( .A1(n18888), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n13525) );
  AOI21_X1 U16998 ( .B1(n9717), .B2(n9846), .A(n13523), .ZN(n18826) );
  NAND2_X1 U16999 ( .A1(n18903), .A2(n18826), .ZN(n13524) );
  OAI211_X1 U17000 ( .C1(n13526), .C2(n18893), .A(n13525), .B(n13524), .ZN(
        P2_U2882) );
  INV_X1 U17001 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13527) );
  NOR2_X1 U17002 ( .A1(n9625), .A2(n13527), .ZN(n13529) );
  OR2_X1 U17003 ( .A1(n9625), .A2(n13528), .ZN(n13595) );
  OAI211_X1 U17004 ( .C1(n13529), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n18899), .B(n13595), .ZN(n13533) );
  OAI21_X1 U17005 ( .B1(n13523), .B2(n13531), .A(n9852), .ZN(n15124) );
  INV_X1 U17006 ( .A(n15124), .ZN(n18814) );
  NAND2_X1 U17007 ( .A1(n18903), .A2(n18814), .ZN(n13532) );
  OAI211_X1 U17008 ( .C1(n18903), .C2(n13534), .A(n13533), .B(n13532), .ZN(
        P2_U2881) );
  INV_X1 U17009 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18950) );
  OAI21_X1 U17010 ( .B1(n13537), .B2(n13536), .A(n13535), .ZN(n18770) );
  OAI222_X1 U17011 ( .A1(n18928), .A2(n14901), .B1(n18926), .B2(n18950), .C1(
        n18936), .C2(n18770), .ZN(P2_U2908) );
  NOR2_X1 U17012 ( .A1(n9625), .A2(n13538), .ZN(n18892) );
  XNOR2_X1 U17013 ( .A(n18892), .B(n18891), .ZN(n13543) );
  OR2_X1 U17014 ( .A1(n13547), .A2(n13539), .ZN(n13541) );
  NAND2_X1 U17015 ( .A1(n13541), .A2(n13540), .ZN(n18788) );
  MUX2_X1 U17016 ( .A(n12324), .B(n18788), .S(n18903), .Z(n13542) );
  OAI21_X1 U17017 ( .B1(n13543), .B2(n18893), .A(n13542), .ZN(P2_U2878) );
  NOR2_X1 U17018 ( .A1(n13544), .A2(n13545), .ZN(n13546) );
  OR2_X1 U17019 ( .A1(n13547), .A2(n13546), .ZN(n18803) );
  NOR2_X1 U17020 ( .A1(n9625), .A2(n13548), .ZN(n13551) );
  INV_X1 U17021 ( .A(n18892), .ZN(n13549) );
  OAI211_X1 U17022 ( .C1(n13551), .C2(n13550), .A(n13549), .B(n18899), .ZN(
        n13553) );
  NAND2_X1 U17023 ( .A1(n18888), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13552) );
  OAI211_X1 U17024 ( .C1(n18803), .C2(n18888), .A(n13553), .B(n13552), .ZN(
        P2_U2879) );
  NOR2_X1 U17025 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13792), .ZN(n13569) );
  XNOR2_X1 U17026 ( .A(n13475), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14752) );
  NOR2_X1 U17027 ( .A1(n13555), .A2(n11186), .ZN(n13556) );
  MUX2_X1 U17028 ( .A(n14744), .B(n13556), .S(n11185), .Z(n13560) );
  INV_X1 U17029 ( .A(n13557), .ZN(n13558) );
  NOR3_X1 U17030 ( .A1(n14745), .A2(n13558), .A3(n14752), .ZN(n13559) );
  AOI211_X1 U17031 ( .C1(n13561), .C2(n14752), .A(n13560), .B(n13559), .ZN(
        n13562) );
  OAI21_X1 U17032 ( .B1(n20678), .B2(n13563), .A(n13562), .ZN(n14751) );
  MUX2_X1 U17033 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14751), .S(
        n13566), .Z(n15584) );
  AOI22_X1 U17034 ( .A1(n13569), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15584), .B2(n13792), .ZN(n13573) );
  MUX2_X1 U17035 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13564), .S(
        n13566), .Z(n15587) );
  AOI22_X1 U17036 ( .A1(n13569), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13792), .B2(n15587), .ZN(n13572) );
  INV_X1 U17037 ( .A(n20159), .ZN(n20407) );
  OR2_X1 U17038 ( .A1(n11468), .A2(n20407), .ZN(n13565) );
  XNOR2_X1 U17039 ( .A(n13565), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19821) );
  AOI21_X1 U17040 ( .B1(n19821), .B2(n15944), .A(n15579), .ZN(n13568) );
  OAI21_X1 U17041 ( .B1(n13566), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13792), .ZN(n13567) );
  OR2_X1 U17042 ( .A1(n13568), .A2(n13567), .ZN(n13571) );
  NAND2_X1 U17043 ( .A1(n13569), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13570) );
  OAI21_X1 U17044 ( .B1(n13573), .B2(n13572), .A(n13574), .ZN(n15596) );
  NAND2_X1 U17045 ( .A1(n13574), .A2(n11191), .ZN(n13575) );
  NAND2_X1 U17046 ( .A1(n15596), .A2(n13575), .ZN(n13580) );
  NAND2_X1 U17047 ( .A1(n13580), .A2(n19770), .ZN(n13577) );
  INV_X1 U17048 ( .A(n15957), .ZN(n13576) );
  NAND2_X1 U17049 ( .A1(n13577), .A2(n13576), .ZN(n13579) );
  NAND2_X1 U17050 ( .A1(n20700), .A2(n13792), .ZN(n20703) );
  NAND2_X1 U17051 ( .A1(n13579), .A2(n20059), .ZN(n20688) );
  NAND2_X1 U17052 ( .A1(n13580), .A2(n15952), .ZN(n15606) );
  INV_X1 U17053 ( .A(n15606), .ZN(n13582) );
  NOR2_X1 U17054 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13792), .ZN(n20682) );
  OAI22_X1 U17055 ( .A1(n11681), .A2(n20377), .B1(n20682), .B2(n20121), .ZN(
        n13581) );
  OAI21_X1 U17056 ( .B1(n13582), .B2(n13581), .A(n20688), .ZN(n13583) );
  OAI21_X1 U17057 ( .B1(n20688), .B2(n20446), .A(n13583), .ZN(P1_U3478) );
  OAI21_X1 U17058 ( .B1(n13587), .B2(n13586), .A(n13585), .ZN(n13861) );
  XNOR2_X1 U17059 ( .A(n13744), .B(n13746), .ZN(n19955) );
  INV_X1 U17060 ( .A(n19854), .ZN(n14392) );
  AOI22_X1 U17061 ( .A1(n19849), .A2(n19955), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14392), .ZN(n13588) );
  OAI21_X1 U17062 ( .B1(n13861), .B2(n14394), .A(n13588), .ZN(P1_U2869) );
  AND2_X1 U17063 ( .A1(n13590), .A2(n13589), .ZN(n18895) );
  XNOR2_X1 U17064 ( .A(n18895), .B(n18884), .ZN(n13594) );
  OAI21_X1 U17065 ( .B1(n13592), .B2(n13591), .A(n13902), .ZN(n18765) );
  MUX2_X1 U17066 ( .A(n10701), .B(n18765), .S(n18903), .Z(n13593) );
  OAI21_X1 U17067 ( .B1(n13594), .B2(n18893), .A(n13593), .ZN(P2_U2876) );
  XNOR2_X1 U17068 ( .A(n13595), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13596) );
  NAND2_X1 U17069 ( .A1(n13596), .A2(n18899), .ZN(n13601) );
  NOR2_X1 U17070 ( .A1(n13530), .A2(n13597), .ZN(n13598) );
  OR2_X1 U17071 ( .A1(n13544), .A2(n13598), .ZN(n16136) );
  INV_X1 U17072 ( .A(n16136), .ZN(n13599) );
  NAND2_X1 U17073 ( .A1(n18903), .A2(n13599), .ZN(n13600) );
  OAI211_X1 U17074 ( .C1(n18903), .C2(n13602), .A(n13601), .B(n13600), .ZN(
        P2_U2880) );
  INV_X1 U17075 ( .A(n19047), .ZN(n13614) );
  NAND2_X1 U17076 ( .A1(n13604), .A2(n13603), .ZN(n13605) );
  AND2_X1 U17077 ( .A1(n13605), .A2(n9921), .ZN(n13961) );
  INV_X1 U17078 ( .A(n13961), .ZN(n19708) );
  NOR2_X1 U17079 ( .A1(n19177), .A2(n19708), .ZN(n13735) );
  AOI21_X1 U17080 ( .B1(n19177), .B2(n19708), .A(n13735), .ZN(n13610) );
  INV_X1 U17081 ( .A(n13606), .ZN(n13607) );
  NAND2_X1 U17082 ( .A1(n13608), .A2(n13607), .ZN(n13609) );
  NAND2_X1 U17083 ( .A1(n13610), .A2(n13609), .ZN(n13737) );
  OAI21_X1 U17084 ( .B1(n13610), .B2(n13609), .A(n13737), .ZN(n13611) );
  NAND2_X1 U17085 ( .A1(n13611), .A2(n16024), .ZN(n13613) );
  AOI22_X1 U17086 ( .A1(n18912), .A2(n19708), .B1(n18921), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13612) );
  OAI211_X1 U17087 ( .C1(n18928), .C2(n13614), .A(n13613), .B(n13612), .ZN(
        P2_U2917) );
  OR2_X1 U17088 ( .A1(n14238), .A2(n13660), .ZN(n13629) );
  NAND2_X1 U17089 ( .A1(n12984), .A2(n13616), .ZN(n13617) );
  INV_X1 U17090 ( .A(n13617), .ZN(n13626) );
  NAND2_X1 U17091 ( .A1(n13618), .A2(n13617), .ZN(n13624) );
  INV_X1 U17092 ( .A(n13619), .ZN(n13621) );
  NAND2_X1 U17093 ( .A1(n10785), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13620) );
  NAND2_X1 U17094 ( .A1(n13621), .A2(n13620), .ZN(n13622) );
  NAND2_X1 U17095 ( .A1(n13656), .A2(n13622), .ZN(n13623) );
  NAND2_X1 U17096 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  AOI21_X1 U17097 ( .B1(n13627), .B2(n13626), .A(n13625), .ZN(n13628) );
  NAND2_X1 U17098 ( .A1(n13629), .A2(n13628), .ZN(n14023) );
  MUX2_X1 U17099 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14023), .S(
        n13654), .Z(n13670) );
  MUX2_X1 U17100 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13630), .S(
        n13654), .Z(n13669) );
  INV_X1 U17101 ( .A(n13631), .ZN(n13637) );
  OAI22_X1 U17102 ( .A1(n13637), .A2(n13634), .B1(n10629), .B2(n13633), .ZN(
        n13635) );
  AOI21_X1 U17103 ( .B1(n13637), .B2(n13636), .A(n13635), .ZN(n19736) );
  INV_X1 U17104 ( .A(n15556), .ZN(n13638) );
  NOR3_X1 U17105 ( .A1(n12821), .A2(n13639), .A3(n13638), .ZN(n13644) );
  INV_X1 U17106 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n13641) );
  AOI21_X1 U17107 ( .B1(n13642), .B2(n13641), .A(n13640), .ZN(n13643) );
  AOI211_X1 U17108 ( .C1(n13646), .C2(n13645), .A(n13644), .B(n13643), .ZN(
        n13647) );
  OAI211_X1 U17109 ( .C1(n13654), .C2(n15561), .A(n19736), .B(n13647), .ZN(
        n13668) );
  INV_X1 U17110 ( .A(n14023), .ZN(n13663) );
  NAND2_X1 U17111 ( .A1(n13656), .A2(n10472), .ZN(n13652) );
  INV_X1 U17112 ( .A(n13648), .ZN(n13649) );
  OR2_X1 U17113 ( .A1(n13650), .A2(n13649), .ZN(n13655) );
  OAI21_X1 U17114 ( .B1(n10826), .B2(n10821), .A(n13655), .ZN(n13651) );
  OAI211_X1 U17115 ( .C1(n13653), .C2(n13660), .A(n13652), .B(n13651), .ZN(
        n14029) );
  OAI21_X1 U17116 ( .B1(n14029), .B2(n19719), .A(n13654), .ZN(n13662) );
  INV_X1 U17117 ( .A(n13655), .ZN(n13658) );
  INV_X1 U17118 ( .A(n13656), .ZN(n13657) );
  MUX2_X1 U17119 ( .A(n13658), .B(n13657), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13659) );
  OAI21_X1 U17120 ( .B1(n18871), .B2(n13660), .A(n13659), .ZN(n14007) );
  AOI211_X1 U17121 ( .C1(n14029), .C2(n19719), .A(n19729), .B(n14007), .ZN(
        n13661) );
  AOI211_X1 U17122 ( .C1(n13663), .C2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n13662), .B(n13661), .ZN(n13664) );
  OAI21_X1 U17123 ( .B1(n13669), .B2(n19704), .A(n13664), .ZN(n13666) );
  NAND2_X1 U17124 ( .A1(n19704), .A2(n19710), .ZN(n19109) );
  INV_X1 U17125 ( .A(n19109), .ZN(n19142) );
  AOI22_X1 U17126 ( .A1(n13669), .A2(n19704), .B1(n13670), .B2(n19142), .ZN(
        n13665) );
  AOI21_X1 U17127 ( .B1(n13666), .B2(n13665), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n13667) );
  AOI211_X1 U17128 ( .C1(n13670), .C2(n13669), .A(n13668), .B(n13667), .ZN(
        n16168) );
  AOI21_X1 U17129 ( .B1(n16168), .B2(n14021), .A(n19751), .ZN(n13675) );
  NOR2_X1 U17130 ( .A1(n13672), .A2(n19549), .ZN(n19742) );
  OAI21_X1 U17131 ( .B1(n13671), .B2(n13673), .A(n19742), .ZN(n13674) );
  NOR2_X1 U17132 ( .A1(n13675), .A2(n13674), .ZN(n16161) );
  OAI21_X1 U17133 ( .B1(n16161), .B2(n19751), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13676) );
  INV_X1 U17134 ( .A(n16158), .ZN(n15623) );
  NAND2_X1 U17135 ( .A1(n13676), .A2(n15623), .ZN(P2_U3593) );
  AOI21_X1 U17136 ( .B1(n13535), .B2(n13677), .A(n13731), .ZN(n15362) );
  INV_X1 U17137 ( .A(n15362), .ZN(n13914) );
  INV_X1 U17138 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18948) );
  OAI222_X1 U17139 ( .A1(n18928), .A2(n14891), .B1(n13914), .B2(n18936), .C1(
        n18948), .C2(n18926), .ZN(P2_U2907) );
  INV_X1 U17140 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13679) );
  AOI22_X1 U17141 ( .A1(n19884), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13678) );
  OAI21_X1 U17142 ( .B1(n13679), .B2(n13692), .A(n13678), .ZN(P1_U2920) );
  INV_X1 U17143 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13681) );
  AOI22_X1 U17144 ( .A1(n19884), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13680) );
  OAI21_X1 U17145 ( .B1(n13681), .B2(n13692), .A(n13680), .ZN(P1_U2919) );
  INV_X1 U17146 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14424) );
  AOI22_X1 U17147 ( .A1(n20709), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13682) );
  OAI21_X1 U17148 ( .B1(n14424), .B2(n13692), .A(n13682), .ZN(P1_U2914) );
  INV_X1 U17149 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13684) );
  AOI22_X1 U17150 ( .A1(n20709), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13683) );
  OAI21_X1 U17151 ( .B1(n13684), .B2(n13692), .A(n13683), .ZN(P1_U2918) );
  INV_X1 U17152 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13686) );
  AOI22_X1 U17153 ( .A1(n20709), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13685) );
  OAI21_X1 U17154 ( .B1(n13686), .B2(n13692), .A(n13685), .ZN(P1_U2917) );
  INV_X1 U17155 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U17156 ( .A1(n20709), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13687) );
  OAI21_X1 U17157 ( .B1(n13688), .B2(n13692), .A(n13687), .ZN(P1_U2916) );
  INV_X1 U17158 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13690) );
  AOI22_X1 U17159 ( .A1(n20709), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13689) );
  OAI21_X1 U17160 ( .B1(n13690), .B2(n13692), .A(n13689), .ZN(P1_U2913) );
  INV_X1 U17161 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U17162 ( .A1(n20709), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13691) );
  OAI21_X1 U17163 ( .B1(n13693), .B2(n13692), .A(n13691), .ZN(P1_U2915) );
  AND2_X1 U17164 ( .A1(n14258), .A2(n15619), .ZN(n13694) );
  OR2_X2 U17165 ( .A1(n13695), .A2(n13694), .ZN(n19920) );
  INV_X1 U17166 ( .A(DATAI_12_), .ZN(n13697) );
  NAND2_X1 U17167 ( .A1(n20007), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13696) );
  OAI21_X1 U17168 ( .B1(n20007), .B2(n13697), .A(n13696), .ZN(n19914) );
  AOI22_X1 U17169 ( .A1(n19922), .A2(n19914), .B1(P1_UWORD_REG_12__SCAN_IN), 
        .B2(n19920), .ZN(n13698) );
  OAI21_X1 U17170 ( .B1(n12111), .B2(n19888), .A(n13698), .ZN(P1_U2949) );
  INV_X1 U17171 ( .A(DATAI_9_), .ZN(n13700) );
  NAND2_X1 U17172 ( .A1(n20007), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13699) );
  OAI21_X1 U17173 ( .B1(n20007), .B2(n13700), .A(n13699), .ZN(n19905) );
  AOI22_X1 U17174 ( .A1(n19922), .A2(n19905), .B1(P1_UWORD_REG_9__SCAN_IN), 
        .B2(n19920), .ZN(n13701) );
  OAI21_X1 U17175 ( .B1(n13702), .B2(n19888), .A(n13701), .ZN(P1_U2946) );
  INV_X1 U17176 ( .A(DATAI_13_), .ZN(n13704) );
  NAND2_X1 U17177 ( .A1(n20007), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13703) );
  OAI21_X1 U17178 ( .B1(n20007), .B2(n13704), .A(n13703), .ZN(n19917) );
  AOI22_X1 U17179 ( .A1(n19922), .A2(n19917), .B1(P1_UWORD_REG_13__SCAN_IN), 
        .B2(n19920), .ZN(n13705) );
  OAI21_X1 U17180 ( .B1(n13706), .B2(n19888), .A(n13705), .ZN(P1_U2950) );
  INV_X1 U17181 ( .A(DATAI_10_), .ZN(n13708) );
  NAND2_X1 U17182 ( .A1(n20007), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13707) );
  OAI21_X1 U17183 ( .B1(n20007), .B2(n13708), .A(n13707), .ZN(n19908) );
  AOI22_X1 U17184 ( .A1(n19922), .A2(n19908), .B1(P1_UWORD_REG_10__SCAN_IN), 
        .B2(n19920), .ZN(n13709) );
  OAI21_X1 U17185 ( .B1(n12067), .B2(n19888), .A(n13709), .ZN(P1_U2947) );
  INV_X1 U17186 ( .A(DATAI_11_), .ZN(n13711) );
  NAND2_X1 U17187 ( .A1(n20007), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13710) );
  OAI21_X1 U17188 ( .B1(n20007), .B2(n13711), .A(n13710), .ZN(n19911) );
  AOI22_X1 U17189 ( .A1(n19922), .A2(n19911), .B1(P1_UWORD_REG_11__SCAN_IN), 
        .B2(n19920), .ZN(n13712) );
  OAI21_X1 U17190 ( .B1(n13713), .B2(n19888), .A(n13712), .ZN(P1_U2948) );
  INV_X1 U17191 ( .A(DATAI_14_), .ZN(n13715) );
  NAND2_X1 U17192 ( .A1(n20007), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13714) );
  OAI21_X1 U17193 ( .B1(n20007), .B2(n13715), .A(n13714), .ZN(n19921) );
  AOI22_X1 U17194 ( .A1(n19922), .A2(n19921), .B1(P1_UWORD_REG_14__SCAN_IN), 
        .B2(n19920), .ZN(n13716) );
  OAI21_X1 U17195 ( .B1(n13717), .B2(n19888), .A(n13716), .ZN(P1_U2951) );
  NAND2_X1 U17196 ( .A1(n20005), .A2(DATAI_2_), .ZN(n13719) );
  NAND2_X1 U17197 ( .A1(n20007), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13718) );
  AND2_X1 U17198 ( .A1(n13719), .A2(n13718), .ZN(n20030) );
  INV_X1 U17199 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20850) );
  OAI222_X1 U17200 ( .A1(n14435), .A2(n13720), .B1(n20030), .B2(n14118), .C1(
        n14437), .C2(n20850), .ZN(P1_U2902) );
  NAND2_X1 U17201 ( .A1(n20005), .A2(DATAI_0_), .ZN(n13722) );
  NAND2_X1 U17202 ( .A1(n20007), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13721) );
  AND2_X1 U17203 ( .A1(n13722), .A2(n13721), .ZN(n20018) );
  INV_X1 U17204 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19887) );
  OAI222_X1 U17205 ( .A1(n14435), .A2(n13809), .B1(n20018), .B2(n14118), .C1(
        n14437), .C2(n19887), .ZN(P1_U2904) );
  INV_X1 U17206 ( .A(DATAI_8_), .ZN(n13724) );
  NAND2_X1 U17207 ( .A1(n20007), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13723) );
  OAI21_X1 U17208 ( .B1(n20007), .B2(n13724), .A(n13723), .ZN(n14415) );
  NAND2_X1 U17209 ( .A1(n19922), .A2(n14415), .ZN(n13728) );
  NAND2_X1 U17210 ( .A1(n19920), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13725) );
  OAI211_X1 U17211 ( .C1(n19888), .C2(n13726), .A(n13728), .B(n13725), .ZN(
        P1_U2945) );
  INV_X1 U17212 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19870) );
  NAND2_X1 U17213 ( .A1(n19920), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13727) );
  OAI211_X1 U17214 ( .C1(n19888), .C2(n19870), .A(n13728), .B(n13727), .ZN(
        P1_U2960) );
  INV_X1 U17215 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19879) );
  INV_X1 U17216 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16256) );
  NAND2_X1 U17217 ( .A1(n20007), .A2(n16256), .ZN(n13729) );
  OAI21_X1 U17218 ( .B1(n20007), .B2(DATAI_3_), .A(n13729), .ZN(n20033) );
  OAI222_X1 U17219 ( .A1(n13861), .A2(n14435), .B1(n14437), .B2(n19879), .C1(
        n20033), .C2(n14118), .ZN(P1_U2901) );
  INV_X1 U17220 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18946) );
  OAI21_X1 U17221 ( .B1(n13731), .B2(n13730), .A(n16119), .ZN(n18758) );
  OAI222_X1 U17222 ( .A1(n18928), .A2(n14884), .B1(n18926), .B2(n18946), .C1(
        n18936), .C2(n18758), .ZN(P2_U2906) );
  OAI21_X1 U17223 ( .B1(n13734), .B2(n13733), .A(n13732), .ZN(n19701) );
  XOR2_X1 U17224 ( .A(n19701), .B(n19320), .Z(n13739) );
  INV_X1 U17225 ( .A(n13735), .ZN(n13736) );
  NAND2_X1 U17226 ( .A1(n13737), .A2(n13736), .ZN(n13738) );
  NAND2_X1 U17227 ( .A1(n13738), .A2(n13739), .ZN(n13778) );
  OAI21_X1 U17228 ( .B1(n13739), .B2(n13738), .A(n13778), .ZN(n13740) );
  NAND2_X1 U17229 ( .A1(n13740), .A2(n16024), .ZN(n13743) );
  INV_X1 U17230 ( .A(n19701), .ZN(n13741) );
  AOI22_X1 U17231 ( .A1(n18912), .A2(n13741), .B1(n18921), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n13742) );
  OAI211_X1 U17232 ( .C1(n14961), .C2(n18928), .A(n13743), .B(n13742), .ZN(
        P2_U2916) );
  XOR2_X1 U17233 ( .A(n13585), .B(n13752), .Z(n19933) );
  INV_X1 U17234 ( .A(n19933), .ZN(n13759) );
  AOI21_X1 U17235 ( .B1(n9777), .B2(n13746), .A(n13745), .ZN(n13748) );
  INV_X1 U17236 ( .A(n13754), .ZN(n13747) );
  NOR2_X1 U17237 ( .A1(n13748), .A2(n13747), .ZN(n19949) );
  AOI22_X1 U17238 ( .A1(n19849), .A2(n19949), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14392), .ZN(n13749) );
  OAI21_X1 U17239 ( .B1(n13759), .B2(n14394), .A(n13749), .ZN(P1_U2868) );
  OAI21_X1 U17240 ( .B1(n13585), .B2(n13752), .A(n13751), .ZN(n13753) );
  AND2_X1 U17241 ( .A1(n13750), .A2(n13753), .ZN(n19816) );
  INV_X1 U17242 ( .A(n19816), .ZN(n13762) );
  AOI21_X1 U17243 ( .B1(n13755), .B2(n13754), .A(n15934), .ZN(n19806) );
  AOI22_X1 U17244 ( .A1(n19806), .A2(n19849), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14392), .ZN(n13756) );
  OAI21_X1 U17245 ( .B1(n13762), .B2(n14394), .A(n13756), .ZN(P1_U2867) );
  INV_X1 U17246 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19877) );
  NAND2_X1 U17247 ( .A1(n20005), .A2(DATAI_4_), .ZN(n13758) );
  NAND2_X1 U17248 ( .A1(n20007), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13757) );
  AND2_X1 U17249 ( .A1(n13758), .A2(n13757), .ZN(n20037) );
  OAI222_X1 U17250 ( .A1(n14435), .A2(n13759), .B1(n14437), .B2(n19877), .C1(
        n20037), .C2(n14118), .ZN(P1_U2900) );
  NAND2_X1 U17251 ( .A1(n20005), .A2(DATAI_5_), .ZN(n13761) );
  NAND2_X1 U17252 ( .A1(n20007), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13760) );
  AND2_X1 U17253 ( .A1(n13761), .A2(n13760), .ZN(n20041) );
  OAI222_X1 U17254 ( .A1(n14435), .A2(n13762), .B1(n20041), .B2(n14118), .C1(
        n14437), .C2(n11704), .ZN(P1_U2899) );
  INV_X1 U17255 ( .A(n9704), .ZN(n13815) );
  XOR2_X1 U17256 ( .A(n13815), .B(n13813), .Z(n13766) );
  INV_X1 U17257 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13764) );
  OAI21_X1 U17258 ( .B1(n13763), .B2(n13904), .A(n13819), .ZN(n16074) );
  MUX2_X1 U17259 ( .A(n13764), .B(n16074), .S(n18903), .Z(n13765) );
  OAI21_X1 U17260 ( .B1(n13766), .B2(n18893), .A(n13765), .ZN(P2_U2874) );
  OAI21_X1 U17261 ( .B1(n13769), .B2(n13768), .A(n13767), .ZN(n13770) );
  INV_X1 U17262 ( .A(n13770), .ZN(n19956) );
  NAND2_X1 U17263 ( .A1(n19956), .A2(n19935), .ZN(n13774) );
  INV_X1 U17264 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13771) );
  NOR2_X1 U17265 ( .A1(n19964), .A2(n13771), .ZN(n19954) );
  NOR2_X1 U17266 ( .A1(n19942), .A2(n13855), .ZN(n13772) );
  AOI211_X1 U17267 ( .C1(n19939), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n19954), .B(n13772), .ZN(n13773) );
  OAI211_X1 U17268 ( .C1(n20006), .C2(n13861), .A(n13774), .B(n13773), .ZN(
        P1_U2996) );
  NAND2_X1 U17269 ( .A1(n19320), .A2(n19701), .ZN(n13777) );
  XNOR2_X1 U17270 ( .A(n13732), .B(n13775), .ZN(n18835) );
  INV_X1 U17271 ( .A(n18835), .ZN(n13776) );
  AOI21_X1 U17272 ( .B1(n13778), .B2(n13777), .A(n13776), .ZN(n18932) );
  INV_X1 U17273 ( .A(n13779), .ZN(n13780) );
  NAND3_X1 U17274 ( .A1(n9715), .A2(n13781), .A3(n13780), .ZN(n13782) );
  NAND2_X1 U17275 ( .A1(n9625), .A2(n13782), .ZN(n18931) );
  XNOR2_X1 U17276 ( .A(n18932), .B(n18931), .ZN(n13786) );
  INV_X1 U17277 ( .A(n18928), .ZN(n18923) );
  OAI22_X1 U17278 ( .A1(n16018), .A2(n18835), .B1(n18926), .B2(n13783), .ZN(
        n13784) );
  AOI21_X1 U17279 ( .B1(n18923), .B2(n19057), .A(n13784), .ZN(n13785) );
  OAI21_X1 U17280 ( .B1(n13786), .B2(n18930), .A(n13785), .ZN(P2_U2915) );
  OR2_X1 U17281 ( .A1(n20780), .A2(n20703), .ZN(n15954) );
  OAI22_X1 U17282 ( .A1(n20702), .A2(n15954), .B1(n15950), .B2(n12120), .ZN(
        n13787) );
  INV_X1 U17283 ( .A(n13788), .ZN(n13789) );
  INV_X1 U17284 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13790) );
  NOR2_X1 U17285 ( .A1(n14450), .A2(n13792), .ZN(n13793) );
  NAND2_X1 U17286 ( .A1(n14251), .A2(n20706), .ZN(n13794) );
  NAND2_X1 U17287 ( .A1(n15779), .A2(n13794), .ZN(n19843) );
  INV_X1 U17288 ( .A(n19843), .ZN(n13860) );
  OR2_X1 U17289 ( .A1(n13795), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13801) );
  INV_X1 U17290 ( .A(n13801), .ZN(n13796) );
  NOR2_X1 U17291 ( .A1(n20012), .A2(n13803), .ZN(n13800) );
  NAND2_X1 U17292 ( .A1(n15659), .A2(n15685), .ZN(n19790) );
  NAND2_X1 U17293 ( .A1(n20025), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13799) );
  AND2_X1 U17294 ( .A1(n20708), .A2(n20771), .ZN(n13797) );
  NOR2_X1 U17295 ( .A1(n13799), .A2(n13797), .ZN(n13798) );
  NAND3_X1 U17296 ( .A1(n13801), .A2(n13800), .A3(n13799), .ZN(n15770) );
  OAI22_X1 U17297 ( .A1(n19994), .A2(n15773), .B1(n13802), .B2(n15770), .ZN(
        n13805) );
  NOR2_X1 U17298 ( .A1(n14257), .A2(n13803), .ZN(n19820) );
  INV_X1 U17299 ( .A(n19820), .ZN(n19841) );
  NOR2_X1 U17300 ( .A1(n20121), .A2(n19841), .ZN(n13804) );
  AOI211_X1 U17301 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n19790), .A(n13805), .B(
        n13804), .ZN(n13808) );
  OAI21_X1 U17302 ( .B1(n19838), .B2(n19837), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13807) );
  OAI211_X1 U17303 ( .C1(n13809), .C2(n13860), .A(n13808), .B(n13807), .ZN(
        P1_U2840) );
  OAI21_X1 U17304 ( .B1(n13810), .B2(n13811), .A(n15305), .ZN(n18731) );
  OAI222_X1 U17305 ( .A1(n18928), .A2(n13812), .B1(n18731), .B2(n18936), .C1(
        n13237), .C2(n18926), .ZN(P2_U2904) );
  INV_X1 U17306 ( .A(n13813), .ZN(n13814) );
  NOR2_X1 U17307 ( .A1(n13815), .A2(n13814), .ZN(n13818) );
  OAI211_X1 U17308 ( .C1(n13818), .C2(n13817), .A(n18899), .B(n13816), .ZN(
        n13825) );
  NAND2_X1 U17309 ( .A1(n13820), .A2(n13819), .ZN(n13823) );
  INV_X1 U17310 ( .A(n13821), .ZN(n13822) );
  NAND2_X1 U17311 ( .A1(n18903), .A2(n18742), .ZN(n13824) );
  OAI211_X1 U17312 ( .C1(n18903), .C2(n13826), .A(n13825), .B(n13824), .ZN(
        P2_U2873) );
  INV_X1 U17313 ( .A(n15659), .ZN(n19830) );
  NAND2_X1 U17314 ( .A1(n19830), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13828) );
  INV_X1 U17315 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20600) );
  AOI22_X1 U17316 ( .A1(n19831), .A2(n20600), .B1(n19832), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13827) );
  OAI211_X1 U17317 ( .C1(n19976), .C2(n15773), .A(n13828), .B(n13827), .ZN(
        n13831) );
  OAI22_X1 U17318 ( .A1(n19818), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13829), .B2(n19841), .ZN(n13830) );
  AOI211_X1 U17319 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19838), .A(
        n13831), .B(n13830), .ZN(n13832) );
  OAI21_X1 U17320 ( .B1(n19947), .B2(n13860), .A(n13832), .ZN(P1_U2839) );
  OAI21_X1 U17321 ( .B1(n13835), .B2(n13834), .A(n13833), .ZN(n15870) );
  OAI22_X1 U17322 ( .A1(n19992), .A2(n13837), .B1(n13838), .B2(n19970), .ZN(
        n13836) );
  NOR2_X1 U17323 ( .A1(n19961), .A2(n19948), .ZN(n13840) );
  INV_X1 U17324 ( .A(n13837), .ZN(n19962) );
  AOI21_X1 U17325 ( .B1(n14661), .B2(n13838), .A(n19981), .ZN(n19975) );
  OAI21_X1 U17326 ( .B1(n19962), .B2(n19992), .A(n19975), .ZN(n19958) );
  AOI21_X1 U17327 ( .B1(n19986), .B2(n14041), .A(n19958), .ZN(n15942) );
  INV_X1 U17328 ( .A(n15942), .ZN(n13839) );
  MUX2_X1 U17329 ( .A(n13840), .B(n13839), .S(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n13841) );
  INV_X1 U17330 ( .A(n13841), .ZN(n13843) );
  AOI22_X1 U17331 ( .A1(n19979), .A2(n19806), .B1(n19977), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n13842) );
  OAI211_X1 U17332 ( .C1(n15870), .C2(n19996), .A(n13843), .B(n13842), .ZN(
        P1_U3026) );
  XOR2_X1 U17333 ( .A(n13750), .B(n13844), .Z(n19851) );
  INV_X1 U17334 ( .A(n19851), .ZN(n13848) );
  NAND2_X1 U17335 ( .A1(n20005), .A2(DATAI_6_), .ZN(n13846) );
  NAND2_X1 U17336 ( .A1(n20007), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13845) );
  AND2_X1 U17337 ( .A1(n13846), .A2(n13845), .ZN(n20045) );
  OAI222_X1 U17338 ( .A1(n14435), .A2(n13848), .B1(n13847), .B2(n14437), .C1(
        n14118), .C2(n20045), .ZN(P1_U2898) );
  NAND2_X1 U17339 ( .A1(n19955), .A2(n19833), .ZN(n13853) );
  OAI221_X1 U17340 ( .B1(n15685), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n15685), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n15659), .ZN(n13851) );
  NOR2_X1 U17341 ( .A1(n15685), .A2(n20600), .ZN(n19835) );
  NAND2_X1 U17342 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n19835), .ZN(n13849) );
  NOR2_X1 U17343 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n13849), .ZN(n13850) );
  AOI21_X1 U17344 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n13851), .A(n13850), .ZN(
        n13852) );
  OAI211_X1 U17345 ( .C1(n13854), .C2(n15770), .A(n13853), .B(n13852), .ZN(
        n13858) );
  OAI22_X1 U17346 ( .A1(n13856), .A2(n19813), .B1(n19818), .B2(n13855), .ZN(
        n13857) );
  AOI211_X1 U17347 ( .C1(n19820), .C2(n20666), .A(n13858), .B(n13857), .ZN(
        n13859) );
  OAI21_X1 U17348 ( .B1(n13861), .B2(n13860), .A(n13859), .ZN(P1_U2837) );
  OR2_X1 U17349 ( .A1(n13863), .A2(n13862), .ZN(n13865) );
  AND2_X1 U17350 ( .A1(n13865), .A2(n13864), .ZN(n19794) );
  INV_X1 U17351 ( .A(n19794), .ZN(n13869) );
  NAND2_X1 U17352 ( .A1(n20005), .A2(DATAI_7_), .ZN(n13867) );
  NAND2_X1 U17353 ( .A1(n20007), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13866) );
  AND2_X1 U17354 ( .A1(n13867), .A2(n13866), .ZN(n20051) );
  INV_X1 U17355 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n19872) );
  OAI222_X1 U17356 ( .A1(n14435), .A2(n13869), .B1(n20051), .B2(n14118), .C1(
        n14437), .C2(n19872), .ZN(P1_U2897) );
  INV_X1 U17357 ( .A(n15936), .ZN(n13873) );
  XNOR2_X1 U17358 ( .A(n13873), .B(n13872), .ZN(n15927) );
  OAI222_X1 U17359 ( .A1(n14394), .A2(n13869), .B1(n13868), .B2(n19854), .C1(
        n14383), .C2(n15927), .ZN(P1_U2865) );
  OAI21_X1 U17360 ( .B1(n10037), .B2(n13870), .A(n9638), .ZN(n14017) );
  AOI21_X1 U17361 ( .B1(n13873), .B2(n13872), .A(n13871), .ZN(n13875) );
  INV_X1 U17362 ( .A(n13917), .ZN(n13874) );
  NOR2_X1 U17363 ( .A1(n13875), .A2(n13874), .ZN(n15921) );
  AOI22_X1 U17364 ( .A1(n15921), .A2(n19849), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14392), .ZN(n13876) );
  OAI21_X1 U17365 ( .B1(n14017), .B2(n14394), .A(n13876), .ZN(P1_U2864) );
  AOI22_X1 U17366 ( .A1(n14086), .A2(n14415), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15801), .ZN(n13877) );
  OAI21_X1 U17367 ( .B1(n14017), .B2(n14435), .A(n13877), .ZN(P1_U2896) );
  INV_X1 U17368 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20612) );
  NAND4_X1 U17369 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19791)
         );
  NAND3_X1 U17370 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n13884) );
  NOR3_X1 U17371 ( .A1(n20612), .A2(n19791), .A3(n13884), .ZN(n13999) );
  OAI21_X1 U17372 ( .B1(n13999), .B2(n15685), .A(n15659), .ZN(n13919) );
  AOI22_X1 U17373 ( .A1(n19833), .A2(n15921), .B1(P1_REIP_REG_8__SCAN_IN), 
        .B2(n13919), .ZN(n13878) );
  OAI211_X1 U17374 ( .C1(n19813), .C2(n13879), .A(n13878), .B(n19964), .ZN(
        n13887) );
  NOR2_X1 U17375 ( .A1(n15685), .A2(n19791), .ZN(n19807) );
  NAND2_X1 U17376 ( .A1(n19807), .A2(n20612), .ZN(n13885) );
  INV_X1 U17377 ( .A(n14013), .ZN(n13882) );
  NOR2_X1 U17378 ( .A1(n15770), .A2(n13880), .ZN(n13881) );
  AOI21_X1 U17379 ( .B1(n19837), .B2(n13882), .A(n13881), .ZN(n13883) );
  OAI21_X1 U17380 ( .B1(n13885), .B2(n13884), .A(n13883), .ZN(n13886) );
  NOR2_X1 U17381 ( .A1(n13887), .A2(n13886), .ZN(n13888) );
  OAI21_X1 U17382 ( .B1(n15779), .B2(n14017), .A(n13888), .ZN(P1_U2832) );
  NAND2_X1 U17383 ( .A1(n13890), .A2(n13889), .ZN(n13892) );
  XNOR2_X1 U17384 ( .A(n13892), .B(n13891), .ZN(n16148) );
  XOR2_X1 U17385 ( .A(n13894), .B(n13893), .Z(n16151) );
  NAND2_X1 U17386 ( .A1(n18822), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16144) );
  OAI21_X1 U17387 ( .B1(n16117), .B2(n20802), .A(n16144), .ZN(n13895) );
  AOI21_X1 U17388 ( .B1(n16108), .B2(n13948), .A(n13895), .ZN(n13896) );
  OAI21_X1 U17389 ( .B1(n13950), .B2(n19026), .A(n13896), .ZN(n13897) );
  AOI21_X1 U17390 ( .B1(n16151), .B2(n16113), .A(n13897), .ZN(n13898) );
  OAI21_X1 U17391 ( .B1(n16148), .B2(n18981), .A(n13898), .ZN(P2_U3011) );
  NOR2_X1 U17392 ( .A1(n10466), .A2(n13899), .ZN(n13900) );
  XNOR2_X1 U17393 ( .A(n13900), .B(n16087), .ZN(n13901) );
  NAND2_X1 U17394 ( .A1(n13901), .A2(n18827), .ZN(n13913) );
  NAND2_X1 U17395 ( .A1(n13903), .A2(n13902), .ZN(n13906) );
  INV_X1 U17396 ( .A(n13904), .ZN(n13905) );
  NOR2_X1 U17397 ( .A1(n18889), .A2(n18870), .ZN(n13910) );
  AOI22_X1 U17398 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n18866), .ZN(n13907) );
  OAI211_X1 U17399 ( .C1(n18774), .C2(n13908), .A(n13907), .B(n18772), .ZN(
        n13909) );
  AOI211_X1 U17400 ( .C1(n13911), .C2(n18865), .A(n13910), .B(n13909), .ZN(
        n13912) );
  OAI211_X1 U17401 ( .C1(n18836), .C2(n13914), .A(n13913), .B(n13912), .ZN(
        P2_U2843) );
  AOI21_X1 U17402 ( .B1(n13915), .B2(n9638), .A(n9685), .ZN(n14039) );
  INV_X1 U17403 ( .A(n14039), .ZN(n13931) );
  NAND2_X1 U17404 ( .A1(n19831), .A2(n13999), .ZN(n14094) );
  AND2_X1 U17405 ( .A1(n13917), .A2(n13916), .ZN(n13918) );
  OR2_X1 U17406 ( .A1(n13918), .A2(n13987), .ZN(n14046) );
  OAI22_X1 U17407 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n14094), .B1(n15773), 
        .B2(n14046), .ZN(n13923) );
  AOI22_X1 U17408 ( .A1(n13919), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_EBX_REG_9__SCAN_IN), .B2(n19832), .ZN(n13920) );
  OAI211_X1 U17409 ( .C1(n19813), .C2(n13921), .A(n13920), .B(n19964), .ZN(
        n13922) );
  AOI211_X1 U17410 ( .C1(n14035), .C2(n19837), .A(n13923), .B(n13922), .ZN(
        n13924) );
  OAI21_X1 U17411 ( .B1(n13931), .B2(n15779), .A(n13924), .ZN(P1_U2831) );
  XNOR2_X1 U17412 ( .A(n13816), .B(n13925), .ZN(n13930) );
  NOR2_X1 U17413 ( .A1(n13927), .A2(n13821), .ZN(n13928) );
  NOR2_X1 U17414 ( .A1(n13926), .A2(n13928), .ZN(n16058) );
  INV_X1 U17415 ( .A(n16058), .ZN(n18730) );
  MUX2_X1 U17416 ( .A(n18724), .B(n18730), .S(n18903), .Z(n13929) );
  OAI21_X1 U17417 ( .B1(n13930), .B2(n18893), .A(n13929), .ZN(P2_U2872) );
  INV_X1 U17418 ( .A(n19905), .ZN(n14410) );
  OAI222_X1 U17419 ( .A1(n13931), .A2(n14435), .B1(n14410), .B2(n14118), .C1(
        n19868), .C2(n14437), .ZN(P1_U2895) );
  OAI222_X1 U17420 ( .A1(n13931), .A2(n14394), .B1(n19854), .B2(n12635), .C1(
        n14046), .C2(n14383), .ZN(P1_U2863) );
  XNOR2_X1 U17421 ( .A(n13933), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13934) );
  XNOR2_X1 U17422 ( .A(n13932), .B(n13934), .ZN(n18979) );
  XOR2_X1 U17423 ( .A(n13936), .B(n13935), .Z(n18978) );
  NOR2_X1 U17424 ( .A1(n15410), .A2(n16156), .ZN(n15444) );
  NOR2_X1 U17425 ( .A1(n10927), .A2(n19017), .ZN(n13937) );
  AOI221_X1 U17426 ( .B1(n15444), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n15435), .C2(n13938), .A(n13937), .ZN(n13942) );
  AOI21_X1 U17427 ( .B1(n13940), .B2(n13939), .A(n13522), .ZN(n18984) );
  NAND2_X1 U17428 ( .A1(n18984), .A2(n19008), .ZN(n13941) );
  OAI211_X1 U17429 ( .C1(n16146), .C2(n18835), .A(n13942), .B(n13941), .ZN(
        n13943) );
  AOI21_X1 U17430 ( .B1(n18978), .B2(n18992), .A(n13943), .ZN(n13944) );
  OAI21_X1 U17431 ( .B1(n18996), .B2(n18979), .A(n13944), .ZN(P2_U3042) );
  INV_X1 U17432 ( .A(n18873), .ZN(n13959) );
  NAND2_X1 U17433 ( .A1(n13945), .A2(n13946), .ZN(n13947) );
  XNOR2_X1 U17434 ( .A(n13948), .B(n13947), .ZN(n13949) );
  NAND2_X1 U17435 ( .A1(n13949), .A2(n18827), .ZN(n13958) );
  INV_X1 U17436 ( .A(n13950), .ZN(n13951) );
  OAI22_X1 U17437 ( .A1(n20802), .A2(n18832), .B1(n18836), .B2(n19701), .ZN(
        n13953) );
  NOR2_X1 U17438 ( .A1(n18774), .A2(n10913), .ZN(n13952) );
  AOI211_X1 U17439 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n18866), .A(n13953), .B(
        n13952), .ZN(n13954) );
  OAI21_X1 U17440 ( .B1(n13955), .B2(n18852), .A(n13954), .ZN(n13956) );
  AOI21_X1 U17441 ( .B1(n13951), .B2(n18840), .A(n13956), .ZN(n13957) );
  OAI211_X1 U17442 ( .C1(n19320), .C2(n13959), .A(n13958), .B(n13957), .ZN(
        P2_U2852) );
  AOI22_X1 U17443 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n18866), .ZN(n13960) );
  OAI21_X1 U17444 ( .B1(n18774), .B2(n14224), .A(n13960), .ZN(n13963) );
  NOR2_X1 U17445 ( .A1(n13961), .A2(n18836), .ZN(n13962) );
  AOI211_X1 U17446 ( .C1(n18865), .C2(n13964), .A(n13963), .B(n13962), .ZN(
        n13965) );
  OAI21_X1 U17447 ( .B1(n14238), .B2(n18870), .A(n13965), .ZN(n13970) );
  INV_X1 U17448 ( .A(n13968), .ZN(n14231) );
  NOR2_X1 U17449 ( .A1(n10466), .A2(n13966), .ZN(n14018) );
  INV_X1 U17450 ( .A(n14018), .ZN(n13967) );
  AOI221_X1 U17451 ( .B1(n14231), .B2(n14018), .C1(n13968), .C2(n13967), .A(
        n18877), .ZN(n13969) );
  AOI211_X1 U17452 ( .C1(n19177), .C2(n18873), .A(n13970), .B(n13969), .ZN(
        n13971) );
  INV_X1 U17453 ( .A(n13971), .ZN(P2_U2853) );
  NAND2_X1 U17454 ( .A1(n13945), .A2(n13972), .ZN(n13973) );
  XNOR2_X1 U17455 ( .A(n15114), .B(n13973), .ZN(n13980) );
  NOR2_X1 U17456 ( .A1(n16138), .A2(n18836), .ZN(n13979) );
  AOI22_X1 U17457 ( .A1(n13974), .A2(n18865), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n18866), .ZN(n13975) );
  OAI211_X1 U17458 ( .C1(n19643), .C2(n18774), .A(n13975), .B(n18772), .ZN(
        n13976) );
  AOI21_X1 U17459 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18874), .A(
        n13976), .ZN(n13977) );
  OAI21_X1 U17460 ( .B1(n18870), .B2(n16136), .A(n13977), .ZN(n13978) );
  AOI211_X1 U17461 ( .C1(n13980), .C2(n18827), .A(n13979), .B(n13978), .ZN(
        n13981) );
  INV_X1 U17462 ( .A(n13981), .ZN(P2_U2848) );
  INV_X1 U17463 ( .A(n13983), .ZN(n13984) );
  OAI21_X1 U17464 ( .B1(n9685), .B2(n13985), .A(n13984), .ZN(n14578) );
  AOI22_X1 U17465 ( .A1(n14086), .A2(n19908), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15801), .ZN(n13986) );
  OAI21_X1 U17466 ( .B1(n14578), .B2(n14435), .A(n13986), .ZN(P1_U2894) );
  INV_X1 U17467 ( .A(n13987), .ZN(n13988) );
  AOI21_X1 U17468 ( .B1(n13989), .B2(n13988), .A(n15781), .ZN(n15910) );
  AOI22_X1 U17469 ( .A1(n15910), .A2(n19849), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14392), .ZN(n13990) );
  OAI21_X1 U17470 ( .B1(n14578), .B2(n14394), .A(n13990), .ZN(P1_U2862) );
  OAI21_X1 U17471 ( .B1(n13991), .B2(n13993), .A(n13992), .ZN(n14979) );
  NAND2_X1 U17472 ( .A1(n15100), .A2(n13994), .ZN(n13995) );
  NAND2_X1 U17473 ( .A1(n15278), .A2(n13995), .ZN(n18708) );
  NOR2_X1 U17474 ( .A1(n18888), .A2(n18708), .ZN(n13996) );
  AOI21_X1 U17475 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n18888), .A(n13996), .ZN(
        n13997) );
  OAI21_X1 U17476 ( .B1(n14979), .B2(n18893), .A(n13997), .ZN(P2_U2870) );
  NOR2_X1 U17477 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n14094), .ZN(n14004) );
  INV_X1 U17478 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13998) );
  OAI22_X1 U17479 ( .A1(n19818), .A2(n14574), .B1(n15770), .B2(n13998), .ZN(
        n14003) );
  INV_X1 U17480 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14001) );
  NAND3_X1 U17481 ( .A1(n13999), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n14213) );
  NOR2_X1 U17482 ( .A1(n19830), .A2(n14213), .ZN(n15745) );
  NOR2_X1 U17483 ( .A1(n19793), .A2(n15745), .ZN(n15786) );
  AOI22_X1 U17484 ( .A1(n19833), .A2(n15910), .B1(P1_REIP_REG_10__SCAN_IN), 
        .B2(n15786), .ZN(n14000) );
  OAI211_X1 U17485 ( .C1(n19813), .C2(n14001), .A(n14000), .B(n19964), .ZN(
        n14002) );
  AOI211_X1 U17486 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n14004), .A(n14003), .B(
        n14002), .ZN(n14005) );
  OAI21_X1 U17487 ( .B1(n15779), .B2(n14578), .A(n14005), .ZN(P1_U2830) );
  INV_X1 U17488 ( .A(n14020), .ZN(n18861) );
  AOI22_X1 U17489 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18861), .B2(n13945), .ZN(n14022) );
  AOI222_X1 U17490 ( .A1(n14007), .A2(n19693), .B1(n14006), .B2(n16163), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n14022), .ZN(n14009) );
  NAND2_X1 U17491 ( .A1(n15559), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14008) );
  OAI21_X1 U17492 ( .B1(n14009), .B2(n15559), .A(n14008), .ZN(P2_U3601) );
  XOR2_X1 U17493 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14011), .Z(
        n14012) );
  XNOR2_X1 U17494 ( .A(n14010), .B(n14012), .ZN(n15923) );
  NAND2_X1 U17495 ( .A1(n15923), .A2(n19935), .ZN(n14016) );
  NOR2_X1 U17496 ( .A1(n19964), .A2(n20612), .ZN(n15920) );
  NOR2_X1 U17497 ( .A1(n19942), .A2(n14013), .ZN(n14014) );
  AOI211_X1 U17498 ( .C1(n19939), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15920), .B(n14014), .ZN(n14015) );
  OAI211_X1 U17499 ( .C1(n20006), .C2(n14017), .A(n14016), .B(n14015), .ZN(
        P1_U2991) );
  OAI21_X1 U17500 ( .B1(n14020), .B2(n14019), .A(n14018), .ZN(n18860) );
  OAI21_X1 U17501 ( .B1(n13945), .B2(n15446), .A(n18860), .ZN(n14026) );
  NOR2_X1 U17502 ( .A1(n14022), .A2(n14021), .ZN(n14027) );
  AOI222_X1 U17503 ( .A1(n14023), .A2(n19693), .B1(n16163), .B2(n19177), .C1(
        n14026), .C2(n14027), .ZN(n14025) );
  NAND2_X1 U17504 ( .A1(n15559), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14024) );
  OAI21_X1 U17505 ( .B1(n14025), .B2(n15559), .A(n14024), .ZN(P2_U3599) );
  INV_X1 U17506 ( .A(n14026), .ZN(n14028) );
  AOI222_X1 U17507 ( .A1(n14029), .A2(n19693), .B1(n16163), .B2(n19715), .C1(
        n14028), .C2(n14027), .ZN(n14032) );
  NAND2_X1 U17508 ( .A1(n15559), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14031) );
  OAI21_X1 U17509 ( .B1(n14032), .B2(n15559), .A(n14031), .ZN(P2_U3600) );
  XNOR2_X1 U17510 ( .A(n14705), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14033) );
  XNOR2_X1 U17511 ( .A(n14034), .B(n14033), .ZN(n14050) );
  NAND2_X1 U17512 ( .A1(n15849), .A2(n14035), .ZN(n14037) );
  INV_X1 U17513 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14036) );
  OR2_X1 U17514 ( .A1(n19964), .A2(n14036), .ZN(n14045) );
  OAI211_X1 U17515 ( .C1(n15823), .C2(n13921), .A(n14037), .B(n14045), .ZN(
        n14038) );
  AOI21_X1 U17516 ( .B1(n14039), .B2(n19934), .A(n14038), .ZN(n14040) );
  OAI21_X1 U17517 ( .B1(n14050), .B2(n19943), .A(n14040), .ZN(P1_U2990) );
  NAND2_X1 U17518 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15937), .ZN(
        n15932) );
  NOR2_X1 U17519 ( .A1(n15919), .A2(n15932), .ZN(n15912) );
  INV_X1 U17520 ( .A(n14661), .ZN(n14730) );
  OAI211_X1 U17521 ( .C1(n14732), .C2(n14730), .A(n14043), .B(n14042), .ZN(
        n14044) );
  AOI21_X1 U17522 ( .B1(n14044), .B2(n19986), .A(n19981), .ZN(n15918) );
  NOR2_X1 U17523 ( .A1(n15918), .A2(n15911), .ZN(n14048) );
  OAI21_X1 U17524 ( .B1(n14046), .B2(n19995), .A(n14045), .ZN(n14047) );
  AOI211_X1 U17525 ( .C1(n15912), .C2(n15911), .A(n14048), .B(n14047), .ZN(
        n14049) );
  OAI21_X1 U17526 ( .B1(n14050), .B2(n19996), .A(n14049), .ZN(P1_U3022) );
  AOI21_X1 U17527 ( .B1(n14055), .B2(n14052), .A(n10032), .ZN(n15843) );
  INV_X1 U17528 ( .A(n15843), .ZN(n14060) );
  AOI22_X1 U17529 ( .A1(n14086), .A2(n19921), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15801), .ZN(n14056) );
  OAI21_X1 U17530 ( .B1(n14060), .B2(n14435), .A(n14056), .ZN(P1_U2890) );
  INV_X1 U17531 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14059) );
  AND2_X1 U17532 ( .A1(n14091), .A2(n14057), .ZN(n14058) );
  OR2_X1 U17533 ( .A1(n14058), .A2(n14111), .ZN(n15759) );
  OAI222_X1 U17534 ( .A1(n14060), .A2(n14394), .B1(n14059), .B2(n19854), .C1(
        n15759), .C2(n14383), .ZN(P1_U2858) );
  OR2_X1 U17535 ( .A1(n13983), .A2(n14062), .ZN(n14063) );
  AND2_X1 U17536 ( .A1(n14061), .A2(n14063), .ZN(n14077) );
  NAND2_X1 U17537 ( .A1(n14077), .A2(n14078), .ZN(n14064) );
  NAND2_X1 U17538 ( .A1(n14064), .A2(n14061), .ZN(n14068) );
  INV_X1 U17539 ( .A(n14068), .ZN(n14066) );
  INV_X1 U17540 ( .A(n14067), .ZN(n14065) );
  NAND2_X1 U17541 ( .A1(n14066), .A2(n14065), .ZN(n14069) );
  NAND2_X1 U17542 ( .A1(n14068), .A2(n14067), .ZN(n14085) );
  INV_X1 U17543 ( .A(n15780), .ZN(n14070) );
  NAND2_X1 U17544 ( .A1(n15781), .A2(n14070), .ZN(n14072) );
  NAND2_X1 U17545 ( .A1(n14072), .A2(n14071), .ZN(n14074) );
  NAND2_X1 U17546 ( .A1(n14074), .A2(n14073), .ZN(n15774) );
  OAI22_X1 U17547 ( .A1(n15774), .A2(n14383), .B1(n15769), .B2(n19854), .ZN(
        n14075) );
  AOI21_X1 U17548 ( .B1(n15847), .B2(n19850), .A(n14075), .ZN(n14076) );
  INV_X1 U17549 ( .A(n14076), .ZN(P1_U2860) );
  XOR2_X1 U17550 ( .A(n14078), .B(n14077), .Z(n15856) );
  INV_X1 U17551 ( .A(n15856), .ZN(n14080) );
  AOI22_X1 U17552 ( .A1(n14086), .A2(n19911), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15801), .ZN(n14079) );
  OAI21_X1 U17553 ( .B1(n14080), .B2(n14435), .A(n14079), .ZN(P1_U2893) );
  INV_X1 U17554 ( .A(n19914), .ZN(n14082) );
  OAI222_X1 U17555 ( .A1(n15778), .A2(n14435), .B1(n14082), .B2(n14118), .C1(
        n14081), .C2(n14437), .ZN(P1_U2892) );
  INV_X1 U17556 ( .A(n14083), .ZN(n14084) );
  AOI21_X1 U17557 ( .B1(n14085), .B2(n14084), .A(n11846), .ZN(n14566) );
  INV_X1 U17558 ( .A(n14566), .ZN(n14088) );
  AOI22_X1 U17559 ( .A1(n14086), .A2(n19917), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15801), .ZN(n14087) );
  OAI21_X1 U17560 ( .B1(n14088), .B2(n14435), .A(n14087), .ZN(P1_U2891) );
  NAND2_X1 U17561 ( .A1(n14073), .A2(n14089), .ZN(n14090) );
  NAND2_X1 U17562 ( .A1(n14091), .A2(n14090), .ZN(n14719) );
  OAI22_X1 U17563 ( .A1(n14719), .A2(n14383), .B1(n14099), .B2(n19854), .ZN(
        n14092) );
  AOI21_X1 U17564 ( .B1(n14566), .B2(n19850), .A(n14092), .ZN(n14093) );
  INV_X1 U17565 ( .A(n14093), .ZN(P1_U2859) );
  INV_X1 U17566 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20619) );
  NAND2_X1 U17567 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14095) );
  NOR2_X1 U17568 ( .A1(n14095), .A2(n14094), .ZN(n15785) );
  NAND2_X1 U17569 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15785), .ZN(n15768) );
  NOR3_X1 U17570 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n20619), .A3(n15768), 
        .ZN(n14105) );
  NAND2_X1 U17571 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14096) );
  INV_X1 U17572 ( .A(n15745), .ZN(n14321) );
  OAI21_X1 U17573 ( .B1(n14096), .B2(n14321), .A(n19790), .ZN(n15767) );
  INV_X1 U17574 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20617) );
  NOR2_X1 U17575 ( .A1(n15773), .A2(n14719), .ZN(n14097) );
  NOR2_X1 U17576 ( .A1(n19977), .A2(n14097), .ZN(n14098) );
  OAI21_X1 U17577 ( .B1(n15770), .B2(n14099), .A(n14098), .ZN(n14100) );
  AOI21_X1 U17578 ( .B1(n19838), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n14100), .ZN(n14103) );
  INV_X1 U17579 ( .A(n14564), .ZN(n14101) );
  NAND2_X1 U17580 ( .A1(n19837), .A2(n14101), .ZN(n14102) );
  OAI211_X1 U17581 ( .C1(n15767), .C2(n20617), .A(n14103), .B(n14102), .ZN(
        n14104) );
  AOI211_X1 U17582 ( .C1(n14566), .C2(n19802), .A(n14105), .B(n14104), .ZN(
        n14106) );
  INV_X1 U17583 ( .A(n14106), .ZN(P1_U2827) );
  INV_X1 U17584 ( .A(n14107), .ZN(n14108) );
  AOI21_X1 U17585 ( .B1(n14109), .B2(n14054), .A(n14108), .ZN(n14553) );
  NOR2_X1 U17586 ( .A1(n14111), .A2(n14110), .ZN(n14112) );
  OR2_X1 U17587 ( .A1(n14389), .A2(n14112), .ZN(n15758) );
  OAI22_X1 U17588 ( .A1(n15758), .A2(n14383), .B1(n14113), .B2(n19854), .ZN(
        n14114) );
  AOI21_X1 U17589 ( .B1(n14553), .B2(n19850), .A(n14114), .ZN(n14115) );
  INV_X1 U17590 ( .A(n14115), .ZN(P1_U2857) );
  INV_X1 U17591 ( .A(n14553), .ZN(n15754) );
  INV_X1 U17592 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19857) );
  NAND2_X1 U17593 ( .A1(n20005), .A2(DATAI_15_), .ZN(n14117) );
  NAND2_X1 U17594 ( .A1(n20007), .A2(BUF1_REG_15__SCAN_IN), .ZN(n14116) );
  AND2_X1 U17595 ( .A1(n14117), .A2(n14116), .ZN(n19928) );
  OAI222_X1 U17596 ( .A1(n15754), .A2(n14435), .B1(n14437), .B2(n19857), .C1(
        n14118), .C2(n19928), .ZN(P1_U2889) );
  OAI21_X1 U17597 ( .B1(n14119), .B2(n14121), .A(n14120), .ZN(n14544) );
  NOR2_X2 U17598 ( .A1(n14123), .A2(n20007), .ZN(n15804) );
  OAI22_X1 U17599 ( .A1(n20026), .A2(n14442), .B1(n14437), .B2(n13681), .ZN(
        n14122) );
  AOI21_X1 U17600 ( .B1(n15804), .B2(DATAI_17_), .A(n14122), .ZN(n14125) );
  NAND2_X1 U17601 ( .A1(n14444), .A2(BUF1_REG_17__SCAN_IN), .ZN(n14124) );
  OAI211_X1 U17602 ( .C1(n14544), .C2(n14435), .A(n14125), .B(n14124), .ZN(
        P1_U2887) );
  INV_X1 U17603 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18409) );
  OAI21_X1 U17604 ( .B1(n18432), .B2(n18572), .A(n18409), .ZN(n14134) );
  NAND2_X1 U17605 ( .A1(n18433), .A2(n14134), .ZN(n18408) );
  NOR2_X1 U17606 ( .A1(n18580), .A2(n18408), .ZN(n14133) );
  INV_X1 U17607 ( .A(n18613), .ZN(n18620) );
  NOR2_X1 U17608 ( .A1(n18620), .A2(n16311), .ZN(n14129) );
  NAND2_X1 U17609 ( .A1(n17971), .A2(n17199), .ZN(n18453) );
  AOI21_X1 U17610 ( .B1(n14129), .B2(n17137), .A(n15628), .ZN(n14130) );
  OAI211_X1 U17611 ( .C1(n15458), .C2(n15460), .A(n14131), .B(n14130), .ZN(
        n18439) );
  NOR2_X1 U17612 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18566), .ZN(n17967) );
  INV_X1 U17613 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16315) );
  NAND3_X1 U17614 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18564)
         );
  NOR2_X1 U17615 ( .A1(n16315), .A2(n18564), .ZN(n14132) );
  MUX2_X1 U17616 ( .A(n14133), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18599), .Z(P3_U3284) );
  NOR2_X1 U17617 ( .A1(n16921), .A2(n14134), .ZN(n17956) );
  OAI221_X1 U17618 ( .B1(n18564), .B2(n17956), .C1(n18564), .C2(n16315), .A(
        n18043), .ZN(n17963) );
  INV_X1 U17619 ( .A(n17963), .ZN(n17959) );
  INV_X1 U17620 ( .A(n17581), .ZN(n17453) );
  NOR2_X1 U17621 ( .A1(n17453), .A2(n18616), .ZN(n15553) );
  AOI21_X1 U17622 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15553), .ZN(n15554) );
  NOR2_X1 U17623 ( .A1(n17959), .A2(n15554), .ZN(n14136) );
  INV_X1 U17624 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18249) );
  NAND2_X1 U17625 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18249), .ZN(n18003) );
  NAND2_X1 U17626 ( .A1(n18003), .A2(n17963), .ZN(n15552) );
  OR2_X1 U17627 ( .A1(n18303), .A2(n15552), .ZN(n14135) );
  MUX2_X1 U17628 ( .A(n14136), .B(n14135), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17629 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16212) );
  XNOR2_X1 U17630 ( .A(n14137), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14465) );
  AOI22_X1 U17631 ( .A1(n12131), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11988), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U17632 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14142) );
  AOI22_X1 U17633 ( .A1(n14138), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13481), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14141) );
  AOI22_X1 U17634 ( .A1(n11370), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14140) );
  NAND4_X1 U17635 ( .A1(n14143), .A2(n14142), .A3(n14141), .A4(n14140), .ZN(
        n14152) );
  AOI22_X1 U17636 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14144), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14150) );
  AOI22_X1 U17637 ( .A1(n14146), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14145), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14149) );
  AOI22_X1 U17638 ( .A1(n11371), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11497), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U17639 ( .A1(n11355), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12058), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14147) );
  NAND4_X1 U17640 ( .A1(n14150), .A2(n14149), .A3(n14148), .A4(n14147), .ZN(
        n14151) );
  NOR2_X1 U17641 ( .A1(n14152), .A2(n14151), .ZN(n14156) );
  NOR2_X1 U17642 ( .A1(n14154), .A2(n14153), .ZN(n14155) );
  XOR2_X1 U17643 ( .A(n14156), .B(n14155), .Z(n14161) );
  AOI21_X1 U17644 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20700), .A(
        n14157), .ZN(n14159) );
  NAND2_X1 U17645 ( .A1(n11685), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n14158) );
  OAI211_X1 U17646 ( .C1(n14161), .C2(n14160), .A(n14159), .B(n14158), .ZN(
        n14162) );
  OAI21_X1 U17647 ( .B1(n12120), .B2(n14465), .A(n14162), .ZN(n14273) );
  AOI22_X1 U17648 ( .A1(n14164), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14163), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14165) );
  NAND2_X1 U17649 ( .A1(n14452), .A2(n10076), .ZN(n14168) );
  AOI22_X1 U17650 ( .A1(n15804), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15801), .ZN(n14167) );
  OAI211_X1 U17651 ( .C1(n15809), .C2(n16212), .A(n14168), .B(n14167), .ZN(
        P1_U2873) );
  AOI21_X1 U17652 ( .B1(n14169), .B2(n15111), .A(n15110), .ZN(n14172) );
  NAND2_X1 U17653 ( .A1(n10088), .A2(n14170), .ZN(n14171) );
  XNOR2_X1 U17654 ( .A(n14172), .B(n14171), .ZN(n14192) );
  NAND2_X1 U17655 ( .A1(n14174), .A2(n9837), .ZN(n14176) );
  NAND2_X1 U17656 ( .A1(n14176), .A2(n14175), .ZN(n14187) );
  NAND3_X1 U17657 ( .A1(n14173), .A2(n14187), .A3(n16152), .ZN(n14186) );
  INV_X1 U17658 ( .A(n18803), .ZN(n14184) );
  OAI22_X1 U17659 ( .A1(n16146), .A2(n18802), .B1(n10998), .B2(n18772), .ZN(
        n14183) );
  NAND2_X1 U17660 ( .A1(n14178), .A2(n14177), .ZN(n16134) );
  OAI21_X1 U17661 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n14179), .ZN(n14180) );
  OAI22_X1 U17662 ( .A1(n14181), .A2(n16134), .B1(n16135), .B2(n14180), .ZN(
        n14182) );
  AOI211_X1 U17663 ( .C1(n14184), .C2(n19008), .A(n14183), .B(n14182), .ZN(
        n14185) );
  OAI211_X1 U17664 ( .C1(n14192), .C2(n16147), .A(n14186), .B(n14185), .ZN(
        P2_U3038) );
  NAND3_X1 U17665 ( .A1(n14173), .A2(n14187), .A3(n16113), .ZN(n14191) );
  NOR2_X1 U17666 ( .A1(n18803), .A2(n19026), .ZN(n14189) );
  OAI22_X1 U17667 ( .A1(n10998), .A2(n18772), .B1(n18989), .B2(n18796), .ZN(
        n14188) );
  AOI211_X1 U17668 ( .C1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18977), .A(
        n14189), .B(n14188), .ZN(n14190) );
  OAI211_X1 U17669 ( .C1(n14192), .C2(n18981), .A(n14191), .B(n14190), .ZN(
        P2_U3006) );
  NAND2_X1 U17670 ( .A1(n14193), .A2(n14989), .ZN(n14196) );
  NOR2_X1 U17671 ( .A1(n14194), .A2(n9662), .ZN(n14195) );
  XNOR2_X1 U17672 ( .A(n14196), .B(n14195), .ZN(n14987) );
  OR3_X1 U17673 ( .A1(n15131), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14197), .ZN(n14198) );
  NAND2_X1 U17674 ( .A1(n18822), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14980) );
  OAI211_X1 U17675 ( .C1(n14199), .C2(n16137), .A(n14198), .B(n14980), .ZN(
        n14200) );
  INV_X1 U17676 ( .A(n14200), .ZN(n14205) );
  NAND2_X1 U17677 ( .A1(n14205), .A2(n14204), .ZN(n14206) );
  OAI21_X1 U17678 ( .B1(n14987), .B2(n16147), .A(n14207), .ZN(P2_U3016) );
  INV_X1 U17679 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14890) );
  AOI22_X1 U17680 ( .A1(n15803), .A2(n19917), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15801), .ZN(n14210) );
  NAND2_X1 U17681 ( .A1(n15804), .A2(DATAI_29_), .ZN(n14209) );
  OAI211_X1 U17682 ( .C1(n15809), .C2(n14890), .A(n14210), .B(n14209), .ZN(
        n14211) );
  INV_X1 U17683 ( .A(n14211), .ZN(n14212) );
  OAI21_X1 U17684 ( .B1(n14208), .B2(n14435), .A(n14212), .ZN(P1_U2875) );
  INV_X1 U17685 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20644) );
  INV_X1 U17686 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20640) );
  INV_X1 U17687 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20633) );
  INV_X1 U17688 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20839) );
  INV_X1 U17689 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20616) );
  NOR3_X1 U17690 ( .A1(n20617), .A2(n20619), .A3(n20616), .ZN(n15762) );
  AND2_X1 U17691 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15762), .ZN(n15744) );
  NAND4_X1 U17692 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(n15744), .ZN(n14322) );
  NOR2_X1 U17693 ( .A1(n14213), .A2(n14322), .ZN(n14320) );
  NAND4_X1 U17694 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14320), .A3(
        P1_REIP_REG_19__SCAN_IN), .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n15707) );
  NOR2_X1 U17695 ( .A1(n20839), .A2(n15707), .ZN(n15696) );
  NAND2_X1 U17696 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15696), .ZN(n15686) );
  NOR2_X1 U17697 ( .A1(n20633), .A2(n15686), .ZN(n15674) );
  NAND2_X1 U17698 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15674), .ZN(n15658) );
  NOR2_X1 U17699 ( .A1(n20640), .A2(n15658), .ZN(n15653) );
  NAND2_X1 U17700 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n15653), .ZN(n15648) );
  NOR2_X1 U17701 ( .A1(n20644), .A2(n15648), .ZN(n14289) );
  NAND2_X1 U17702 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n14289), .ZN(n14264) );
  NOR2_X1 U17703 ( .A1(n19830), .A2(n14264), .ZN(n14263) );
  NOR2_X1 U17704 ( .A1(n14263), .A2(n19793), .ZN(n14295) );
  NOR3_X1 U17705 ( .A1(n15685), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14264), 
        .ZN(n14214) );
  AOI21_X1 U17706 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(n19832), .A(n14214), .ZN(
        n14217) );
  NAND2_X1 U17707 ( .A1(n19837), .A2(n14215), .ZN(n14216) );
  OAI211_X1 U17708 ( .C1(n19813), .C2(n14218), .A(n14217), .B(n14216), .ZN(
        n14221) );
  OAI21_X1 U17709 ( .B1(n14296), .B2(n14219), .A(n14277), .ZN(n14590) );
  NOR2_X1 U17710 ( .A1(n14590), .A2(n15773), .ZN(n14220) );
  AOI211_X1 U17711 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14295), .A(n14221), 
        .B(n14220), .ZN(n14222) );
  OAI21_X1 U17712 ( .B1(n14208), .B2(n15779), .A(n14222), .ZN(P1_U2811) );
  INV_X1 U17713 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14223) );
  OAI222_X1 U17714 ( .A1(n14394), .A2(n14208), .B1(n14223), .B2(n19854), .C1(
        n14590), .C2(n14383), .ZN(P1_U2843) );
  INV_X1 U17715 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14225) );
  OAI22_X1 U17716 ( .A1(n16117), .A2(n14225), .B1(n14224), .B2(n19017), .ZN(
        n14230) );
  OAI21_X1 U17717 ( .B1(n14228), .B2(n14227), .A(n14226), .ZN(n18997) );
  NOR2_X1 U17718 ( .A1(n18997), .A2(n18980), .ZN(n14229) );
  AOI211_X1 U17719 ( .C1(n16108), .C2(n14231), .A(n14230), .B(n14229), .ZN(
        n14237) );
  INV_X1 U17720 ( .A(n14232), .ZN(n14235) );
  INV_X1 U17721 ( .A(n14233), .ZN(n14234) );
  NAND2_X1 U17722 ( .A1(n14235), .A2(n14234), .ZN(n18990) );
  NAND3_X1 U17723 ( .A1(n16112), .A2(n18991), .A3(n18990), .ZN(n14236) );
  OAI211_X1 U17724 ( .C1(n19026), .C2(n14238), .A(n14237), .B(n14236), .ZN(
        P2_U3012) );
  NAND2_X1 U17725 ( .A1(n14240), .A2(n14239), .ZN(n14241) );
  AND2_X1 U17726 ( .A1(n14242), .A2(n14241), .ZN(n14244) );
  MUX2_X1 U17727 ( .A(n14244), .B(n14243), .S(n14252), .Z(n14249) );
  INV_X1 U17728 ( .A(n14245), .ZN(n14247) );
  NAND2_X1 U17729 ( .A1(n14247), .A2(n14246), .ZN(n14248) );
  NAND2_X1 U17730 ( .A1(n14249), .A2(n14248), .ZN(n14250) );
  NAND2_X1 U17731 ( .A1(n14250), .A2(n11310), .ZN(n15592) );
  INV_X1 U17732 ( .A(n15592), .ZN(n14261) );
  OR2_X1 U17733 ( .A1(n14252), .A2(n14251), .ZN(n14256) );
  INV_X1 U17734 ( .A(n14253), .ZN(n14254) );
  NAND2_X1 U17735 ( .A1(n14254), .A2(n12700), .ZN(n14255) );
  NAND2_X1 U17736 ( .A1(n14256), .A2(n14255), .ZN(n19764) );
  NAND2_X1 U17737 ( .A1(n14258), .A2(n14257), .ZN(n14259) );
  AOI21_X1 U17738 ( .B1(n14259), .B2(n15620), .A(n15619), .ZN(n20705) );
  OR2_X1 U17739 ( .A1(n19764), .A2(n20705), .ZN(n15593) );
  AND2_X1 U17740 ( .A1(n15593), .A2(n14260), .ZN(n19771) );
  MUX2_X1 U17741 ( .A(P1_MORE_REG_SCAN_IN), .B(n14261), .S(n19771), .Z(
        P1_U3484) );
  NAND2_X1 U17742 ( .A1(n14452), .A2(n19802), .ZN(n14270) );
  INV_X1 U17743 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20647) );
  INV_X1 U17744 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14463) );
  NOR2_X1 U17745 ( .A1(n20647), .A2(n14463), .ZN(n14262) );
  AOI21_X1 U17746 ( .B1(n14263), .B2(n14262), .A(n19793), .ZN(n14280) );
  INV_X1 U17747 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14328) );
  NAND2_X1 U17748 ( .A1(n19838), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14267) );
  NOR3_X1 U17749 ( .A1(n15685), .A2(n14264), .A3(n20647), .ZN(n14281) );
  INV_X1 U17750 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14265) );
  NAND3_X1 U17751 ( .A1(n14281), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n14265), 
        .ZN(n14266) );
  OAI211_X1 U17752 ( .C1(n14328), .C2(n15770), .A(n14267), .B(n14266), .ZN(
        n14268) );
  AOI21_X1 U17753 ( .B1(n14280), .B2(P1_REIP_REG_31__SCAN_IN), .A(n14268), 
        .ZN(n14269) );
  OAI211_X1 U17754 ( .C1(n14329), .C2(n15773), .A(n14270), .B(n14269), .ZN(
        P1_U2809) );
  AOI21_X1 U17755 ( .B1(n14273), .B2(n14272), .A(n14271), .ZN(n14467) );
  INV_X1 U17756 ( .A(n14467), .ZN(n14400) );
  INV_X1 U17757 ( .A(n14274), .ZN(n14275) );
  AOI22_X1 U17758 ( .A1(n14277), .A2(n14276), .B1(n14275), .B2(n14296), .ZN(
        n14279) );
  OAI21_X1 U17759 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14281), .A(n14280), 
        .ZN(n14283) );
  AOI22_X1 U17760 ( .A1(n19838), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n19832), .ZN(n14282) );
  OAI211_X1 U17761 ( .C1(n14465), .C2(n19818), .A(n14283), .B(n14282), .ZN(
        n14284) );
  AOI21_X1 U17762 ( .B1(n14584), .B2(n19833), .A(n14284), .ZN(n14285) );
  OAI21_X1 U17763 ( .B1(n14400), .B2(n15779), .A(n14285), .ZN(P1_U2810) );
  INV_X1 U17764 ( .A(n14479), .ZN(n14333) );
  NOR2_X1 U17765 ( .A1(n19818), .A2(n14477), .ZN(n14294) );
  INV_X1 U17766 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14288) );
  NAND3_X1 U17767 ( .A1(n19831), .A2(n14289), .A3(n14288), .ZN(n14291) );
  NAND2_X1 U17768 ( .A1(n19832), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14290) );
  OAI211_X1 U17769 ( .C1(n19813), .C2(n14292), .A(n14291), .B(n14290), .ZN(
        n14293) );
  AOI211_X1 U17770 ( .C1(n14295), .C2(P1_REIP_REG_28__SCAN_IN), .A(n14294), 
        .B(n14293), .ZN(n14299) );
  AOI21_X1 U17771 ( .B1(n14297), .B2(n14302), .A(n14296), .ZN(n14595) );
  NAND2_X1 U17772 ( .A1(n14595), .A2(n19833), .ZN(n14298) );
  OAI211_X1 U17773 ( .C1(n14333), .C2(n15779), .A(n14299), .B(n14298), .ZN(
        P1_U2812) );
  NAND2_X1 U17774 ( .A1(n14614), .A2(n14300), .ZN(n14301) );
  NAND2_X1 U17775 ( .A1(n14302), .A2(n14301), .ZN(n14604) );
  NAND2_X1 U17776 ( .A1(n14488), .A2(n19802), .ZN(n14311) );
  NOR3_X1 U17777 ( .A1(n15648), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n15685), 
        .ZN(n14306) );
  AOI21_X1 U17778 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(n19832), .A(n14306), .ZN(
        n14307) );
  OAI21_X1 U17779 ( .B1(n19813), .B2(n14486), .A(n14307), .ZN(n14309) );
  OAI21_X1 U17780 ( .B1(n19830), .B2(n15648), .A(n19790), .ZN(n15650) );
  NOR2_X1 U17781 ( .A1(n15650), .A2(n20644), .ZN(n14308) );
  AOI211_X1 U17782 ( .C1(n19837), .C2(n14484), .A(n14309), .B(n14308), .ZN(
        n14310) );
  OAI211_X1 U17783 ( .C1(n15773), .C2(n14604), .A(n14311), .B(n14310), .ZN(
        P1_U2813) );
  AOI21_X1 U17784 ( .B1(n14315), .B2(n14313), .A(n14314), .ZN(n14532) );
  INV_X1 U17785 ( .A(n14532), .ZN(n14436) );
  AND2_X1 U17786 ( .A1(n14376), .A2(n14316), .ZN(n14317) );
  OR2_X1 U17787 ( .A1(n14317), .A2(n14654), .ZN(n14677) );
  INV_X1 U17788 ( .A(n14677), .ZN(n14326) );
  AOI21_X1 U17789 ( .B1(n19832), .B2(P1_EBX_REG_19__SCAN_IN), .A(n19977), .ZN(
        n14319) );
  NAND2_X1 U17790 ( .A1(n19837), .A2(n14529), .ZN(n14318) );
  OAI211_X1 U17791 ( .C1(n19813), .C2(n11933), .A(n14319), .B(n14318), .ZN(
        n14325) );
  INV_X1 U17792 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20630) );
  INV_X1 U17793 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20628) );
  NOR2_X1 U17794 ( .A1(n20630), .A2(n20628), .ZN(n15716) );
  AND2_X1 U17795 ( .A1(n19831), .A2(n14320), .ZN(n15725) );
  OAI21_X1 U17796 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15725), .ZN(n14323) );
  OAI21_X1 U17797 ( .B1(n14322), .B2(n14321), .A(n19790), .ZN(n15739) );
  OAI22_X1 U17798 ( .A1(n15716), .A2(n14323), .B1(n20630), .B2(n15739), .ZN(
        n14324) );
  AOI211_X1 U17799 ( .C1(n14326), .C2(n19833), .A(n14325), .B(n14324), .ZN(
        n14327) );
  OAI21_X1 U17800 ( .B1(n14436), .B2(n15779), .A(n14327), .ZN(P1_U2821) );
  OAI22_X1 U17801 ( .A1(n14329), .A2(n14383), .B1(n19854), .B2(n14328), .ZN(
        P1_U2841) );
  INV_X1 U17802 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14331) );
  OAI222_X1 U17803 ( .A1(n14394), .A2(n14400), .B1(n14331), .B2(n19854), .C1(
        n14330), .C2(n14383), .ZN(P1_U2842) );
  AOI22_X1 U17804 ( .A1(n14595), .A2(n19849), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14392), .ZN(n14332) );
  OAI21_X1 U17805 ( .B1(n14333), .B2(n14394), .A(n14332), .ZN(P1_U2844) );
  INV_X1 U17806 ( .A(n14488), .ZN(n14335) );
  OAI222_X1 U17807 ( .A1(n14394), .A2(n14335), .B1(n14334), .B2(n19854), .C1(
        n14604), .C2(n14383), .ZN(P1_U2845) );
  OR2_X1 U17808 ( .A1(n14337), .A2(n14338), .ZN(n14339) );
  NAND2_X1 U17809 ( .A1(n14336), .A2(n14339), .ZN(n15668) );
  NOR2_X1 U17810 ( .A1(n14347), .A2(n14340), .ZN(n14341) );
  OR2_X1 U17811 ( .A1(n14612), .A2(n14341), .ZN(n15672) );
  OAI22_X1 U17812 ( .A1(n15672), .A2(n14383), .B1(n15661), .B2(n19854), .ZN(
        n14342) );
  INV_X1 U17813 ( .A(n14342), .ZN(n14343) );
  OAI21_X1 U17814 ( .B1(n15668), .B2(n14394), .A(n14343), .ZN(P1_U2847) );
  NOR2_X1 U17815 ( .A1(n14344), .A2(n14345), .ZN(n14346) );
  OR2_X1 U17816 ( .A1(n14337), .A2(n14346), .ZN(n14414) );
  AOI21_X1 U17817 ( .B1(n14348), .B2(n14355), .A(n14347), .ZN(n15679) );
  AOI22_X1 U17818 ( .A1(n15679), .A2(n19849), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14392), .ZN(n14349) );
  OAI21_X1 U17819 ( .B1(n14414), .B2(n14394), .A(n14349), .ZN(P1_U2848) );
  INV_X1 U17820 ( .A(n14350), .ZN(n14351) );
  AOI21_X1 U17821 ( .B1(n14352), .B2(n14351), .A(n14344), .ZN(n14420) );
  NAND2_X1 U17822 ( .A1(n14361), .A2(n14353), .ZN(n14354) );
  NAND2_X1 U17823 ( .A1(n14355), .A2(n14354), .ZN(n15689) );
  OAI22_X1 U17824 ( .A1(n15689), .A2(n14383), .B1(n14356), .B2(n19854), .ZN(
        n14357) );
  AOI21_X1 U17825 ( .B1(n14420), .B2(n19850), .A(n14357), .ZN(n14358) );
  INV_X1 U17826 ( .A(n14358), .ZN(P1_U2849) );
  OR2_X1 U17827 ( .A1(n14368), .A2(n14359), .ZN(n14360) );
  NAND2_X1 U17828 ( .A1(n14361), .A2(n14360), .ZN(n15703) );
  INV_X1 U17829 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15698) );
  AOI21_X1 U17830 ( .B1(n14363), .B2(n14362), .A(n14350), .ZN(n15813) );
  INV_X1 U17831 ( .A(n15813), .ZN(n14428) );
  OAI222_X1 U17832 ( .A1(n15703), .A2(n14383), .B1(n15698), .B2(n19854), .C1(
        n14428), .C2(n14394), .ZN(P1_U2850) );
  OAI21_X1 U17833 ( .B1(n14364), .B2(n14365), .A(n14362), .ZN(n15710) );
  NOR2_X1 U17834 ( .A1(n14656), .A2(n14366), .ZN(n14367) );
  OR2_X1 U17835 ( .A1(n14368), .A2(n14367), .ZN(n15709) );
  OAI22_X1 U17836 ( .A1(n15709), .A2(n14383), .B1(n14369), .B2(n19854), .ZN(
        n14370) );
  INV_X1 U17837 ( .A(n14370), .ZN(n14371) );
  OAI21_X1 U17838 ( .B1(n15710), .B2(n14394), .A(n14371), .ZN(P1_U2851) );
  OAI22_X1 U17839 ( .A1(n14677), .A2(n14383), .B1(n20863), .B2(n19854), .ZN(
        n14372) );
  AOI21_X1 U17840 ( .B1(n14532), .B2(n19850), .A(n14372), .ZN(n14373) );
  INV_X1 U17841 ( .A(n14373), .ZN(P1_U2853) );
  NAND2_X1 U17842 ( .A1(n14382), .A2(n14374), .ZN(n14375) );
  NAND2_X1 U17843 ( .A1(n14376), .A2(n14375), .ZN(n15889) );
  INV_X1 U17844 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14379) );
  NAND2_X1 U17845 ( .A1(n14120), .A2(n14377), .ZN(n14378) );
  NAND2_X1 U17846 ( .A1(n14313), .A2(n14378), .ZN(n15827) );
  OAI222_X1 U17847 ( .A1(n15889), .A2(n14383), .B1(n14379), .B2(n19854), .C1(
        n15827), .C2(n14394), .ZN(P1_U2854) );
  INV_X1 U17848 ( .A(n14544), .ZN(n15736) );
  NAND2_X1 U17849 ( .A1(n14391), .A2(n14380), .ZN(n14381) );
  NAND2_X1 U17850 ( .A1(n14382), .A2(n14381), .ZN(n15734) );
  OAI22_X1 U17851 ( .A1(n15734), .A2(n14383), .B1(n15731), .B2(n19854), .ZN(
        n14384) );
  AOI21_X1 U17852 ( .B1(n15736), .B2(n19850), .A(n14384), .ZN(n14385) );
  INV_X1 U17853 ( .A(n14385), .ZN(P1_U2855) );
  AND2_X1 U17854 ( .A1(n14107), .A2(n14386), .ZN(n14387) );
  NOR2_X1 U17855 ( .A1(n14119), .A2(n14387), .ZN(n15838) );
  INV_X1 U17856 ( .A(n15838), .ZN(n14447) );
  OR2_X1 U17857 ( .A1(n14389), .A2(n14388), .ZN(n14390) );
  AND2_X1 U17858 ( .A1(n14391), .A2(n14390), .ZN(n15898) );
  AOI22_X1 U17859 ( .A1(n15898), .A2(n19849), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14392), .ZN(n14393) );
  OAI21_X1 U17860 ( .B1(n14447), .B2(n14394), .A(n14393), .ZN(P1_U2856) );
  AOI22_X1 U17861 ( .A1(n15803), .A2(n19921), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n15801), .ZN(n14396) );
  NAND2_X1 U17862 ( .A1(n15804), .A2(DATAI_30_), .ZN(n14395) );
  OAI211_X1 U17863 ( .C1(n15809), .C2(n14397), .A(n14396), .B(n14395), .ZN(
        n14398) );
  INV_X1 U17864 ( .A(n14398), .ZN(n14399) );
  OAI21_X1 U17865 ( .B1(n14400), .B2(n14435), .A(n14399), .ZN(P1_U2874) );
  INV_X1 U17866 ( .A(n14435), .ZN(n15805) );
  NAND2_X1 U17867 ( .A1(n14479), .A2(n15805), .ZN(n14404) );
  AOI22_X1 U17868 ( .A1(n15803), .A2(n19914), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n15801), .ZN(n14403) );
  NAND2_X1 U17869 ( .A1(n14444), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14402) );
  NAND2_X1 U17870 ( .A1(n15804), .A2(DATAI_28_), .ZN(n14401) );
  NAND4_X1 U17871 ( .A1(n14404), .A2(n14403), .A3(n14402), .A4(n14401), .ZN(
        P1_U2876) );
  NAND2_X1 U17872 ( .A1(n14488), .A2(n15805), .ZN(n14408) );
  AOI22_X1 U17873 ( .A1(n15803), .A2(n19911), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15801), .ZN(n14407) );
  NAND2_X1 U17874 ( .A1(n14444), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14406) );
  NAND2_X1 U17875 ( .A1(n15804), .A2(DATAI_27_), .ZN(n14405) );
  NAND4_X1 U17876 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        P1_U2877) );
  NAND2_X1 U17877 ( .A1(n15801), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n14409) );
  OAI21_X1 U17878 ( .B1(n14442), .B2(n14410), .A(n14409), .ZN(n14411) );
  AOI21_X1 U17879 ( .B1(n15804), .B2(DATAI_25_), .A(n14411), .ZN(n14413) );
  NAND2_X1 U17880 ( .A1(n14444), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14412) );
  OAI211_X1 U17881 ( .C1(n15668), .C2(n14435), .A(n14413), .B(n14412), .ZN(
        P1_U2879) );
  NAND2_X1 U17882 ( .A1(n15680), .A2(n15805), .ZN(n14419) );
  AOI22_X1 U17883 ( .A1(n15803), .A2(n14415), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n15801), .ZN(n14418) );
  NAND2_X1 U17884 ( .A1(n14444), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14417) );
  NAND2_X1 U17885 ( .A1(n15804), .A2(DATAI_24_), .ZN(n14416) );
  NAND4_X1 U17886 ( .A1(n14419), .A2(n14418), .A3(n14417), .A4(n14416), .ZN(
        P1_U2880) );
  INV_X1 U17887 ( .A(n14420), .ZN(n15690) );
  OAI22_X1 U17888 ( .A1(n20051), .A2(n14442), .B1(n14437), .B2(n13690), .ZN(
        n14421) );
  AOI21_X1 U17889 ( .B1(n15804), .B2(DATAI_23_), .A(n14421), .ZN(n14423) );
  NAND2_X1 U17890 ( .A1(n14444), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14422) );
  OAI211_X1 U17891 ( .C1(n15690), .C2(n14435), .A(n14423), .B(n14422), .ZN(
        P1_U2881) );
  OAI22_X1 U17892 ( .A1(n20045), .A2(n14442), .B1(n14437), .B2(n14424), .ZN(
        n14425) );
  AOI21_X1 U17893 ( .B1(n15804), .B2(DATAI_22_), .A(n14425), .ZN(n14427) );
  NAND2_X1 U17894 ( .A1(n14444), .A2(BUF1_REG_22__SCAN_IN), .ZN(n14426) );
  OAI211_X1 U17895 ( .C1(n14428), .C2(n14435), .A(n14427), .B(n14426), .ZN(
        P1_U2882) );
  OAI22_X1 U17896 ( .A1(n20041), .A2(n14442), .B1(n14437), .B2(n13693), .ZN(
        n14429) );
  AOI21_X1 U17897 ( .B1(n15804), .B2(DATAI_21_), .A(n14429), .ZN(n14431) );
  NAND2_X1 U17898 ( .A1(n14444), .A2(BUF1_REG_21__SCAN_IN), .ZN(n14430) );
  OAI211_X1 U17899 ( .C1(n15710), .C2(n14435), .A(n14431), .B(n14430), .ZN(
        P1_U2883) );
  OAI22_X1 U17900 ( .A1(n14442), .A2(n20033), .B1(n14437), .B2(n13686), .ZN(
        n14432) );
  AOI21_X1 U17901 ( .B1(n15804), .B2(DATAI_19_), .A(n14432), .ZN(n14434) );
  NAND2_X1 U17902 ( .A1(n14444), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14433) );
  OAI211_X1 U17903 ( .C1(n14436), .C2(n14435), .A(n14434), .B(n14433), .ZN(
        P1_U2885) );
  OAI22_X1 U17904 ( .A1(n20030), .A2(n14442), .B1(n14437), .B2(n13684), .ZN(
        n14438) );
  AOI21_X1 U17905 ( .B1(n15804), .B2(DATAI_18_), .A(n14438), .ZN(n14440) );
  NAND2_X1 U17906 ( .A1(n14444), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14439) );
  OAI211_X1 U17907 ( .C1(n15827), .C2(n14435), .A(n14440), .B(n14439), .ZN(
        P1_U2886) );
  NAND2_X1 U17908 ( .A1(n15801), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n14441) );
  OAI21_X1 U17909 ( .B1(n14442), .B2(n20018), .A(n14441), .ZN(n14443) );
  AOI21_X1 U17910 ( .B1(n15804), .B2(DATAI_16_), .A(n14443), .ZN(n14446) );
  NAND2_X1 U17911 ( .A1(n14444), .A2(BUF1_REG_16__SCAN_IN), .ZN(n14445) );
  OAI211_X1 U17912 ( .C1(n14447), .C2(n14435), .A(n14446), .B(n14445), .ZN(
        P1_U2888) );
  NAND2_X1 U17913 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14448) );
  OAI211_X1 U17914 ( .C1(n19942), .C2(n14450), .A(n14449), .B(n14448), .ZN(
        n14451) );
  AOI21_X1 U17915 ( .B1(n14452), .B2(n19934), .A(n14451), .ZN(n14453) );
  OAI21_X1 U17916 ( .B1(n14454), .B2(n19943), .A(n14453), .ZN(P1_U2968) );
  INV_X1 U17917 ( .A(n14455), .ZN(n14457) );
  NOR2_X1 U17918 ( .A1(n14705), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14456) );
  NAND2_X1 U17919 ( .A1(n14457), .A2(n14456), .ZN(n14461) );
  NAND3_X1 U17920 ( .A1(n14461), .A2(n14462), .A3(n14458), .ZN(n14459) );
  OAI211_X1 U17921 ( .C1(n14462), .C2(n14461), .A(n14460), .B(n14459), .ZN(
        n14585) );
  NOR2_X1 U17922 ( .A1(n19964), .A2(n14463), .ZN(n14583) );
  AOI21_X1 U17923 ( .B1(n19939), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14583), .ZN(n14464) );
  OAI21_X1 U17924 ( .B1(n19942), .B2(n14465), .A(n14464), .ZN(n14466) );
  AOI21_X1 U17925 ( .B1(n14467), .B2(n19934), .A(n14466), .ZN(n14468) );
  OAI21_X1 U17926 ( .B1(n19943), .B2(n14585), .A(n14468), .ZN(P1_U2969) );
  INV_X1 U17927 ( .A(n14469), .ZN(n14490) );
  NAND2_X1 U17928 ( .A1(n14539), .A2(n14471), .ZN(n14491) );
  NAND3_X1 U17929 ( .A1(n14470), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14491), .ZN(n14472) );
  OAI21_X1 U17930 ( .B1(n14490), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14472), .ZN(n14474) );
  MUX2_X1 U17931 ( .A(n11616), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n14539), .Z(n14473) );
  NAND2_X1 U17932 ( .A1(n14474), .A2(n14473), .ZN(n14475) );
  XOR2_X1 U17933 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14475), .Z(
        n14601) );
  NAND2_X1 U17934 ( .A1(n19977), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U17935 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14476) );
  OAI211_X1 U17936 ( .C1(n19942), .C2(n14477), .A(n14596), .B(n14476), .ZN(
        n14478) );
  AOI21_X1 U17937 ( .B1(n14479), .B2(n19934), .A(n14478), .ZN(n14480) );
  OAI21_X1 U17938 ( .B1(n19943), .B2(n14601), .A(n14480), .ZN(P1_U2971) );
  MUX2_X1 U17939 ( .A(n14482), .B(n14481), .S(n9634), .Z(n14483) );
  XNOR2_X1 U17940 ( .A(n14483), .B(n11616), .ZN(n14609) );
  NAND2_X1 U17941 ( .A1(n15849), .A2(n14484), .ZN(n14485) );
  OR2_X1 U17942 ( .A1(n19964), .A2(n20644), .ZN(n14602) );
  OAI211_X1 U17943 ( .C1(n15823), .C2(n14486), .A(n14485), .B(n14602), .ZN(
        n14487) );
  AOI21_X1 U17944 ( .B1(n14488), .B2(n19934), .A(n14487), .ZN(n14489) );
  OAI21_X1 U17945 ( .B1(n19943), .B2(n14609), .A(n14489), .ZN(P1_U2972) );
  INV_X1 U17946 ( .A(n14470), .ZN(n14509) );
  OAI21_X1 U17947 ( .B1(n9634), .B2(n14509), .A(n14490), .ZN(n14492) );
  NAND2_X1 U17948 ( .A1(n14492), .A2(n14491), .ZN(n14493) );
  XOR2_X1 U17949 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14493), .Z(
        n14620) );
  NAND2_X1 U17950 ( .A1(n14336), .A2(n14494), .ZN(n14495) );
  AND2_X1 U17951 ( .A1(n14496), .A2(n14495), .ZN(n15798) );
  INV_X1 U17952 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14497) );
  OR2_X1 U17953 ( .A1(n19964), .A2(n14497), .ZN(n14617) );
  NAND2_X1 U17954 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14498) );
  OAI211_X1 U17955 ( .C1(n19942), .C2(n15657), .A(n14617), .B(n14498), .ZN(
        n14499) );
  AOI21_X1 U17956 ( .B1(n15798), .B2(n19934), .A(n14499), .ZN(n14500) );
  OAI21_X1 U17957 ( .B1(n14620), .B2(n19943), .A(n14500), .ZN(P1_U2973) );
  NAND2_X1 U17958 ( .A1(n14501), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14510) );
  NOR2_X1 U17959 ( .A1(n14510), .A2(n14512), .ZN(n14504) );
  NOR2_X1 U17960 ( .A1(n14502), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14503) );
  MUX2_X1 U17961 ( .A(n14504), .B(n14503), .S(n9634), .Z(n14505) );
  XNOR2_X1 U17962 ( .A(n14505), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14628) );
  OR2_X1 U17963 ( .A1(n19964), .A2(n20640), .ZN(n14624) );
  OAI21_X1 U17964 ( .B1(n15823), .B2(n15662), .A(n14624), .ZN(n14507) );
  NOR2_X1 U17965 ( .A1(n15668), .A2(n20006), .ZN(n14506) );
  AOI211_X1 U17966 ( .C1(n15849), .C2(n15666), .A(n14507), .B(n14506), .ZN(
        n14508) );
  OAI21_X1 U17967 ( .B1(n19943), .B2(n14628), .A(n14508), .ZN(P1_U2974) );
  NAND2_X1 U17968 ( .A1(n14509), .A2(n9634), .ZN(n14511) );
  MUX2_X1 U17969 ( .A(n9634), .B(n14511), .S(n14510), .Z(n14513) );
  XNOR2_X1 U17970 ( .A(n14513), .B(n14512), .ZN(n14635) );
  INV_X1 U17971 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n15677) );
  NOR2_X1 U17972 ( .A1(n19964), .A2(n15677), .ZN(n14630) );
  AOI21_X1 U17973 ( .B1(n19939), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14630), .ZN(n14514) );
  OAI21_X1 U17974 ( .B1(n19942), .B2(n15683), .A(n14514), .ZN(n14515) );
  AOI21_X1 U17975 ( .B1(n15680), .B2(n19934), .A(n14515), .ZN(n14516) );
  OAI21_X1 U17976 ( .B1(n14635), .B2(n19943), .A(n14516), .ZN(P1_U2975) );
  XNOR2_X1 U17977 ( .A(n14705), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14517) );
  XNOR2_X1 U17978 ( .A(n14470), .B(n14517), .ZN(n14643) );
  OAI22_X1 U17979 ( .A1(n15823), .A2(n15695), .B1(n19964), .B2(n20633), .ZN(
        n14519) );
  NOR2_X1 U17980 ( .A1(n15690), .A2(n20006), .ZN(n14518) );
  AOI211_X1 U17981 ( .C1(n15849), .C2(n15692), .A(n14519), .B(n14518), .ZN(
        n14520) );
  OAI21_X1 U17982 ( .B1(n14643), .B2(n19943), .A(n14520), .ZN(P1_U2976) );
  NOR2_X1 U17983 ( .A1(n14521), .A2(n9634), .ZN(n14650) );
  OAI22_X1 U17984 ( .A1(n14650), .A2(n9669), .B1(n9634), .B2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14522) );
  XNOR2_X1 U17985 ( .A(n14522), .B(n11611), .ZN(n14649) );
  NAND2_X1 U17986 ( .A1(n19977), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14645) );
  OAI21_X1 U17987 ( .B1(n15823), .B2(n15715), .A(n14645), .ZN(n14524) );
  NOR2_X1 U17988 ( .A1(n15710), .A2(n20006), .ZN(n14523) );
  AOI211_X1 U17989 ( .C1(n15849), .C2(n15712), .A(n14524), .B(n14523), .ZN(
        n14525) );
  OAI21_X1 U17990 ( .B1(n19943), .B2(n14649), .A(n14525), .ZN(P1_U2978) );
  NOR2_X1 U17991 ( .A1(n14705), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14527) );
  MUX2_X1 U17992 ( .A(n14539), .B(n14527), .S(n14526), .Z(n14528) );
  XNOR2_X1 U17993 ( .A(n14528), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14681) );
  NAND2_X1 U17994 ( .A1(n15849), .A2(n14529), .ZN(n14530) );
  NAND2_X1 U17995 ( .A1(n19977), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14675) );
  OAI211_X1 U17996 ( .C1(n15823), .C2(n11933), .A(n14530), .B(n14675), .ZN(
        n14531) );
  AOI21_X1 U17997 ( .B1(n14532), .B2(n19934), .A(n14531), .ZN(n14533) );
  OAI21_X1 U17998 ( .B1(n19943), .B2(n14681), .A(n14533), .ZN(P1_U2980) );
  NAND2_X1 U17999 ( .A1(n14534), .A2(n14535), .ZN(n14703) );
  NAND3_X1 U18000 ( .A1(n14703), .A2(n14702), .A3(n14536), .ZN(n14538) );
  OAI21_X1 U18001 ( .B1(n14539), .B2(n15895), .A(n14549), .ZN(n15835) );
  NAND2_X1 U18002 ( .A1(n15835), .A2(n14540), .ZN(n15832) );
  MUX2_X1 U18003 ( .A(n15835), .B(n15832), .S(n14541), .Z(n14542) );
  XNOR2_X1 U18004 ( .A(n14542), .B(n14682), .ZN(n14694) );
  NAND2_X1 U18005 ( .A1(n19977), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n14690) );
  OAI21_X1 U18006 ( .B1(n15823), .B2(n14543), .A(n14690), .ZN(n14546) );
  NOR2_X1 U18007 ( .A1(n14544), .A2(n20006), .ZN(n14545) );
  AOI211_X1 U18008 ( .C1(n15849), .C2(n15733), .A(n14546), .B(n14545), .ZN(
        n14547) );
  OAI21_X1 U18009 ( .B1(n14694), .B2(n19943), .A(n14547), .ZN(P1_U2982) );
  XNOR2_X1 U18010 ( .A(n14705), .B(n15895), .ZN(n14548) );
  XNOR2_X1 U18011 ( .A(n14549), .B(n14548), .ZN(n14699) );
  AOI22_X1 U18012 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14550) );
  OAI21_X1 U18013 ( .B1(n19942), .B2(n14551), .A(n14550), .ZN(n14552) );
  AOI21_X1 U18014 ( .B1(n14553), .B2(n19934), .A(n14552), .ZN(n14554) );
  OAI21_X1 U18015 ( .B1(n14699), .B2(n19943), .A(n14554), .ZN(P1_U2984) );
  INV_X1 U18016 ( .A(n14555), .ZN(n14556) );
  OR2_X1 U18017 ( .A1(n14534), .A2(n14556), .ZN(n14558) );
  NAND2_X1 U18018 ( .A1(n14558), .A2(n14557), .ZN(n14728) );
  NAND2_X1 U18019 ( .A1(n14559), .A2(n14560), .ZN(n14727) );
  NAND2_X1 U18020 ( .A1(n14725), .A2(n14560), .ZN(n14562) );
  XNOR2_X1 U18021 ( .A(n14562), .B(n14561), .ZN(n14724) );
  AOI22_X1 U18022 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14563) );
  OAI21_X1 U18023 ( .B1(n19942), .B2(n14564), .A(n14563), .ZN(n14565) );
  AOI21_X1 U18024 ( .B1(n14566), .B2(n19934), .A(n14565), .ZN(n14567) );
  OAI21_X1 U18025 ( .B1(n14724), .B2(n19943), .A(n14567), .ZN(P1_U2986) );
  XOR2_X1 U18026 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n14534), .Z(
        n14570) );
  NAND2_X1 U18027 ( .A1(n14568), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14569) );
  MUX2_X1 U18028 ( .A(n14570), .B(n14569), .S(n9634), .Z(n14572) );
  NOR3_X1 U18029 ( .A1(n14568), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14705), .ZN(n15853) );
  INV_X1 U18030 ( .A(n15853), .ZN(n14571) );
  NAND2_X1 U18031 ( .A1(n14572), .A2(n14571), .ZN(n15914) );
  NAND2_X1 U18032 ( .A1(n15914), .A2(n19935), .ZN(n14577) );
  INV_X1 U18033 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14573) );
  NOR2_X1 U18034 ( .A1(n19964), .A2(n14573), .ZN(n15909) );
  NOR2_X1 U18035 ( .A1(n19942), .A2(n14574), .ZN(n14575) );
  AOI211_X1 U18036 ( .C1(n19939), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15909), .B(n14575), .ZN(n14576) );
  OAI211_X1 U18037 ( .C1(n20006), .C2(n14578), .A(n14577), .B(n14576), .ZN(
        P1_U2989) );
  INV_X1 U18038 ( .A(n14579), .ZN(n14581) );
  AOI21_X1 U18039 ( .B1(n14587), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14580) );
  NOR2_X1 U18040 ( .A1(n14581), .A2(n14580), .ZN(n14582) );
  INV_X1 U18041 ( .A(n14586), .ZN(n14592) );
  NAND2_X1 U18042 ( .A1(n14587), .A2(n9767), .ZN(n14588) );
  OAI211_X1 U18043 ( .C1(n14590), .C2(n19995), .A(n14589), .B(n14588), .ZN(
        n14591) );
  AOI21_X1 U18044 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14592), .A(
        n14591), .ZN(n14593) );
  OAI21_X1 U18045 ( .B1(n14594), .B2(n19996), .A(n14593), .ZN(P1_U3002) );
  XNOR2_X1 U18046 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14598) );
  NAND2_X1 U18047 ( .A1(n14595), .A2(n19979), .ZN(n14597) );
  OAI211_X1 U18048 ( .C1(n14603), .C2(n14598), .A(n14597), .B(n14596), .ZN(
        n14599) );
  AOI21_X1 U18049 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14607), .A(
        n14599), .ZN(n14600) );
  OAI21_X1 U18050 ( .B1(n14601), .B2(n19996), .A(n14600), .ZN(P1_U3003) );
  OAI21_X1 U18051 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14603), .A(
        n14602), .ZN(n14606) );
  NOR2_X1 U18052 ( .A1(n14604), .A2(n19995), .ZN(n14605) );
  AOI211_X1 U18053 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14607), .A(
        n14606), .B(n14605), .ZN(n14608) );
  OAI21_X1 U18054 ( .B1(n14609), .B2(n19996), .A(n14608), .ZN(P1_U3004) );
  INV_X1 U18055 ( .A(n14610), .ZN(n14626) );
  OR2_X1 U18056 ( .A1(n14612), .A2(n14611), .ZN(n14613) );
  NAND2_X1 U18057 ( .A1(n14614), .A2(n14613), .ZN(n15789) );
  OAI211_X1 U18058 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n14622), .B(n14615), .ZN(
        n14616) );
  OAI211_X1 U18059 ( .C1(n15789), .C2(n19995), .A(n14617), .B(n14616), .ZN(
        n14618) );
  AOI21_X1 U18060 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14626), .A(
        n14618), .ZN(n14619) );
  OAI21_X1 U18061 ( .B1(n14620), .B2(n19996), .A(n14619), .ZN(P1_U3005) );
  NAND2_X1 U18062 ( .A1(n14622), .A2(n14621), .ZN(n14623) );
  OAI211_X1 U18063 ( .C1(n15672), .C2(n19995), .A(n14624), .B(n14623), .ZN(
        n14625) );
  AOI21_X1 U18064 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14626), .A(
        n14625), .ZN(n14627) );
  OAI21_X1 U18065 ( .B1(n14628), .B2(n19996), .A(n14627), .ZN(P1_U3006) );
  NOR3_X1 U18066 ( .A1(n14638), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n14639), .ZN(n14629) );
  AOI211_X1 U18067 ( .C1(n15679), .C2(n19979), .A(n14630), .B(n14629), .ZN(
        n14634) );
  OAI21_X1 U18068 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n19970), .A(
        n14631), .ZN(n14632) );
  NAND2_X1 U18069 ( .A1(n14632), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14633) );
  OAI211_X1 U18070 ( .C1(n14635), .C2(n19996), .A(n14634), .B(n14633), .ZN(
        P1_U3007) );
  INV_X1 U18071 ( .A(n15689), .ZN(n14641) );
  NAND2_X1 U18072 ( .A1(n19977), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14636) );
  OAI221_X1 U18073 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14639), 
        .C1(n14638), .C2(n14637), .A(n14636), .ZN(n14640) );
  AOI21_X1 U18074 ( .B1(n14641), .B2(n19979), .A(n14640), .ZN(n14642) );
  OAI21_X1 U18075 ( .B1(n14643), .B2(n19996), .A(n14642), .ZN(P1_U3008) );
  INV_X1 U18076 ( .A(n14644), .ZN(n15874) );
  NAND2_X1 U18077 ( .A1(n15874), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14646) );
  OAI211_X1 U18078 ( .C1(n15709), .C2(n19995), .A(n14646), .B(n14645), .ZN(
        n14647) );
  AOI21_X1 U18079 ( .B1(n15878), .B2(n11611), .A(n14647), .ZN(n14648) );
  OAI21_X1 U18080 ( .B1(n14649), .B2(n19996), .A(n14648), .ZN(P1_U3010) );
  AOI21_X1 U18081 ( .B1(n14651), .B2(n9634), .A(n14650), .ZN(n14652) );
  XNOR2_X1 U18082 ( .A(n14652), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15820) );
  INV_X1 U18083 ( .A(n15820), .ZN(n14673) );
  NOR2_X1 U18084 ( .A1(n14654), .A2(n14653), .ZN(n14655) );
  OR2_X1 U18085 ( .A1(n14656), .A2(n14655), .ZN(n15793) );
  INV_X1 U18086 ( .A(n15793), .ZN(n14671) );
  INV_X1 U18087 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14663) );
  AND2_X1 U18088 ( .A1(n14663), .A2(n14657), .ZN(n14679) );
  NAND3_X1 U18089 ( .A1(n19991), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n14717), .ZN(n14659) );
  NAND2_X1 U18090 ( .A1(n14659), .A2(n14658), .ZN(n14683) );
  INV_X1 U18091 ( .A(n14660), .ZN(n14666) );
  OAI21_X1 U18092 ( .B1(n14663), .B2(n14662), .A(n14661), .ZN(n14665) );
  OAI211_X1 U18093 ( .C1(n14666), .C2(n19992), .A(n14665), .B(n14664), .ZN(
        n14674) );
  AOI21_X1 U18094 ( .B1(n14679), .B2(n14683), .A(n14674), .ZN(n14667) );
  NAND2_X1 U18095 ( .A1(n19977), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15821) );
  OAI221_X1 U18096 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14669), 
        .C1(n14668), .C2(n14667), .A(n15821), .ZN(n14670) );
  AOI21_X1 U18097 ( .B1(n14671), .B2(n19979), .A(n14670), .ZN(n14672) );
  OAI21_X1 U18098 ( .B1(n14673), .B2(n19996), .A(n14672), .ZN(P1_U3011) );
  NAND2_X1 U18099 ( .A1(n14674), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14676) );
  OAI211_X1 U18100 ( .C1(n14677), .C2(n19995), .A(n14676), .B(n14675), .ZN(
        n14678) );
  AOI21_X1 U18101 ( .B1(n14713), .B2(n14679), .A(n14678), .ZN(n14680) );
  OAI21_X1 U18102 ( .B1(n14681), .B2(n19996), .A(n14680), .ZN(P1_U3012) );
  NAND2_X1 U18103 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15896) );
  NAND3_X1 U18104 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n14713), .ZN(n15894) );
  INV_X1 U18105 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14682) );
  OAI21_X1 U18106 ( .B1(n15896), .B2(n15894), .A(n14682), .ZN(n14692) );
  INV_X1 U18107 ( .A(n15884), .ZN(n14689) );
  AND2_X1 U18108 ( .A1(n14711), .A2(n14683), .ZN(n14720) );
  NAND2_X1 U18109 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14717), .ZN(
        n14684) );
  AND2_X1 U18110 ( .A1(n20001), .A2(n14684), .ZN(n14716) );
  NAND2_X1 U18111 ( .A1(n19991), .A2(n14685), .ZN(n14686) );
  OAI21_X1 U18112 ( .B1(n14687), .B2(n19992), .A(n14686), .ZN(n14688) );
  OR3_X1 U18113 ( .A1(n19981), .A2(n14716), .A3(n14688), .ZN(n14722) );
  OR2_X1 U18114 ( .A1(n14720), .A2(n14722), .ZN(n14710) );
  AOI21_X1 U18115 ( .B1(n14704), .B2(n19986), .A(n14710), .ZN(n15902) );
  OAI21_X1 U18116 ( .B1(n15922), .B2(n14689), .A(n15902), .ZN(n15890) );
  OAI21_X1 U18117 ( .B1(n15734), .B2(n19995), .A(n14690), .ZN(n14691) );
  AOI21_X1 U18118 ( .B1(n14692), .B2(n15890), .A(n14691), .ZN(n14693) );
  OAI21_X1 U18119 ( .B1(n14694), .B2(n19996), .A(n14693), .ZN(P1_U3014) );
  INV_X1 U18120 ( .A(n15758), .ZN(n14697) );
  NAND2_X1 U18121 ( .A1(n19977), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14695) );
  OAI221_X1 U18122 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15894), 
        .C1(n15895), .C2(n15902), .A(n14695), .ZN(n14696) );
  AOI21_X1 U18123 ( .B1(n14697), .B2(n19979), .A(n14696), .ZN(n14698) );
  OAI21_X1 U18124 ( .B1(n14699), .B2(n19996), .A(n14698), .ZN(P1_U3016) );
  INV_X1 U18125 ( .A(n14700), .ZN(n14701) );
  AOI21_X1 U18126 ( .B1(n14703), .B2(n14702), .A(n14701), .ZN(n14707) );
  XNOR2_X1 U18127 ( .A(n14705), .B(n14704), .ZN(n14706) );
  XNOR2_X1 U18128 ( .A(n14707), .B(n14706), .ZN(n15846) );
  INV_X1 U18129 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14708) );
  OAI22_X1 U18130 ( .A1(n15759), .A2(n19995), .B1(n19964), .B2(n14708), .ZN(
        n14709) );
  AOI21_X1 U18131 ( .B1(n14710), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n14709), .ZN(n14715) );
  NOR2_X1 U18132 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14711), .ZN(
        n14712) );
  NAND2_X1 U18133 ( .A1(n14713), .A2(n14712), .ZN(n14714) );
  OAI211_X1 U18134 ( .C1(n15846), .C2(n19996), .A(n14715), .B(n14714), .ZN(
        P1_U3017) );
  AOI22_X1 U18135 ( .A1(n19977), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n14717), 
        .B2(n14716), .ZN(n14718) );
  OAI21_X1 U18136 ( .B1(n14719), .B2(n19995), .A(n14718), .ZN(n14721) );
  AOI211_X1 U18137 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n14722), .A(
        n14721), .B(n14720), .ZN(n14723) );
  OAI21_X1 U18138 ( .B1(n14724), .B2(n19996), .A(n14723), .ZN(P1_U3018) );
  INV_X1 U18139 ( .A(n14725), .ZN(n14726) );
  AOI21_X1 U18140 ( .B1(n14728), .B2(n14727), .A(n14726), .ZN(n15852) );
  NAND3_X1 U18141 ( .A1(n14729), .A2(n15937), .A3(n20856), .ZN(n14741) );
  INV_X1 U18142 ( .A(n14735), .ZN(n14731) );
  AOI21_X1 U18143 ( .B1(n14732), .B2(n14731), .A(n14730), .ZN(n14733) );
  AOI211_X1 U18144 ( .C1(n19968), .C2(n14734), .A(n14733), .B(n19981), .ZN(
        n15908) );
  NOR2_X1 U18145 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14735), .ZN(
        n15904) );
  NAND2_X1 U18146 ( .A1(n15904), .A2(n14736), .ZN(n14737) );
  AOI21_X1 U18147 ( .B1(n15908), .B2(n14737), .A(n20856), .ZN(n14739) );
  OAI22_X1 U18148 ( .A1(n15774), .A2(n19995), .B1(n20619), .B2(n19964), .ZN(
        n14738) );
  NOR2_X1 U18149 ( .A1(n14739), .A2(n14738), .ZN(n14740) );
  OAI211_X1 U18150 ( .C1(n15852), .C2(n19996), .A(n14741), .B(n14740), .ZN(
        P1_U3019) );
  INV_X1 U18151 ( .A(n13829), .ZN(n20687) );
  NOR3_X1 U18152 ( .A1(n14742), .A2(n13475), .A3(n11191), .ZN(n14743) );
  AOI211_X1 U18153 ( .C1(n20687), .C2(n14745), .A(n14744), .B(n14743), .ZN(
        n15580) );
  INV_X1 U18154 ( .A(n15945), .ZN(n14758) );
  AOI22_X1 U18155 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19987), .B2(n12737), .ZN(
        n14756) );
  INV_X1 U18156 ( .A(n14756), .ZN(n14747) );
  NOR2_X1 U18157 ( .A1(n13792), .A2(n20798), .ZN(n14755) );
  NOR3_X1 U18158 ( .A1(n11191), .A2(n13475), .A3(n15599), .ZN(n14746) );
  AOI21_X1 U18159 ( .B1(n14747), .B2(n14755), .A(n14746), .ZN(n14748) );
  OAI21_X1 U18160 ( .B1(n15580), .B2(n14758), .A(n14748), .ZN(n14750) );
  INV_X1 U18161 ( .A(n14749), .ZN(n15948) );
  MUX2_X1 U18162 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14750), .S(
        n15948), .Z(P1_U3473) );
  INV_X1 U18163 ( .A(n14751), .ZN(n14759) );
  INV_X1 U18164 ( .A(n14752), .ZN(n14754) );
  AOI22_X1 U18165 ( .A1(n14756), .A2(n14755), .B1(n14754), .B2(n14753), .ZN(
        n14757) );
  OAI21_X1 U18166 ( .B1(n14759), .B2(n14758), .A(n14757), .ZN(n14760) );
  MUX2_X1 U18167 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14760), .S(
        n15948), .Z(P1_U3472) );
  OR2_X1 U18168 ( .A1(n14762), .A2(n14761), .ZN(n14763) );
  NAND2_X1 U18169 ( .A1(n14764), .A2(n14763), .ZN(n15136) );
  OAI21_X1 U18170 ( .B1(n14894), .B2(n14766), .A(n14765), .ZN(n15133) );
  AOI22_X1 U18171 ( .A1(n14767), .A2(n18865), .B1(P2_REIP_REG_29__SCAN_IN), 
        .B2(n18867), .ZN(n14769) );
  AOI22_X1 U18172 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n18866), .ZN(n14768) );
  OAI211_X1 U18173 ( .C1(n15133), .C2(n18836), .A(n14769), .B(n14768), .ZN(
        n14772) );
  NOR2_X1 U18174 ( .A1(n14772), .A2(n14771), .ZN(n14773) );
  OAI21_X1 U18175 ( .B1(n15136), .B2(n18870), .A(n14773), .ZN(P2_U2826) );
  INV_X1 U18176 ( .A(n12480), .ZN(n14774) );
  AOI21_X1 U18177 ( .B1(n14775), .B2(n14850), .A(n14774), .ZN(n15153) );
  INV_X1 U18178 ( .A(n15153), .ZN(n14786) );
  OAI21_X1 U18179 ( .B1(n14911), .B2(n14776), .A(n14893), .ZN(n15159) );
  INV_X1 U18180 ( .A(n14777), .ZN(n14778) );
  AOI22_X1 U18181 ( .A1(n14778), .A2(n18865), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18874), .ZN(n14780) );
  AOI22_X1 U18182 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n18867), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n18866), .ZN(n14779) );
  OAI211_X1 U18183 ( .C1(n15159), .C2(n18836), .A(n14780), .B(n14779), .ZN(
        n14784) );
  AOI211_X1 U18184 ( .C1(n15004), .C2(n14782), .A(n14781), .B(n18877), .ZN(
        n14783) );
  NOR2_X1 U18185 ( .A1(n14784), .A2(n14783), .ZN(n14785) );
  OAI21_X1 U18186 ( .B1(n14786), .B2(n18870), .A(n14785), .ZN(P2_U2828) );
  AND2_X1 U18187 ( .A1(n14861), .A2(n14787), .ZN(n14788) );
  OR2_X1 U18188 ( .A1(n14788), .A2(n14848), .ZN(n16036) );
  INV_X1 U18189 ( .A(n14789), .ZN(n14790) );
  OAI21_X1 U18190 ( .B1(n14930), .B2(n14791), .A(n14790), .ZN(n15183) );
  OAI22_X1 U18191 ( .A1(n14793), .A2(n18852), .B1(n14792), .B2(n18774), .ZN(
        n14794) );
  INV_X1 U18192 ( .A(n14794), .ZN(n14796) );
  AOI22_X1 U18193 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n18866), .ZN(n14795) );
  OAI211_X1 U18194 ( .C1(n15183), .C2(n18836), .A(n14796), .B(n14795), .ZN(
        n14800) );
  AOI211_X1 U18195 ( .C1(n16031), .C2(n14798), .A(n14797), .B(n18877), .ZN(
        n14799) );
  NOR2_X1 U18196 ( .A1(n14800), .A2(n14799), .ZN(n14801) );
  OAI21_X1 U18197 ( .B1(n16036), .B2(n18870), .A(n14801), .ZN(P2_U2830) );
  AOI211_X1 U18198 ( .C1(n14804), .C2(n14803), .A(n14802), .B(n18877), .ZN(
        n14806) );
  INV_X1 U18199 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16009) );
  INV_X1 U18200 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19663) );
  OAI22_X1 U18201 ( .A1(n18837), .A2(n16009), .B1(n19663), .B2(n18774), .ZN(
        n14805) );
  AOI211_X1 U18202 ( .C1(n18874), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14806), .B(n14805), .ZN(n14813) );
  XOR2_X1 U18203 ( .A(n14807), .B(n14808), .Z(n15217) );
  INV_X1 U18204 ( .A(n14809), .ZN(n14810) );
  OAI21_X1 U18205 ( .B1(n14811), .B2(n9859), .A(n14810), .ZN(n15222) );
  INV_X1 U18206 ( .A(n15222), .ZN(n16006) );
  AOI22_X1 U18207 ( .A1(n15217), .A2(n18863), .B1(n16006), .B2(n18840), .ZN(
        n14812) );
  OAI211_X1 U18208 ( .C1(n14814), .C2(n18852), .A(n14813), .B(n14812), .ZN(
        P2_U2833) );
  INV_X1 U18209 ( .A(n14815), .ZN(n14829) );
  OAI21_X1 U18210 ( .B1(n14818), .B2(n14816), .A(n14817), .ZN(n16046) );
  OAI21_X1 U18211 ( .B1(n14819), .B2(n15634), .A(n14807), .ZN(n15236) );
  INV_X1 U18212 ( .A(n15236), .ZN(n14820) );
  AOI22_X1 U18213 ( .A1(n18866), .A2(P2_EBX_REG_21__SCAN_IN), .B1(n18863), 
        .B2(n14820), .ZN(n14821) );
  OAI21_X1 U18214 ( .B1(n16046), .B2(n18870), .A(n14821), .ZN(n14828) );
  NAND3_X1 U18215 ( .A1(n18827), .A2(n13945), .A3(n14822), .ZN(n18665) );
  NAND2_X1 U18216 ( .A1(n18827), .A2(n14823), .ZN(n14825) );
  AOI22_X1 U18217 ( .A1(P2_REIP_REG_21__SCAN_IN), .A2(n18867), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18874), .ZN(n14824) );
  OAI221_X1 U18218 ( .B1(n16040), .B2(n18665), .C1(n14826), .C2(n14825), .A(
        n14824), .ZN(n14827) );
  AOI211_X1 U18219 ( .C1(n18865), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        n14830) );
  INV_X1 U18220 ( .A(n14830), .ZN(P2_U2834) );
  OR2_X1 U18221 ( .A1(n14832), .A2(n14831), .ZN(n14883) );
  NAND3_X1 U18222 ( .A1(n14883), .A2(n14833), .A3(n18899), .ZN(n14835) );
  NAND2_X1 U18223 ( .A1(n18888), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14834) );
  OAI211_X1 U18224 ( .C1(n18888), .C2(n15136), .A(n14835), .B(n14834), .ZN(
        P2_U2858) );
  NAND2_X1 U18225 ( .A1(n14837), .A2(n14836), .ZN(n14838) );
  XOR2_X1 U18226 ( .A(n14839), .B(n14838), .Z(n14900) );
  NOR2_X1 U18227 ( .A1(n18888), .A2(n15966), .ZN(n14840) );
  AOI21_X1 U18228 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n18888), .A(n14840), .ZN(
        n14841) );
  OAI21_X1 U18229 ( .B1(n14900), .B2(n18893), .A(n14841), .ZN(P2_U2859) );
  OAI21_X1 U18230 ( .B1(n14842), .B2(n14844), .A(n14843), .ZN(n14907) );
  NAND2_X1 U18231 ( .A1(n18888), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14846) );
  NAND2_X1 U18232 ( .A1(n15153), .A2(n18903), .ZN(n14845) );
  OAI211_X1 U18233 ( .C1(n14907), .C2(n18893), .A(n14846), .B(n14845), .ZN(
        P2_U2860) );
  OR2_X1 U18234 ( .A1(n14848), .A2(n14847), .ZN(n14849) );
  NAND2_X1 U18235 ( .A1(n14850), .A2(n14849), .ZN(n15980) );
  AOI21_X1 U18236 ( .B1(n14853), .B2(n14852), .A(n14851), .ZN(n14908) );
  NAND2_X1 U18237 ( .A1(n14908), .A2(n18899), .ZN(n14855) );
  NAND2_X1 U18238 ( .A1(n18888), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14854) );
  OAI211_X1 U18239 ( .C1(n15980), .C2(n18888), .A(n14855), .B(n14854), .ZN(
        P2_U2861) );
  AOI21_X1 U18240 ( .B1(n9702), .B2(n14857), .A(n14856), .ZN(n14928) );
  NAND2_X1 U18241 ( .A1(n14928), .A2(n18899), .ZN(n14864) );
  INV_X1 U18242 ( .A(n14858), .ZN(n14860) );
  NAND2_X1 U18243 ( .A1(n14860), .A2(n14859), .ZN(n14862) );
  AND2_X1 U18244 ( .A1(n14862), .A2(n14861), .ZN(n15991) );
  NAND2_X1 U18245 ( .A1(n18903), .A2(n15991), .ZN(n14863) );
  OAI211_X1 U18246 ( .C1(n18903), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        P2_U2863) );
  AOI21_X1 U18247 ( .B1(n14868), .B2(n14867), .A(n14866), .ZN(n14938) );
  NAND2_X1 U18248 ( .A1(n14938), .A2(n18899), .ZN(n14871) );
  INV_X1 U18249 ( .A(n15208), .ZN(n14869) );
  NAND2_X1 U18250 ( .A1(n18903), .A2(n14869), .ZN(n14870) );
  OAI211_X1 U18251 ( .C1(n18903), .C2(n11161), .A(n14871), .B(n14870), .ZN(
        P2_U2864) );
  OAI21_X1 U18252 ( .B1(n14872), .B2(n14874), .A(n14873), .ZN(n14958) );
  OR2_X1 U18253 ( .A1(n14958), .A2(n18893), .ZN(n14876) );
  INV_X1 U18254 ( .A(n16046), .ZN(n15234) );
  NAND2_X1 U18255 ( .A1(n18903), .A2(n15234), .ZN(n14875) );
  OAI211_X1 U18256 ( .C1(n18903), .C2(n9950), .A(n14876), .B(n14875), .ZN(
        P2_U2866) );
  OAI21_X1 U18257 ( .B1(n14877), .B2(n15279), .A(n15060), .ZN(n18684) );
  AOI21_X1 U18258 ( .B1(n14880), .B2(n14878), .A(n14879), .ZN(n14959) );
  NAND2_X1 U18259 ( .A1(n14959), .A2(n18899), .ZN(n14882) );
  NAND2_X1 U18260 ( .A1(n18888), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14881) );
  OAI211_X1 U18261 ( .C1(n18684), .C2(n18888), .A(n14882), .B(n14881), .ZN(
        P2_U2868) );
  NAND3_X1 U18262 ( .A1(n14883), .A2(n14833), .A3(n16024), .ZN(n14889) );
  NOR2_X1 U18263 ( .A1(n16017), .A2(n14884), .ZN(n14887) );
  OAI22_X1 U18264 ( .A1(n16018), .A2(n15133), .B1(n18926), .B2(n14885), .ZN(
        n14886) );
  AOI211_X1 U18265 ( .C1(BUF2_REG_29__SCAN_IN), .C2(n18908), .A(n14887), .B(
        n14886), .ZN(n14888) );
  OAI211_X1 U18266 ( .C1(n14918), .C2(n14890), .A(n14889), .B(n14888), .ZN(
        P2_U2890) );
  OAI22_X1 U18267 ( .A1(n16017), .A2(n14891), .B1(n18926), .B2(n20796), .ZN(
        n14897) );
  AND2_X1 U18268 ( .A1(n14893), .A2(n14892), .ZN(n14895) );
  OR2_X1 U18269 ( .A1(n14895), .A2(n14894), .ZN(n15965) );
  NOR2_X1 U18270 ( .A1(n16018), .A2(n15965), .ZN(n14896) );
  AOI211_X1 U18271 ( .C1(BUF1_REG_28__SCAN_IN), .C2(n18909), .A(n14897), .B(
        n14896), .ZN(n14899) );
  NAND2_X1 U18272 ( .A1(n18908), .A2(BUF2_REG_28__SCAN_IN), .ZN(n14898) );
  OAI211_X1 U18273 ( .C1(n14900), .C2(n18930), .A(n14899), .B(n14898), .ZN(
        P2_U2891) );
  NOR2_X1 U18274 ( .A1(n16017), .A2(n14901), .ZN(n14904) );
  OAI22_X1 U18275 ( .A1(n16018), .A2(n15159), .B1(n18926), .B2(n14902), .ZN(
        n14903) );
  AOI211_X1 U18276 ( .C1(BUF2_REG_27__SCAN_IN), .C2(n18908), .A(n14904), .B(
        n14903), .ZN(n14906) );
  NAND2_X1 U18277 ( .A1(n18909), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14905) );
  OAI211_X1 U18278 ( .C1(n14907), .C2(n18930), .A(n14906), .B(n14905), .ZN(
        P2_U2892) );
  INV_X1 U18279 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n14917) );
  NAND2_X1 U18280 ( .A1(n14908), .A2(n16024), .ZN(n14916) );
  NOR2_X1 U18281 ( .A1(n14789), .A2(n14909), .ZN(n14910) );
  NOR2_X1 U18282 ( .A1(n14911), .A2(n14910), .ZN(n15978) );
  AOI22_X1 U18283 ( .A1(n18912), .A2(n15978), .B1(n18921), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n14912) );
  OAI21_X1 U18284 ( .B1(n14913), .B2(n16017), .A(n14912), .ZN(n14914) );
  AOI21_X1 U18285 ( .B1(n18908), .B2(BUF2_REG_26__SCAN_IN), .A(n14914), .ZN(
        n14915) );
  OAI211_X1 U18286 ( .C1(n14918), .C2(n14917), .A(n14916), .B(n14915), .ZN(
        P2_U2893) );
  OAI21_X1 U18287 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n16003) );
  OAI22_X1 U18288 ( .A1(n16017), .A2(n14923), .B1(n18926), .B2(n14922), .ZN(
        n14925) );
  NOR2_X1 U18289 ( .A1(n16018), .A2(n15183), .ZN(n14924) );
  AOI211_X1 U18290 ( .C1(BUF1_REG_25__SCAN_IN), .C2(n18909), .A(n14925), .B(
        n14924), .ZN(n14927) );
  NAND2_X1 U18291 ( .A1(n18908), .A2(BUF2_REG_25__SCAN_IN), .ZN(n14926) );
  OAI211_X1 U18292 ( .C1(n16003), .C2(n18930), .A(n14927), .B(n14926), .ZN(
        P2_U2894) );
  INV_X1 U18293 ( .A(n18908), .ZN(n14968) );
  INV_X1 U18294 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n14937) );
  NAND2_X1 U18295 ( .A1(n14928), .A2(n16024), .ZN(n14936) );
  OAI22_X1 U18296 ( .A1(n16017), .A2(n14929), .B1(n18926), .B2(n11128), .ZN(
        n14934) );
  INV_X1 U18297 ( .A(n14930), .ZN(n14931) );
  OAI21_X1 U18298 ( .B1(n14932), .B2(n13214), .A(n14931), .ZN(n15989) );
  NOR2_X1 U18299 ( .A1(n16018), .A2(n15989), .ZN(n14933) );
  AOI211_X1 U18300 ( .C1(BUF1_REG_24__SCAN_IN), .C2(n18909), .A(n14934), .B(
        n14933), .ZN(n14935) );
  OAI211_X1 U18301 ( .C1(n14968), .C2(n14937), .A(n14936), .B(n14935), .ZN(
        P2_U2895) );
  INV_X1 U18302 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n14944) );
  NAND2_X1 U18303 ( .A1(n14938), .A2(n16024), .ZN(n14943) );
  OAI22_X1 U18304 ( .A1(n16017), .A2(n14939), .B1(n18926), .B2(n11126), .ZN(
        n14941) );
  NOR2_X1 U18305 ( .A1(n16018), .A2(n15204), .ZN(n14940) );
  AOI211_X1 U18306 ( .C1(BUF1_REG_23__SCAN_IN), .C2(n18909), .A(n14941), .B(
        n14940), .ZN(n14942) );
  OAI211_X1 U18307 ( .C1(n14968), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        P2_U2896) );
  INV_X1 U18308 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n14953) );
  AOI21_X1 U18309 ( .B1(n14945), .B2(n14873), .A(n13020), .ZN(n16007) );
  NAND2_X1 U18310 ( .A1(n16007), .A2(n16024), .ZN(n14952) );
  OAI22_X1 U18311 ( .A1(n16017), .A2(n14947), .B1(n18926), .B2(n14946), .ZN(
        n14950) );
  INV_X1 U18312 ( .A(n15217), .ZN(n14948) );
  NOR2_X1 U18313 ( .A1(n16018), .A2(n14948), .ZN(n14949) );
  AOI211_X1 U18314 ( .C1(BUF1_REG_22__SCAN_IN), .C2(n18909), .A(n14950), .B(
        n14949), .ZN(n14951) );
  OAI211_X1 U18315 ( .C1(n14968), .C2(n14953), .A(n14952), .B(n14951), .ZN(
        P2_U2897) );
  OAI22_X1 U18316 ( .A1(n16017), .A2(n18927), .B1(n18926), .B2(n20852), .ZN(
        n14955) );
  NOR2_X1 U18317 ( .A1(n16018), .A2(n15236), .ZN(n14954) );
  AOI211_X1 U18318 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n18909), .A(n14955), .B(
        n14954), .ZN(n14957) );
  NAND2_X1 U18319 ( .A1(n18908), .A2(BUF2_REG_21__SCAN_IN), .ZN(n14956) );
  OAI211_X1 U18320 ( .C1(n14958), .C2(n18930), .A(n14957), .B(n14956), .ZN(
        P2_U2898) );
  INV_X1 U18321 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14967) );
  NAND2_X1 U18322 ( .A1(n14959), .A2(n16024), .ZN(n14966) );
  OAI22_X1 U18323 ( .A1(n16017), .A2(n14961), .B1(n18926), .B2(n14960), .ZN(
        n14964) );
  OAI21_X1 U18324 ( .B1(n14962), .B2(n15271), .A(n15632), .ZN(n18683) );
  NOR2_X1 U18325 ( .A1(n16018), .A2(n18683), .ZN(n14963) );
  AOI211_X1 U18326 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n18909), .A(n14964), .B(
        n14963), .ZN(n14965) );
  OAI211_X1 U18327 ( .C1(n14968), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        P2_U2900) );
  OAI21_X1 U18328 ( .B1(n14969), .B2(n14971), .A(n14970), .ZN(n18707) );
  OAI22_X1 U18329 ( .A1(n16017), .A2(n14973), .B1(n18926), .B2(n14972), .ZN(
        n14974) );
  AOI21_X1 U18330 ( .B1(n18909), .B2(BUF1_REG_17__SCAN_IN), .A(n14974), .ZN(
        n14976) );
  NAND2_X1 U18331 ( .A1(n18908), .A2(BUF2_REG_17__SCAN_IN), .ZN(n14975) );
  OAI211_X1 U18332 ( .C1(n18707), .C2(n16018), .A(n14976), .B(n14975), .ZN(
        n14977) );
  INV_X1 U18333 ( .A(n14977), .ZN(n14978) );
  OAI21_X1 U18334 ( .B1(n18930), .B2(n14979), .A(n14978), .ZN(P2_U2902) );
  INV_X1 U18335 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14981) );
  OAI21_X1 U18336 ( .B1(n16117), .B2(n14981), .A(n14980), .ZN(n14982) );
  OAI21_X1 U18337 ( .B1(n14987), .B2(n18981), .A(n14986), .ZN(P2_U2984) );
  NAND2_X1 U18338 ( .A1(n14989), .A2(n14988), .ZN(n14991) );
  XOR2_X1 U18339 ( .A(n14991), .B(n14990), .Z(n15141) );
  AOI21_X1 U18340 ( .B1(n15128), .B2(n12552), .A(n14992), .ZN(n15139) );
  NAND2_X1 U18341 ( .A1(n14993), .A2(n16108), .ZN(n14995) );
  NOR2_X1 U18342 ( .A1(n18772), .A2(n19673), .ZN(n15129) );
  AOI21_X1 U18343 ( .B1(n18977), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15129), .ZN(n14994) );
  OAI211_X1 U18344 ( .C1(n15136), .C2(n19026), .A(n14995), .B(n14994), .ZN(
        n14996) );
  AOI21_X1 U18345 ( .B1(n15139), .B2(n16113), .A(n14996), .ZN(n14997) );
  OAI21_X1 U18346 ( .B1(n15141), .B2(n18981), .A(n14997), .ZN(P2_U2985) );
  NAND2_X1 U18347 ( .A1(n14998), .A2(n20763), .ZN(n15152) );
  NAND2_X1 U18348 ( .A1(n15152), .A2(n16112), .ZN(n15006) );
  NAND2_X1 U18349 ( .A1(n15153), .A2(n18985), .ZN(n14999) );
  NAND2_X1 U18350 ( .A1(n18822), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15154) );
  OAI211_X1 U18351 ( .C1(n16117), .C2(n15000), .A(n14999), .B(n15154), .ZN(
        n15003) );
  NOR3_X1 U18352 ( .A1(n15160), .A2(n12479), .A3(n18980), .ZN(n15002) );
  OAI21_X1 U18353 ( .B1(n15165), .B2(n15006), .A(n15005), .ZN(P2_U2987) );
  NAND2_X1 U18354 ( .A1(n15007), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15027) );
  NAND2_X1 U18355 ( .A1(n15027), .A2(n15008), .ZN(n15022) );
  OR2_X1 U18356 ( .A1(n15007), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15024) );
  NAND2_X1 U18357 ( .A1(n15022), .A2(n15024), .ZN(n15178) );
  INV_X1 U18358 ( .A(n15177), .ZN(n15009) );
  OAI21_X1 U18359 ( .B1(n15178), .B2(n15009), .A(n15011), .ZN(n15010) );
  MUX2_X1 U18360 ( .A(n15011), .B(n15010), .S(n15176), .Z(n15012) );
  NAND2_X1 U18361 ( .A1(n15012), .A2(n12534), .ZN(n15175) );
  NAND2_X1 U18362 ( .A1(n15014), .A2(n15166), .ZN(n15015) );
  AND2_X1 U18363 ( .A1(n15001), .A2(n15015), .ZN(n15173) );
  NOR2_X1 U18364 ( .A1(n18772), .A2(n15016), .ZN(n15167) );
  NOR2_X1 U18365 ( .A1(n19026), .A2(n15980), .ZN(n15017) );
  AOI211_X1 U18366 ( .C1(n18977), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15167), .B(n15017), .ZN(n15018) );
  OAI21_X1 U18367 ( .B1(n15019), .B2(n18989), .A(n15018), .ZN(n15020) );
  AOI21_X1 U18368 ( .B1(n15173), .B2(n16113), .A(n15020), .ZN(n15021) );
  OAI21_X1 U18369 ( .B1(n15175), .B2(n18981), .A(n15021), .ZN(P2_U2988) );
  INV_X1 U18370 ( .A(n15178), .ZN(n15028) );
  INV_X1 U18371 ( .A(n15022), .ZN(n15025) );
  AOI21_X1 U18372 ( .B1(n15025), .B2(n15024), .A(n15023), .ZN(n15026) );
  AOI21_X1 U18373 ( .B1(n15028), .B2(n15027), .A(n15026), .ZN(n15192) );
  NAND2_X1 U18374 ( .A1(n15192), .A2(n16112), .ZN(n15036) );
  AOI22_X1 U18375 ( .A1(n18985), .A2(n15991), .B1(n18977), .B2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15035) );
  AND2_X1 U18376 ( .A1(n15038), .A2(n15195), .ZN(n15030) );
  NOR2_X1 U18377 ( .A1(n15029), .A2(n15030), .ZN(n15200) );
  NAND2_X1 U18378 ( .A1(n15200), .A2(n16113), .ZN(n15034) );
  OAI22_X1 U18379 ( .A1(n11127), .A2(n18772), .B1(n18989), .B2(n15031), .ZN(
        n15032) );
  INV_X1 U18380 ( .A(n15032), .ZN(n15033) );
  NAND4_X1 U18381 ( .A1(n15036), .A2(n15035), .A3(n15034), .A4(n15033), .ZN(
        P2_U2990) );
  NOR2_X1 U18382 ( .A1(n15037), .A2(n15218), .ZN(n15051) );
  OAI21_X1 U18383 ( .B1(n15051), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15038), .ZN(n15214) );
  NOR2_X1 U18384 ( .A1(n19026), .A2(n15208), .ZN(n15041) );
  OAI22_X1 U18385 ( .A1(n15039), .A2(n16117), .B1(n11125), .B2(n18772), .ZN(
        n15040) );
  AOI211_X1 U18386 ( .C1(n15042), .C2(n16108), .A(n15041), .B(n15040), .ZN(
        n15046) );
  XOR2_X1 U18387 ( .A(n15043), .B(n15044), .Z(n15211) );
  NAND2_X1 U18388 ( .A1(n15211), .A2(n16112), .ZN(n15045) );
  OAI211_X1 U18389 ( .C1(n15214), .C2(n18980), .A(n15046), .B(n15045), .ZN(
        P2_U2991) );
  NAND2_X1 U18390 ( .A1(n15048), .A2(n15047), .ZN(n15050) );
  XOR2_X1 U18391 ( .A(n15050), .B(n9612), .Z(n15226) );
  INV_X1 U18392 ( .A(n15051), .ZN(n15216) );
  NAND2_X1 U18393 ( .A1(n15037), .A2(n15218), .ZN(n15215) );
  NAND3_X1 U18394 ( .A1(n15216), .A2(n16113), .A3(n15215), .ZN(n15056) );
  NOR2_X1 U18395 ( .A1(n19026), .A2(n15222), .ZN(n15054) );
  OAI22_X1 U18396 ( .A1(n19663), .A2(n19017), .B1(n18989), .B2(n15052), .ZN(
        n15053) );
  AOI211_X1 U18397 ( .C1(n18977), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15054), .B(n15053), .ZN(n15055) );
  OAI211_X1 U18398 ( .C1(n15226), .C2(n18981), .A(n15056), .B(n15055), .ZN(
        P2_U2992) );
  OAI21_X1 U18399 ( .B1(n15057), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15058), .ZN(n15639) );
  INV_X1 U18400 ( .A(n15059), .ZN(n18669) );
  NAND2_X1 U18401 ( .A1(n15061), .A2(n15060), .ZN(n15063) );
  INV_X1 U18402 ( .A(n14816), .ZN(n15062) );
  NAND2_X1 U18403 ( .A1(n15063), .A2(n15062), .ZN(n18671) );
  NAND2_X1 U18404 ( .A1(n18822), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15645) );
  NAND2_X1 U18405 ( .A1(n18977), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15064) );
  OAI211_X1 U18406 ( .C1(n19026), .C2(n18671), .A(n15645), .B(n15064), .ZN(
        n15080) );
  INV_X1 U18407 ( .A(n15230), .ZN(n15074) );
  INV_X1 U18408 ( .A(n15065), .ZN(n15070) );
  AOI21_X2 U18409 ( .B1(n15070), .B2(n15069), .A(n15319), .ZN(n15098) );
  OAI21_X1 U18410 ( .B1(n15075), .B2(n15074), .A(n15076), .ZN(n15078) );
  NAND2_X1 U18411 ( .A1(n15078), .A2(n15229), .ZN(n15640) );
  NOR2_X1 U18412 ( .A1(n15640), .A2(n18981), .ZN(n15079) );
  OAI21_X1 U18413 ( .B1(n15639), .B2(n18980), .A(n15081), .ZN(P2_U2994) );
  INV_X1 U18414 ( .A(n18702), .ZN(n15096) );
  BUF_X1 U18415 ( .A(n15082), .Z(n15083) );
  AND2_X1 U18416 ( .A1(n15314), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15084) );
  NAND2_X1 U18417 ( .A1(n15358), .A2(n15084), .ZN(n15316) );
  OAI211_X1 U18418 ( .C1(n15291), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16113), .B(n15263), .ZN(n15095) );
  INV_X1 U18419 ( .A(n15097), .ZN(n15086) );
  NOR2_X1 U18420 ( .A1(n15087), .A2(n15086), .ZN(n15091) );
  NOR2_X1 U18421 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  XNOR2_X1 U18422 ( .A(n15091), .B(n15090), .ZN(n15297) );
  NAND2_X1 U18423 ( .A1(n18822), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15294) );
  OAI21_X1 U18424 ( .B1(n16117), .B2(n18703), .A(n15294), .ZN(n15093) );
  NOR2_X1 U18425 ( .A1(n19026), .A2(n18708), .ZN(n15092) );
  AOI211_X1 U18426 ( .C1(n16112), .C2(n15297), .A(n15093), .B(n15092), .ZN(
        n15094) );
  OAI211_X1 U18427 ( .C1(n18989), .C2(n15096), .A(n15095), .B(n15094), .ZN(
        P2_U2997) );
  OAI21_X1 U18428 ( .B1(n15099), .B2(n15098), .A(n15097), .ZN(n15307) );
  INV_X1 U18429 ( .A(n15316), .ZN(n15301) );
  OAI211_X1 U18430 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15301), .A(
        n9742), .B(n16113), .ZN(n15106) );
  INV_X1 U18431 ( .A(n18715), .ZN(n15104) );
  OAI21_X1 U18432 ( .B1(n13926), .B2(n15101), .A(n15100), .ZN(n18880) );
  NAND2_X1 U18433 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18977), .ZN(
        n15102) );
  NAND2_X1 U18434 ( .A1(n18822), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15308) );
  OAI211_X1 U18435 ( .C1(n19026), .C2(n18880), .A(n15102), .B(n15308), .ZN(
        n15103) );
  AOI21_X1 U18436 ( .B1(n16108), .B2(n15104), .A(n15103), .ZN(n15105) );
  OAI211_X1 U18437 ( .C1(n15307), .C2(n18981), .A(n15106), .B(n15105), .ZN(
        P2_U2998) );
  XOR2_X1 U18438 ( .A(n9839), .B(n15108), .Z(n15109) );
  XNOR2_X1 U18439 ( .A(n15107), .B(n15109), .ZN(n16143) );
  NAND2_X1 U18440 ( .A1(n12320), .A2(n15111), .ZN(n15112) );
  XNOR2_X1 U18441 ( .A(n14169), .B(n15112), .ZN(n16141) );
  OAI22_X1 U18442 ( .A1(n15113), .A2(n16117), .B1(n19643), .B2(n18772), .ZN(
        n15117) );
  INV_X1 U18443 ( .A(n15114), .ZN(n15115) );
  OAI22_X1 U18444 ( .A1(n18989), .A2(n15115), .B1(n19026), .B2(n16136), .ZN(
        n15116) );
  AOI211_X1 U18445 ( .C1(n16141), .C2(n16112), .A(n15117), .B(n15116), .ZN(
        n15118) );
  OAI21_X1 U18446 ( .B1(n18980), .B2(n16143), .A(n15118), .ZN(P2_U3007) );
  XNOR2_X1 U18447 ( .A(n15119), .B(n15120), .ZN(n15428) );
  OAI21_X1 U18448 ( .B1(n15122), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15121), .ZN(n15123) );
  INV_X1 U18449 ( .A(n15123), .ZN(n15420) );
  OAI22_X1 U18450 ( .A1(n19641), .A2(n19017), .B1(n18989), .B2(n18812), .ZN(
        n15126) );
  OAI22_X1 U18451 ( .A1(n19026), .A2(n15124), .B1(n16117), .B2(n9823), .ZN(
        n15125) );
  AOI211_X1 U18452 ( .C1(n15420), .C2(n16113), .A(n15126), .B(n15125), .ZN(
        n15127) );
  OAI21_X1 U18453 ( .B1(n18981), .B2(n15428), .A(n15127), .ZN(P2_U3008) );
  INV_X1 U18454 ( .A(n15131), .ZN(n15156) );
  NAND2_X1 U18455 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15130) );
  AOI21_X1 U18456 ( .B1(n15156), .B2(n15130), .A(n15162), .ZN(n15145) );
  NOR2_X1 U18457 ( .A1(n15145), .A2(n15128), .ZN(n15138) );
  INV_X1 U18458 ( .A(n15129), .ZN(n15132) );
  OAI211_X1 U18459 ( .C1(n16146), .C2(n15133), .A(n15132), .B(n10074), .ZN(
        n15134) );
  INV_X1 U18460 ( .A(n15134), .ZN(n15135) );
  OAI21_X1 U18461 ( .B1(n16137), .B2(n15136), .A(n15135), .ZN(n15137) );
  OAI21_X1 U18462 ( .B1(n15141), .B2(n16147), .A(n15140), .ZN(P2_U3017) );
  NAND2_X1 U18463 ( .A1(n15142), .A2(n18992), .ZN(n15150) );
  OAI21_X1 U18464 ( .B1(n16146), .B2(n15965), .A(n15143), .ZN(n15147) );
  AOI21_X1 U18465 ( .B1(n15156), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15144) );
  NOR2_X1 U18466 ( .A1(n15145), .A2(n15144), .ZN(n15146) );
  AOI211_X1 U18467 ( .C1(n19008), .C2(n15148), .A(n15147), .B(n15146), .ZN(
        n15149) );
  OAI211_X1 U18468 ( .C1(n18996), .C2(n15151), .A(n15150), .B(n15149), .ZN(
        P2_U3018) );
  NAND2_X1 U18469 ( .A1(n15152), .A2(n18992), .ZN(n15164) );
  NAND2_X1 U18470 ( .A1(n19008), .A2(n15153), .ZN(n15158) );
  INV_X1 U18471 ( .A(n15154), .ZN(n15155) );
  AOI21_X1 U18472 ( .B1(n15156), .B2(n20763), .A(n15155), .ZN(n15157) );
  OAI211_X1 U18473 ( .C1(n16146), .C2(n15159), .A(n15158), .B(n15157), .ZN(
        n15161) );
  OAI21_X1 U18474 ( .B1(n15165), .B2(n15164), .A(n15163), .ZN(P2_U3019) );
  NOR2_X1 U18475 ( .A1(n15188), .A2(n15166), .ZN(n15172) );
  NAND2_X1 U18476 ( .A1(n18993), .A2(n15978), .ZN(n15170) );
  XNOR2_X1 U18477 ( .A(n15166), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15168) );
  AOI21_X1 U18478 ( .B1(n15181), .B2(n15168), .A(n15167), .ZN(n15169) );
  OAI211_X1 U18479 ( .C1(n15980), .C2(n16137), .A(n15170), .B(n15169), .ZN(
        n15171) );
  AOI211_X1 U18480 ( .C1(n15173), .C2(n16152), .A(n15172), .B(n15171), .ZN(
        n15174) );
  OAI21_X1 U18481 ( .B1(n15175), .B2(n16147), .A(n15174), .ZN(P2_U3020) );
  NAND2_X1 U18482 ( .A1(n15177), .A2(n15176), .ZN(n15179) );
  XOR2_X1 U18483 ( .A(n15179), .B(n15178), .Z(n16033) );
  INV_X1 U18484 ( .A(n16033), .ZN(n15191) );
  INV_X1 U18485 ( .A(n15029), .ZN(n15180) );
  AOI21_X1 U18486 ( .B1(n15187), .B2(n15180), .A(n15013), .ZN(n16032) );
  INV_X1 U18487 ( .A(n16036), .ZN(n15185) );
  AOI22_X1 U18488 ( .A1(n15181), .A2(n15187), .B1(n18822), .B2(
        P2_REIP_REG_25__SCAN_IN), .ZN(n15182) );
  OAI21_X1 U18489 ( .B1(n16146), .B2(n15183), .A(n15182), .ZN(n15184) );
  AOI21_X1 U18490 ( .B1(n19008), .B2(n15185), .A(n15184), .ZN(n15186) );
  OAI21_X1 U18491 ( .B1(n15188), .B2(n15187), .A(n15186), .ZN(n15189) );
  AOI21_X1 U18492 ( .B1(n16032), .B2(n16152), .A(n15189), .ZN(n15190) );
  OAI21_X1 U18493 ( .B1(n15191), .B2(n16147), .A(n15190), .ZN(P2_U3021) );
  INV_X1 U18494 ( .A(n15192), .ZN(n15202) );
  AOI21_X1 U18495 ( .B1(n15195), .B2(n15194), .A(n15193), .ZN(n15197) );
  NOR2_X1 U18496 ( .A1(n18772), .A2(n11127), .ZN(n15196) );
  AOI211_X1 U18497 ( .C1(n19008), .C2(n15991), .A(n15197), .B(n15196), .ZN(
        n15198) );
  OAI21_X1 U18498 ( .B1(n16146), .B2(n15989), .A(n15198), .ZN(n15199) );
  AOI21_X1 U18499 ( .B1(n15200), .B2(n16152), .A(n15199), .ZN(n15201) );
  OAI21_X1 U18500 ( .B1(n15202), .B2(n16147), .A(n15201), .ZN(P2_U3022) );
  OAI22_X1 U18501 ( .A1(n15293), .A2(n15203), .B1(n15410), .B2(n15409), .ZN(
        n15240) );
  NOR2_X1 U18502 ( .A1(n16146), .A2(n15204), .ZN(n15210) );
  XNOR2_X1 U18503 ( .A(n15205), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15206) );
  AOI22_X1 U18504 ( .A1(n18822), .A2(P2_REIP_REG_23__SCAN_IN), .B1(n15219), 
        .B2(n15206), .ZN(n15207) );
  OAI21_X1 U18505 ( .B1(n16137), .B2(n15208), .A(n15207), .ZN(n15209) );
  AOI211_X1 U18506 ( .C1(n15240), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15210), .B(n15209), .ZN(n15213) );
  NAND2_X1 U18507 ( .A1(n15211), .A2(n18992), .ZN(n15212) );
  OAI211_X1 U18508 ( .C1(n15214), .C2(n18996), .A(n15213), .B(n15212), .ZN(
        P2_U3023) );
  NAND3_X1 U18509 ( .A1(n15216), .A2(n16152), .A3(n15215), .ZN(n15225) );
  NAND2_X1 U18510 ( .A1(n18993), .A2(n15217), .ZN(n15221) );
  AOI22_X1 U18511 ( .A1(n18822), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n15219), 
        .B2(n15218), .ZN(n15220) );
  OAI211_X1 U18512 ( .C1(n15222), .C2(n16137), .A(n15221), .B(n15220), .ZN(
        n15223) );
  AOI21_X1 U18513 ( .B1(n15240), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15223), .ZN(n15224) );
  OAI211_X1 U18514 ( .C1(n15226), .C2(n16147), .A(n15225), .B(n15224), .ZN(
        P2_U3024) );
  NAND2_X1 U18515 ( .A1(n15058), .A2(n15227), .ZN(n15228) );
  AND2_X1 U18516 ( .A1(n15037), .A2(n15228), .ZN(n16041) );
  INV_X1 U18517 ( .A(n16041), .ZN(n15243) );
  NAND2_X1 U18518 ( .A1(n15230), .A2(n15229), .ZN(n15233) );
  NAND2_X1 U18519 ( .A1(n16043), .A2(n18992), .ZN(n15242) );
  NOR2_X1 U18520 ( .A1(n19661), .A2(n19017), .ZN(n16039) );
  AOI21_X1 U18521 ( .B1(n19008), .B2(n15234), .A(n16039), .ZN(n15235) );
  OAI21_X1 U18522 ( .B1(n16146), .B2(n15236), .A(n15235), .ZN(n15239) );
  NOR2_X1 U18523 ( .A1(n15237), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15238) );
  AOI211_X1 U18524 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15240), .A(
        n15239), .B(n15238), .ZN(n15241) );
  OAI211_X1 U18525 ( .C1(n15243), .C2(n18996), .A(n15242), .B(n15241), .ZN(
        P2_U3025) );
  AND2_X1 U18526 ( .A1(n15244), .A2(n15259), .ZN(n15245) );
  NOR2_X1 U18527 ( .A1(n15057), .A2(n15245), .ZN(n16048) );
  INV_X1 U18528 ( .A(n16048), .ZN(n15262) );
  INV_X1 U18529 ( .A(n15246), .ZN(n15248) );
  NAND2_X1 U18530 ( .A1(n15248), .A2(n15247), .ZN(n15251) );
  INV_X1 U18531 ( .A(n15249), .ZN(n15269) );
  AOI21_X1 U18532 ( .B1(n15267), .B2(n15269), .A(n15265), .ZN(n15250) );
  XNOR2_X1 U18533 ( .A(n15251), .B(n15250), .ZN(n16049) );
  NAND2_X1 U18534 ( .A1(n16049), .A2(n18992), .ZN(n15261) );
  NAND2_X1 U18535 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15252) );
  INV_X1 U18536 ( .A(n15413), .ZN(n15287) );
  NOR2_X1 U18537 ( .A1(n15412), .A2(n15287), .ZN(n15394) );
  AOI21_X1 U18538 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15409), .A(
        n15410), .ZN(n15395) );
  AOI21_X1 U18539 ( .B1(n15252), .B2(n15394), .A(n15395), .ZN(n15371) );
  OAI21_X1 U18540 ( .B1(n15314), .B2(n15293), .A(n15371), .ZN(n15333) );
  AOI21_X1 U18541 ( .B1(n15253), .B2(n15452), .A(n15333), .ZN(n15274) );
  INV_X1 U18542 ( .A(n15274), .ZN(n15254) );
  AOI21_X1 U18543 ( .B1(n15452), .B2(n15275), .A(n15254), .ZN(n15637) );
  INV_X1 U18544 ( .A(n18683), .ZN(n15256) );
  OAI22_X1 U18545 ( .A1(n16137), .A2(n18684), .B1(n20834), .B2(n18772), .ZN(
        n15255) );
  AOI21_X1 U18546 ( .B1(n18993), .B2(n15256), .A(n15255), .ZN(n15257) );
  OAI21_X1 U18547 ( .B1(n15637), .B2(n15259), .A(n15257), .ZN(n15258) );
  AOI21_X1 U18548 ( .B1(n15643), .B2(n15259), .A(n15258), .ZN(n15260) );
  OAI211_X1 U18549 ( .C1(n15262), .C2(n18996), .A(n15261), .B(n15260), .ZN(
        P2_U3027) );
  NAND2_X1 U18550 ( .A1(n15263), .A2(n15275), .ZN(n15264) );
  NAND2_X1 U18551 ( .A1(n15264), .A2(n15244), .ZN(n16052) );
  INV_X1 U18552 ( .A(n15265), .ZN(n15266) );
  NAND2_X1 U18553 ( .A1(n15267), .A2(n15266), .ZN(n15268) );
  XNOR2_X1 U18554 ( .A(n15269), .B(n15268), .ZN(n16053) );
  INV_X1 U18555 ( .A(n16053), .ZN(n15270) );
  NAND2_X1 U18556 ( .A1(n15270), .A2(n18992), .ZN(n15286) );
  AOI21_X1 U18557 ( .B1(n14970), .B2(n15272), .A(n15271), .ZN(n18696) );
  NAND2_X1 U18558 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n18839), .ZN(n15273) );
  OAI221_X1 U18559 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15276), 
        .C1(n15275), .C2(n15274), .A(n15273), .ZN(n15283) );
  NAND2_X1 U18560 ( .A1(n15278), .A2(n15277), .ZN(n15281) );
  INV_X1 U18561 ( .A(n15279), .ZN(n15280) );
  INV_X1 U18562 ( .A(n18695), .ZN(n16016) );
  NOR2_X1 U18563 ( .A1(n16137), .A2(n16016), .ZN(n15282) );
  OR2_X1 U18564 ( .A1(n15283), .A2(n15282), .ZN(n15284) );
  AOI21_X1 U18565 ( .B1(n18696), .B2(n18993), .A(n15284), .ZN(n15285) );
  OAI211_X1 U18566 ( .C1(n16052), .C2(n18996), .A(n15286), .B(n15285), .ZN(
        P2_U3028) );
  NOR2_X1 U18567 ( .A1(n15288), .A2(n15287), .ZN(n15327) );
  NOR2_X1 U18568 ( .A1(n15289), .A2(n15315), .ZN(n15290) );
  AOI22_X1 U18569 ( .A1(n15291), .A2(n16152), .B1(n15327), .B2(n15290), .ZN(
        n15300) );
  INV_X1 U18570 ( .A(n19000), .ZN(n15292) );
  OAI21_X1 U18571 ( .B1(n16137), .B2(n18708), .A(n15294), .ZN(n15296) );
  NOR2_X1 U18572 ( .A1(n18707), .A2(n16146), .ZN(n15295) );
  AOI211_X1 U18573 ( .C1(n18992), .C2(n15297), .A(n15296), .B(n15295), .ZN(
        n15298) );
  OAI211_X1 U18574 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n15300), .A(
        n15299), .B(n15298), .ZN(P2_U3029) );
  AOI22_X1 U18575 ( .A1(n15301), .A2(n16152), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15327), .ZN(n15313) );
  INV_X1 U18576 ( .A(n15302), .ZN(n15303) );
  NAND2_X1 U18577 ( .A1(n15303), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15312) );
  AND2_X1 U18578 ( .A1(n15305), .A2(n15304), .ZN(n15306) );
  NOR2_X1 U18579 ( .A1(n14969), .A2(n15306), .ZN(n18913) );
  NOR2_X1 U18580 ( .A1(n15307), .A2(n16147), .ZN(n15310) );
  OAI21_X1 U18581 ( .B1(n16137), .B2(n18880), .A(n15308), .ZN(n15309) );
  AOI211_X1 U18582 ( .C1(n18913), .C2(n18993), .A(n15310), .B(n15309), .ZN(
        n15311) );
  OAI211_X1 U18583 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15313), .A(
        n15312), .B(n15311), .ZN(P2_U3030) );
  NAND2_X1 U18584 ( .A1(n15358), .A2(n15314), .ZN(n16066) );
  NAND2_X1 U18585 ( .A1(n16066), .A2(n15315), .ZN(n15317) );
  NAND2_X1 U18586 ( .A1(n15317), .A2(n15316), .ZN(n16057) );
  NOR2_X1 U18587 ( .A1(n15319), .A2(n15318), .ZN(n15326) );
  INV_X1 U18588 ( .A(n15320), .ZN(n15324) );
  OAI21_X1 U18589 ( .B1(n15337), .B2(n15322), .A(n15066), .ZN(n16065) );
  OR2_X1 U18590 ( .A1(n15323), .A2(n15324), .ZN(n16064) );
  NOR2_X1 U18591 ( .A1(n16065), .A2(n16064), .ZN(n16063) );
  NOR2_X1 U18592 ( .A1(n15324), .A2(n16063), .ZN(n15325) );
  XOR2_X1 U18593 ( .A(n15326), .B(n15325), .Z(n16060) );
  NAND2_X1 U18594 ( .A1(n16060), .A2(n18992), .ZN(n15335) );
  INV_X1 U18595 ( .A(n15327), .ZN(n15330) );
  NOR2_X1 U18596 ( .A1(n10711), .A2(n18772), .ZN(n15328) );
  AOI21_X1 U18597 ( .B1(n19008), .B2(n16058), .A(n15328), .ZN(n15329) );
  OAI21_X1 U18598 ( .B1(n15330), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15329), .ZN(n15332) );
  NOR2_X1 U18599 ( .A1(n18731), .A2(n16146), .ZN(n15331) );
  AOI211_X1 U18600 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15333), .A(
        n15332), .B(n15331), .ZN(n15334) );
  OAI211_X1 U18601 ( .C1(n16057), .C2(n18996), .A(n15335), .B(n15334), .ZN(
        P2_U3031) );
  NOR2_X1 U18602 ( .A1(n15337), .A2(n15336), .ZN(n15340) );
  NAND2_X1 U18603 ( .A1(n15066), .A2(n15338), .ZN(n15339) );
  XNOR2_X1 U18604 ( .A(n15340), .B(n15339), .ZN(n16076) );
  INV_X1 U18605 ( .A(n16076), .ZN(n15350) );
  NAND2_X1 U18606 ( .A1(n15358), .A2(n16120), .ZN(n16068) );
  INV_X1 U18607 ( .A(n16068), .ZN(n15342) );
  AOI21_X1 U18608 ( .B1(n15358), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15341) );
  NOR2_X1 U18609 ( .A1(n15342), .A2(n15341), .ZN(n16075) );
  NAND3_X1 U18610 ( .A1(n15343), .A2(n15413), .A3(n15364), .ZN(n15360) );
  NAND2_X1 U18611 ( .A1(n15371), .A2(n15360), .ZN(n16127) );
  NAND2_X1 U18612 ( .A1(n15343), .A2(n15413), .ZN(n16122) );
  NOR2_X1 U18613 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16122), .ZN(
        n16128) );
  INV_X1 U18614 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19651) );
  NOR2_X1 U18615 ( .A1(n19651), .A2(n18772), .ZN(n15344) );
  AOI21_X1 U18616 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16128), .A(
        n15344), .ZN(n15345) );
  OAI21_X1 U18617 ( .B1(n16137), .B2(n16074), .A(n15345), .ZN(n15346) );
  AOI21_X1 U18618 ( .B1(n16127), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15346), .ZN(n15347) );
  OAI21_X1 U18619 ( .B1(n18758), .B2(n16146), .A(n15347), .ZN(n15348) );
  AOI21_X1 U18620 ( .B1(n16075), .B2(n16152), .A(n15348), .ZN(n15349) );
  OAI21_X1 U18621 ( .B1(n15350), .B2(n16147), .A(n15349), .ZN(P2_U3033) );
  INV_X1 U18622 ( .A(n15351), .ZN(n15352) );
  NAND2_X1 U18623 ( .A1(n15353), .A2(n15352), .ZN(n15357) );
  NOR2_X1 U18624 ( .A1(n15355), .A2(n15336), .ZN(n15356) );
  XNOR2_X1 U18625 ( .A(n15357), .B(n15356), .ZN(n16081) );
  XNOR2_X1 U18626 ( .A(n9745), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16080) );
  NAND2_X1 U18627 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18822), .ZN(n15359) );
  OAI211_X1 U18628 ( .C1(n16137), .C2(n18889), .A(n15360), .B(n15359), .ZN(
        n15361) );
  AOI21_X1 U18629 ( .B1(n15362), .B2(n18993), .A(n15361), .ZN(n15363) );
  OAI21_X1 U18630 ( .B1(n15371), .B2(n15364), .A(n15363), .ZN(n15365) );
  AOI21_X1 U18631 ( .B1(n16080), .B2(n16152), .A(n15365), .ZN(n15366) );
  OAI21_X1 U18632 ( .B1(n16081), .B2(n16147), .A(n15366), .ZN(P2_U3034) );
  OAI21_X1 U18633 ( .B1(n16104), .B2(n15393), .A(n15367), .ZN(n15368) );
  NAND2_X1 U18634 ( .A1(n15368), .A2(n9745), .ZN(n16088) );
  INV_X1 U18635 ( .A(n18770), .ZN(n15374) );
  INV_X1 U18636 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15369) );
  OAI22_X1 U18637 ( .A1(n16137), .A2(n18765), .B1(n18772), .B2(n15369), .ZN(
        n15373) );
  AOI21_X1 U18638 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15394), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15370) );
  NOR2_X1 U18639 ( .A1(n15371), .A2(n15370), .ZN(n15372) );
  AOI211_X1 U18640 ( .C1(n18993), .C2(n15374), .A(n15373), .B(n15372), .ZN(
        n15383) );
  NAND2_X1 U18641 ( .A1(n15376), .A2(n15375), .ZN(n15381) );
  INV_X1 U18642 ( .A(n15377), .ZN(n15379) );
  OR2_X1 U18643 ( .A1(n15379), .A2(n15378), .ZN(n15380) );
  XNOR2_X1 U18644 ( .A(n15381), .B(n15380), .ZN(n16089) );
  NAND2_X1 U18645 ( .A1(n16089), .A2(n18992), .ZN(n15382) );
  OAI211_X1 U18646 ( .C1(n16088), .C2(n18996), .A(n15383), .B(n15382), .ZN(
        P2_U3035) );
  XNOR2_X1 U18647 ( .A(n16104), .B(n15393), .ZN(n16097) );
  INV_X1 U18648 ( .A(n15384), .ZN(n15404) );
  OR2_X1 U18649 ( .A1(n15385), .A2(n15404), .ZN(n15389) );
  AND2_X1 U18650 ( .A1(n15387), .A2(n15386), .ZN(n15388) );
  XNOR2_X1 U18651 ( .A(n15389), .B(n15388), .ZN(n16096) );
  INV_X1 U18652 ( .A(n16096), .ZN(n15402) );
  XNOR2_X1 U18653 ( .A(n15391), .B(n15390), .ZN(n18925) );
  NOR2_X1 U18654 ( .A1(n11030), .A2(n18772), .ZN(n15392) );
  AOI221_X1 U18655 ( .B1(n15395), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n15394), .C2(n15393), .A(n15392), .ZN(n15400) );
  NAND2_X1 U18656 ( .A1(n15396), .A2(n13540), .ZN(n15398) );
  INV_X1 U18657 ( .A(n13591), .ZN(n15397) );
  AND2_X1 U18658 ( .A1(n15398), .A2(n15397), .ZN(n18897) );
  NAND2_X1 U18659 ( .A1(n19008), .A2(n18897), .ZN(n15399) );
  OAI211_X1 U18660 ( .C1(n16146), .C2(n18925), .A(n15400), .B(n15399), .ZN(
        n15401) );
  AOI21_X1 U18661 ( .B1(n15402), .B2(n18992), .A(n15401), .ZN(n15403) );
  OAI21_X1 U18662 ( .B1(n16097), .B2(n18996), .A(n15403), .ZN(P2_U3036) );
  NOR2_X1 U18663 ( .A1(n15405), .A2(n15404), .ZN(n15407) );
  XOR2_X1 U18664 ( .A(n15407), .B(n15406), .Z(n16102) );
  INV_X1 U18665 ( .A(n16101), .ZN(n15408) );
  NAND3_X1 U18666 ( .A1(n15408), .A2(n16152), .A3(n16104), .ZN(n15419) );
  NOR2_X1 U18667 ( .A1(n15410), .A2(n15409), .ZN(n15414) );
  INV_X1 U18668 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19646) );
  NOR2_X1 U18669 ( .A1(n19646), .A2(n18772), .ZN(n15411) );
  AOI221_X1 U18670 ( .B1(n15414), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n15413), .C2(n15412), .A(n15411), .ZN(n15415) );
  INV_X1 U18671 ( .A(n15415), .ZN(n15417) );
  OAI22_X1 U18672 ( .A1(n18789), .A2(n16146), .B1(n16137), .B2(n18788), .ZN(
        n15416) );
  NOR2_X1 U18673 ( .A1(n15417), .A2(n15416), .ZN(n15418) );
  OAI211_X1 U18674 ( .C1(n16102), .C2(n16147), .A(n15419), .B(n15418), .ZN(
        P2_U3037) );
  NAND2_X1 U18675 ( .A1(n15420), .A2(n16152), .ZN(n15427) );
  INV_X1 U18676 ( .A(n16134), .ZN(n15425) );
  AOI22_X1 U18677 ( .A1(n19008), .A2(n18814), .B1(n18822), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n15421) );
  OAI21_X1 U18678 ( .B1(n18818), .B2(n16146), .A(n15421), .ZN(n15424) );
  INV_X1 U18679 ( .A(n15435), .ZN(n15422) );
  NOR3_X1 U18680 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15422), .A3(
        n15434), .ZN(n15423) );
  AOI211_X1 U18681 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15425), .A(
        n15424), .B(n15423), .ZN(n15426) );
  OAI211_X1 U18682 ( .C1(n15428), .C2(n16147), .A(n15427), .B(n15426), .ZN(
        P2_U3040) );
  XNOR2_X1 U18683 ( .A(n15429), .B(n15430), .ZN(n16110) );
  OAI21_X1 U18684 ( .B1(n15433), .B2(n15432), .A(n15431), .ZN(n18935) );
  OAI211_X1 U18685 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n15435), .B(n15434), .ZN(n15437) );
  AOI22_X1 U18686 ( .A1(n19008), .A2(n18826), .B1(n18822), .B2(
        P2_REIP_REG_5__SCAN_IN), .ZN(n15436) );
  OAI211_X1 U18687 ( .C1(n18935), .C2(n16146), .A(n15437), .B(n15436), .ZN(
        n15443) );
  NAND2_X1 U18688 ( .A1(n15439), .A2(n15438), .ZN(n15440) );
  XOR2_X1 U18689 ( .A(n15441), .B(n15440), .Z(n16109) );
  NOR2_X1 U18690 ( .A1(n16109), .A2(n18996), .ZN(n15442) );
  AOI211_X1 U18691 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15444), .A(
        n15443), .B(n15442), .ZN(n15445) );
  OAI21_X1 U18692 ( .B1(n16147), .B2(n16110), .A(n15445), .ZN(P2_U3041) );
  OAI22_X1 U18693 ( .A1(n16147), .A2(n15447), .B1(n19004), .B2(n15446), .ZN(
        n15448) );
  AOI211_X1 U18694 ( .C1(n18993), .C2(n19717), .A(n15449), .B(n15448), .ZN(
        n15455) );
  OAI22_X1 U18695 ( .A1(n15450), .A2(n18996), .B1(n16137), .B2(n18853), .ZN(
        n15451) );
  INV_X1 U18696 ( .A(n15451), .ZN(n15454) );
  OAI211_X1 U18697 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15452), .B(n19001), .ZN(n15453) );
  NAND3_X1 U18698 ( .A1(n15455), .A2(n15454), .A3(n15453), .ZN(P2_U3045) );
  INV_X1 U18699 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16683) );
  INV_X1 U18700 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16681) );
  NAND4_X1 U18701 ( .A1(n17999), .A2(n17983), .A3(n15457), .A4(n15456), .ZN(
        n15459) );
  INV_X1 U18702 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n15462) );
  NAND2_X1 U18703 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16664) );
  INV_X1 U18704 ( .A(n16664), .ZN(n16973) );
  AND2_X1 U18705 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n16973), .ZN(n16965) );
  NAND3_X1 U18706 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n16965), .ZN(n16960) );
  INV_X1 U18707 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16949) );
  INV_X1 U18708 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16956) );
  NOR4_X1 U18709 ( .A1(n16949), .A2(n16589), .A3(n16956), .A4(n16896), .ZN(
        n15461) );
  NAND4_X1 U18710 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(n15461), .ZN(n16883) );
  NOR3_X1 U18711 ( .A1(n15462), .A2(n16960), .A3(n16883), .ZN(n15549) );
  NAND2_X1 U18712 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16869), .ZN(n16868) );
  NAND2_X1 U18713 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16843), .ZN(n16817) );
  NOR2_X2 U18714 ( .A1(n16475), .A2(n16817), .ZN(n16831) );
  NAND2_X1 U18715 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16831), .ZN(n16814) );
  NOR2_X1 U18716 ( .A1(n17032), .A2(n16773), .ZN(n16775) );
  NAND2_X1 U18717 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16775), .ZN(n16762) );
  NAND2_X1 U18718 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16744), .ZN(n16738) );
  NOR2_X2 U18719 ( .A1(n16683), .A2(n16738), .ZN(n16743) );
  INV_X1 U18720 ( .A(n16728), .ZN(n16733) );
  NAND2_X1 U18721 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16733), .ZN(n15536) );
  NOR2_X2 U18722 ( .A1(n17999), .A2(n16978), .ZN(n16982) );
  INV_X1 U18723 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16685) );
  NOR3_X1 U18724 ( .A1(n16685), .A2(n16684), .A3(n16728), .ZN(n16722) );
  NOR2_X1 U18725 ( .A1(n16982), .A2(n16722), .ZN(n16723) );
  AOI22_X1 U18726 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U18727 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16919), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15465) );
  AOI22_X1 U18728 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9600), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15464) );
  AOI22_X1 U18729 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15463) );
  NAND4_X1 U18730 ( .A1(n15466), .A2(n15465), .A3(n15464), .A4(n15463), .ZN(
        n15472) );
  AOI22_X1 U18731 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U18732 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15469) );
  AOI22_X1 U18733 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15468) );
  AOI22_X1 U18734 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15467) );
  NAND4_X1 U18735 ( .A1(n15470), .A2(n15469), .A3(n15468), .A4(n15467), .ZN(
        n15471) );
  NOR2_X1 U18736 ( .A1(n15472), .A2(n15471), .ZN(n15534) );
  AOI22_X1 U18737 ( .A1(n16921), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U18738 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15475) );
  AOI22_X1 U18739 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15474) );
  AOI22_X1 U18740 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9609), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15473) );
  NAND4_X1 U18741 ( .A1(n15476), .A2(n15475), .A3(n15474), .A4(n15473), .ZN(
        n15482) );
  AOI22_X1 U18742 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15480) );
  AOI22_X1 U18743 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15479) );
  AOI22_X1 U18744 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U18745 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16919), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15477) );
  NAND4_X1 U18746 ( .A1(n15480), .A2(n15479), .A3(n15478), .A4(n15477), .ZN(
        n15481) );
  NOR2_X1 U18747 ( .A1(n15482), .A2(n15481), .ZN(n16730) );
  AOI22_X1 U18748 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16920), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15486) );
  AOI22_X1 U18749 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n16932), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15485) );
  AOI22_X1 U18750 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n16919), .ZN(n15484) );
  AOI22_X1 U18751 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n16819), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n9609), .ZN(n15483) );
  NAND4_X1 U18752 ( .A1(n15486), .A2(n15485), .A3(n15484), .A4(n15483), .ZN(
        n15492) );
  AOI22_X1 U18753 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9608), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n9600), .ZN(n15490) );
  AOI22_X1 U18754 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n15537), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15489) );
  AOI22_X1 U18755 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10299), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n15538), .ZN(n15488) );
  AOI22_X1 U18756 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n16933), .ZN(n15487) );
  NAND4_X1 U18757 ( .A1(n15490), .A2(n15489), .A3(n15488), .A4(n15487), .ZN(
        n15491) );
  NOR2_X1 U18758 ( .A1(n15492), .A2(n15491), .ZN(n16740) );
  AOI22_X1 U18759 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15502) );
  AOI22_X1 U18760 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15501) );
  AOI22_X1 U18761 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9604), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15493) );
  OAI21_X1 U18762 ( .B1(n10094), .B2(n20816), .A(n15493), .ZN(n15499) );
  AOI22_X1 U18763 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15497) );
  AOI22_X1 U18764 ( .A1(n16939), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15496) );
  AOI22_X1 U18765 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15495) );
  AOI22_X1 U18766 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15494) );
  NAND4_X1 U18767 ( .A1(n15497), .A2(n15496), .A3(n15495), .A4(n15494), .ZN(
        n15498) );
  AOI211_X1 U18768 ( .C1(n15537), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n15499), .B(n15498), .ZN(n15500) );
  NAND3_X1 U18769 ( .A1(n15502), .A2(n15501), .A3(n15500), .ZN(n16746) );
  AOI22_X1 U18770 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15512) );
  AOI22_X1 U18771 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15511) );
  AOI22_X1 U18772 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9609), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15503) );
  OAI21_X1 U18773 ( .B1(n16804), .B2(n16953), .A(n15503), .ZN(n15509) );
  AOI22_X1 U18774 ( .A1(n10311), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15507) );
  AOI22_X1 U18775 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16931), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15506) );
  AOI22_X1 U18776 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15505) );
  AOI22_X1 U18777 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15504) );
  NAND4_X1 U18778 ( .A1(n15507), .A2(n15506), .A3(n15505), .A4(n15504), .ZN(
        n15508) );
  AOI211_X1 U18779 ( .C1(n15537), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n15509), .B(n15508), .ZN(n15510) );
  NAND3_X1 U18780 ( .A1(n15512), .A2(n15511), .A3(n15510), .ZN(n16747) );
  NAND2_X1 U18781 ( .A1(n16746), .A2(n16747), .ZN(n16745) );
  NOR2_X1 U18782 ( .A1(n16740), .A2(n16745), .ZN(n16739) );
  AOI22_X1 U18783 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U18784 ( .A1(n16921), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15521) );
  AOI22_X1 U18785 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15513) );
  OAI21_X1 U18786 ( .B1(n16705), .B2(n16976), .A(n15513), .ZN(n15519) );
  AOI22_X1 U18787 ( .A1(n15538), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15517) );
  AOI22_X1 U18788 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15516) );
  AOI22_X1 U18789 ( .A1(n10150), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15515) );
  AOI22_X1 U18790 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9609), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15514) );
  NAND4_X1 U18791 ( .A1(n15517), .A2(n15516), .A3(n15515), .A4(n15514), .ZN(
        n15518) );
  AOI211_X1 U18792 ( .C1(n16914), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n15519), .B(n15518), .ZN(n15520) );
  NAND3_X1 U18793 ( .A1(n15522), .A2(n15521), .A3(n15520), .ZN(n16735) );
  NAND2_X1 U18794 ( .A1(n16739), .A2(n16735), .ZN(n16734) );
  NOR2_X1 U18795 ( .A1(n16730), .A2(n16734), .ZN(n16729) );
  AOI22_X1 U18796 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15533) );
  AOI22_X1 U18797 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15532) );
  INV_X1 U18798 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U18799 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15523) );
  OAI21_X1 U18800 ( .B1(n16705), .B2(n16967), .A(n15523), .ZN(n15530) );
  AOI22_X1 U18801 ( .A1(n16940), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15528) );
  AOI22_X1 U18802 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U18803 ( .A1(n16939), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15526) );
  AOI22_X1 U18804 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15525) );
  NAND4_X1 U18805 ( .A1(n15528), .A2(n15527), .A3(n15526), .A4(n15525), .ZN(
        n15529) );
  AOI211_X1 U18806 ( .C1(n15537), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n15530), .B(n15529), .ZN(n15531) );
  NAND3_X1 U18807 ( .A1(n15533), .A2(n15532), .A3(n15531), .ZN(n16726) );
  NAND2_X1 U18808 ( .A1(n16729), .A2(n16726), .ZN(n16725) );
  NOR2_X1 U18809 ( .A1(n15534), .A2(n16725), .ZN(n16720) );
  AOI21_X1 U18810 ( .B1(n15534), .B2(n16725), .A(n16720), .ZN(n17002) );
  AOI22_X1 U18811 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16723), .B1(n17002), 
        .B2(n16982), .ZN(n15535) );
  OAI21_X1 U18812 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15536), .A(n15535), .ZN(
        P3_U2675) );
  AOI22_X1 U18813 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9604), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U18814 ( .A1(n16939), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15541) );
  AOI22_X1 U18815 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15540) );
  AOI22_X1 U18816 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15539) );
  NAND4_X1 U18817 ( .A1(n15542), .A2(n15541), .A3(n15540), .A4(n15539), .ZN(
        n15548) );
  AOI22_X1 U18818 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15546) );
  AOI22_X1 U18819 ( .A1(n10311), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15545) );
  AOI22_X1 U18820 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10143), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15544) );
  AOI22_X1 U18821 ( .A1(n16921), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15543) );
  NAND4_X1 U18822 ( .A1(n15546), .A2(n15545), .A3(n15544), .A4(n15543), .ZN(
        n15547) );
  NOR2_X1 U18823 ( .A1(n15548), .A2(n15547), .ZN(n17080) );
  NAND3_X1 U18824 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16969), .A3(n16884), 
        .ZN(n15551) );
  NOR2_X1 U18825 ( .A1(n17032), .A2(n16978), .ZN(n16981) );
  NAND3_X1 U18826 ( .A1(n15549), .A2(n16981), .A3(n16518), .ZN(n15550) );
  OAI211_X1 U18827 ( .C1(n17080), .C2(n16969), .A(n15551), .B(n15550), .ZN(
        P3_U2690) );
  NAND2_X1 U18828 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18133) );
  AOI221_X1 U18829 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18133), .C1(n15553), 
        .C2(n18133), .A(n15552), .ZN(n17962) );
  NOR2_X1 U18830 ( .A1(n15554), .A2(n18423), .ZN(n15555) );
  OAI21_X1 U18831 ( .B1(n15555), .B2(n18303), .A(n17963), .ZN(n17960) );
  AOI22_X1 U18832 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17962), .B1(
        n17960), .B2(n18442), .ZN(P3_U2865) );
  NAND4_X1 U18833 ( .A1(n15557), .A2(n12747), .A3(n19693), .A4(n15556), .ZN(
        n15558) );
  OR2_X1 U18834 ( .A1(n15559), .A2(n15558), .ZN(n15560) );
  OAI21_X1 U18835 ( .B1(n15562), .B2(n15561), .A(n15560), .ZN(P2_U3595) );
  NOR2_X1 U18836 ( .A1(n17951), .A2(n17690), .ZN(n17863) );
  INV_X1 U18837 ( .A(n15563), .ZN(n15564) );
  NOR2_X1 U18838 ( .A1(n15565), .A2(n15564), .ZN(n17657) );
  NAND4_X1 U18839 ( .A1(n15566), .A2(n17934), .A3(n17268), .A4(n17657), .ZN(
        n16198) );
  OAI21_X1 U18840 ( .B1(n17930), .B2(n16187), .A(n16198), .ZN(n15567) );
  AOI21_X1 U18841 ( .B1(n15568), .B2(n17863), .A(n15567), .ZN(n15613) );
  INV_X1 U18842 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16190) );
  INV_X1 U18843 ( .A(n17897), .ZN(n17855) );
  NAND2_X1 U18844 ( .A1(n17934), .A2(n17855), .ZN(n17936) );
  NOR2_X1 U18845 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17936), .ZN(
        n15570) );
  AOI22_X1 U18846 ( .A1(n16170), .A2(n17863), .B1(n16169), .B2(n17947), .ZN(
        n15569) );
  INV_X1 U18847 ( .A(n15569), .ZN(n15615) );
  AOI211_X1 U18848 ( .C1(n17950), .C2(n15571), .A(n15570), .B(n15615), .ZN(
        n15576) );
  OAI21_X1 U18849 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15573), .A(
        n15572), .ZN(n15574) );
  INV_X1 U18850 ( .A(n15574), .ZN(n16193) );
  AOI22_X1 U18851 ( .A1(n17877), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n17862), 
        .B2(n16193), .ZN(n15575) );
  OAI221_X1 U18852 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15613), 
        .C1(n16190), .C2(n15576), .A(n15575), .ZN(P3_U2833) );
  NOR3_X1 U18853 ( .A1(n15578), .A2(n15577), .A3(n20446), .ZN(n15581) );
  NAND2_X1 U18854 ( .A1(n15581), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15583) );
  OAI22_X1 U18855 ( .A1(n15581), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n15580), .B2(n15579), .ZN(n15582) );
  NAND2_X1 U18856 ( .A1(n15583), .A2(n15582), .ZN(n15586) );
  INV_X1 U18857 ( .A(n15584), .ZN(n15585) );
  AOI222_X1 U18858 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15586), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15585), .C1(n15586), 
        .C2(n15585), .ZN(n15588) );
  AOI222_X1 U18859 ( .A1(n15588), .A2(n20673), .B1(n15588), .B2(n15587), .C1(
        n20673), .C2(n15587), .ZN(n15589) );
  OR2_X1 U18860 ( .A1(n15589), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n15598) );
  NOR2_X1 U18861 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15594) );
  INV_X1 U18862 ( .A(n15590), .ZN(n15591) );
  OAI211_X1 U18863 ( .C1(n15594), .C2(n15593), .A(n15592), .B(n15591), .ZN(
        n15595) );
  NOR2_X1 U18864 ( .A1(n15596), .A2(n15595), .ZN(n15597) );
  NOR3_X1 U18865 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20703), .A3(n15599), 
        .ZN(n15609) );
  NAND2_X1 U18866 ( .A1(n15600), .A2(n20771), .ZN(n15603) );
  OAI21_X1 U18867 ( .B1(n15601), .B2(n20708), .A(n20582), .ZN(n15602) );
  OAI21_X1 U18868 ( .B1(n15604), .B2(n15603), .A(n15602), .ZN(n15951) );
  INV_X1 U18869 ( .A(n15610), .ZN(n15605) );
  OAI21_X1 U18870 ( .B1(n15951), .B2(n15605), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n15956) );
  OAI211_X1 U18871 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20708), .A(n15606), 
        .B(n15954), .ZN(n15607) );
  OAI22_X1 U18872 ( .A1(n15950), .A2(n15951), .B1(n15956), .B2(n15607), .ZN(
        n15608) );
  OAI22_X1 U18873 ( .A1(n15610), .A2(n19763), .B1(n15609), .B2(n15608), .ZN(
        P1_U3161) );
  OAI21_X1 U18874 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15612), .A(
        n15611), .ZN(n16181) );
  OR2_X1 U18875 ( .A1(n15613), .A2(n16190), .ZN(n15617) );
  AOI221_X1 U18876 ( .B1(n17897), .B2(n15614), .C1(n16178), .C2(n15614), .A(
        n17877), .ZN(n16203) );
  NOR2_X1 U18877 ( .A1(n16203), .A2(n15615), .ZN(n15616) );
  MUX2_X1 U18878 ( .A(n15617), .B(n15616), .S(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n15618) );
  NAND2_X1 U18879 ( .A1(n17877), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16171) );
  OAI211_X1 U18880 ( .C1(n17807), .C2(n16181), .A(n15618), .B(n16171), .ZN(
        P3_U2832) );
  INV_X1 U18881 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20599) );
  INV_X1 U18882 ( .A(HOLD), .ZN(n20585) );
  NOR2_X1 U18883 ( .A1(n20599), .A2(n20585), .ZN(n15622) );
  AOI22_X1 U18884 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15621) );
  NAND2_X1 U18885 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15619), .ZN(n20593) );
  OAI211_X1 U18886 ( .C1(n15622), .C2(n15621), .A(n15620), .B(n20593), .ZN(
        P1_U3195) );
  AND2_X1 U18887 ( .A1(n19875), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OAI221_X1 U18888 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n19692), .C1(n19751), 
        .C2(n19618), .A(n19549), .ZN(n19616) );
  OAI211_X1 U18889 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(
        P2_STATE2_REG_1__SCAN_IN), .A(n15623), .B(n19616), .ZN(n15624) );
  INV_X1 U18890 ( .A(n15624), .ZN(P2_U3178) );
  AOI221_X1 U18891 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16158), .C1(n19732), .C2(
        n16158), .A(n19554), .ZN(n19727) );
  INV_X1 U18892 ( .A(n19727), .ZN(n19728) );
  NOR2_X1 U18893 ( .A1(n15625), .A2(n19728), .ZN(P2_U3047) );
  NOR2_X1 U18894 ( .A1(n18619), .A2(n17138), .ZN(n15626) );
  NOR2_X1 U18895 ( .A1(n18418), .A2(n17123), .ZN(n17133) );
  AOI22_X1 U18896 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17133), .B1(n17130), .B2(
        P3_EAX_REG_0__SCAN_IN), .ZN(n15630) );
  NOR2_X1 U18897 ( .A1(n17130), .A2(n17032), .ZN(n17129) );
  INV_X1 U18898 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17197) );
  NAND2_X1 U18899 ( .A1(n17129), .A2(n17197), .ZN(n15629) );
  OAI211_X1 U18900 ( .C1(n15631), .C2(n17125), .A(n15630), .B(n15629), .ZN(
        P3_U2735) );
  NAND2_X1 U18901 ( .A1(n15633), .A2(n15632), .ZN(n15635) );
  NAND2_X1 U18902 ( .A1(n15635), .A2(n9932), .ZN(n18670) );
  OAI22_X1 U18903 ( .A1(n15637), .A2(n15636), .B1(n16146), .B2(n18670), .ZN(
        n15638) );
  INV_X1 U18904 ( .A(n15638), .ZN(n15647) );
  OAI222_X1 U18905 ( .A1(n18671), .A2(n16137), .B1(n15640), .B2(n16147), .C1(
        n15639), .C2(n18996), .ZN(n15641) );
  INV_X1 U18906 ( .A(n15641), .ZN(n15646) );
  OAI211_X1 U18907 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15643), .B(n15642), .ZN(
        n15644) );
  NAND4_X1 U18908 ( .A1(n15647), .A2(n15646), .A3(n15645), .A4(n15644), .ZN(
        P2_U3026) );
  AND2_X1 U18909 ( .A1(n15648), .A2(n19831), .ZN(n15652) );
  AOI22_X1 U18910 ( .A1(n19838), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n19832), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n15649) );
  OAI21_X1 U18911 ( .B1(n15650), .B2(n14497), .A(n15649), .ZN(n15651) );
  AOI21_X1 U18912 ( .B1(n15653), .B2(n15652), .A(n15651), .ZN(n15656) );
  NOR2_X1 U18913 ( .A1(n15789), .A2(n15773), .ZN(n15654) );
  AOI21_X1 U18914 ( .B1(n15798), .B2(n19802), .A(n15654), .ZN(n15655) );
  OAI211_X1 U18915 ( .C1(n15657), .C2(n19818), .A(n15656), .B(n15655), .ZN(
        P1_U2814) );
  NOR2_X1 U18916 ( .A1(n15685), .A2(n15658), .ZN(n15665) );
  NAND2_X1 U18917 ( .A1(n15659), .A2(n15674), .ZN(n15660) );
  NAND2_X1 U18918 ( .A1(n19790), .A2(n15660), .ZN(n15684) );
  OAI21_X1 U18919 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n15685), .A(n15684), 
        .ZN(n15664) );
  OAI22_X1 U18920 ( .A1(n19813), .A2(n15662), .B1(n15661), .B2(n15770), .ZN(
        n15663) );
  AOI221_X1 U18921 ( .B1(n15665), .B2(n20640), .C1(n15664), .C2(
        P1_REIP_REG_25__SCAN_IN), .A(n15663), .ZN(n15671) );
  INV_X1 U18922 ( .A(n15666), .ZN(n15667) );
  OAI22_X1 U18923 ( .A1(n15668), .A2(n15779), .B1(n15667), .B2(n19818), .ZN(
        n15669) );
  INV_X1 U18924 ( .A(n15669), .ZN(n15670) );
  OAI211_X1 U18925 ( .C1(n15773), .C2(n15672), .A(n15671), .B(n15670), .ZN(
        P1_U2815) );
  NOR2_X1 U18926 ( .A1(n15685), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15673) );
  AOI22_X1 U18927 ( .A1(n15674), .A2(n15673), .B1(n19832), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n15676) );
  NAND2_X1 U18928 ( .A1(n19838), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15675) );
  OAI211_X1 U18929 ( .C1(n15684), .C2(n15677), .A(n15676), .B(n15675), .ZN(
        n15678) );
  INV_X1 U18930 ( .A(n15678), .ZN(n15682) );
  AOI22_X1 U18931 ( .A1(n15680), .A2(n19802), .B1(n15679), .B2(n19833), .ZN(
        n15681) );
  OAI211_X1 U18932 ( .C1(n15683), .C2(n19818), .A(n15682), .B(n15681), .ZN(
        P1_U2816) );
  INV_X1 U18933 ( .A(n15684), .ZN(n15688) );
  OAI21_X1 U18934 ( .B1(n15686), .B2(n15685), .A(n20633), .ZN(n15687) );
  AOI22_X1 U18935 ( .A1(n15688), .A2(n15687), .B1(n19832), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n15694) );
  OAI22_X1 U18936 ( .A1(n15690), .A2(n15779), .B1(n15689), .B2(n15773), .ZN(
        n15691) );
  AOI21_X1 U18937 ( .B1(n15692), .B2(n19837), .A(n15691), .ZN(n15693) );
  OAI211_X1 U18938 ( .C1(n15695), .C2(n19813), .A(n15694), .B(n15693), .ZN(
        P1_U2817) );
  OAI21_X1 U18939 ( .B1(n19830), .B2(n15707), .A(n19790), .ZN(n15717) );
  NAND2_X1 U18940 ( .A1(n19831), .A2(n20839), .ZN(n15706) );
  INV_X1 U18941 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20635) );
  AOI21_X1 U18942 ( .B1(n15717), .B2(n15706), .A(n20635), .ZN(n15702) );
  NAND2_X1 U18943 ( .A1(n19831), .A2(n15696), .ZN(n15697) );
  NOR2_X1 U18944 ( .A1(n15697), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15701) );
  INV_X1 U18945 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15699) );
  OAI22_X1 U18946 ( .A1(n19813), .A2(n15699), .B1(n15770), .B2(n15698), .ZN(
        n15700) );
  NOR3_X1 U18947 ( .A1(n15702), .A2(n15701), .A3(n15700), .ZN(n15705) );
  INV_X1 U18948 ( .A(n15703), .ZN(n15876) );
  AOI22_X1 U18949 ( .A1(n15813), .A2(n19802), .B1(n19833), .B2(n15876), .ZN(
        n15704) );
  OAI211_X1 U18950 ( .C1(n15816), .C2(n19818), .A(n15705), .B(n15704), .ZN(
        P1_U2818) );
  OAI22_X1 U18951 ( .A1(n15717), .A2(n20839), .B1(n15707), .B2(n15706), .ZN(
        n15708) );
  AOI21_X1 U18952 ( .B1(n19832), .B2(P1_EBX_REG_21__SCAN_IN), .A(n15708), .ZN(
        n15714) );
  OAI22_X1 U18953 ( .A1(n15710), .A2(n15779), .B1(n15709), .B2(n15773), .ZN(
        n15711) );
  AOI21_X1 U18954 ( .B1(n15712), .B2(n19837), .A(n15711), .ZN(n15713) );
  OAI211_X1 U18955 ( .C1(n15715), .C2(n19813), .A(n15714), .B(n15713), .ZN(
        P1_U2819) );
  AOI21_X1 U18956 ( .B1(n15716), .B2(n15725), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15718) );
  OAI22_X1 U18957 ( .A1(n15718), .A2(n15717), .B1(n20822), .B2(n15770), .ZN(
        n15719) );
  AOI21_X1 U18958 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19838), .A(
        n15719), .ZN(n15724) );
  NOR2_X1 U18959 ( .A1(n14314), .A2(n15720), .ZN(n15721) );
  OR2_X1 U18960 ( .A1(n14364), .A2(n15721), .ZN(n15818) );
  OAI22_X1 U18961 ( .A1(n15818), .A2(n15779), .B1(n15773), .B2(n15793), .ZN(
        n15722) );
  INV_X1 U18962 ( .A(n15722), .ZN(n15723) );
  OAI211_X1 U18963 ( .C1(n15817), .C2(n19818), .A(n15724), .B(n15723), .ZN(
        P1_U2820) );
  AOI22_X1 U18964 ( .A1(n15725), .A2(n20628), .B1(n19832), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n15726) );
  OAI21_X1 U18965 ( .B1(n20628), .B2(n15739), .A(n15726), .ZN(n15727) );
  AOI211_X1 U18966 ( .C1(n19838), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19977), .B(n15727), .ZN(n15730) );
  OAI22_X1 U18967 ( .A1(n15827), .A2(n15779), .B1(n15773), .B2(n15889), .ZN(
        n15728) );
  INV_X1 U18968 ( .A(n15728), .ZN(n15729) );
  OAI211_X1 U18969 ( .C1(n15831), .C2(n19818), .A(n15730), .B(n15729), .ZN(
        P1_U2822) );
  INV_X1 U18970 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20623) );
  NAND2_X1 U18971 ( .A1(n15744), .A2(n15785), .ZN(n15746) );
  NOR2_X1 U18972 ( .A1(n20623), .A2(n15746), .ZN(n15741) );
  AOI21_X1 U18973 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n15741), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n15740) );
  OAI22_X1 U18974 ( .A1(n19813), .A2(n14543), .B1(n15731), .B2(n15770), .ZN(
        n15732) );
  AOI211_X1 U18975 ( .C1(n19837), .C2(n15733), .A(n19977), .B(n15732), .ZN(
        n15738) );
  INV_X1 U18976 ( .A(n15734), .ZN(n15735) );
  AOI22_X1 U18977 ( .A1(n15736), .A2(n19802), .B1(n15735), .B2(n19833), .ZN(
        n15737) );
  OAI211_X1 U18978 ( .C1(n15740), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        P1_U2823) );
  INV_X1 U18979 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20625) );
  AOI22_X1 U18980 ( .A1(n15741), .A2(n20625), .B1(n19832), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n15742) );
  OAI21_X1 U18981 ( .B1(n15841), .B2(n19818), .A(n15742), .ZN(n15743) );
  AOI211_X1 U18982 ( .C1(n19838), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19977), .B(n15743), .ZN(n15749) );
  AOI22_X1 U18983 ( .A1(n15838), .A2(n19802), .B1(n19833), .B2(n15898), .ZN(
        n15748) );
  AOI21_X1 U18984 ( .B1(n15745), .B2(n15744), .A(n19793), .ZN(n15761) );
  NOR2_X1 U18985 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15746), .ZN(n15751) );
  OAI21_X1 U18986 ( .B1(n15761), .B2(n15751), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15747) );
  NAND3_X1 U18987 ( .A1(n15749), .A2(n15748), .A3(n15747), .ZN(P1_U2824) );
  AOI21_X1 U18988 ( .B1(n19832), .B2(P1_EBX_REG_15__SCAN_IN), .A(n19977), .ZN(
        n15750) );
  OAI21_X1 U18989 ( .B1(n19813), .B2(n11864), .A(n15750), .ZN(n15752) );
  AOI211_X1 U18990 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15761), .A(n15752), 
        .B(n15751), .ZN(n15753) );
  OAI21_X1 U18991 ( .B1(n15754), .B2(n15779), .A(n15753), .ZN(n15755) );
  AOI21_X1 U18992 ( .B1(n15756), .B2(n19837), .A(n15755), .ZN(n15757) );
  OAI21_X1 U18993 ( .B1(n15773), .B2(n15758), .A(n15757), .ZN(P1_U2825) );
  INV_X1 U18994 ( .A(n15759), .ZN(n15760) );
  AOI22_X1 U18995 ( .A1(n15760), .A2(n19833), .B1(n19832), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n15766) );
  AOI21_X1 U18996 ( .B1(n19838), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n19977), .ZN(n15765) );
  AOI22_X1 U18997 ( .A1(n15843), .A2(n19802), .B1(n19837), .B2(n15842), .ZN(
        n15764) );
  OAI221_X1 U18998 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n15762), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(n15785), .A(n15761), .ZN(n15763) );
  NAND4_X1 U18999 ( .A1(n15766), .A2(n15765), .A3(n15764), .A4(n15763), .ZN(
        P1_U2826) );
  AOI21_X1 U19000 ( .B1(n20619), .B2(n15768), .A(n15767), .ZN(n15776) );
  NOR2_X1 U19001 ( .A1(n15770), .A2(n15769), .ZN(n15771) );
  AOI211_X1 U19002 ( .C1(n19838), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n19977), .B(n15771), .ZN(n15772) );
  OAI21_X1 U19003 ( .B1(n15774), .B2(n15773), .A(n15772), .ZN(n15775) );
  AOI211_X1 U19004 ( .C1(n19837), .C2(n15848), .A(n15776), .B(n15775), .ZN(
        n15777) );
  OAI21_X1 U19005 ( .B1(n15779), .B2(n15778), .A(n15777), .ZN(P1_U2828) );
  INV_X1 U19006 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15783) );
  XNOR2_X1 U19007 ( .A(n15781), .B(n15780), .ZN(n15903) );
  AOI22_X1 U19008 ( .A1(n15903), .A2(n19833), .B1(n19832), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15782) );
  OAI211_X1 U19009 ( .C1(n19813), .C2(n15783), .A(n15782), .B(n19964), .ZN(
        n15784) );
  AOI221_X1 U19010 ( .B1(n15786), .B2(P1_REIP_REG_11__SCAN_IN), .C1(n15785), 
        .C2(n20616), .A(n15784), .ZN(n15788) );
  NAND2_X1 U19011 ( .A1(n19802), .A2(n15856), .ZN(n15787) );
  OAI211_X1 U19012 ( .C1(n19818), .C2(n15859), .A(n15788), .B(n15787), .ZN(
        P1_U2829) );
  NOR2_X1 U19013 ( .A1(n15789), .A2(n14383), .ZN(n15790) );
  AOI21_X1 U19014 ( .B1(n15798), .B2(n19850), .A(n15790), .ZN(n15791) );
  OAI21_X1 U19015 ( .B1(n19854), .B2(n15792), .A(n15791), .ZN(P1_U2846) );
  OAI22_X1 U19016 ( .A1(n15818), .A2(n14394), .B1(n15793), .B2(n14383), .ZN(
        n15794) );
  INV_X1 U19017 ( .A(n15794), .ZN(n15795) );
  OAI21_X1 U19018 ( .B1(n19854), .B2(n20822), .A(n15795), .ZN(P1_U2852) );
  AOI22_X1 U19019 ( .A1(n15856), .A2(n19850), .B1(n19849), .B2(n15903), .ZN(
        n15796) );
  OAI21_X1 U19020 ( .B1(n19854), .B2(n15797), .A(n15796), .ZN(P1_U2861) );
  AOI22_X1 U19021 ( .A1(n15803), .A2(n19908), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n15801), .ZN(n15800) );
  AOI22_X1 U19022 ( .A1(n15798), .A2(n15805), .B1(n15804), .B2(DATAI_26_), 
        .ZN(n15799) );
  OAI211_X1 U19023 ( .C1(n15809), .C2(n14917), .A(n15800), .B(n15799), .ZN(
        P1_U2878) );
  INV_X1 U19024 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16231) );
  INV_X1 U19025 ( .A(n20037), .ZN(n15802) );
  AOI22_X1 U19026 ( .A1(n15803), .A2(n15802), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n15801), .ZN(n15808) );
  INV_X1 U19027 ( .A(n15818), .ZN(n15806) );
  AOI22_X1 U19028 ( .A1(n15806), .A2(n15805), .B1(n15804), .B2(DATAI_20_), 
        .ZN(n15807) );
  OAI211_X1 U19029 ( .C1(n15809), .C2(n16231), .A(n15808), .B(n15807), .ZN(
        P1_U2884) );
  AOI22_X1 U19030 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15815) );
  NAND2_X1 U19031 ( .A1(n15811), .A2(n15810), .ZN(n15812) );
  XNOR2_X1 U19032 ( .A(n15812), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15875) );
  AOI22_X1 U19033 ( .A1(n15813), .A2(n19934), .B1(n19935), .B2(n15875), .ZN(
        n15814) );
  OAI211_X1 U19034 ( .C1(n19942), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        P1_U2977) );
  INV_X1 U19035 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15824) );
  OAI22_X1 U19036 ( .A1(n15818), .A2(n20006), .B1(n15817), .B2(n19942), .ZN(
        n15819) );
  AOI21_X1 U19037 ( .B1(n15820), .B2(n19935), .A(n15819), .ZN(n15822) );
  OAI211_X1 U19038 ( .C1(n15824), .C2(n15823), .A(n15822), .B(n15821), .ZN(
        P1_U2979) );
  AOI22_X1 U19039 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n15830) );
  OAI21_X1 U19040 ( .B1(n15826), .B2(n15825), .A(n14526), .ZN(n15883) );
  OAI22_X1 U19041 ( .A1(n15883), .A2(n19943), .B1(n15827), .B2(n20006), .ZN(
        n15828) );
  INV_X1 U19042 ( .A(n15828), .ZN(n15829) );
  OAI211_X1 U19043 ( .C1(n19942), .C2(n15831), .A(n15830), .B(n15829), .ZN(
        P1_U2981) );
  AOI22_X1 U19044 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15840) );
  INV_X1 U19045 ( .A(n15832), .ZN(n15837) );
  AOI21_X1 U19046 ( .B1(n15835), .B2(n15834), .A(n15833), .ZN(n15836) );
  NOR2_X1 U19047 ( .A1(n15837), .A2(n15836), .ZN(n15899) );
  AOI22_X1 U19048 ( .A1(n15899), .A2(n19935), .B1(n19934), .B2(n15838), .ZN(
        n15839) );
  OAI211_X1 U19049 ( .C1(n19942), .C2(n15841), .A(n15840), .B(n15839), .ZN(
        P1_U2983) );
  AOI22_X1 U19050 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15845) );
  AOI22_X1 U19051 ( .A1(n15843), .A2(n19934), .B1(n15849), .B2(n15842), .ZN(
        n15844) );
  OAI211_X1 U19052 ( .C1(n15846), .C2(n19943), .A(n15845), .B(n15844), .ZN(
        P1_U2985) );
  AOI22_X1 U19053 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15851) );
  AOI22_X1 U19054 ( .A1(n15849), .A2(n15848), .B1(n19934), .B2(n15847), .ZN(
        n15850) );
  OAI211_X1 U19055 ( .C1(n15852), .C2(n19943), .A(n15851), .B(n15850), .ZN(
        P1_U2987) );
  AOI22_X1 U19056 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15858) );
  NOR3_X1 U19057 ( .A1(n14534), .A2(n9634), .A3(n15917), .ZN(n15854) );
  NOR2_X1 U19058 ( .A1(n15854), .A2(n15853), .ZN(n15855) );
  XOR2_X1 U19059 ( .A(n12643), .B(n15855), .Z(n15905) );
  AOI22_X1 U19060 ( .A1(n19935), .A2(n15905), .B1(n19934), .B2(n15856), .ZN(
        n15857) );
  OAI211_X1 U19061 ( .C1(n19942), .C2(n15859), .A(n15858), .B(n15857), .ZN(
        P1_U2988) );
  AOI22_X1 U19062 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15863) );
  XNOR2_X1 U19063 ( .A(n15860), .B(n15861), .ZN(n15929) );
  AOI22_X1 U19064 ( .A1(n15929), .A2(n19935), .B1(n19934), .B2(n19794), .ZN(
        n15862) );
  OAI211_X1 U19065 ( .C1(n19942), .C2(n19797), .A(n15863), .B(n15862), .ZN(
        P1_U2992) );
  AOI22_X1 U19066 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15869) );
  NAND2_X1 U19067 ( .A1(n15865), .A2(n15864), .ZN(n15866) );
  NAND2_X1 U19068 ( .A1(n15867), .A2(n15866), .ZN(n15938) );
  AOI22_X1 U19069 ( .A1(n15938), .A2(n19935), .B1(n19934), .B2(n19851), .ZN(
        n15868) );
  OAI211_X1 U19070 ( .C1(n19942), .C2(n19805), .A(n15869), .B(n15868), .ZN(
        P1_U2993) );
  AOI22_X1 U19071 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15873) );
  INV_X1 U19072 ( .A(n15870), .ZN(n15871) );
  AOI22_X1 U19073 ( .A1(n15871), .A2(n19935), .B1(n19934), .B2(n19816), .ZN(
        n15872) );
  OAI211_X1 U19074 ( .C1(n19942), .C2(n19819), .A(n15873), .B(n15872), .ZN(
        P1_U2994) );
  AOI22_X1 U19075 ( .A1(n15875), .A2(n19957), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15874), .ZN(n15882) );
  NAND2_X1 U19076 ( .A1(n19977), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15881) );
  NAND2_X1 U19077 ( .A1(n15876), .A2(n19979), .ZN(n15880) );
  OAI211_X1 U19078 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15878), .B(n15877), .ZN(
        n15879) );
  NAND4_X1 U19079 ( .A1(n15882), .A2(n15881), .A3(n15880), .A4(n15879), .ZN(
        P1_U3009) );
  INV_X1 U19080 ( .A(n15883), .ZN(n15888) );
  NOR3_X1 U19081 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15884), .A3(
        n15894), .ZN(n15886) );
  NOR2_X1 U19082 ( .A1(n19964), .A2(n20628), .ZN(n15885) );
  OR2_X1 U19083 ( .A1(n15886), .A2(n15885), .ZN(n15887) );
  AOI21_X1 U19084 ( .B1(n15888), .B2(n19957), .A(n15887), .ZN(n15893) );
  INV_X1 U19085 ( .A(n15889), .ZN(n15891) );
  AOI22_X1 U19086 ( .A1(n15891), .A2(n19979), .B1(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15890), .ZN(n15892) );
  NAND2_X1 U19087 ( .A1(n15893), .A2(n15892), .ZN(P1_U3013) );
  AOI21_X1 U19088 ( .B1(n15895), .B2(n9765), .A(n15894), .ZN(n15897) );
  AOI22_X1 U19089 ( .A1(n19977), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n15897), 
        .B2(n15896), .ZN(n15901) );
  AOI22_X1 U19090 ( .A1(n15899), .A2(n19957), .B1(n19979), .B2(n15898), .ZN(
        n15900) );
  OAI211_X1 U19091 ( .C1(n15902), .C2(n9765), .A(n15901), .B(n15900), .ZN(
        P1_U3015) );
  AOI22_X1 U19092 ( .A1(n15903), .A2(n19979), .B1(n19977), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15907) );
  AOI22_X1 U19093 ( .A1(n15905), .A2(n19957), .B1(n15937), .B2(n15904), .ZN(
        n15906) );
  OAI211_X1 U19094 ( .C1(n15908), .C2(n12643), .A(n15907), .B(n15906), .ZN(
        P1_U3020) );
  AOI21_X1 U19095 ( .B1(n15910), .B2(n19979), .A(n15909), .ZN(n15916) );
  AOI22_X1 U19096 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n15911), .B2(n15917), .ZN(
        n15913) );
  AOI22_X1 U19097 ( .A1(n15914), .A2(n19957), .B1(n15913), .B2(n15912), .ZN(
        n15915) );
  OAI211_X1 U19098 ( .C1(n15918), .C2(n15917), .A(n15916), .B(n15915), .ZN(
        P1_U3021) );
  OAI21_X1 U19099 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15919), .ZN(n15926) );
  AOI21_X1 U19100 ( .B1(n15921), .B2(n19979), .A(n15920), .ZN(n15925) );
  OAI21_X1 U19101 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15922), .A(
        n15942), .ZN(n15928) );
  AOI22_X1 U19102 ( .A1(n15923), .A2(n19957), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n15928), .ZN(n15924) );
  OAI211_X1 U19103 ( .C1(n15932), .C2(n15926), .A(n15925), .B(n15924), .ZN(
        P1_U3023) );
  INV_X1 U19104 ( .A(n15927), .ZN(n19785) );
  AOI22_X1 U19105 ( .A1(n19785), .A2(n19979), .B1(n19977), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n15931) );
  AOI22_X1 U19106 ( .A1(n15929), .A2(n19957), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15928), .ZN(n15930) );
  OAI211_X1 U19107 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n15932), .A(
        n15931), .B(n15930), .ZN(P1_U3024) );
  OR2_X1 U19108 ( .A1(n15934), .A2(n15933), .ZN(n15935) );
  AND2_X1 U19109 ( .A1(n15936), .A2(n15935), .ZN(n19848) );
  AOI22_X1 U19110 ( .A1(n19979), .A2(n19848), .B1(n19977), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15940) );
  AOI22_X1 U19111 ( .A1(n15938), .A2(n19957), .B1(n15937), .B2(n15941), .ZN(
        n15939) );
  OAI211_X1 U19112 ( .C1(n15942), .C2(n15941), .A(n15940), .B(n15939), .ZN(
        P1_U3025) );
  NAND4_X1 U19113 ( .A1(n19821), .A2(n15945), .A3(n15944), .A4(n15943), .ZN(
        n15946) );
  OAI21_X1 U19114 ( .B1(n15948), .B2(n15947), .A(n15946), .ZN(P1_U3468) );
  NAND4_X1 U19115 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20700), .A4(n20708), .ZN(n15949) );
  OAI21_X1 U19116 ( .B1(n15950), .B2(n20771), .A(n15949), .ZN(n20581) );
  OAI21_X1 U19117 ( .B1(n15952), .B2(n20581), .A(n15951), .ZN(n15953) );
  OAI211_X1 U19118 ( .C1(n20703), .C2(n20708), .A(n15954), .B(n15953), .ZN(
        n15955) );
  AOI21_X1 U19119 ( .B1(n13792), .B2(n15956), .A(n15955), .ZN(P1_U3162) );
  INV_X1 U19120 ( .A(n15956), .ZN(n20584) );
  OAI21_X1 U19121 ( .B1(n20584), .B2(n20780), .A(n15957), .ZN(P1_U3466) );
  AOI22_X1 U19122 ( .A1(n15958), .A2(n18865), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n18867), .ZN(n15964) );
  AOI22_X1 U19123 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n15959), .ZN(n15963) );
  AOI22_X1 U19124 ( .A1(n16001), .A2(n18840), .B1(n18863), .B2(n18904), .ZN(
        n15962) );
  NAND3_X1 U19125 ( .A1(n18827), .A2(n15960), .A3(n13945), .ZN(n15961) );
  NAND4_X1 U19126 ( .A1(n15964), .A2(n15963), .A3(n15962), .A4(n15961), .ZN(
        P2_U2824) );
  OAI22_X1 U19127 ( .A1(n15966), .A2(n18870), .B1(n15965), .B2(n18836), .ZN(
        n15967) );
  INV_X1 U19128 ( .A(n15967), .ZN(n15976) );
  AOI211_X1 U19129 ( .C1(n15970), .C2(n15969), .A(n15968), .B(n18877), .ZN(
        n15974) );
  AOI22_X1 U19130 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n18867), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n18866), .ZN(n15971) );
  OAI21_X1 U19131 ( .B1(n15972), .B2(n18852), .A(n15971), .ZN(n15973) );
  AOI211_X1 U19132 ( .C1(n18874), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15974), .B(n15973), .ZN(n15975) );
  NAND2_X1 U19133 ( .A1(n15976), .A2(n15975), .ZN(P2_U2827) );
  AOI22_X1 U19134 ( .A1(n15977), .A2(n18865), .B1(P2_REIP_REG_26__SCAN_IN), 
        .B2(n18867), .ZN(n15988) );
  AOI22_X1 U19135 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n18866), .ZN(n15987) );
  INV_X1 U19136 ( .A(n15978), .ZN(n15979) );
  OAI22_X1 U19137 ( .A1(n15980), .A2(n18870), .B1(n15979), .B2(n18836), .ZN(
        n15981) );
  INV_X1 U19138 ( .A(n15981), .ZN(n15986) );
  AOI21_X1 U19139 ( .B1(n15983), .B2(n9701), .A(n15982), .ZN(n15984) );
  NAND2_X1 U19140 ( .A1(n18827), .A2(n15984), .ZN(n15985) );
  NAND4_X1 U19141 ( .A1(n15988), .A2(n15987), .A3(n15986), .A4(n15985), .ZN(
        P2_U2829) );
  INV_X1 U19142 ( .A(n15989), .ZN(n15990) );
  AOI22_X1 U19143 ( .A1(n15991), .A2(n18840), .B1(n15990), .B2(n18863), .ZN(
        n16000) );
  AOI211_X1 U19144 ( .C1(n15994), .C2(n15993), .A(n15992), .B(n18877), .ZN(
        n15998) );
  AOI22_X1 U19145 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n18867), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n18866), .ZN(n15995) );
  OAI21_X1 U19146 ( .B1(n15996), .B2(n18852), .A(n15995), .ZN(n15997) );
  AOI211_X1 U19147 ( .C1(n18874), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15998), .B(n15997), .ZN(n15999) );
  NAND2_X1 U19148 ( .A1(n16000), .A2(n15999), .ZN(P2_U2831) );
  OAI22_X1 U19149 ( .A1(n18888), .A2(n16001), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n18903), .ZN(n16002) );
  INV_X1 U19150 ( .A(n16002), .ZN(P2_U2856) );
  INV_X1 U19151 ( .A(n16003), .ZN(n16004) );
  AOI22_X1 U19152 ( .A1(n16004), .A2(n18899), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n18888), .ZN(n16005) );
  OAI21_X1 U19153 ( .B1(n18888), .B2(n16036), .A(n16005), .ZN(P2_U2862) );
  AOI22_X1 U19154 ( .A1(n16007), .A2(n18899), .B1(n18903), .B2(n16006), .ZN(
        n16008) );
  OAI21_X1 U19155 ( .B1(n18903), .B2(n16009), .A(n16008), .ZN(P2_U2865) );
  NOR2_X1 U19156 ( .A1(n14879), .A2(n16010), .ZN(n16011) );
  OR2_X1 U19157 ( .A1(n14872), .A2(n16011), .ZN(n16019) );
  OAI22_X1 U19158 ( .A1(n16019), .A2(n18893), .B1(n18888), .B2(n18671), .ZN(
        n16012) );
  INV_X1 U19159 ( .A(n16012), .ZN(n16013) );
  OAI21_X1 U19160 ( .B1(n18903), .B2(n11159), .A(n16013), .ZN(P2_U2867) );
  AOI21_X1 U19161 ( .B1(n16014), .B2(n13992), .A(n10014), .ZN(n16025) );
  AOI22_X1 U19162 ( .A1(n16025), .A2(n18899), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n18888), .ZN(n16015) );
  OAI21_X1 U19163 ( .B1(n18888), .B2(n16016), .A(n16015), .ZN(P2_U2869) );
  INV_X1 U19164 ( .A(n16017), .ZN(n18907) );
  AOI22_X1 U19165 ( .A1(n18907), .A2(n19057), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n18921), .ZN(n16023) );
  AOI22_X1 U19166 ( .A1(n18909), .A2(BUF1_REG_20__SCAN_IN), .B1(n18908), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16022) );
  OAI22_X1 U19167 ( .A1(n16019), .A2(n18930), .B1(n16018), .B2(n18670), .ZN(
        n16020) );
  INV_X1 U19168 ( .A(n16020), .ZN(n16021) );
  NAND3_X1 U19169 ( .A1(n16023), .A2(n16022), .A3(n16021), .ZN(P2_U2899) );
  AOI22_X1 U19170 ( .A1(n18907), .A2(n19047), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n18921), .ZN(n16028) );
  AOI22_X1 U19171 ( .A1(n18909), .A2(BUF1_REG_18__SCAN_IN), .B1(n18908), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16027) );
  AOI22_X1 U19172 ( .A1(n18696), .A2(n18912), .B1(n16025), .B2(n16024), .ZN(
        n16026) );
  NAND3_X1 U19173 ( .A1(n16028), .A2(n16027), .A3(n16026), .ZN(P2_U2901) );
  OAI22_X1 U19174 ( .A1(n14792), .A2(n18772), .B1(n16029), .B2(n16117), .ZN(
        n16030) );
  AOI21_X1 U19175 ( .B1(n16108), .B2(n16031), .A(n16030), .ZN(n16035) );
  AOI22_X1 U19176 ( .A1(n16033), .A2(n16112), .B1(n16032), .B2(n16113), .ZN(
        n16034) );
  OAI211_X1 U19177 ( .C1(n19026), .C2(n16036), .A(n16035), .B(n16034), .ZN(
        P2_U2989) );
  NOR2_X1 U19178 ( .A1(n16037), .A2(n16117), .ZN(n16038) );
  AOI211_X1 U19179 ( .C1(n16108), .C2(n16040), .A(n16039), .B(n16038), .ZN(
        n16045) );
  OAI211_X1 U19180 ( .C1(n19026), .C2(n16046), .A(n16045), .B(n16044), .ZN(
        P2_U2993) );
  OAI22_X1 U19181 ( .A1(n20750), .A2(n16117), .B1(n20834), .B2(n19017), .ZN(
        n16047) );
  AOI21_X1 U19182 ( .B1(n16108), .B2(n18679), .A(n16047), .ZN(n16051) );
  AOI22_X1 U19183 ( .A1(n16049), .A2(n16112), .B1(n16113), .B2(n16048), .ZN(
        n16050) );
  OAI211_X1 U19184 ( .C1(n19026), .C2(n18684), .A(n16051), .B(n16050), .ZN(
        P2_U2995) );
  AOI22_X1 U19185 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18977), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18839), .ZN(n16056) );
  OAI22_X1 U19186 ( .A1(n16053), .A2(n18981), .B1(n18980), .B2(n16052), .ZN(
        n16054) );
  AOI21_X1 U19187 ( .B1(n18985), .B2(n18695), .A(n16054), .ZN(n16055) );
  OAI211_X1 U19188 ( .C1(n18989), .C2(n18690), .A(n16056), .B(n16055), .ZN(
        P2_U2996) );
  AOI22_X1 U19189 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n18839), .B1(n16108), 
        .B2(n18729), .ZN(n16062) );
  INV_X1 U19190 ( .A(n16057), .ZN(n16059) );
  AOI222_X1 U19191 ( .A1(n16060), .A2(n16112), .B1(n16113), .B2(n16059), .C1(
        n18985), .C2(n16058), .ZN(n16061) );
  OAI211_X1 U19192 ( .C1(n18736), .C2(n16117), .A(n16062), .B(n16061), .ZN(
        P2_U2999) );
  AOI22_X1 U19193 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18977), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18839), .ZN(n16073) );
  AOI21_X1 U19194 ( .B1(n16065), .B2(n16064), .A(n16063), .ZN(n16124) );
  INV_X1 U19195 ( .A(n16066), .ZN(n16067) );
  AOI21_X1 U19196 ( .B1(n16069), .B2(n16068), .A(n16067), .ZN(n16125) );
  INV_X1 U19197 ( .A(n16125), .ZN(n16070) );
  OAI22_X1 U19198 ( .A1(n16124), .A2(n18981), .B1(n18980), .B2(n16070), .ZN(
        n16071) );
  AOI21_X1 U19199 ( .B1(n18985), .B2(n18742), .A(n16071), .ZN(n16072) );
  OAI211_X1 U19200 ( .C1(n18989), .C2(n18738), .A(n16073), .B(n16072), .ZN(
        P2_U3000) );
  AOI22_X1 U19201 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n18839), .B1(n16108), 
        .B2(n18755), .ZN(n16078) );
  INV_X1 U19202 ( .A(n16074), .ZN(n18754) );
  AOI222_X1 U19203 ( .A1(n16076), .A2(n16112), .B1(n16075), .B2(n16113), .C1(
        n18985), .C2(n18754), .ZN(n16077) );
  OAI211_X1 U19204 ( .C1(n16079), .C2(n16117), .A(n16078), .B(n16077), .ZN(
        P2_U3001) );
  AOI22_X1 U19205 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18977), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18839), .ZN(n16086) );
  INV_X1 U19206 ( .A(n16080), .ZN(n16082) );
  OAI22_X1 U19207 ( .A1(n16082), .A2(n18980), .B1(n16081), .B2(n18981), .ZN(
        n16083) );
  AOI21_X1 U19208 ( .B1(n18985), .B2(n16084), .A(n16083), .ZN(n16085) );
  OAI211_X1 U19209 ( .C1(n18989), .C2(n16087), .A(n16086), .B(n16085), .ZN(
        P2_U3002) );
  AOI22_X1 U19210 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18839), .B1(n16108), 
        .B2(n18764), .ZN(n16094) );
  OR2_X1 U19211 ( .A1(n16088), .A2(n18980), .ZN(n16091) );
  NAND2_X1 U19212 ( .A1(n16089), .A2(n16112), .ZN(n16090) );
  OAI211_X1 U19213 ( .C1(n19026), .C2(n18765), .A(n16091), .B(n16090), .ZN(
        n16092) );
  INV_X1 U19214 ( .A(n16092), .ZN(n16093) );
  OAI211_X1 U19215 ( .C1(n16095), .C2(n16117), .A(n16094), .B(n16093), .ZN(
        P2_U3003) );
  AOI22_X1 U19216 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18977), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18839), .ZN(n16100) );
  OAI22_X1 U19217 ( .A1(n16097), .A2(n18980), .B1(n16096), .B2(n18981), .ZN(
        n16098) );
  AOI21_X1 U19218 ( .B1(n18985), .B2(n18897), .A(n16098), .ZN(n16099) );
  OAI211_X1 U19219 ( .C1(n18989), .C2(n18777), .A(n16100), .B(n16099), .ZN(
        P2_U3004) );
  AOI22_X1 U19220 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18839), .B1(n16108), 
        .B2(n18787), .ZN(n16107) );
  NOR2_X1 U19221 ( .A1(n16101), .A2(n18980), .ZN(n16105) );
  OAI22_X1 U19222 ( .A1(n16102), .A2(n18981), .B1(n19026), .B2(n18788), .ZN(
        n16103) );
  AOI21_X1 U19223 ( .B1(n16105), .B2(n16104), .A(n16103), .ZN(n16106) );
  OAI211_X1 U19224 ( .C1(n18794), .C2(n16117), .A(n16107), .B(n16106), .ZN(
        P2_U3005) );
  AOI22_X1 U19225 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18839), .B1(n16108), 
        .B2(n18825), .ZN(n16116) );
  INV_X1 U19226 ( .A(n16109), .ZN(n16114) );
  INV_X1 U19227 ( .A(n16110), .ZN(n16111) );
  AOI222_X1 U19228 ( .A1(n16114), .A2(n16113), .B1(n18985), .B2(n18826), .C1(
        n16112), .C2(n16111), .ZN(n16115) );
  OAI211_X1 U19229 ( .C1(n20762), .C2(n16117), .A(n16116), .B(n16115), .ZN(
        P2_U3009) );
  AOI21_X1 U19230 ( .B1(n16119), .B2(n16118), .A(n13810), .ZN(n18917) );
  INV_X1 U19231 ( .A(n16120), .ZN(n16121) );
  NOR3_X1 U19232 ( .A1(n16122), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16121), .ZN(n16123) );
  AOI21_X1 U19233 ( .B1(n18917), .B2(n18993), .A(n16123), .ZN(n16132) );
  INV_X1 U19234 ( .A(n16124), .ZN(n16126) );
  AOI222_X1 U19235 ( .A1(n16126), .A2(n18992), .B1(n19008), .B2(n18742), .C1(
        n16152), .C2(n16125), .ZN(n16131) );
  NAND2_X1 U19236 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n18839), .ZN(n16130) );
  OAI21_X1 U19237 ( .B1(n16128), .B2(n16127), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16129) );
  NAND4_X1 U19238 ( .A1(n16132), .A2(n16131), .A3(n16130), .A4(n16129), .ZN(
        P2_U3032) );
  NAND2_X1 U19239 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n18839), .ZN(n16133) );
  OAI221_X1 U19240 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16135), .C1(
        n9839), .C2(n16134), .A(n16133), .ZN(n16140) );
  OAI22_X1 U19241 ( .A1(n16138), .A2(n16146), .B1(n16137), .B2(n16136), .ZN(
        n16139) );
  AOI211_X1 U19242 ( .C1(n16141), .C2(n18992), .A(n16140), .B(n16139), .ZN(
        n16142) );
  OAI21_X1 U19243 ( .B1(n18996), .B2(n16143), .A(n16142), .ZN(P2_U3039) );
  NAND2_X1 U19244 ( .A1(n19008), .A2(n13951), .ZN(n16145) );
  OAI211_X1 U19245 ( .C1(n16146), .C2(n19701), .A(n16145), .B(n16144), .ZN(
        n16150) );
  NOR2_X1 U19246 ( .A1(n16148), .A2(n16147), .ZN(n16149) );
  AOI211_X1 U19247 ( .C1(n16152), .C2(n16151), .A(n16150), .B(n16149), .ZN(
        n16153) );
  OAI221_X1 U19248 ( .B1(n16156), .B2(n16155), .C1(n16156), .C2(n16154), .A(
        n16153), .ZN(P2_U3043) );
  AOI21_X1 U19249 ( .B1(n16159), .B2(n16158), .A(n16157), .ZN(n16166) );
  INV_X1 U19250 ( .A(n16161), .ZN(n16160) );
  OAI21_X1 U19251 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19747), .A(n16160), 
        .ZN(n19611) );
  NAND2_X1 U19252 ( .A1(n16161), .A2(n19618), .ZN(n19615) );
  OAI21_X1 U19253 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16163), .A(n16162), 
        .ZN(n16164) );
  AOI22_X1 U19254 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19611), .B1(n19615), 
        .B2(n16164), .ZN(n16165) );
  OAI211_X1 U19255 ( .C1(n16168), .C2(n16167), .A(n16166), .B(n16165), .ZN(
        P2_U3176) );
  NAND2_X1 U19256 ( .A1(n9632), .A2(n16169), .ZN(n16186) );
  NAND2_X1 U19257 ( .A1(n17529), .A2(n16170), .ZN(n16188) );
  AOI21_X1 U19258 ( .B1(n16186), .B2(n16188), .A(n16177), .ZN(n16176) );
  INV_X1 U19259 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16173) );
  OAI221_X1 U19260 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16174), .C1(
        n16173), .C2(n16172), .A(n16171), .ZN(n16175) );
  AOI211_X1 U19261 ( .C1(n17475), .C2(n16330), .A(n16176), .B(n16175), .ZN(
        n16180) );
  NOR2_X2 U19262 ( .A1(n17300), .A2(n17422), .ZN(n17328) );
  NAND4_X1 U19263 ( .A1(n16178), .A2(n17268), .A3(n17328), .A4(n16177), .ZN(
        n16179) );
  OAI211_X1 U19264 ( .C1(n16181), .C2(n17470), .A(n16180), .B(n16179), .ZN(
        P3_U2800) );
  INV_X2 U19265 ( .A(n17835), .ZN(n17940) );
  OAI21_X1 U19266 ( .B1(n17991), .B2(n16183), .A(n16182), .ZN(n16184) );
  AOI22_X1 U19267 ( .A1(n17940), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n16185), 
        .B2(n16184), .ZN(n16197) );
  AOI21_X1 U19268 ( .B1(n16187), .B2(n16190), .A(n16186), .ZN(n16192) );
  AOI21_X1 U19269 ( .B1(n16190), .B2(n16189), .A(n16188), .ZN(n16191) );
  AOI211_X1 U19270 ( .C1(n16193), .C2(n17533), .A(n16192), .B(n16191), .ZN(
        n16196) );
  OAI21_X1 U19271 ( .B1(n17475), .B2(n16194), .A(n16343), .ZN(n16195) );
  NAND3_X1 U19272 ( .A1(n16197), .A2(n16196), .A3(n16195), .ZN(P3_U2801) );
  OAI22_X1 U19273 ( .A1(n16200), .A2(n17936), .B1(n16199), .B2(n16198), .ZN(
        n16201) );
  AOI211_X1 U19274 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16203), .A(
        n16202), .B(n16201), .ZN(n16207) );
  AOI22_X1 U19275 ( .A1(n17863), .A2(n16205), .B1(n17947), .B2(n16204), .ZN(
        n16206) );
  OAI211_X1 U19276 ( .C1(n16208), .C2(n17807), .A(n16207), .B(n16206), .ZN(
        P3_U2831) );
  NOR3_X1 U19277 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16210) );
  NOR4_X1 U19278 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16209) );
  INV_X2 U19279 ( .A(n16298), .ZN(U215) );
  NAND4_X1 U19280 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16210), .A3(n16209), .A4(
        U215), .ZN(U213) );
  INV_X1 U19281 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n18937) );
  INV_X2 U19282 ( .A(U214), .ZN(n16261) );
  NOR2_X1 U19283 ( .A1(n16261), .A2(n16211), .ZN(n16251) );
  INV_X1 U19284 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16301) );
  OAI222_X1 U19285 ( .A1(U212), .A2(n18937), .B1(n16263), .B2(n16212), .C1(
        U214), .C2(n16301), .ZN(U216) );
  AOI222_X1 U19286 ( .A1(n16260), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16251), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16261), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n16213) );
  INV_X1 U19287 ( .A(n16213), .ZN(U217) );
  AOI22_X1 U19288 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16260), .ZN(n16214) );
  OAI21_X1 U19289 ( .B1(n14890), .B2(n16263), .A(n16214), .ZN(U218) );
  INV_X1 U19290 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16216) );
  AOI22_X1 U19291 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16260), .ZN(n16215) );
  OAI21_X1 U19292 ( .B1(n16216), .B2(n16263), .A(n16215), .ZN(U219) );
  INV_X1 U19293 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16218) );
  AOI22_X1 U19294 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16260), .ZN(n16217) );
  OAI21_X1 U19295 ( .B1(n16218), .B2(n16263), .A(n16217), .ZN(U220) );
  AOI22_X1 U19296 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16260), .ZN(n16219) );
  OAI21_X1 U19297 ( .B1(n14917), .B2(n16263), .A(n16219), .ZN(U221) );
  INV_X1 U19298 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16221) );
  AOI22_X1 U19299 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16260), .ZN(n16220) );
  OAI21_X1 U19300 ( .B1(n16221), .B2(n16263), .A(n16220), .ZN(U222) );
  INV_X1 U19301 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16223) );
  AOI22_X1 U19302 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16260), .ZN(n16222) );
  OAI21_X1 U19303 ( .B1(n16223), .B2(n16263), .A(n16222), .ZN(U223) );
  INV_X1 U19304 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16225) );
  AOI22_X1 U19305 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16260), .ZN(n16224) );
  OAI21_X1 U19306 ( .B1(n16225), .B2(n16263), .A(n16224), .ZN(U224) );
  INV_X1 U19307 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16227) );
  AOI22_X1 U19308 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16260), .ZN(n16226) );
  OAI21_X1 U19309 ( .B1(n16227), .B2(n16263), .A(n16226), .ZN(U225) );
  INV_X1 U19310 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16229) );
  AOI22_X1 U19311 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16260), .ZN(n16228) );
  OAI21_X1 U19312 ( .B1(n16229), .B2(n16263), .A(n16228), .ZN(U226) );
  AOI22_X1 U19313 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16260), .ZN(n16230) );
  OAI21_X1 U19314 ( .B1(n16231), .B2(n16263), .A(n16230), .ZN(U227) );
  INV_X1 U19315 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16233) );
  AOI22_X1 U19316 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16260), .ZN(n16232) );
  OAI21_X1 U19317 ( .B1(n16233), .B2(n16263), .A(n16232), .ZN(U228) );
  INV_X1 U19318 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16235) );
  AOI22_X1 U19319 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16260), .ZN(n16234) );
  OAI21_X1 U19320 ( .B1(n16235), .B2(n16263), .A(n16234), .ZN(U229) );
  INV_X1 U19321 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16237) );
  AOI22_X1 U19322 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16260), .ZN(n16236) );
  OAI21_X1 U19323 ( .B1(n16237), .B2(n16263), .A(n16236), .ZN(U230) );
  INV_X1 U19324 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16239) );
  AOI22_X1 U19325 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16260), .ZN(n16238) );
  OAI21_X1 U19326 ( .B1(n16239), .B2(n16263), .A(n16238), .ZN(U231) );
  INV_X1 U19327 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n20768) );
  AOI22_X1 U19328 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16251), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16260), .ZN(n16240) );
  OAI21_X1 U19329 ( .B1(n20768), .B2(U214), .A(n16240), .ZN(U232) );
  INV_X1 U19330 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16279) );
  AOI22_X1 U19331 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16251), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16261), .ZN(n16241) );
  OAI21_X1 U19332 ( .B1(n16279), .B2(U212), .A(n16241), .ZN(U233) );
  INV_X1 U19333 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16278) );
  AOI22_X1 U19334 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16251), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16261), .ZN(n16242) );
  OAI21_X1 U19335 ( .B1(n16278), .B2(U212), .A(n16242), .ZN(U234) );
  INV_X1 U19336 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16277) );
  AOI22_X1 U19337 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16251), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16261), .ZN(n16243) );
  OAI21_X1 U19338 ( .B1(n16277), .B2(U212), .A(n16243), .ZN(U235) );
  INV_X1 U19339 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16276) );
  AOI22_X1 U19340 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16251), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16261), .ZN(n16244) );
  OAI21_X1 U19341 ( .B1(n16276), .B2(U212), .A(n16244), .ZN(U236) );
  AOI22_X1 U19342 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16260), .ZN(n16245) );
  OAI21_X1 U19343 ( .B1(n16246), .B2(n16263), .A(n16245), .ZN(U237) );
  INV_X1 U19344 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16274) );
  AOI22_X1 U19345 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16251), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16261), .ZN(n16247) );
  OAI21_X1 U19346 ( .B1(n16274), .B2(U212), .A(n16247), .ZN(U238) );
  INV_X1 U19347 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16273) );
  AOI22_X1 U19348 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n16251), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16261), .ZN(n16248) );
  OAI21_X1 U19349 ( .B1(n16273), .B2(U212), .A(n16248), .ZN(U239) );
  INV_X1 U19350 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16272) );
  AOI22_X1 U19351 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16251), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16261), .ZN(n16249) );
  OAI21_X1 U19352 ( .B1(n16272), .B2(U212), .A(n16249), .ZN(U240) );
  INV_X1 U19353 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16271) );
  AOI22_X1 U19354 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16251), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16261), .ZN(n16250) );
  OAI21_X1 U19355 ( .B1(n16271), .B2(U212), .A(n16250), .ZN(U241) );
  INV_X1 U19356 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16270) );
  AOI22_X1 U19357 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16251), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16261), .ZN(n16252) );
  OAI21_X1 U19358 ( .B1(n16270), .B2(U212), .A(n16252), .ZN(U242) );
  AOI22_X1 U19359 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16260), .ZN(n16253) );
  OAI21_X1 U19360 ( .B1(n16254), .B2(n16263), .A(n16253), .ZN(U243) );
  AOI22_X1 U19361 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16260), .ZN(n16255) );
  OAI21_X1 U19362 ( .B1(n16256), .B2(n16263), .A(n16255), .ZN(U244) );
  AOI22_X1 U19363 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16260), .ZN(n16257) );
  OAI21_X1 U19364 ( .B1(n16258), .B2(n16263), .A(n16257), .ZN(U245) );
  INV_X1 U19365 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20766) );
  AOI22_X1 U19366 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16260), .ZN(n16259) );
  OAI21_X1 U19367 ( .B1(n20766), .B2(n16263), .A(n16259), .ZN(U246) );
  AOI22_X1 U19368 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16261), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16260), .ZN(n16262) );
  OAI21_X1 U19369 ( .B1(n16264), .B2(n16263), .A(n16262), .ZN(U247) );
  INV_X1 U19370 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16265) );
  AOI22_X1 U19371 ( .A1(n16298), .A2(n16265), .B1(n17964), .B2(U215), .ZN(U251) );
  OAI22_X1 U19372 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16298), .ZN(n16266) );
  INV_X1 U19373 ( .A(n16266), .ZN(U252) );
  INV_X1 U19374 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16267) );
  AOI22_X1 U19375 ( .A1(n16298), .A2(n16267), .B1(n17974), .B2(U215), .ZN(U253) );
  INV_X1 U19376 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16268) );
  INV_X1 U19377 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n17978) );
  AOI22_X1 U19378 ( .A1(n16298), .A2(n16268), .B1(n17978), .B2(U215), .ZN(U254) );
  INV_X1 U19379 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16269) );
  AOI22_X1 U19380 ( .A1(n16298), .A2(n16269), .B1(n17982), .B2(U215), .ZN(U255) );
  INV_X1 U19381 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n17987) );
  AOI22_X1 U19382 ( .A1(n16296), .A2(n16270), .B1(n17987), .B2(U215), .ZN(U256) );
  INV_X1 U19383 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n17992) );
  AOI22_X1 U19384 ( .A1(n16298), .A2(n16271), .B1(n17992), .B2(U215), .ZN(U257) );
  INV_X1 U19385 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n17996) );
  AOI22_X1 U19386 ( .A1(n16298), .A2(n16272), .B1(n17996), .B2(U215), .ZN(U258) );
  INV_X1 U19387 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U19388 ( .A1(n16298), .A2(n16273), .B1(n17230), .B2(U215), .ZN(U259) );
  INV_X1 U19389 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U19390 ( .A1(n16296), .A2(n16274), .B1(n17232), .B2(U215), .ZN(U260) );
  INV_X1 U19391 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16275) );
  INV_X1 U19392 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U19393 ( .A1(n16298), .A2(n16275), .B1(n17234), .B2(U215), .ZN(U261) );
  INV_X1 U19394 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U19395 ( .A1(n16296), .A2(n16276), .B1(n17236), .B2(U215), .ZN(U262) );
  INV_X1 U19396 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U19397 ( .A1(n16298), .A2(n16277), .B1(n17238), .B2(U215), .ZN(U263) );
  INV_X1 U19398 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U19399 ( .A1(n16298), .A2(n16278), .B1(n17243), .B2(U215), .ZN(U264) );
  AOI22_X1 U19400 ( .A1(n16296), .A2(n16279), .B1(n13175), .B2(U215), .ZN(U265) );
  OAI22_X1 U19401 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16298), .ZN(n16280) );
  INV_X1 U19402 ( .A(n16280), .ZN(U266) );
  OAI22_X1 U19403 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16298), .ZN(n16281) );
  INV_X1 U19404 ( .A(n16281), .ZN(U267) );
  OAI22_X1 U19405 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16298), .ZN(n16282) );
  INV_X1 U19406 ( .A(n16282), .ZN(U268) );
  OAI22_X1 U19407 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16298), .ZN(n16283) );
  INV_X1 U19408 ( .A(n16283), .ZN(U269) );
  OAI22_X1 U19409 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16298), .ZN(n16284) );
  INV_X1 U19410 ( .A(n16284), .ZN(U270) );
  OAI22_X1 U19411 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16298), .ZN(n16285) );
  INV_X1 U19412 ( .A(n16285), .ZN(U271) );
  INV_X1 U19413 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16286) );
  INV_X1 U19414 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n17986) );
  AOI22_X1 U19415 ( .A1(n16298), .A2(n16286), .B1(n17986), .B2(U215), .ZN(U272) );
  INV_X1 U19416 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16287) );
  AOI22_X1 U19417 ( .A1(n16298), .A2(n16287), .B1(n14953), .B2(U215), .ZN(U273) );
  OAI22_X1 U19418 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16298), .ZN(n16288) );
  INV_X1 U19419 ( .A(n16288), .ZN(U274) );
  OAI22_X1 U19420 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16296), .ZN(n16289) );
  INV_X1 U19421 ( .A(n16289), .ZN(U275) );
  OAI22_X1 U19422 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16296), .ZN(n16290) );
  INV_X1 U19423 ( .A(n16290), .ZN(U276) );
  OAI22_X1 U19424 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16296), .ZN(n16291) );
  INV_X1 U19425 ( .A(n16291), .ZN(U277) );
  OAI22_X1 U19426 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16296), .ZN(n16292) );
  INV_X1 U19427 ( .A(n16292), .ZN(U278) );
  INV_X1 U19428 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16294) );
  INV_X1 U19429 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U19430 ( .A1(n16298), .A2(n16294), .B1(n17007), .B2(U215), .ZN(U279) );
  OAI22_X1 U19431 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16296), .ZN(n16295) );
  INV_X1 U19432 ( .A(n16295), .ZN(U280) );
  OAI22_X1 U19433 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16296), .ZN(n16297) );
  INV_X1 U19434 ( .A(n16297), .ZN(U281) );
  OAI22_X1 U19435 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n16298), .ZN(n16299) );
  INV_X1 U19436 ( .A(n16299), .ZN(U282) );
  INV_X1 U19437 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16300) );
  AOI222_X1 U19438 ( .A1(n16301), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n18937), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16300), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16302) );
  INV_X2 U19439 ( .A(n16304), .ZN(n16303) );
  INV_X1 U19440 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18509) );
  INV_X1 U19441 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19648) );
  AOI22_X1 U19442 ( .A1(n16303), .A2(n18509), .B1(n19648), .B2(n16304), .ZN(
        U347) );
  INV_X1 U19443 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18507) );
  INV_X1 U19444 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19647) );
  AOI22_X1 U19445 ( .A1(n16303), .A2(n18507), .B1(n19647), .B2(n16304), .ZN(
        U348) );
  INV_X1 U19446 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18504) );
  INV_X1 U19447 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19645) );
  AOI22_X1 U19448 ( .A1(n16303), .A2(n18504), .B1(n19645), .B2(n16304), .ZN(
        U349) );
  INV_X1 U19449 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18503) );
  INV_X1 U19450 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19644) );
  AOI22_X1 U19451 ( .A1(n16303), .A2(n18503), .B1(n19644), .B2(n16304), .ZN(
        U350) );
  INV_X1 U19452 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18501) );
  INV_X1 U19453 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19642) );
  AOI22_X1 U19454 ( .A1(n16303), .A2(n18501), .B1(n19642), .B2(n16304), .ZN(
        U351) );
  INV_X1 U19455 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18499) );
  INV_X1 U19456 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19640) );
  AOI22_X1 U19457 ( .A1(n16303), .A2(n18499), .B1(n19640), .B2(n16304), .ZN(
        U352) );
  INV_X1 U19458 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18497) );
  INV_X1 U19459 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19639) );
  AOI22_X1 U19460 ( .A1(n16303), .A2(n18497), .B1(n19639), .B2(n16304), .ZN(
        U353) );
  INV_X1 U19461 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18495) );
  AOI22_X1 U19462 ( .A1(n16303), .A2(n18495), .B1(n19638), .B2(n16304), .ZN(
        U354) );
  INV_X1 U19463 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18550) );
  INV_X1 U19464 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U19465 ( .A1(n16303), .A2(n18550), .B1(n20840), .B2(n16304), .ZN(
        U355) );
  INV_X1 U19466 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18548) );
  INV_X1 U19467 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19674) );
  AOI22_X1 U19468 ( .A1(n16303), .A2(n18548), .B1(n19674), .B2(n16304), .ZN(
        U356) );
  INV_X1 U19469 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18545) );
  INV_X1 U19470 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19672) );
  AOI22_X1 U19471 ( .A1(n16303), .A2(n18545), .B1(n19672), .B2(n16304), .ZN(
        U357) );
  INV_X1 U19472 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18544) );
  INV_X1 U19473 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19669) );
  AOI22_X1 U19474 ( .A1(n16303), .A2(n18544), .B1(n19669), .B2(n16304), .ZN(
        U358) );
  INV_X1 U19475 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18542) );
  INV_X1 U19476 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19668) );
  AOI22_X1 U19477 ( .A1(n16303), .A2(n18542), .B1(n19668), .B2(n16304), .ZN(
        U359) );
  INV_X1 U19478 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18540) );
  INV_X1 U19479 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19667) );
  AOI22_X1 U19480 ( .A1(n16303), .A2(n18540), .B1(n19667), .B2(n16304), .ZN(
        U360) );
  INV_X1 U19481 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18537) );
  INV_X1 U19482 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19666) );
  AOI22_X1 U19483 ( .A1(n16303), .A2(n18537), .B1(n19666), .B2(n16304), .ZN(
        U361) );
  INV_X1 U19484 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18534) );
  INV_X1 U19485 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19665) );
  AOI22_X1 U19486 ( .A1(n16303), .A2(n18534), .B1(n19665), .B2(n16304), .ZN(
        U362) );
  INV_X1 U19487 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18533) );
  INV_X1 U19488 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19664) );
  AOI22_X1 U19489 ( .A1(n16303), .A2(n18533), .B1(n19664), .B2(n16304), .ZN(
        U363) );
  INV_X1 U19490 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18531) );
  INV_X1 U19491 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U19492 ( .A1(n16303), .A2(n18531), .B1(n19662), .B2(n16304), .ZN(
        U364) );
  INV_X1 U19493 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18493) );
  INV_X1 U19494 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19637) );
  AOI22_X1 U19495 ( .A1(n16303), .A2(n18493), .B1(n19637), .B2(n16304), .ZN(
        U365) );
  INV_X1 U19496 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18529) );
  INV_X1 U19497 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19660) );
  AOI22_X1 U19498 ( .A1(n16303), .A2(n18529), .B1(n19660), .B2(n16304), .ZN(
        U366) );
  INV_X1 U19499 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18527) );
  INV_X1 U19500 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19659) );
  AOI22_X1 U19501 ( .A1(n16303), .A2(n18527), .B1(n19659), .B2(n16304), .ZN(
        U367) );
  INV_X1 U19502 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18525) );
  INV_X1 U19503 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19658) );
  AOI22_X1 U19504 ( .A1(n16303), .A2(n18525), .B1(n19658), .B2(n16304), .ZN(
        U368) );
  INV_X1 U19505 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18523) );
  INV_X1 U19506 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19657) );
  AOI22_X1 U19507 ( .A1(n16303), .A2(n18523), .B1(n19657), .B2(n16304), .ZN(
        U369) );
  INV_X1 U19508 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18521) );
  INV_X1 U19509 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19655) );
  AOI22_X1 U19510 ( .A1(n16303), .A2(n18521), .B1(n19655), .B2(n16304), .ZN(
        U370) );
  INV_X1 U19511 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18519) );
  INV_X1 U19512 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19654) );
  AOI22_X1 U19513 ( .A1(n16303), .A2(n18519), .B1(n19654), .B2(n16304), .ZN(
        U371) );
  INV_X1 U19514 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18516) );
  INV_X1 U19515 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19653) );
  AOI22_X1 U19516 ( .A1(n16303), .A2(n18516), .B1(n19653), .B2(n16304), .ZN(
        U372) );
  INV_X1 U19517 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18515) );
  INV_X1 U19518 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19652) );
  AOI22_X1 U19519 ( .A1(n16303), .A2(n18515), .B1(n19652), .B2(n16304), .ZN(
        U373) );
  INV_X1 U19520 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18512) );
  INV_X1 U19521 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U19522 ( .A1(n16303), .A2(n18512), .B1(n19650), .B2(n16304), .ZN(
        U374) );
  INV_X1 U19523 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18511) );
  INV_X1 U19524 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19649) );
  AOI22_X1 U19525 ( .A1(n16303), .A2(n18511), .B1(n19649), .B2(n16304), .ZN(
        U375) );
  INV_X1 U19526 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18491) );
  INV_X1 U19527 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19635) );
  AOI22_X1 U19528 ( .A1(n16303), .A2(n18491), .B1(n19635), .B2(n16304), .ZN(
        U376) );
  INV_X1 U19529 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16305) );
  NAND2_X1 U19530 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18490), .ZN(n18480) );
  AOI22_X1 U19531 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18480), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18488), .ZN(n18563) );
  OAI21_X1 U19532 ( .B1(n18488), .B2(n16305), .A(n9594), .ZN(P3_U2633) );
  OAI21_X1 U19533 ( .B1(n16313), .B2(n17200), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16306) );
  OAI21_X1 U19534 ( .B1(n16307), .B2(n17621), .A(n16306), .ZN(P3_U2634) );
  AOI21_X1 U19535 ( .B1(n18488), .B2(n18490), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16308) );
  AOI22_X1 U19536 ( .A1(n18610), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16308), 
        .B2(n18629), .ZN(P3_U2635) );
  INV_X1 U19537 ( .A(BS16), .ZN(n18645) );
  AOI21_X1 U19538 ( .B1(n18474), .B2(n18645), .A(n9594), .ZN(n18559) );
  INV_X1 U19539 ( .A(n18559), .ZN(n18561) );
  OAI21_X1 U19540 ( .B1(n18563), .B2(n16309), .A(n18561), .ZN(P3_U2636) );
  INV_X1 U19541 ( .A(n16310), .ZN(n16312) );
  NOR3_X1 U19542 ( .A1(n16313), .A2(n16312), .A3(n16311), .ZN(n18406) );
  NOR2_X1 U19543 ( .A1(n18406), .A2(n18459), .ZN(n18611) );
  OAI21_X1 U19544 ( .B1(n18611), .B2(n16315), .A(n16314), .ZN(P3_U2637) );
  NOR4_X1 U19545 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16319) );
  NOR4_X1 U19546 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16318) );
  NOR4_X1 U19547 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16317) );
  NOR4_X1 U19548 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16316) );
  NAND4_X1 U19549 ( .A1(n16319), .A2(n16318), .A3(n16317), .A4(n16316), .ZN(
        n16325) );
  NOR4_X1 U19550 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16323) );
  AOI211_X1 U19551 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16322) );
  NOR4_X1 U19552 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16321) );
  NOR4_X1 U19553 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16320) );
  NAND4_X1 U19554 ( .A1(n16323), .A2(n16322), .A3(n16321), .A4(n16320), .ZN(
        n16324) );
  NOR2_X1 U19555 ( .A1(n16325), .A2(n16324), .ZN(n18604) );
  INV_X1 U19556 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18557) );
  NOR3_X1 U19557 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16327) );
  OAI21_X1 U19558 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16327), .A(n18604), .ZN(
        n16326) );
  OAI21_X1 U19559 ( .B1(n18604), .B2(n18557), .A(n16326), .ZN(P3_U2638) );
  INV_X1 U19560 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18600) );
  INV_X1 U19561 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18562) );
  AOI21_X1 U19562 ( .B1(n18600), .B2(n18562), .A(n16327), .ZN(n16328) );
  INV_X1 U19563 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18554) );
  INV_X1 U19564 ( .A(n18604), .ZN(n18607) );
  AOI22_X1 U19565 ( .A1(n18604), .A2(n16328), .B1(n18554), .B2(n18607), .ZN(
        P3_U2639) );
  XNOR2_X1 U19566 ( .A(n16330), .B(n16329), .ZN(n16337) );
  NAND2_X1 U19567 ( .A1(n16631), .A2(n16331), .ZN(n16339) );
  INV_X1 U19568 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18551) );
  OAI22_X1 U19569 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16339), .B1(n16338), 
        .B2(n18551), .ZN(n16332) );
  AOI211_X1 U19570 ( .C1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n9591), .A(
        n16333), .B(n16332), .ZN(n16336) );
  OAI21_X1 U19571 ( .B1(n16662), .B2(n16334), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16335) );
  OAI211_X1 U19572 ( .C1(n18467), .C2(n16337), .A(n16336), .B(n16335), .ZN(
        P3_U2641) );
  NAND3_X1 U19573 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16362), .ZN(n16349) );
  AOI22_X1 U19574 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n9591), .B1(
        n16662), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16348) );
  INV_X1 U19575 ( .A(n16338), .ZN(n16346) );
  INV_X1 U19576 ( .A(n16350), .ZN(n16340) );
  AOI21_X1 U19577 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16340), .A(n16339), .ZN(
        n16345) );
  AOI211_X1 U19578 ( .C1(n16343), .C2(n16342), .A(n16341), .B(n16571), .ZN(
        n16344) );
  AOI211_X1 U19579 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16346), .A(n16345), 
        .B(n16344), .ZN(n16347) );
  AOI22_X1 U19580 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n9591), .B1(
        n16662), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16358) );
  AOI211_X1 U19581 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16364), .A(n16350), .B(
        n16673), .ZN(n16354) );
  AOI211_X1 U19582 ( .C1(n16352), .C2(n16351), .A(n9664), .B(n16571), .ZN(
        n16353) );
  AOI211_X1 U19583 ( .C1(n16363), .C2(P3_REIP_REG_28__SCAN_IN), .A(n16354), 
        .B(n16353), .ZN(n16357) );
  NAND2_X1 U19584 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16355) );
  OAI211_X1 U19585 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16362), .B(n16355), .ZN(n16356) );
  NAND3_X1 U19586 ( .A1(n16358), .A2(n16357), .A3(n16356), .ZN(P3_U2643) );
  AOI22_X1 U19587 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n9591), .B1(
        n16662), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16367) );
  INV_X1 U19588 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18543) );
  AOI211_X1 U19589 ( .C1(n17276), .C2(n16360), .A(n16359), .B(n16571), .ZN(
        n16361) );
  AOI221_X1 U19590 ( .B1(n16363), .B2(P3_REIP_REG_27__SCAN_IN), .C1(n16362), 
        .C2(n18543), .A(n16361), .ZN(n16366) );
  OAI211_X1 U19591 ( .C1(n16368), .C2(n16684), .A(n16631), .B(n16364), .ZN(
        n16365) );
  NAND3_X1 U19592 ( .A1(n16367), .A2(n16366), .A3(n16365), .ZN(P3_U2644) );
  AOI211_X1 U19593 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16369), .A(n16368), .B(
        n16673), .ZN(n16375) );
  AOI211_X1 U19594 ( .C1(n16371), .C2(n9658), .A(n16370), .B(n16571), .ZN(
        n16374) );
  INV_X1 U19595 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16372) );
  OAI22_X1 U19596 ( .A1(n17281), .A2(n16659), .B1(n16674), .B2(n16372), .ZN(
        n16373) );
  NOR3_X1 U19597 ( .A1(n16375), .A2(n16374), .A3(n16373), .ZN(n16376) );
  OAI221_X1 U19598 ( .B1(n16378), .B2(n18541), .C1(n16378), .C2(n16377), .A(
        n16376), .ZN(P3_U2645) );
  AOI21_X1 U19599 ( .B1(n16631), .B2(n16379), .A(n16662), .ZN(n16389) );
  NOR2_X1 U19600 ( .A1(n16379), .A2(n16673), .ZN(n16393) );
  AOI22_X1 U19601 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n9591), .B1(
        n16393), .B2(n16388), .ZN(n16387) );
  AOI211_X1 U19602 ( .C1(n16382), .C2(n16381), .A(n16380), .B(n16571), .ZN(
        n16383) );
  AOI221_X1 U19603 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n16385), .C1(n16384), 
        .C2(n16385), .A(n16383), .ZN(n16386) );
  OAI211_X1 U19604 ( .C1(n16389), .C2(n16388), .A(n16387), .B(n16386), .ZN(
        P3_U2646) );
  INV_X1 U19605 ( .A(n16397), .ZN(n16390) );
  AOI21_X1 U19606 ( .B1(n16646), .B2(n16390), .A(n16676), .ZN(n16401) );
  INV_X1 U19607 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18536) );
  AOI22_X1 U19608 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n9591), .B1(
        n16662), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16400) );
  AOI211_X1 U19609 ( .C1(n17310), .C2(n16392), .A(n16391), .B(n16571), .ZN(
        n16396) );
  INV_X1 U19610 ( .A(n16393), .ZN(n16394) );
  AOI21_X1 U19611 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16407), .A(n16394), .ZN(
        n16395) );
  AOI211_X1 U19612 ( .C1(n16398), .C2(n16397), .A(n16396), .B(n16395), .ZN(
        n16399) );
  OAI211_X1 U19613 ( .C1(n16401), .C2(n18536), .A(n16400), .B(n16399), .ZN(
        P3_U2647) );
  AOI221_X1 U19614 ( .B1(n16666), .B2(n18535), .C1(n16402), .C2(n18535), .A(
        n16401), .ZN(n16406) );
  AOI211_X1 U19615 ( .C1(n17321), .C2(n16404), .A(n16403), .B(n16571), .ZN(
        n16405) );
  AOI211_X1 U19616 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16662), .A(n16406), .B(
        n16405), .ZN(n16409) );
  OAI211_X1 U19617 ( .C1(n16414), .C2(n16682), .A(n16631), .B(n16407), .ZN(
        n16408) );
  OAI211_X1 U19618 ( .C1(n16659), .C2(n17324), .A(n16409), .B(n16408), .ZN(
        P3_U2648) );
  AOI221_X1 U19619 ( .B1(n18530), .B2(n16646), .C1(n16420), .C2(n16646), .A(
        n16676), .ZN(n16419) );
  INV_X1 U19620 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18532) );
  NOR2_X1 U19621 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16666), .ZN(n16410) );
  AOI22_X1 U19622 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n9591), .B1(
        n16411), .B2(n16410), .ZN(n16418) );
  AOI211_X1 U19623 ( .C1(n17334), .C2(n16413), .A(n16412), .B(n16571), .ZN(
        n16416) );
  AOI211_X1 U19624 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16427), .A(n16414), .B(
        n16673), .ZN(n16415) );
  AOI211_X1 U19625 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16662), .A(n16416), .B(
        n16415), .ZN(n16417) );
  OAI211_X1 U19626 ( .C1(n16419), .C2(n18532), .A(n16418), .B(n16417), .ZN(
        P3_U2649) );
  INV_X1 U19627 ( .A(n16420), .ZN(n16423) );
  NOR2_X1 U19628 ( .A1(n16666), .A2(n16423), .ZN(n16435) );
  OR2_X1 U19629 ( .A1(n16676), .A2(n16435), .ZN(n16437) );
  AOI211_X1 U19630 ( .C1(n17353), .C2(n16422), .A(n16421), .B(n16571), .ZN(
        n16426) );
  NAND3_X1 U19631 ( .A1(n16646), .A2(n16423), .A3(n18530), .ZN(n16424) );
  OAI21_X1 U19632 ( .B1(n16659), .B2(n20869), .A(n16424), .ZN(n16425) );
  AOI211_X1 U19633 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16437), .A(n16426), 
        .B(n16425), .ZN(n16429) );
  OAI211_X1 U19634 ( .C1(n16433), .C2(n16774), .A(n16631), .B(n16427), .ZN(
        n16428) );
  OAI211_X1 U19635 ( .C1(n16774), .C2(n16674), .A(n16429), .B(n16428), .ZN(
        P3_U2650) );
  AOI211_X1 U19636 ( .C1(n17371), .C2(n16431), .A(n16430), .B(n16571), .ZN(
        n16432) );
  AOI21_X1 U19637 ( .B1(n9591), .B2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16432), .ZN(n16440) );
  AOI211_X1 U19638 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16441), .A(n16433), .B(
        n16673), .ZN(n16434) );
  AOI21_X1 U19639 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16662), .A(n16434), .ZN(
        n16439) );
  AOI22_X1 U19640 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16437), .B1(n16436), 
        .B2(n16435), .ZN(n16438) );
  NAND3_X1 U19641 ( .A1(n16440), .A2(n16439), .A3(n16438), .ZN(P3_U2651) );
  AOI21_X1 U19642 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16458), .A(n16673), .ZN(
        n16442) );
  AOI22_X1 U19643 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n9591), .B1(
        n16442), .B2(n16441), .ZN(n16452) );
  INV_X1 U19644 ( .A(n16463), .ZN(n17378) );
  INV_X1 U19645 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U19646 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16463), .B1(
        n17378), .B2(n17391), .ZN(n17388) );
  AOI21_X1 U19647 ( .B1(n16454), .B2(n17388), .A(n16603), .ZN(n16444) );
  NOR2_X1 U19648 ( .A1(n17391), .A2(n16463), .ZN(n16443) );
  OAI21_X1 U19649 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16443), .A(
        n17330), .ZN(n17383) );
  XNOR2_X1 U19650 ( .A(n16444), .B(n17383), .ZN(n16445) );
  AOI22_X1 U19651 ( .A1(n16662), .A2(P3_EBX_REG_19__SCAN_IN), .B1(n16650), 
        .B2(n16445), .ZN(n16451) );
  INV_X1 U19652 ( .A(n16448), .ZN(n16447) );
  NOR2_X1 U19653 ( .A1(n16676), .A2(n16446), .ZN(n16502) );
  AOI21_X1 U19654 ( .B1(n16447), .B2(n16502), .A(n16479), .ZN(n16471) );
  NAND4_X1 U19655 ( .A1(n16646), .A2(n16501), .A3(P3_REIP_REG_14__SCAN_IN), 
        .A4(P3_REIP_REG_13__SCAN_IN), .ZN(n16492) );
  NOR2_X1 U19656 ( .A1(n16448), .A2(n16492), .ZN(n16457) );
  XNOR2_X1 U19657 ( .A(P3_REIP_REG_19__SCAN_IN), .B(n18524), .ZN(n16449) );
  AOI22_X1 U19658 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16471), .B1(n16457), 
        .B2(n16449), .ZN(n16450) );
  NAND4_X1 U19659 ( .A1(n16452), .A2(n16451), .A3(n16450), .A4(n17835), .ZN(
        P3_U2652) );
  NAND2_X1 U19660 ( .A1(n16454), .A2(n17388), .ZN(n16453) );
  OAI211_X1 U19661 ( .C1(n16454), .C2(n17388), .A(n16650), .B(n16453), .ZN(
        n16455) );
  OAI211_X1 U19662 ( .C1(n17391), .C2(n16659), .A(n17950), .B(n16455), .ZN(
        n16456) );
  AOI221_X1 U19663 ( .B1(n16471), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16457), 
        .C2(n18524), .A(n16456), .ZN(n16461) );
  OAI211_X1 U19664 ( .C1(n16459), .C2(n16462), .A(n16631), .B(n16458), .ZN(
        n16460) );
  OAI211_X1 U19665 ( .C1(n16462), .C2(n16674), .A(n16461), .B(n16460), .ZN(
        P3_U2653) );
  NAND2_X1 U19666 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16476) );
  NOR3_X1 U19667 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16476), .A3(n16492), 
        .ZN(n16470) );
  NAND2_X1 U19668 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17398), .ZN(
        n16480) );
  INV_X1 U19669 ( .A(n16480), .ZN(n16464) );
  OAI21_X1 U19670 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16464), .A(
        n16463), .ZN(n17399) );
  NOR2_X1 U19671 ( .A1(n17617), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16651) );
  AOI21_X1 U19672 ( .B1(n17398), .B2(n16651), .A(n16603), .ZN(n16465) );
  INV_X1 U19673 ( .A(n16465), .ZN(n16467) );
  AOI21_X1 U19674 ( .B1(n17399), .B2(n16467), .A(n18467), .ZN(n16466) );
  OAI21_X1 U19675 ( .B1(n17399), .B2(n16467), .A(n16466), .ZN(n16468) );
  OAI211_X1 U19676 ( .C1(n9723), .C2(n16659), .A(n17950), .B(n16468), .ZN(
        n16469) );
  AOI211_X1 U19677 ( .C1(n16471), .C2(P3_REIP_REG_17__SCAN_IN), .A(n16470), 
        .B(n16469), .ZN(n16474) );
  OAI211_X1 U19678 ( .C1(n16477), .C2(n16475), .A(n16631), .B(n16472), .ZN(
        n16473) );
  OAI211_X1 U19679 ( .C1(n16475), .C2(n16674), .A(n16474), .B(n16473), .ZN(
        P3_U2654) );
  OAI21_X1 U19680 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), 
        .A(n16476), .ZN(n16486) );
  AOI211_X1 U19681 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16494), .A(n16477), .B(
        n16673), .ZN(n16478) );
  AOI21_X1 U19682 ( .B1(n9591), .B2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16478), .ZN(n16485) );
  NOR2_X1 U19683 ( .A1(n16479), .A2(n16502), .ZN(n16504) );
  INV_X1 U19684 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16842) );
  OAI21_X1 U19685 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16487), .A(
        n16480), .ZN(n17418) );
  NAND2_X1 U19686 ( .A1(n10414), .A2(n16481), .ZN(n16488) );
  XNOR2_X1 U19687 ( .A(n17418), .B(n16488), .ZN(n16482) );
  OAI22_X1 U19688 ( .A1(n16674), .A2(n16842), .B1(n18467), .B2(n16482), .ZN(
        n16483) );
  AOI211_X1 U19689 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n16504), .A(n17940), 
        .B(n16483), .ZN(n16484) );
  OAI211_X1 U19690 ( .C1(n16492), .C2(n16486), .A(n16485), .B(n16484), .ZN(
        P3_U2655) );
  AOI21_X1 U19691 ( .B1(n17425), .B2(n17411), .A(n16487), .ZN(n17424) );
  NOR3_X1 U19692 ( .A1(n17424), .A2(n18467), .A3(n16488), .ZN(n16489) );
  AOI211_X1 U19693 ( .C1(n16662), .C2(P3_EBX_REG_15__SCAN_IN), .A(n17940), .B(
        n16489), .ZN(n16491) );
  NOR2_X1 U19694 ( .A1(n10414), .A2(n16571), .ZN(n16620) );
  AOI21_X1 U19695 ( .B1(n10414), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18467), .ZN(n16669) );
  OAI211_X1 U19696 ( .C1(n16620), .C2(n17425), .A(n17424), .B(n16669), .ZN(
        n16490) );
  OAI211_X1 U19697 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n16492), .A(n16491), 
        .B(n16490), .ZN(n16493) );
  AOI21_X1 U19698 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16504), .A(n16493), 
        .ZN(n16497) );
  OAI211_X1 U19699 ( .C1(n16498), .C2(n16495), .A(n16631), .B(n16494), .ZN(
        n16496) );
  OAI211_X1 U19700 ( .C1(n16659), .C2(n17425), .A(n16497), .B(n16496), .ZN(
        P3_U2656) );
  AOI22_X1 U19701 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n9591), .B1(
        n16662), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16507) );
  OAI21_X1 U19702 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16509), .A(
        n17411), .ZN(n17438) );
  INV_X1 U19703 ( .A(n17456), .ZN(n16523) );
  NAND2_X1 U19704 ( .A1(n16675), .A2(n16523), .ZN(n16524) );
  OAI21_X1 U19705 ( .B1(n17460), .B2(n16524), .A(n10414), .ZN(n16511) );
  XOR2_X1 U19706 ( .A(n17438), .B(n16511), .Z(n16500) );
  AOI211_X1 U19707 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16517), .A(n16498), .B(
        n16673), .ZN(n16499) );
  AOI21_X1 U19708 ( .B1(n16500), .B2(n16650), .A(n16499), .ZN(n16506) );
  NAND2_X1 U19709 ( .A1(n16646), .A2(n16501), .ZN(n16515) );
  NOR2_X1 U19710 ( .A1(n16502), .A2(n16515), .ZN(n16503) );
  AOI22_X1 U19711 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16504), .B1(
        P3_REIP_REG_13__SCAN_IN), .B2(n16503), .ZN(n16505) );
  NAND4_X1 U19712 ( .A1(n16507), .A2(n16506), .A3(n16505), .A4(n17835), .ZN(
        P3_U2657) );
  INV_X1 U19713 ( .A(n16508), .ZN(n16528) );
  INV_X1 U19714 ( .A(n16676), .ZN(n16552) );
  OAI21_X1 U19715 ( .B1(n16528), .B2(n16666), .A(n16552), .ZN(n16536) );
  NOR2_X1 U19716 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16666), .ZN(n16527) );
  NAND2_X1 U19717 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16523), .ZN(
        n16510) );
  AOI21_X1 U19718 ( .B1(n17463), .B2(n16510), .A(n16509), .ZN(n17468) );
  NOR3_X1 U19719 ( .A1(n17468), .A2(n16571), .A3(n16511), .ZN(n16512) );
  AOI211_X1 U19720 ( .C1(n16662), .C2(P3_EBX_REG_13__SCAN_IN), .A(n17877), .B(
        n16512), .ZN(n16514) );
  OAI211_X1 U19721 ( .C1(n16603), .C2(n17463), .A(n17468), .B(n16669), .ZN(
        n16513) );
  OAI211_X1 U19722 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16515), .A(n16514), 
        .B(n16513), .ZN(n16516) );
  AOI221_X1 U19723 ( .B1(n16536), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16527), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16516), .ZN(n16520) );
  OAI211_X1 U19724 ( .C1(n16521), .C2(n16518), .A(n16631), .B(n16517), .ZN(
        n16519) );
  OAI211_X1 U19725 ( .C1(n16659), .C2(n17463), .A(n16520), .B(n16519), .ZN(
        P3_U2658) );
  AOI211_X1 U19726 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16537), .A(n16521), .B(
        n16673), .ZN(n16522) );
  AOI21_X1 U19727 ( .B1(n9591), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16522), .ZN(n16531) );
  AOI22_X1 U19728 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16523), .B1(
        n17456), .B2(n17477), .ZN(n17474) );
  AND2_X1 U19729 ( .A1(n16524), .A2(n10414), .ZN(n16525) );
  XOR2_X1 U19730 ( .A(n17474), .B(n16525), .Z(n16526) );
  AOI22_X1 U19731 ( .A1(n16662), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16650), 
        .B2(n16526), .ZN(n16530) );
  AOI22_X1 U19732 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16536), .B1(n16528), 
        .B2(n16527), .ZN(n16529) );
  NAND4_X1 U19733 ( .A1(n16531), .A2(n16530), .A3(n16529), .A4(n17835), .ZN(
        P3_U2659) );
  AND3_X1 U19734 ( .A1(n17487), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        n16592), .ZN(n16544) );
  OAI21_X1 U19735 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16544), .A(
        n17456), .ZN(n17488) );
  INV_X1 U19736 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17499) );
  NAND3_X1 U19737 ( .A1(n16532), .A2(n17487), .A3(n16651), .ZN(n16543) );
  OAI21_X1 U19738 ( .B1(n17499), .B2(n16543), .A(n10414), .ZN(n16546) );
  XOR2_X1 U19739 ( .A(n17488), .B(n16546), .Z(n16533) );
  AOI22_X1 U19740 ( .A1(n16662), .A2(P3_EBX_REG_11__SCAN_IN), .B1(n16650), 
        .B2(n16533), .ZN(n16541) );
  NAND2_X1 U19741 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16534) );
  NAND2_X1 U19742 ( .A1(n16646), .A2(n16568), .ZN(n16551) );
  INV_X1 U19743 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18510) );
  OAI21_X1 U19744 ( .B1(n16534), .B2(n16551), .A(n18510), .ZN(n16535) );
  AOI22_X1 U19745 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n9591), .B1(
        n16536), .B2(n16535), .ZN(n16540) );
  OAI211_X1 U19746 ( .C1(n16542), .C2(n16538), .A(n16631), .B(n16537), .ZN(
        n16539) );
  NAND4_X1 U19747 ( .A1(n16541), .A2(n16540), .A3(n17835), .A4(n16539), .ZN(
        P3_U2660) );
  AOI22_X1 U19748 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n9591), .B1(
        n16662), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n16555) );
  INV_X1 U19749 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18506) );
  NOR3_X1 U19750 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18506), .A3(n16551), 
        .ZN(n16550) );
  AOI211_X1 U19751 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16564), .A(n16542), .B(
        n16673), .ZN(n16549) );
  INV_X1 U19752 ( .A(n16543), .ZN(n16561) );
  NOR2_X1 U19753 ( .A1(n16561), .A2(n16603), .ZN(n16547) );
  NAND2_X1 U19754 ( .A1(n17487), .A2(n16592), .ZN(n16556) );
  AOI21_X1 U19755 ( .B1(n17499), .B2(n16556), .A(n16544), .ZN(n17501) );
  INV_X1 U19756 ( .A(n17501), .ZN(n16545) );
  AOI221_X1 U19757 ( .B1(n16547), .B2(n17501), .C1(n16546), .C2(n16545), .A(
        n18467), .ZN(n16548) );
  NOR4_X1 U19758 ( .A1(n17940), .A2(n16550), .A3(n16549), .A4(n16548), .ZN(
        n16554) );
  NOR2_X1 U19759 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16551), .ZN(n16563) );
  OAI21_X1 U19760 ( .B1(n16568), .B2(n16666), .A(n16552), .ZN(n16575) );
  OAI21_X1 U19761 ( .B1(n16563), .B2(n16575), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16553) );
  NAND3_X1 U19762 ( .A1(n16555), .A2(n16554), .A3(n16553), .ZN(P3_U2661) );
  NOR2_X1 U19763 ( .A1(n16603), .A2(n18467), .ZN(n16661) );
  NAND3_X1 U19764 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16532), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16581) );
  NOR2_X1 U19765 ( .A1(n17526), .A2(n16581), .ZN(n16570) );
  OAI21_X1 U19766 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16570), .A(
        n16556), .ZN(n17514) );
  NOR2_X1 U19767 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18467), .ZN(
        n16557) );
  AOI22_X1 U19768 ( .A1(n16661), .A2(n17514), .B1(n16570), .B2(n16557), .ZN(
        n16560) );
  INV_X1 U19769 ( .A(n17514), .ZN(n16558) );
  AOI22_X1 U19770 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n9591), .B1(
        n16558), .B2(n16620), .ZN(n16559) );
  OAI211_X1 U19771 ( .C1(n16561), .C2(n16560), .A(n16559), .B(n17835), .ZN(
        n16562) );
  AOI211_X1 U19772 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n16575), .A(n16563), .B(
        n16562), .ZN(n16566) );
  OAI211_X1 U19773 ( .C1(n16569), .C2(n16567), .A(n16631), .B(n16564), .ZN(
        n16565) );
  OAI211_X1 U19774 ( .C1(n16567), .C2(n16674), .A(n16566), .B(n16565), .ZN(
        P3_U2662) );
  OR2_X1 U19775 ( .A1(n16666), .A2(n16568), .ZN(n16578) );
  AOI22_X1 U19776 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n9591), .B1(
        n16662), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n16577) );
  AOI211_X1 U19777 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16588), .A(n16569), .B(
        n16673), .ZN(n16574) );
  OAI21_X1 U19778 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16581), .A(
        n10414), .ZN(n16582) );
  AOI21_X1 U19779 ( .B1(n17526), .B2(n16581), .A(n16570), .ZN(n17532) );
  XOR2_X1 U19780 ( .A(n16582), .B(n17532), .Z(n16572) );
  OAI21_X1 U19781 ( .B1(n16572), .B2(n16571), .A(n17835), .ZN(n16573) );
  AOI211_X1 U19782 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n16575), .A(n16574), .B(
        n16573), .ZN(n16576) );
  OAI211_X1 U19783 ( .C1(n16579), .C2(n16578), .A(n16577), .B(n16576), .ZN(
        P3_U2663) );
  INV_X1 U19784 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18502) );
  AND3_X1 U19785 ( .A1(n16646), .A2(n16580), .A3(n18502), .ZN(n16587) );
  AOI21_X1 U19786 ( .B1(n16532), .B2(n16651), .A(n16603), .ZN(n16593) );
  OAI21_X1 U19787 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16592), .A(
        n16581), .ZN(n17545) );
  INV_X1 U19788 ( .A(n17545), .ZN(n16583) );
  AOI221_X1 U19789 ( .B1(n16593), .B2(n16583), .C1(n16582), .C2(n17545), .A(
        n18467), .ZN(n16586) );
  AOI221_X1 U19790 ( .B1(n18500), .B2(n16646), .C1(n16602), .C2(n16646), .A(
        n16676), .ZN(n16584) );
  OAI22_X1 U19791 ( .A1(n16584), .A2(n18502), .B1(n16674), .B2(n16589), .ZN(
        n16585) );
  NOR4_X1 U19792 ( .A1(n17940), .A2(n16587), .A3(n16586), .A4(n16585), .ZN(
        n16591) );
  OAI211_X1 U19793 ( .C1(n16597), .C2(n16589), .A(n16631), .B(n16588), .ZN(
        n16590) );
  OAI211_X1 U19794 ( .C1(n16659), .C2(n20781), .A(n16591), .B(n16590), .ZN(
        P3_U2664) );
  AOI21_X1 U19795 ( .B1(n16646), .B2(n16602), .A(n16676), .ZN(n16608) );
  AOI21_X1 U19796 ( .B1(n17555), .B2(n16604), .A(n16592), .ZN(n17558) );
  NAND2_X1 U19797 ( .A1(n16650), .A2(n16593), .ZN(n16595) );
  OAI211_X1 U19798 ( .C1(n16620), .C2(n17555), .A(n17558), .B(n16669), .ZN(
        n16594) );
  OAI21_X1 U19799 ( .B1(n17558), .B2(n16595), .A(n16594), .ZN(n16596) );
  AOI211_X1 U19800 ( .C1(n16662), .C2(P3_EBX_REG_6__SCAN_IN), .A(n17877), .B(
        n16596), .ZN(n16601) );
  NOR3_X1 U19801 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16666), .A3(n16602), .ZN(
        n16599) );
  AOI211_X1 U19802 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16612), .A(n16597), .B(
        n16673), .ZN(n16598) );
  AOI211_X1 U19803 ( .C1(n9591), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16599), .B(n16598), .ZN(n16600) );
  OAI211_X1 U19804 ( .C1(n16608), .C2(n18500), .A(n16601), .B(n16600), .ZN(
        P3_U2665) );
  INV_X1 U19805 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16615) );
  AND2_X1 U19806 ( .A1(n16602), .A2(n16646), .ZN(n16610) );
  INV_X1 U19807 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18498) );
  AOI21_X1 U19808 ( .B1(n17567), .B2(n16651), .A(n16603), .ZN(n16619) );
  NAND2_X1 U19809 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17567), .ZN(
        n16618) );
  INV_X1 U19810 ( .A(n16618), .ZN(n16605) );
  OAI21_X1 U19811 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16605), .A(
        n16604), .ZN(n17570) );
  XNOR2_X1 U19812 ( .A(n16619), .B(n17570), .ZN(n16606) );
  AOI22_X1 U19813 ( .A1(n16662), .A2(P3_EBX_REG_5__SCAN_IN), .B1(n16650), .B2(
        n16606), .ZN(n16607) );
  OAI211_X1 U19814 ( .C1(n16608), .C2(n18498), .A(n16607), .B(n17950), .ZN(
        n16609) );
  AOI21_X1 U19815 ( .B1(n16611), .B2(n16610), .A(n16609), .ZN(n16614) );
  OAI211_X1 U19816 ( .C1(n16616), .C2(n16896), .A(n16631), .B(n16612), .ZN(
        n16613) );
  OAI211_X1 U19817 ( .C1(n16659), .C2(n16615), .A(n16614), .B(n16613), .ZN(
        P3_U2666) );
  AOI21_X1 U19818 ( .B1(n16646), .B2(n16629), .A(n16676), .ZN(n16643) );
  AOI22_X1 U19819 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n9591), .B1(
        n16662), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16628) );
  AOI211_X1 U19820 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16630), .A(n16616), .B(
        n16673), .ZN(n16626) );
  NOR3_X1 U19821 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16666), .A3(n16629), .ZN(
        n16625) );
  INV_X1 U19822 ( .A(n17582), .ZN(n16617) );
  NOR2_X1 U19823 ( .A1(n16617), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17575) );
  NOR2_X1 U19824 ( .A1(n17617), .A2(n16617), .ZN(n16633) );
  OAI21_X1 U19825 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16633), .A(
        n16618), .ZN(n17585) );
  AOI22_X1 U19826 ( .A1(n16651), .A2(n17575), .B1(n16619), .B2(n17585), .ZN(
        n16621) );
  INV_X1 U19827 ( .A(n16620), .ZN(n16654) );
  OAI22_X1 U19828 ( .A1(n16621), .A2(n18467), .B1(n17585), .B2(n16654), .ZN(
        n16624) );
  NAND2_X1 U19829 ( .A1(n17968), .A2(n18634), .ZN(n18637) );
  OAI221_X1 U19830 ( .B1(n18637), .B2(n16622), .C1(n18637), .C2(n18409), .A(
        n17835), .ZN(n16623) );
  NOR4_X1 U19831 ( .A1(n16626), .A2(n16625), .A3(n16624), .A4(n16623), .ZN(
        n16627) );
  OAI211_X1 U19832 ( .C1(n16643), .C2(n18496), .A(n16628), .B(n16627), .ZN(
        P3_U2667) );
  INV_X1 U19833 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18494) );
  INV_X1 U19834 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18492) );
  NOR2_X1 U19835 ( .A1(n18600), .A2(n18492), .ZN(n16648) );
  AND2_X1 U19836 ( .A1(n16629), .A2(n16646), .ZN(n16641) );
  OAI22_X1 U19837 ( .A1(n16634), .A2(n16659), .B1(n16674), .B2(n16632), .ZN(
        n16640) );
  INV_X1 U19838 ( .A(n18432), .ZN(n18413) );
  NAND2_X1 U19839 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18413), .ZN(
        n18415) );
  AOI21_X1 U19840 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18415), .A(
        n16819), .ZN(n18567) );
  OAI211_X1 U19841 ( .C1(n16644), .C2(n16632), .A(n16631), .B(n16630), .ZN(
        n16638) );
  NAND2_X1 U19842 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16649) );
  AOI21_X1 U19843 ( .B1(n16634), .B2(n16649), .A(n16633), .ZN(n16635) );
  INV_X1 U19844 ( .A(n16635), .ZN(n17594) );
  OAI21_X1 U19845 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16649), .A(
        n10414), .ZN(n16653) );
  AOI21_X1 U19846 ( .B1(n17594), .B2(n16653), .A(n18467), .ZN(n16636) );
  OAI21_X1 U19847 ( .B1(n17594), .B2(n16653), .A(n16636), .ZN(n16637) );
  OAI211_X1 U19848 ( .C1(n18567), .C2(n18637), .A(n16638), .B(n16637), .ZN(
        n16639) );
  AOI211_X1 U19849 ( .C1(n16648), .C2(n16641), .A(n16640), .B(n16639), .ZN(
        n16642) );
  OAI21_X1 U19850 ( .B1(n16643), .B2(n18494), .A(n16642), .ZN(P3_U2668) );
  OR2_X1 U19851 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n16665) );
  AOI211_X1 U19852 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16665), .A(n16644), .B(
        n16673), .ZN(n16645) );
  AOI21_X1 U19853 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n16662), .A(n16645), .ZN(
        n16658) );
  OAI21_X1 U19854 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16646), .ZN(n16647) );
  NAND2_X1 U19855 ( .A1(n18584), .A2(n18429), .ZN(n18412) );
  OAI21_X1 U19856 ( .B1(n18432), .B2(n18598), .A(n18412), .ZN(n18578) );
  OAI22_X1 U19857 ( .A1(n16648), .A2(n16647), .B1(n18637), .B2(n18578), .ZN(
        n16656) );
  OAI21_X1 U19858 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16649), .ZN(n17604) );
  OAI21_X1 U19859 ( .B1(n16651), .B2(n17604), .A(n16650), .ZN(n16652) );
  OAI22_X1 U19860 ( .A1(n17604), .A2(n16654), .B1(n16653), .B2(n16652), .ZN(
        n16655) );
  AOI211_X1 U19861 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n16676), .A(n16656), .B(
        n16655), .ZN(n16657) );
  OAI211_X1 U19862 ( .C1(n17608), .C2(n16659), .A(n16658), .B(n16657), .ZN(
        P3_U2669) );
  AOI21_X1 U19863 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16661), .A(
        n9591), .ZN(n16672) );
  AOI22_X1 U19864 ( .A1(n16662), .A2(P3_EBX_REG_1__SCAN_IN), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n16676), .ZN(n16671) );
  NAND2_X1 U19865 ( .A1(n18429), .A2(n16663), .ZN(n18585) );
  NOR2_X1 U19866 ( .A1(n18585), .A2(n18637), .ZN(n16668) );
  NAND2_X1 U19867 ( .A1(n16665), .A2(n16664), .ZN(n16977) );
  OAI22_X1 U19868 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16666), .B1(n16673), 
        .B2(n16977), .ZN(n16667) );
  AOI211_X1 U19869 ( .C1(n17617), .C2(n16669), .A(n16668), .B(n16667), .ZN(
        n16670) );
  OAI211_X1 U19870 ( .C1(n16672), .C2(n17617), .A(n16671), .B(n16670), .ZN(
        P3_U2670) );
  INV_X1 U19871 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n16984) );
  AOI21_X1 U19872 ( .B1(n16674), .B2(n16673), .A(n16984), .ZN(n16678) );
  NOR3_X1 U19873 ( .A1(n18632), .A2(n16676), .A3(n16675), .ZN(n16677) );
  AOI211_X1 U19874 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n16679), .A(n16678), .B(
        n16677), .ZN(n16680) );
  OAI21_X1 U19875 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18637), .A(
        n16680), .ZN(P3_U2671) );
  NOR4_X1 U19876 ( .A1(n16683), .A2(n16682), .A3(n16681), .A4(n16774), .ZN(
        n16687) );
  NOR4_X1 U19877 ( .A1(n16721), .A2(n16685), .A3(n16684), .A4(n16773), .ZN(
        n16686) );
  NAND4_X1 U19878 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16687), .A4(n16686), .ZN(n16690) );
  NOR2_X1 U19879 ( .A1(n16691), .A2(n16690), .ZN(n16717) );
  NAND2_X1 U19880 ( .A1(n16969), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16689) );
  NAND2_X1 U19881 ( .A1(n16717), .A2(n17999), .ZN(n16688) );
  OAI22_X1 U19882 ( .A1(n16717), .A2(n16689), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16688), .ZN(P3_U2672) );
  NAND2_X1 U19883 ( .A1(n16691), .A2(n16690), .ZN(n16692) );
  NAND2_X1 U19884 ( .A1(n16692), .A2(n16969), .ZN(n16716) );
  AOI22_X1 U19885 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16696) );
  AOI22_X1 U19886 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16695) );
  AOI22_X1 U19887 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16694) );
  AOI22_X1 U19888 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9608), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16693) );
  NAND4_X1 U19889 ( .A1(n16696), .A2(n16695), .A3(n16694), .A4(n16693), .ZN(
        n16703) );
  AOI22_X1 U19890 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16701) );
  AOI22_X1 U19891 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16920), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16700) );
  AOI22_X1 U19892 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16699) );
  AOI22_X1 U19893 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16698) );
  NAND4_X1 U19894 ( .A1(n16701), .A2(n16700), .A3(n16699), .A4(n16698), .ZN(
        n16702) );
  NOR2_X1 U19895 ( .A1(n16703), .A2(n16702), .ZN(n16715) );
  AOI22_X1 U19896 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16940), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16714) );
  AOI22_X1 U19897 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16713) );
  AOI22_X1 U19898 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16704) );
  OAI21_X1 U19899 ( .B1(n16705), .B2(n16959), .A(n16704), .ZN(n16711) );
  AOI22_X1 U19900 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16709) );
  AOI22_X1 U19901 ( .A1(n16819), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16708) );
  AOI22_X1 U19902 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16707) );
  AOI22_X1 U19903 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16706) );
  NAND4_X1 U19904 ( .A1(n16709), .A2(n16708), .A3(n16707), .A4(n16706), .ZN(
        n16710) );
  AOI211_X1 U19905 ( .C1(n16914), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n16711), .B(n16710), .ZN(n16712) );
  NAND3_X1 U19906 ( .A1(n16714), .A2(n16713), .A3(n16712), .ZN(n16719) );
  NAND2_X1 U19907 ( .A1(n16720), .A2(n16719), .ZN(n16718) );
  XNOR2_X1 U19908 ( .A(n16715), .B(n16718), .ZN(n16997) );
  OAI22_X1 U19909 ( .A1(n16717), .A2(n16716), .B1(n16997), .B2(n16969), .ZN(
        P3_U2673) );
  OAI21_X1 U19910 ( .B1(n16720), .B2(n16719), .A(n16718), .ZN(n17001) );
  AOI22_X1 U19911 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16723), .B1(n16722), 
        .B2(n16721), .ZN(n16724) );
  OAI21_X1 U19912 ( .B1(n17001), .B2(n16969), .A(n16724), .ZN(P3_U2674) );
  OAI21_X1 U19913 ( .B1(n16729), .B2(n16726), .A(n16725), .ZN(n17011) );
  NAND3_X1 U19914 ( .A1(n16728), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n16969), 
        .ZN(n16727) );
  OAI221_X1 U19915 ( .B1(n16728), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n16969), 
        .C2(n17011), .A(n16727), .ZN(P3_U2676) );
  AOI21_X1 U19916 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16969), .A(n16737), .ZN(
        n16732) );
  AOI21_X1 U19917 ( .B1(n16730), .B2(n16734), .A(n16729), .ZN(n17012) );
  INV_X1 U19918 ( .A(n17012), .ZN(n16731) );
  OAI22_X1 U19919 ( .A1(n16733), .A2(n16732), .B1(n16969), .B2(n16731), .ZN(
        P3_U2677) );
  AOI21_X1 U19920 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16969), .A(n16743), .ZN(
        n16736) );
  OAI21_X1 U19921 ( .B1(n16739), .B2(n16735), .A(n16734), .ZN(n17020) );
  OAI22_X1 U19922 ( .A1(n16737), .A2(n16736), .B1(n16969), .B2(n17020), .ZN(
        P3_U2678) );
  INV_X1 U19923 ( .A(n16738), .ZN(n16749) );
  AOI21_X1 U19924 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16969), .A(n16749), .ZN(
        n16742) );
  AOI21_X1 U19925 ( .B1(n16740), .B2(n16745), .A(n16739), .ZN(n17021) );
  INV_X1 U19926 ( .A(n17021), .ZN(n16741) );
  OAI22_X1 U19927 ( .A1(n16743), .A2(n16742), .B1(n16969), .B2(n16741), .ZN(
        P3_U2679) );
  AOI21_X1 U19928 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n16969), .A(n16744), .ZN(
        n16748) );
  OAI21_X1 U19929 ( .B1(n16747), .B2(n16746), .A(n16745), .ZN(n17030) );
  OAI22_X1 U19930 ( .A1(n16749), .A2(n16748), .B1(n16969), .B2(n17030), .ZN(
        P3_U2680) );
  AOI22_X1 U19931 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16753) );
  AOI22_X1 U19932 ( .A1(n16819), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16752) );
  AOI22_X1 U19933 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16751) );
  AOI22_X1 U19934 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16750) );
  NAND4_X1 U19935 ( .A1(n16753), .A2(n16752), .A3(n16751), .A4(n16750), .ZN(
        n16760) );
  AOI22_X1 U19936 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9600), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16758) );
  AOI22_X1 U19937 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16920), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16757) );
  AOI22_X1 U19938 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16754), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16756) );
  AOI22_X1 U19939 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16939), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16755) );
  NAND4_X1 U19940 ( .A1(n16758), .A2(n16757), .A3(n16756), .A4(n16755), .ZN(
        n16759) );
  NOR2_X1 U19941 ( .A1(n16760), .A2(n16759), .ZN(n17033) );
  NAND3_X1 U19942 ( .A1(n16762), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n16969), 
        .ZN(n16761) );
  OAI221_X1 U19943 ( .B1(n16762), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n16969), 
        .C2(n17033), .A(n16761), .ZN(P3_U2681) );
  AOI22_X1 U19944 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16940), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16766) );
  AOI22_X1 U19945 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16765) );
  AOI22_X1 U19946 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16764) );
  AOI22_X1 U19947 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16763) );
  NAND4_X1 U19948 ( .A1(n16766), .A2(n16765), .A3(n16764), .A4(n16763), .ZN(
        n16772) );
  AOI22_X1 U19949 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16770) );
  AOI22_X1 U19950 ( .A1(n16919), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16769) );
  AOI22_X1 U19951 ( .A1(n16819), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16768) );
  AOI22_X1 U19952 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16767) );
  NAND4_X1 U19953 ( .A1(n16770), .A2(n16769), .A3(n16768), .A4(n16767), .ZN(
        n16771) );
  NOR2_X1 U19954 ( .A1(n16772), .A2(n16771), .ZN(n17039) );
  AND2_X1 U19955 ( .A1(n16969), .A2(n16773), .ZN(n16787) );
  AOI22_X1 U19956 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16787), .B1(n16775), 
        .B2(n16774), .ZN(n16776) );
  OAI21_X1 U19957 ( .B1(n17039), .B2(n16969), .A(n16776), .ZN(P3_U2682) );
  AOI22_X1 U19958 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16940), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16786) );
  AOI22_X1 U19959 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16785) );
  AOI22_X1 U19960 ( .A1(n15538), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16777) );
  OAI21_X1 U19961 ( .B1(n16804), .B2(n16967), .A(n16777), .ZN(n16783) );
  AOI22_X1 U19962 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9608), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16781) );
  AOI22_X1 U19963 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16780) );
  AOI22_X1 U19964 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16779) );
  AOI22_X1 U19965 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16778) );
  NAND4_X1 U19966 ( .A1(n16781), .A2(n16780), .A3(n16779), .A4(n16778), .ZN(
        n16782) );
  AOI211_X1 U19967 ( .C1(n9609), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n16783), .B(n16782), .ZN(n16784) );
  NAND3_X1 U19968 ( .A1(n16786), .A2(n16785), .A3(n16784), .ZN(n17044) );
  INV_X1 U19969 ( .A(n17044), .ZN(n16789) );
  OAI21_X1 U19970 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16802), .A(n16787), .ZN(
        n16788) );
  OAI21_X1 U19971 ( .B1(n16789), .B2(n16969), .A(n16788), .ZN(P3_U2683) );
  OAI21_X1 U19972 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16790), .A(n16969), .ZN(
        n16801) );
  AOI22_X1 U19973 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16794) );
  AOI22_X1 U19974 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16919), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16793) );
  AOI22_X1 U19975 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16792) );
  AOI22_X1 U19976 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16791) );
  NAND4_X1 U19977 ( .A1(n16794), .A2(n16793), .A3(n16792), .A4(n16791), .ZN(
        n16800) );
  AOI22_X1 U19978 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16920), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16798) );
  AOI22_X1 U19979 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16797) );
  AOI22_X1 U19980 ( .A1(n16940), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16796) );
  AOI22_X1 U19981 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16795) );
  NAND4_X1 U19982 ( .A1(n16798), .A2(n16797), .A3(n16796), .A4(n16795), .ZN(
        n16799) );
  NOR2_X1 U19983 ( .A1(n16800), .A2(n16799), .ZN(n17052) );
  OAI22_X1 U19984 ( .A1(n16802), .A2(n16801), .B1(n17052), .B2(n16969), .ZN(
        P3_U2684) );
  AOI22_X1 U19985 ( .A1(n16819), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16813) );
  AOI22_X1 U19986 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16812) );
  AOI22_X1 U19987 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16803) );
  OAI21_X1 U19988 ( .B1(n16804), .B2(n16976), .A(n16803), .ZN(n16810) );
  AOI22_X1 U19989 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9604), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16808) );
  AOI22_X1 U19990 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16807) );
  AOI22_X1 U19991 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16806) );
  AOI22_X1 U19992 ( .A1(n16939), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16805) );
  NAND4_X1 U19993 ( .A1(n16808), .A2(n16807), .A3(n16806), .A4(n16805), .ZN(
        n16809) );
  AOI211_X1 U19994 ( .C1(n16914), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n16810), .B(n16809), .ZN(n16811) );
  NAND3_X1 U19995 ( .A1(n16813), .A2(n16812), .A3(n16811), .ZN(n17053) );
  INV_X1 U19996 ( .A(n17053), .ZN(n16816) );
  OAI21_X1 U19997 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16831), .A(n16814), .ZN(
        n16815) );
  AOI22_X1 U19998 ( .A1(n16982), .A2(n16816), .B1(n16815), .B2(n16969), .ZN(
        P3_U2685) );
  INV_X1 U19999 ( .A(n16817), .ZN(n16818) );
  OAI21_X1 U20000 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16818), .A(n16969), .ZN(
        n16830) );
  AOI22_X1 U20001 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16823) );
  AOI22_X1 U20002 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n16819), .B1(
        n9604), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16822) );
  AOI22_X1 U20003 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n16920), .ZN(n16821) );
  AOI22_X1 U20004 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n9609), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9600), .ZN(n16820) );
  NAND4_X1 U20005 ( .A1(n16823), .A2(n16822), .A3(n16821), .A4(n16820), .ZN(
        n16829) );
  AOI22_X1 U20006 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n15538), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n10299), .ZN(n16827) );
  AOI22_X1 U20007 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n16933), .ZN(n16826) );
  AOI22_X1 U20008 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n16919), .ZN(n16825) );
  AOI22_X1 U20009 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n16871), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16824) );
  NAND4_X1 U20010 ( .A1(n16827), .A2(n16826), .A3(n16825), .A4(n16824), .ZN(
        n16828) );
  NOR2_X1 U20011 ( .A1(n16829), .A2(n16828), .ZN(n17063) );
  OAI22_X1 U20012 ( .A1(n16831), .A2(n16830), .B1(n17063), .B2(n16969), .ZN(
        P3_U2686) );
  AOI22_X1 U20013 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16835) );
  AOI22_X1 U20014 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U20015 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16920), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16833) );
  AOI22_X1 U20016 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9609), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16832) );
  NAND4_X1 U20017 ( .A1(n16835), .A2(n16834), .A3(n16833), .A4(n16832), .ZN(
        n16841) );
  AOI22_X1 U20018 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16839) );
  AOI22_X1 U20019 ( .A1(n10311), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16838) );
  AOI22_X1 U20020 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16837) );
  AOI22_X1 U20021 ( .A1(n16939), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16836) );
  NAND4_X1 U20022 ( .A1(n16839), .A2(n16838), .A3(n16837), .A4(n16836), .ZN(
        n16840) );
  NOR2_X1 U20023 ( .A1(n16841), .A2(n16840), .ZN(n17069) );
  NOR2_X1 U20024 ( .A1(n16982), .A2(n16843), .ZN(n16855) );
  OAI222_X1 U20025 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17999), .B1(
        P3_EBX_REG_16__SCAN_IN), .B2(n16843), .C1(n16855), .C2(n16842), .ZN(
        n16844) );
  OAI21_X1 U20026 ( .B1(n17069), .B2(n16969), .A(n16844), .ZN(P3_U2687) );
  AOI22_X1 U20027 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16848) );
  AOI22_X1 U20028 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16920), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16847) );
  AOI22_X1 U20029 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9608), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16846) );
  AOI22_X1 U20030 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16845) );
  NAND4_X1 U20031 ( .A1(n16848), .A2(n16847), .A3(n16846), .A4(n16845), .ZN(
        n16854) );
  AOI22_X1 U20032 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16919), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16852) );
  AOI22_X1 U20033 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16851) );
  AOI22_X1 U20034 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16850) );
  AOI22_X1 U20035 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16849) );
  NAND4_X1 U20036 ( .A1(n16852), .A2(n16851), .A3(n16850), .A4(n16849), .ZN(
        n16853) );
  NOR2_X1 U20037 ( .A1(n16854), .A2(n16853), .ZN(n17073) );
  INV_X1 U20038 ( .A(n16868), .ZN(n16856) );
  OAI21_X1 U20039 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16856), .A(n16855), .ZN(
        n16857) );
  OAI21_X1 U20040 ( .B1(n17073), .B2(n16969), .A(n16857), .ZN(P3_U2688) );
  AOI22_X1 U20041 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16919), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U20042 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16860) );
  AOI22_X1 U20043 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16920), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20044 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16858) );
  NAND4_X1 U20045 ( .A1(n16861), .A2(n16860), .A3(n16859), .A4(n16858), .ZN(
        n16867) );
  AOI22_X1 U20046 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16865) );
  AOI22_X1 U20047 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16864) );
  AOI22_X1 U20048 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16863) );
  AOI22_X1 U20049 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16862) );
  NAND4_X1 U20050 ( .A1(n16865), .A2(n16864), .A3(n16863), .A4(n16862), .ZN(
        n16866) );
  NOR2_X1 U20051 ( .A1(n16867), .A2(n16866), .ZN(n17078) );
  OAI221_X1 U20052 ( .B1(n16869), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n17999), 
        .C2(n16978), .A(n16868), .ZN(n16870) );
  OAI21_X1 U20053 ( .B1(n17078), .B2(n16969), .A(n16870), .ZN(P3_U2689) );
  AOI22_X1 U20054 ( .A1(n16921), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16919), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16875) );
  AOI22_X1 U20055 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16874) );
  AOI22_X1 U20056 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9604), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16873) );
  AOI22_X1 U20057 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16872) );
  NAND4_X1 U20058 ( .A1(n16875), .A2(n16874), .A3(n16873), .A4(n16872), .ZN(
        n16882) );
  AOI22_X1 U20059 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16880) );
  AOI22_X1 U20060 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20061 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16878) );
  AOI22_X1 U20062 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16877) );
  NAND4_X1 U20063 ( .A1(n16880), .A2(n16879), .A3(n16878), .A4(n16877), .ZN(
        n16881) );
  NOR2_X1 U20064 ( .A1(n16882), .A2(n16881), .ZN(n17083) );
  NOR3_X1 U20065 ( .A1(n16978), .A2(n16960), .A3(n16883), .ZN(n16898) );
  OAI211_X1 U20066 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16898), .A(n16884), .B(
        n16969), .ZN(n16885) );
  OAI21_X1 U20067 ( .B1(n17083), .B2(n16969), .A(n16885), .ZN(P3_U2691) );
  AOI22_X1 U20068 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U20069 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16888) );
  AOI22_X1 U20070 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20071 ( .A1(n10311), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16886) );
  NAND4_X1 U20072 ( .A1(n16889), .A2(n16888), .A3(n16887), .A4(n16886), .ZN(
        n16895) );
  AOI22_X1 U20073 ( .A1(n16940), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20074 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16892) );
  AOI22_X1 U20075 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16939), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20076 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16890) );
  NAND4_X1 U20077 ( .A1(n16893), .A2(n16892), .A3(n16891), .A4(n16890), .ZN(
        n16894) );
  NOR2_X1 U20078 ( .A1(n16895), .A2(n16894), .ZN(n17086) );
  NOR3_X1 U20079 ( .A1(n16896), .A2(n16978), .A3(n16960), .ZN(n16957) );
  NAND3_X1 U20080 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(n16957), .ZN(n16952) );
  NOR2_X1 U20081 ( .A1(n16949), .A2(n16952), .ZN(n16929) );
  NAND2_X1 U20082 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16929), .ZN(n16928) );
  INV_X1 U20083 ( .A(n16928), .ZN(n16910) );
  AND2_X1 U20084 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16910), .ZN(n16912) );
  OAI21_X1 U20085 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n16912), .A(n16969), .ZN(
        n16897) );
  OAI22_X1 U20086 ( .A1(n17086), .A2(n16969), .B1(n16898), .B2(n16897), .ZN(
        P3_U2692) );
  AOI22_X1 U20087 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20088 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16919), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16901) );
  AOI22_X1 U20089 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16921), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16900) );
  AOI22_X1 U20090 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16899) );
  NAND4_X1 U20091 ( .A1(n16902), .A2(n16901), .A3(n16900), .A4(n16899), .ZN(
        n16909) );
  AOI22_X1 U20092 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16907) );
  AOI22_X1 U20093 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10144), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16906) );
  AOI22_X1 U20094 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16905) );
  AOI22_X1 U20095 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16904) );
  NAND4_X1 U20096 ( .A1(n16907), .A2(n16906), .A3(n16905), .A4(n16904), .ZN(
        n16908) );
  NOR2_X1 U20097 ( .A1(n16909), .A2(n16908), .ZN(n17092) );
  OAI21_X1 U20098 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n16910), .A(n16969), .ZN(
        n16911) );
  OAI22_X1 U20099 ( .A1(n17092), .A2(n16969), .B1(n16912), .B2(n16911), .ZN(
        P3_U2693) );
  AOI22_X1 U20100 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n15538), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n9600), .ZN(n16918) );
  AOI22_X1 U20101 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n16913), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16917) );
  AOI22_X1 U20102 ( .A1(n16939), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16916) );
  AOI22_X1 U20103 ( .A1(n16914), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16915) );
  NAND4_X1 U20104 ( .A1(n16918), .A2(n16917), .A3(n16916), .A4(n16915), .ZN(
        n16927) );
  AOI22_X1 U20105 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n16919), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16925) );
  AOI22_X1 U20106 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9604), .ZN(n16924) );
  AOI22_X1 U20107 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U20108 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n16921), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n16933), .ZN(n16922) );
  NAND4_X1 U20109 ( .A1(n16925), .A2(n16924), .A3(n16923), .A4(n16922), .ZN(
        n16926) );
  NOR2_X1 U20110 ( .A1(n16927), .A2(n16926), .ZN(n17093) );
  OAI21_X1 U20111 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n16929), .A(n16928), .ZN(
        n16930) );
  AOI22_X1 U20112 ( .A1(n16982), .A2(n17093), .B1(n16930), .B2(n16969), .ZN(
        P3_U2694) );
  AOI22_X1 U20113 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15538), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16937) );
  AOI22_X1 U20114 ( .A1(n16920), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16936) );
  AOI22_X1 U20115 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U20116 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9609), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16934) );
  NAND4_X1 U20117 ( .A1(n16937), .A2(n16936), .A3(n16935), .A4(n16934), .ZN(
        n16947) );
  AOI22_X1 U20118 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16945) );
  AOI22_X1 U20119 ( .A1(n15524), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16938), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16944) );
  AOI22_X1 U20120 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10299), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20121 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9604), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16942) );
  NAND4_X1 U20122 ( .A1(n16945), .A2(n16944), .A3(n16943), .A4(n16942), .ZN(
        n16946) );
  NOR2_X1 U20123 ( .A1(n16947), .A2(n16946), .ZN(n17101) );
  INV_X1 U20124 ( .A(n16952), .ZN(n16948) );
  OAI33_X1 U20125 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17032), .A3(n16952), .B1(
        n16949), .B2(n16982), .B3(n16948), .ZN(n16950) );
  INV_X1 U20126 ( .A(n16950), .ZN(n16951) );
  OAI21_X1 U20127 ( .B1(n17101), .B2(n16969), .A(n16951), .ZN(P3_U2695) );
  AOI21_X1 U20128 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n16957), .A(
        P3_EBX_REG_7__SCAN_IN), .ZN(n16955) );
  NAND2_X1 U20129 ( .A1(n16969), .A2(n16952), .ZN(n16954) );
  OAI22_X1 U20130 ( .A1(n16955), .A2(n16954), .B1(n16953), .B2(n16969), .ZN(
        P3_U2696) );
  INV_X1 U20131 ( .A(n16957), .ZN(n16961) );
  AOI22_X1 U20132 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16961), .B1(n16957), .B2(
        n16956), .ZN(n16958) );
  AOI22_X1 U20133 ( .A1(n16982), .A2(n16959), .B1(n16958), .B2(n16969), .ZN(
        P3_U2697) );
  NOR2_X1 U20134 ( .A1(n16978), .A2(n16960), .ZN(n16962) );
  OAI21_X1 U20135 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n16962), .A(n16961), .ZN(
        n16963) );
  AOI22_X1 U20136 ( .A1(n16982), .A2(n16964), .B1(n16963), .B2(n16969), .ZN(
        P3_U2698) );
  AND2_X1 U20137 ( .A1(n16965), .A2(n16981), .ZN(n16974) );
  NAND2_X1 U20138 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16974), .ZN(n16968) );
  NAND3_X1 U20139 ( .A1(n16968), .A2(P3_EBX_REG_4__SCAN_IN), .A3(n16969), .ZN(
        n16966) );
  OAI221_X1 U20140 ( .B1(n16968), .B2(P3_EBX_REG_4__SCAN_IN), .C1(n16969), 
        .C2(n16967), .A(n16966), .ZN(P3_U2699) );
  INV_X1 U20141 ( .A(n16968), .ZN(n16972) );
  AOI21_X1 U20142 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n16969), .A(n16974), .ZN(
        n16971) );
  OAI22_X1 U20143 ( .A1(n16972), .A2(n16971), .B1(n16970), .B2(n16969), .ZN(
        P3_U2700) );
  AOI211_X1 U20144 ( .C1(n16982), .C2(n16976), .A(n16975), .B(n16974), .ZN(
        P3_U2701) );
  INV_X1 U20145 ( .A(n16977), .ZN(n16979) );
  AOI222_X1 U20146 ( .A1(n16981), .A2(n16979), .B1(P3_EBX_REG_1__SCAN_IN), 
        .B2(n16978), .C1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .C2(n16982), .ZN(
        n16980) );
  INV_X1 U20147 ( .A(n16980), .ZN(P3_U2702) );
  AOI22_X1 U20148 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n16982), .B1(
        n16981), .B2(n16984), .ZN(n16983) );
  OAI21_X1 U20149 ( .B1(n16985), .B2(n16984), .A(n16983), .ZN(P3_U2703) );
  INV_X1 U20150 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17144) );
  INV_X1 U20151 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17148) );
  INV_X1 U20152 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17154) );
  INV_X1 U20153 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17250) );
  INV_X1 U20154 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17180) );
  NAND3_X1 U20155 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .ZN(n17102) );
  NAND4_X1 U20156 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_1__SCAN_IN), .ZN(n16986) );
  NOR3_X1 U20157 ( .A1(n17197), .A2(n17102), .A3(n16986), .ZN(n17105) );
  NAND2_X1 U20158 ( .A1(n17105), .A2(n16987), .ZN(n17098) );
  INV_X1 U20159 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17245) );
  INV_X1 U20160 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17170) );
  INV_X1 U20161 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17172) );
  INV_X1 U20162 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17178) );
  NOR4_X1 U20163 ( .A1(n17245), .A2(n17170), .A3(n17172), .A4(n17178), .ZN(
        n16988) );
  INV_X1 U20164 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17156) );
  INV_X1 U20165 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17158) );
  NOR2_X1 U20166 ( .A1(n17156), .A2(n17158), .ZN(n16989) );
  NAND4_X1 U20167 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n16989), .ZN(n17031) );
  NAND2_X1 U20168 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17027), .ZN(n17026) );
  NAND2_X1 U20169 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17023), .ZN(n17022) );
  NAND2_X1 U20170 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17003), .ZN(n16998) );
  NAND2_X1 U20171 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n16994), .ZN(n16993) );
  NAND2_X1 U20172 ( .A1(n16993), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n16991) );
  NOR2_X2 U20173 ( .A1(n17993), .A2(n17123), .ZN(n17064) );
  NAND2_X1 U20174 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17064), .ZN(n16990) );
  OAI221_X1 U20175 ( .B1(n16993), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n16991), 
        .C2(n17097), .A(n16990), .ZN(P3_U2704) );
  NOR2_X1 U20176 ( .A1(n16992), .A2(n17123), .ZN(n17065) );
  AOI22_X1 U20177 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17065), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17064), .ZN(n16996) );
  OAI211_X1 U20178 ( .C1(n16994), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17123), .B(
        n16993), .ZN(n16995) );
  OAI211_X1 U20179 ( .C1(n16997), .C2(n17125), .A(n16996), .B(n16995), .ZN(
        P3_U2705) );
  AOI22_X1 U20180 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17065), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17064), .ZN(n17000) );
  OAI211_X1 U20181 ( .C1(n17003), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17123), .B(
        n16998), .ZN(n16999) );
  OAI211_X1 U20182 ( .C1(n17001), .C2(n17125), .A(n17000), .B(n16999), .ZN(
        P3_U2706) );
  INV_X1 U20183 ( .A(n17064), .ZN(n17038) );
  AOI22_X1 U20184 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17065), .B1(n17132), .B2(
        n17002), .ZN(n17006) );
  AOI211_X1 U20185 ( .C1(n17144), .C2(n17008), .A(n17003), .B(n17097), .ZN(
        n17004) );
  INV_X1 U20186 ( .A(n17004), .ZN(n17005) );
  OAI211_X1 U20187 ( .C1(n17038), .C2(n17007), .A(n17006), .B(n17005), .ZN(
        P3_U2707) );
  AOI22_X1 U20188 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17065), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17064), .ZN(n17010) );
  OAI211_X1 U20189 ( .C1(n9686), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17123), .B(
        n17008), .ZN(n17009) );
  OAI211_X1 U20190 ( .C1(n17011), .C2(n17125), .A(n17010), .B(n17009), .ZN(
        P3_U2708) );
  AOI22_X1 U20191 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17064), .B1(n17132), .B2(
        n17012), .ZN(n17015) );
  AOI211_X1 U20192 ( .C1(n17148), .C2(n17016), .A(n9686), .B(n17097), .ZN(
        n17013) );
  INV_X1 U20193 ( .A(n17013), .ZN(n17014) );
  OAI211_X1 U20194 ( .C1(n17058), .C2(n17234), .A(n17015), .B(n17014), .ZN(
        P3_U2709) );
  AOI22_X1 U20195 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17065), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17064), .ZN(n17019) );
  OAI211_X1 U20196 ( .C1(n17017), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17123), .B(
        n17016), .ZN(n17018) );
  OAI211_X1 U20197 ( .C1(n17020), .C2(n17125), .A(n17019), .B(n17018), .ZN(
        P3_U2710) );
  AOI22_X1 U20198 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17064), .B1(n17132), .B2(
        n17021), .ZN(n17025) );
  OAI211_X1 U20199 ( .C1(n17023), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17123), .B(
        n17022), .ZN(n17024) );
  OAI211_X1 U20200 ( .C1(n17058), .C2(n17230), .A(n17025), .B(n17024), .ZN(
        P3_U2711) );
  AOI22_X1 U20201 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17065), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17064), .ZN(n17029) );
  OAI211_X1 U20202 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17027), .A(n17123), .B(
        n17026), .ZN(n17028) );
  OAI211_X1 U20203 ( .C1(n17030), .C2(n17125), .A(n17029), .B(n17028), .ZN(
        P3_U2712) );
  INV_X1 U20204 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17160) );
  NOR2_X1 U20205 ( .A1(n17032), .A2(n17066), .ZN(n17060) );
  NAND2_X1 U20206 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17060), .ZN(n17059) );
  NAND2_X1 U20207 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17055), .ZN(n17054) );
  NAND2_X1 U20208 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17048), .ZN(n17045) );
  INV_X1 U20209 ( .A(n17045), .ZN(n17041) );
  NOR2_X1 U20210 ( .A1(n17097), .A2(n17041), .ZN(n17042) );
  AOI21_X1 U20211 ( .B1(n17129), .B2(n17156), .A(n17042), .ZN(n17037) );
  NOR4_X1 U20212 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17032), .A3(n17066), .A4(
        n17031), .ZN(n17035) );
  OAI22_X1 U20213 ( .A1(n17033), .A2(n17125), .B1(n14953), .B2(n17038), .ZN(
        n17034) );
  AOI211_X1 U20214 ( .C1(n17065), .C2(BUF2_REG_6__SCAN_IN), .A(n17035), .B(
        n17034), .ZN(n17036) );
  OAI21_X1 U20215 ( .B1(n17037), .B2(n17154), .A(n17036), .ZN(P3_U2713) );
  OAI22_X1 U20216 ( .A1(n17039), .A2(n17125), .B1(n17986), .B2(n17038), .ZN(
        n17040) );
  AOI221_X1 U20217 ( .B1(n17042), .B2(P3_EAX_REG_21__SCAN_IN), .C1(n17041), 
        .C2(n17156), .A(n17040), .ZN(n17043) );
  OAI21_X1 U20218 ( .B1(n17987), .B2(n17058), .A(n17043), .ZN(P3_U2714) );
  AOI22_X1 U20219 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17064), .B1(n17132), .B2(
        n17044), .ZN(n17047) );
  OAI211_X1 U20220 ( .C1(n17048), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17123), .B(
        n17045), .ZN(n17046) );
  OAI211_X1 U20221 ( .C1(n17058), .C2(n17982), .A(n17047), .B(n17046), .ZN(
        P3_U2715) );
  AOI22_X1 U20222 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17065), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17064), .ZN(n17051) );
  AOI211_X1 U20223 ( .C1(n17160), .C2(n17054), .A(n17048), .B(n17097), .ZN(
        n17049) );
  INV_X1 U20224 ( .A(n17049), .ZN(n17050) );
  OAI211_X1 U20225 ( .C1(n17052), .C2(n17125), .A(n17051), .B(n17050), .ZN(
        P3_U2716) );
  AOI22_X1 U20226 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17064), .B1(n17132), .B2(
        n17053), .ZN(n17057) );
  OAI211_X1 U20227 ( .C1(n17055), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17123), .B(
        n17054), .ZN(n17056) );
  OAI211_X1 U20228 ( .C1(n17058), .C2(n17974), .A(n17057), .B(n17056), .ZN(
        P3_U2717) );
  AOI22_X1 U20229 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17065), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17064), .ZN(n17062) );
  OAI211_X1 U20230 ( .C1(n17060), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17123), .B(
        n17059), .ZN(n17061) );
  OAI211_X1 U20231 ( .C1(n17063), .C2(n17125), .A(n17062), .B(n17061), .ZN(
        P3_U2718) );
  AOI22_X1 U20232 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17065), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17064), .ZN(n17068) );
  OAI211_X1 U20233 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17070), .A(n17123), .B(
        n17066), .ZN(n17067) );
  OAI211_X1 U20234 ( .C1(n17069), .C2(n17125), .A(n17068), .B(n17067), .ZN(
        P3_U2719) );
  AOI211_X1 U20235 ( .C1(n17250), .C2(n17075), .A(n17097), .B(n17070), .ZN(
        n17071) );
  AOI21_X1 U20236 ( .B1(n17133), .B2(BUF2_REG_15__SCAN_IN), .A(n17071), .ZN(
        n17072) );
  OAI21_X1 U20237 ( .B1(n17073), .B2(n17125), .A(n17072), .ZN(P3_U2720) );
  NAND2_X1 U20238 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .ZN(n17074) );
  NAND3_X1 U20239 ( .A1(n17999), .A2(n17096), .A3(P3_EAX_REG_9__SCAN_IN), .ZN(
        n17089) );
  NOR2_X1 U20240 ( .A1(n17074), .A2(n17089), .ZN(n17088) );
  NAND2_X1 U20241 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17088), .ZN(n17079) );
  NOR2_X1 U20242 ( .A1(n17170), .A2(n17079), .ZN(n17082) );
  OAI211_X1 U20243 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17082), .A(n17123), .B(
        n17075), .ZN(n17077) );
  NAND2_X1 U20244 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17133), .ZN(n17076) );
  OAI211_X1 U20245 ( .C1(n17078), .C2(n17125), .A(n17077), .B(n17076), .ZN(
        P3_U2721) );
  INV_X1 U20246 ( .A(n17079), .ZN(n17085) );
  AOI21_X1 U20247 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17123), .A(n17085), .ZN(
        n17081) );
  OAI222_X1 U20248 ( .A1(n17128), .A2(n17243), .B1(n17082), .B2(n17081), .C1(
        n17125), .C2(n17080), .ZN(P3_U2722) );
  AOI21_X1 U20249 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17123), .A(n17088), .ZN(
        n17084) );
  OAI222_X1 U20250 ( .A1(n17128), .A2(n17238), .B1(n17085), .B2(n17084), .C1(
        n17125), .C2(n17083), .ZN(P3_U2723) );
  INV_X1 U20251 ( .A(n17089), .ZN(n17095) );
  AOI22_X1 U20252 ( .A1(n17095), .A2(P3_EAX_REG_10__SCAN_IN), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n17123), .ZN(n17087) );
  OAI222_X1 U20253 ( .A1(n17128), .A2(n17236), .B1(n17088), .B2(n17087), .C1(
        n17125), .C2(n17086), .ZN(P3_U2724) );
  INV_X1 U20254 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17176) );
  AOI221_X1 U20255 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n17095), .C1(n17176), 
        .C2(n17089), .A(n17097), .ZN(n17090) );
  AOI21_X1 U20256 ( .B1(n17133), .B2(BUF2_REG_10__SCAN_IN), .A(n17090), .ZN(
        n17091) );
  OAI21_X1 U20257 ( .B1(n17092), .B2(n17125), .A(n17091), .ZN(P3_U2725) );
  AOI22_X1 U20258 ( .A1(n17999), .A2(n17096), .B1(P3_EAX_REG_9__SCAN_IN), .B2(
        n17123), .ZN(n17094) );
  OAI222_X1 U20259 ( .A1(n17128), .A2(n17232), .B1(n17095), .B2(n17094), .C1(
        n17125), .C2(n17093), .ZN(P3_U2726) );
  AOI211_X1 U20260 ( .C1(n17180), .C2(n17098), .A(n17097), .B(n17096), .ZN(
        n17099) );
  AOI21_X1 U20261 ( .B1(n17133), .B2(BUF2_REG_8__SCAN_IN), .A(n17099), .ZN(
        n17100) );
  OAI21_X1 U20262 ( .B1(n17101), .B2(n17125), .A(n17100), .ZN(P3_U2727) );
  INV_X1 U20263 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17192) );
  NAND3_X1 U20264 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(n17129), .ZN(n17121) );
  NOR2_X1 U20265 ( .A1(n17192), .A2(n17121), .ZN(n17127) );
  NAND2_X1 U20266 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17127), .ZN(n17114) );
  NOR2_X1 U20267 ( .A1(n17102), .A2(n17114), .ZN(n17110) );
  AOI21_X1 U20268 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17123), .A(n17110), .ZN(
        n17106) );
  AOI22_X1 U20269 ( .A1(n17133), .A2(BUF2_REG_7__SCAN_IN), .B1(n17132), .B2(
        n17103), .ZN(n17104) );
  OAI221_X1 U20270 ( .B1(n17106), .B2(n17105), .C1(n17106), .C2(n17129), .A(
        n17104), .ZN(P3_U2728) );
  NAND2_X1 U20271 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n17107) );
  NOR2_X1 U20272 ( .A1(n17107), .A2(n17114), .ZN(n17113) );
  AOI21_X1 U20273 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17123), .A(n17113), .ZN(
        n17109) );
  OAI222_X1 U20274 ( .A1(n17992), .A2(n17128), .B1(n17110), .B2(n17109), .C1(
        n17125), .C2(n17108), .ZN(P3_U2729) );
  INV_X1 U20275 ( .A(n17114), .ZN(n17120) );
  AOI22_X1 U20276 ( .A1(n17120), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n17123), .ZN(n17112) );
  OAI222_X1 U20277 ( .A1(n17987), .A2(n17128), .B1(n17113), .B2(n17112), .C1(
        n17125), .C2(n17111), .ZN(P3_U2730) );
  INV_X1 U20278 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17188) );
  NOR2_X1 U20279 ( .A1(n17188), .A2(n17114), .ZN(n17117) );
  AOI21_X1 U20280 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17123), .A(n17120), .ZN(
        n17116) );
  OAI222_X1 U20281 ( .A1(n17982), .A2(n17128), .B1(n17117), .B2(n17116), .C1(
        n17125), .C2(n17115), .ZN(P3_U2731) );
  AOI21_X1 U20282 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17123), .A(n17127), .ZN(
        n17119) );
  OAI222_X1 U20283 ( .A1(n17978), .A2(n17128), .B1(n17120), .B2(n17119), .C1(
        n17125), .C2(n17118), .ZN(P3_U2732) );
  INV_X1 U20284 ( .A(n17121), .ZN(n17122) );
  AOI21_X1 U20285 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17123), .A(n17122), .ZN(
        n17126) );
  OAI222_X1 U20286 ( .A1(n17974), .A2(n17128), .B1(n17127), .B2(n17126), .C1(
        n17125), .C2(n17124), .ZN(P3_U2733) );
  NAND2_X1 U20287 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17129), .ZN(n17136) );
  INV_X1 U20288 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17221) );
  AOI21_X1 U20289 ( .B1(n17999), .B2(n17197), .A(n17130), .ZN(n17135) );
  AOI22_X1 U20290 ( .A1(n17133), .A2(BUF2_REG_1__SCAN_IN), .B1(n17132), .B2(
        n17131), .ZN(n17134) );
  OAI221_X1 U20291 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17136), .C1(n17221), 
        .C2(n17135), .A(n17134), .ZN(P3_U2734) );
  NOR2_X2 U20292 ( .A1(n18577), .A2(n18472), .ZN(n18614) );
  NOR2_X4 U20293 ( .A1(n18614), .A2(n17139), .ZN(n17182) );
  AND2_X1 U20294 ( .A1(n17182), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20295 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20296 ( .A1(n18614), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17140) );
  OAI21_X1 U20297 ( .B1(n17218), .B2(n17165), .A(n17140), .ZN(P3_U2737) );
  INV_X1 U20298 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20299 ( .A1(n18614), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17141) );
  OAI21_X1 U20300 ( .B1(n17142), .B2(n17165), .A(n17141), .ZN(P3_U2738) );
  AOI22_X1 U20301 ( .A1(n18614), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17143) );
  OAI21_X1 U20302 ( .B1(n17144), .B2(n17165), .A(n17143), .ZN(P3_U2739) );
  INV_X1 U20303 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U20304 ( .A1(n18614), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17145) );
  OAI21_X1 U20305 ( .B1(n17146), .B2(n17165), .A(n17145), .ZN(P3_U2740) );
  AOI22_X1 U20306 ( .A1(n18614), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17147) );
  OAI21_X1 U20307 ( .B1(n17148), .B2(n17165), .A(n17147), .ZN(P3_U2741) );
  INV_X1 U20308 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20815) );
  AOI22_X1 U20309 ( .A1(n18614), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17149) );
  OAI21_X1 U20310 ( .B1(n20815), .B2(n17165), .A(n17149), .ZN(P3_U2742) );
  INV_X1 U20311 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20312 ( .A1(n18614), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17150) );
  OAI21_X1 U20313 ( .B1(n17151), .B2(n17165), .A(n17150), .ZN(P3_U2743) );
  INV_X1 U20314 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20315 ( .A1(n18614), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17152) );
  OAI21_X1 U20316 ( .B1(n17210), .B2(n17165), .A(n17152), .ZN(P3_U2744) );
  AOI22_X1 U20317 ( .A1(n17194), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17153) );
  OAI21_X1 U20318 ( .B1(n17154), .B2(n17165), .A(n17153), .ZN(P3_U2745) );
  AOI22_X1 U20319 ( .A1(n17194), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17155) );
  OAI21_X1 U20320 ( .B1(n17156), .B2(n17165), .A(n17155), .ZN(P3_U2746) );
  AOI22_X1 U20321 ( .A1(n17194), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17157) );
  OAI21_X1 U20322 ( .B1(n17158), .B2(n17165), .A(n17157), .ZN(P3_U2747) );
  AOI22_X1 U20323 ( .A1(n17194), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17159) );
  OAI21_X1 U20324 ( .B1(n17160), .B2(n17165), .A(n17159), .ZN(P3_U2748) );
  INV_X1 U20325 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20326 ( .A1(n17194), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17161) );
  OAI21_X1 U20327 ( .B1(n17162), .B2(n17165), .A(n17161), .ZN(P3_U2749) );
  INV_X1 U20328 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20329 ( .A1(n17194), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17163) );
  OAI21_X1 U20330 ( .B1(n17203), .B2(n17165), .A(n17163), .ZN(P3_U2750) );
  INV_X1 U20331 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20332 ( .A1(n17194), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17164) );
  OAI21_X1 U20333 ( .B1(n17166), .B2(n17165), .A(n17164), .ZN(P3_U2751) );
  AOI22_X1 U20334 ( .A1(n17194), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17167) );
  OAI21_X1 U20335 ( .B1(n17250), .B2(n17196), .A(n17167), .ZN(P3_U2752) );
  AOI22_X1 U20336 ( .A1(n17194), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17168) );
  OAI21_X1 U20337 ( .B1(n17245), .B2(n17196), .A(n17168), .ZN(P3_U2753) );
  AOI22_X1 U20338 ( .A1(n17194), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17169) );
  OAI21_X1 U20339 ( .B1(n17170), .B2(n17196), .A(n17169), .ZN(P3_U2754) );
  AOI22_X1 U20340 ( .A1(n17194), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17171) );
  OAI21_X1 U20341 ( .B1(n17172), .B2(n17196), .A(n17171), .ZN(P3_U2755) );
  INV_X1 U20342 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20343 ( .A1(n17194), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17173) );
  OAI21_X1 U20344 ( .B1(n17174), .B2(n17196), .A(n17173), .ZN(P3_U2756) );
  AOI22_X1 U20345 ( .A1(n17194), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17175) );
  OAI21_X1 U20346 ( .B1(n17176), .B2(n17196), .A(n17175), .ZN(P3_U2757) );
  AOI22_X1 U20347 ( .A1(n17194), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17177) );
  OAI21_X1 U20348 ( .B1(n17178), .B2(n17196), .A(n17177), .ZN(P3_U2758) );
  AOI22_X1 U20349 ( .A1(n17194), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17179) );
  OAI21_X1 U20350 ( .B1(n17180), .B2(n17196), .A(n17179), .ZN(P3_U2759) );
  INV_X1 U20351 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20352 ( .A1(n17194), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17181) );
  OAI21_X1 U20353 ( .B1(n17228), .B2(n17196), .A(n17181), .ZN(P3_U2760) );
  INV_X1 U20354 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20355 ( .A1(n17194), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17183) );
  OAI21_X1 U20356 ( .B1(n17184), .B2(n17196), .A(n17183), .ZN(P3_U2761) );
  INV_X1 U20357 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17186) );
  AOI22_X1 U20358 ( .A1(n17194), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17185) );
  OAI21_X1 U20359 ( .B1(n17186), .B2(n17196), .A(n17185), .ZN(P3_U2762) );
  AOI22_X1 U20360 ( .A1(n17194), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17187) );
  OAI21_X1 U20361 ( .B1(n17188), .B2(n17196), .A(n17187), .ZN(P3_U2763) );
  INV_X1 U20362 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20363 ( .A1(n17194), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17189) );
  OAI21_X1 U20364 ( .B1(n17190), .B2(n17196), .A(n17189), .ZN(P3_U2764) );
  AOI22_X1 U20365 ( .A1(n17194), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17191) );
  OAI21_X1 U20366 ( .B1(n17192), .B2(n17196), .A(n17191), .ZN(P3_U2765) );
  AOI22_X1 U20367 ( .A1(n17194), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17193) );
  OAI21_X1 U20368 ( .B1(n17221), .B2(n17196), .A(n17193), .ZN(P3_U2766) );
  AOI22_X1 U20369 ( .A1(n17194), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17195) );
  OAI21_X1 U20370 ( .B1(n17197), .B2(n17196), .A(n17195), .ZN(P3_U2767) );
  OAI211_X1 U20371 ( .C1(n18613), .C2(n17971), .A(n17199), .B(n17198), .ZN(
        n17246) );
  AOI22_X1 U20372 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17239), .ZN(n17201) );
  OAI21_X1 U20373 ( .B1(n17964), .B2(n17242), .A(n17201), .ZN(P3_U2768) );
  AOI22_X1 U20374 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17247), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17239), .ZN(n17202) );
  OAI21_X1 U20375 ( .B1(n17203), .B2(n17249), .A(n17202), .ZN(P3_U2769) );
  AOI22_X1 U20376 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17239), .ZN(n17204) );
  OAI21_X1 U20377 ( .B1(n17974), .B2(n17242), .A(n17204), .ZN(P3_U2770) );
  AOI22_X1 U20378 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17239), .ZN(n17205) );
  OAI21_X1 U20379 ( .B1(n17978), .B2(n17242), .A(n17205), .ZN(P3_U2771) );
  AOI22_X1 U20380 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17239), .ZN(n17206) );
  OAI21_X1 U20381 ( .B1(n17982), .B2(n17242), .A(n17206), .ZN(P3_U2772) );
  AOI22_X1 U20382 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17239), .ZN(n17207) );
  OAI21_X1 U20383 ( .B1(n17987), .B2(n17242), .A(n17207), .ZN(P3_U2773) );
  AOI22_X1 U20384 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17239), .ZN(n17208) );
  OAI21_X1 U20385 ( .B1(n17992), .B2(n17242), .A(n17208), .ZN(P3_U2774) );
  AOI22_X1 U20386 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17247), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17239), .ZN(n17209) );
  OAI21_X1 U20387 ( .B1(n17210), .B2(n17249), .A(n17209), .ZN(P3_U2775) );
  AOI22_X1 U20388 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17239), .ZN(n17211) );
  OAI21_X1 U20389 ( .B1(n17230), .B2(n17242), .A(n17211), .ZN(P3_U2776) );
  AOI22_X1 U20390 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17239), .ZN(n17212) );
  OAI21_X1 U20391 ( .B1(n17232), .B2(n17242), .A(n17212), .ZN(P3_U2777) );
  AOI22_X1 U20392 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17239), .ZN(n17213) );
  OAI21_X1 U20393 ( .B1(n17234), .B2(n17242), .A(n17213), .ZN(P3_U2778) );
  AOI22_X1 U20394 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17239), .ZN(n17214) );
  OAI21_X1 U20395 ( .B1(n17236), .B2(n17242), .A(n17214), .ZN(P3_U2779) );
  AOI22_X1 U20396 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17239), .ZN(n17215) );
  OAI21_X1 U20397 ( .B1(n17238), .B2(n17242), .A(n17215), .ZN(P3_U2780) );
  AOI22_X1 U20398 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17240), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17239), .ZN(n17216) );
  OAI21_X1 U20399 ( .B1(n17243), .B2(n17242), .A(n17216), .ZN(P3_U2781) );
  AOI22_X1 U20400 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17247), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17239), .ZN(n17217) );
  OAI21_X1 U20401 ( .B1(n17218), .B2(n17249), .A(n17217), .ZN(P3_U2782) );
  AOI22_X1 U20402 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17239), .ZN(n17219) );
  OAI21_X1 U20403 ( .B1(n17964), .B2(n17242), .A(n17219), .ZN(P3_U2783) );
  AOI22_X1 U20404 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17247), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17239), .ZN(n17220) );
  OAI21_X1 U20405 ( .B1(n17221), .B2(n17249), .A(n17220), .ZN(P3_U2784) );
  AOI22_X1 U20406 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17246), .ZN(n17222) );
  OAI21_X1 U20407 ( .B1(n17974), .B2(n17242), .A(n17222), .ZN(P3_U2785) );
  AOI22_X1 U20408 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17246), .ZN(n17223) );
  OAI21_X1 U20409 ( .B1(n17978), .B2(n17242), .A(n17223), .ZN(P3_U2786) );
  AOI22_X1 U20410 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17246), .ZN(n17224) );
  OAI21_X1 U20411 ( .B1(n17982), .B2(n17242), .A(n17224), .ZN(P3_U2787) );
  AOI22_X1 U20412 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17246), .ZN(n17225) );
  OAI21_X1 U20413 ( .B1(n17987), .B2(n17242), .A(n17225), .ZN(P3_U2788) );
  AOI22_X1 U20414 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17246), .ZN(n17226) );
  OAI21_X1 U20415 ( .B1(n17992), .B2(n17242), .A(n17226), .ZN(P3_U2789) );
  AOI22_X1 U20416 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17247), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17246), .ZN(n17227) );
  OAI21_X1 U20417 ( .B1(n17228), .B2(n17249), .A(n17227), .ZN(P3_U2790) );
  AOI22_X1 U20418 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17246), .ZN(n17229) );
  OAI21_X1 U20419 ( .B1(n17230), .B2(n17242), .A(n17229), .ZN(P3_U2791) );
  AOI22_X1 U20420 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17246), .ZN(n17231) );
  OAI21_X1 U20421 ( .B1(n17232), .B2(n17242), .A(n17231), .ZN(P3_U2792) );
  AOI22_X1 U20422 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17239), .ZN(n17233) );
  OAI21_X1 U20423 ( .B1(n17234), .B2(n17242), .A(n17233), .ZN(P3_U2793) );
  AOI22_X1 U20424 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17239), .ZN(n17235) );
  OAI21_X1 U20425 ( .B1(n17236), .B2(n17242), .A(n17235), .ZN(P3_U2794) );
  AOI22_X1 U20426 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17239), .ZN(n17237) );
  OAI21_X1 U20427 ( .B1(n17238), .B2(n17242), .A(n17237), .ZN(P3_U2795) );
  AOI22_X1 U20428 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17240), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17239), .ZN(n17241) );
  OAI21_X1 U20429 ( .B1(n17243), .B2(n17242), .A(n17241), .ZN(P3_U2796) );
  AOI22_X1 U20430 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17247), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17246), .ZN(n17244) );
  OAI21_X1 U20431 ( .B1(n17245), .B2(n17249), .A(n17244), .ZN(P3_U2797) );
  AOI22_X1 U20432 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17247), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17246), .ZN(n17248) );
  OAI21_X1 U20433 ( .B1(n17250), .B2(n17249), .A(n17248), .ZN(P3_U2798) );
  INV_X1 U20434 ( .A(n17333), .ZN(n17364) );
  NAND2_X1 U20435 ( .A1(n17457), .A2(n17251), .ZN(n17252) );
  OAI211_X1 U20436 ( .C1(n17253), .C2(n17581), .A(n17622), .B(n17252), .ZN(
        n17286) );
  AOI21_X1 U20437 ( .B1(n17364), .B2(n17281), .A(n17286), .ZN(n17278) );
  NAND3_X1 U20438 ( .A1(n17253), .A2(n9726), .A3(n17294), .ZN(n17277) );
  AOI21_X1 U20439 ( .B1(n17278), .B2(n17277), .A(n9727), .ZN(n17256) );
  INV_X1 U20440 ( .A(n17294), .ZN(n17459) );
  NOR3_X1 U20441 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17459), .A3(
        n17254), .ZN(n17255) );
  AOI211_X1 U20442 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17877), .A(n17256), 
        .B(n17255), .ZN(n17266) );
  INV_X1 U20443 ( .A(n17257), .ZN(n17264) );
  NOR2_X1 U20444 ( .A1(n9632), .A2(n17529), .ZN(n17372) );
  OAI22_X1 U20445 ( .A1(n17628), .A2(n17626), .B1(n17638), .B2(n17494), .ZN(
        n17287) );
  NOR2_X1 U20446 ( .A1(n17627), .A2(n17287), .ZN(n17275) );
  NOR3_X1 U20447 ( .A1(n17372), .A2(n17275), .A3(n12521), .ZN(n17260) );
  OAI211_X1 U20448 ( .C1(n17417), .C2(n17267), .A(n17266), .B(n17265), .ZN(
        P3_U2802) );
  NOR2_X1 U20449 ( .A1(n17950), .A2(n18543), .ZN(n17643) );
  OAI21_X1 U20450 ( .B1(n17271), .B2(n17270), .A(n17428), .ZN(n17272) );
  INV_X1 U20451 ( .A(n17272), .ZN(n17273) );
  OR2_X1 U20452 ( .A1(n17646), .A2(n17470), .ZN(n17274) );
  AOI21_X1 U20453 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17280), .A(
        n17279), .ZN(n17655) );
  OAI21_X1 U20454 ( .B1(n17282), .B2(n17991), .A(n17281), .ZN(n17285) );
  AOI21_X1 U20455 ( .B1(n17417), .B2(n17333), .A(n17283), .ZN(n17284) );
  NOR2_X1 U20456 ( .A1(n17950), .A2(n18541), .ZN(n17652) );
  AOI211_X1 U20457 ( .C1(n17286), .C2(n17285), .A(n17284), .B(n17652), .ZN(
        n17289) );
  NAND2_X1 U20458 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17658), .ZN(
        n17635) );
  NOR2_X1 U20459 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17635), .ZN(
        n17647) );
  AOI22_X1 U20460 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17287), .B1(
        n17328), .B2(n17647), .ZN(n17288) );
  OAI211_X1 U20461 ( .C1(n17655), .C2(n17470), .A(n17289), .B(n17288), .ZN(
        P3_U2804) );
  OAI21_X1 U20462 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17291), .A(
        n17290), .ZN(n17668) );
  OAI21_X1 U20463 ( .B1(n17295), .B2(n17991), .A(n17622), .ZN(n17292) );
  AOI21_X1 U20464 ( .B1(n17457), .B2(n17293), .A(n17292), .ZN(n17323) );
  OAI21_X1 U20465 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18472), .A(
        n17323), .ZN(n17314) );
  INV_X1 U20466 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n20866) );
  NAND2_X1 U20467 ( .A1(n17295), .A2(n17294), .ZN(n17312) );
  AOI221_X1 U20468 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n20866), .C2(n17296), .A(
        n17312), .ZN(n17299) );
  OAI22_X1 U20469 ( .A1(n17835), .A2(n18539), .B1(n17417), .B2(n17297), .ZN(
        n17298) );
  AOI211_X1 U20470 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17314), .A(
        n17299), .B(n17298), .ZN(n17307) );
  NOR3_X1 U20471 ( .A1(n17771), .A2(n17300), .A3(n17635), .ZN(n17301) );
  AOI21_X1 U20472 ( .B1(n17302), .B2(n17659), .A(n17301), .ZN(n17665) );
  AOI21_X1 U20473 ( .B1(n17304), .B2(n17428), .A(n17303), .ZN(n17305) );
  XNOR2_X1 U20474 ( .A(n17305), .B(n17659), .ZN(n17664) );
  AOI22_X1 U20475 ( .A1(n9632), .A2(n17665), .B1(n17533), .B2(n17664), .ZN(
        n17306) );
  OAI211_X1 U20476 ( .C1(n17494), .C2(n17668), .A(n17307), .B(n17306), .ZN(
        P3_U2805) );
  AOI21_X1 U20477 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17309), .A(
        n17308), .ZN(n17683) );
  NOR2_X1 U20478 ( .A1(n17950), .A2(n18536), .ZN(n17679) );
  INV_X1 U20479 ( .A(n17310), .ZN(n17311) );
  OAI22_X1 U20480 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17312), .B1(
        n17417), .B2(n17311), .ZN(n17313) );
  AOI211_X1 U20481 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17314), .A(
        n17679), .B(n17313), .ZN(n17317) );
  INV_X1 U20482 ( .A(n17315), .ZN(n17669) );
  OAI22_X1 U20483 ( .A1(n17670), .A2(n17626), .B1(n17669), .B2(n17494), .ZN(
        n17327) );
  NOR2_X1 U20484 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n20785), .ZN(
        n17681) );
  AOI22_X1 U20485 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17327), .B1(
        n17328), .B2(n17681), .ZN(n17316) );
  OAI211_X1 U20486 ( .C1(n17683), .C2(n17470), .A(n17317), .B(n17316), .ZN(
        P3_U2806) );
  AOI22_X1 U20487 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17428), .B1(
        n17318), .B2(n17340), .ZN(n17319) );
  NAND2_X1 U20488 ( .A1(n17362), .A2(n17319), .ZN(n17320) );
  XNOR2_X1 U20489 ( .A(n17320), .B(n20785), .ZN(n17688) );
  NOR2_X1 U20490 ( .A1(n17459), .A2(n17332), .ZN(n17357) );
  NAND2_X1 U20491 ( .A1(n17335), .A2(n17357), .ZN(n17325) );
  AOI22_X1 U20492 ( .A1(n17877), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17475), 
        .B2(n17321), .ZN(n17322) );
  OAI221_X1 U20493 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17325), .C1(
        n17324), .C2(n17323), .A(n17322), .ZN(n17326) );
  AOI221_X1 U20494 ( .B1(n17328), .B2(n20785), .C1(n17327), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17326), .ZN(n17329) );
  OAI21_X1 U20495 ( .B1(n17470), .B2(n17688), .A(n17329), .ZN(P3_U2807) );
  INV_X1 U20496 ( .A(n17622), .ZN(n17589) );
  AND2_X1 U20497 ( .A1(n17330), .A2(n17457), .ZN(n17331) );
  AOI211_X1 U20498 ( .C1(n17453), .C2(n17332), .A(n17589), .B(n17331), .ZN(
        n17365) );
  OAI21_X1 U20499 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17333), .A(
        n17365), .ZN(n17356) );
  AOI22_X1 U20500 ( .A1(n17475), .A2(n17334), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17356), .ZN(n17348) );
  AOI21_X1 U20501 ( .B1(n20869), .B2(n17336), .A(n17335), .ZN(n17337) );
  AOI22_X1 U20502 ( .A1(n17877), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17357), 
        .B2(n17337), .ZN(n17347) );
  NOR2_X1 U20503 ( .A1(n17338), .A2(n17341), .ZN(n17695) );
  NOR2_X1 U20504 ( .A1(n17691), .A2(n17494), .ZN(n17423) );
  AOI21_X1 U20505 ( .B1(n9632), .B2(n17771), .A(n17423), .ZN(n17421) );
  OAI21_X1 U20506 ( .B1(n17372), .B2(n17695), .A(n17421), .ZN(n17359) );
  INV_X1 U20507 ( .A(n17362), .ZN(n17339) );
  AOI221_X1 U20508 ( .B1(n17341), .B2(n17340), .C1(n17349), .C2(n17340), .A(
        n17339), .ZN(n17342) );
  XOR2_X1 U20509 ( .A(n17342), .B(n17700), .Z(n17706) );
  INV_X1 U20510 ( .A(n17706), .ZN(n17343) );
  AOI22_X1 U20511 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17359), .B1(
        n17533), .B2(n17343), .ZN(n17346) );
  INV_X1 U20512 ( .A(n17422), .ZN(n17344) );
  NAND3_X1 U20513 ( .A1(n17344), .A2(n17695), .A3(n17700), .ZN(n17345) );
  NAND4_X1 U20514 ( .A1(n17348), .A2(n17347), .A3(n17346), .A4(n17345), .ZN(
        P3_U2808) );
  INV_X1 U20515 ( .A(n17358), .ZN(n17713) );
  INV_X1 U20516 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17707) );
  NOR3_X1 U20517 ( .A1(n17707), .A2(n17428), .A3(n17349), .ZN(n17375) );
  INV_X1 U20518 ( .A(n17394), .ZN(n17376) );
  AOI22_X1 U20519 ( .A1(n17713), .A2(n17375), .B1(n17376), .B2(n17350), .ZN(
        n17352) );
  XNOR2_X1 U20520 ( .A(n17352), .B(n17351), .ZN(n17717) );
  AOI22_X1 U20521 ( .A1(n17877), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17475), 
        .B2(n17353), .ZN(n17354) );
  INV_X1 U20522 ( .A(n17354), .ZN(n17355) );
  AOI221_X1 U20523 ( .B1(n17357), .B2(n20869), .C1(n17356), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17355), .ZN(n17361) );
  NOR2_X1 U20524 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17358), .ZN(
        n17709) );
  NAND2_X1 U20525 ( .A1(n17738), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17630) );
  NOR2_X1 U20526 ( .A1(n17422), .A2(n17630), .ZN(n17386) );
  AOI22_X1 U20527 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17359), .B1(
        n17709), .B2(n17386), .ZN(n17360) );
  OAI211_X1 U20528 ( .C1(n17717), .C2(n17470), .A(n17361), .B(n17360), .ZN(
        P3_U2809) );
  OAI221_X1 U20529 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17393), 
        .C1(n17730), .C2(n17375), .A(n17362), .ZN(n17363) );
  XOR2_X1 U20530 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17363), .Z(
        n17728) );
  INV_X1 U20531 ( .A(n17605), .ZN(n17370) );
  INV_X1 U20532 ( .A(n10407), .ZN(n17367) );
  AOI221_X1 U20533 ( .B1(n17367), .B2(n17366), .C1(n17991), .C2(n17366), .A(
        n17365), .ZN(n17369) );
  INV_X1 U20534 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18528) );
  NOR2_X1 U20535 ( .A1(n17950), .A2(n18528), .ZN(n17368) );
  AOI211_X1 U20536 ( .C1(n17371), .C2(n17370), .A(n17369), .B(n17368), .ZN(
        n17374) );
  NOR2_X1 U20537 ( .A1(n17730), .A2(n17630), .ZN(n17721) );
  OAI21_X1 U20538 ( .B1(n17372), .B2(n17721), .A(n17421), .ZN(n17385) );
  NOR2_X1 U20539 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17730), .ZN(
        n17718) );
  AOI22_X1 U20540 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17385), .B1(
        n17386), .B2(n17718), .ZN(n17373) );
  OAI211_X1 U20541 ( .C1(n17470), .C2(n17728), .A(n17374), .B(n17373), .ZN(
        P3_U2810) );
  AOI21_X1 U20542 ( .B1(n17376), .B2(n17393), .A(n17375), .ZN(n17377) );
  XNOR2_X1 U20543 ( .A(n17377), .B(n17730), .ZN(n17734) );
  AOI21_X1 U20544 ( .B1(n17453), .B2(n17379), .A(n17589), .ZN(n17400) );
  OAI21_X1 U20545 ( .B1(n17378), .B2(n18472), .A(n17400), .ZN(n17390) );
  AOI22_X1 U20546 ( .A1(n17877), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17390), .ZN(n17382) );
  NOR2_X1 U20547 ( .A1(n17459), .A2(n17379), .ZN(n17392) );
  OAI211_X1 U20548 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17392), .B(n17380), .ZN(n17381) );
  OAI211_X1 U20549 ( .C1(n17383), .C2(n17417), .A(n17382), .B(n17381), .ZN(
        n17384) );
  AOI221_X1 U20550 ( .B1(n17386), .B2(n17730), .C1(n17385), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17384), .ZN(n17387) );
  OAI21_X1 U20551 ( .B1(n17734), .B2(n17470), .A(n17387), .ZN(P3_U2811) );
  NAND2_X1 U20552 ( .A1(n17738), .A2(n17707), .ZN(n17746) );
  OAI22_X1 U20553 ( .A1(n17835), .A2(n18524), .B1(n17417), .B2(n17388), .ZN(
        n17389) );
  AOI221_X1 U20554 ( .B1(n17392), .B2(n17391), .C1(n17390), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17389), .ZN(n17397) );
  OAI21_X1 U20555 ( .B1(n17738), .B2(n17422), .A(n17421), .ZN(n17405) );
  AOI21_X1 U20556 ( .B1(n17531), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17393), .ZN(n17395) );
  XNOR2_X1 U20557 ( .A(n17395), .B(n17394), .ZN(n17742) );
  AOI22_X1 U20558 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17405), .B1(
        n17533), .B2(n17742), .ZN(n17396) );
  OAI211_X1 U20559 ( .C1(n17422), .C2(n17746), .A(n17397), .B(n17396), .ZN(
        P3_U2812) );
  NAND2_X1 U20560 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17747), .ZN(
        n17753) );
  AOI21_X1 U20561 ( .B1(n17398), .B2(n18344), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17401) );
  OAI22_X1 U20562 ( .A1(n17401), .A2(n17400), .B1(n17605), .B2(n17399), .ZN(
        n17402) );
  AOI21_X1 U20563 ( .B1(n17940), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17402), 
        .ZN(n17407) );
  OAI21_X1 U20564 ( .B1(n17404), .B2(n17747), .A(n17403), .ZN(n17750) );
  AOI22_X1 U20565 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17405), .B1(
        n17533), .B2(n17750), .ZN(n17406) );
  OAI211_X1 U20566 ( .C1(n17422), .C2(n17753), .A(n17407), .B(n17406), .ZN(
        P3_U2813) );
  AOI21_X1 U20567 ( .B1(n17531), .B2(n17409), .A(n17408), .ZN(n17410) );
  XNOR2_X1 U20568 ( .A(n17410), .B(n17762), .ZN(n17759) );
  INV_X1 U20569 ( .A(n17411), .ZN(n17412) );
  AOI21_X1 U20570 ( .B1(n17453), .B2(n17413), .A(n17589), .ZN(n17440) );
  OAI21_X1 U20571 ( .B1(n17412), .B2(n18472), .A(n17440), .ZN(n17427) );
  AOI22_X1 U20572 ( .A1(n17877), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17427), .ZN(n17416) );
  NOR2_X1 U20573 ( .A1(n17459), .A2(n17413), .ZN(n17426) );
  OAI211_X1 U20574 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17426), .B(n17414), .ZN(n17415) );
  OAI211_X1 U20575 ( .C1(n17418), .C2(n17417), .A(n17416), .B(n17415), .ZN(
        n17419) );
  AOI21_X1 U20576 ( .B1(n17533), .B2(n17759), .A(n17419), .ZN(n17420) );
  OAI221_X1 U20577 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17422), 
        .C1(n17762), .C2(n17421), .A(n17420), .ZN(P3_U2814) );
  INV_X1 U20578 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17774) );
  NAND2_X1 U20579 ( .A1(n17757), .A2(n17495), .ZN(n17441) );
  NAND2_X1 U20580 ( .A1(n17774), .A2(n17441), .ZN(n17768) );
  AOI22_X1 U20581 ( .A1(n17475), .A2(n17424), .B1(n17423), .B2(n17768), .ZN(
        n17434) );
  AOI22_X1 U20582 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17427), .B1(
        n17426), .B2(n17425), .ZN(n17433) );
  INV_X1 U20583 ( .A(n17780), .ZN(n17784) );
  NOR2_X1 U20584 ( .A1(n17428), .A2(n17818), .ZN(n17511) );
  INV_X1 U20585 ( .A(n17511), .ZN(n17503) );
  NOR2_X1 U20586 ( .A1(n17784), .A2(n17503), .ZN(n17442) );
  NOR2_X1 U20587 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17809), .ZN(
        n17796) );
  INV_X1 U20588 ( .A(n17796), .ZN(n17465) );
  OAI221_X1 U20589 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17443), 
        .C1(n20872), .C2(n17442), .A(n17465), .ZN(n17429) );
  XNOR2_X1 U20590 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17429), .ZN(
        n17776) );
  NOR2_X1 U20591 ( .A1(n17430), .A2(n17626), .ZN(n17431) );
  NOR2_X1 U20592 ( .A1(n17820), .A2(n17784), .ZN(n17802) );
  NAND3_X1 U20593 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n17802), .ZN(n17435) );
  NAND2_X1 U20594 ( .A1(n17774), .A2(n17435), .ZN(n17770) );
  AOI22_X1 U20595 ( .A1(n17533), .A2(n17776), .B1(n17431), .B2(n17770), .ZN(
        n17432) );
  NAND2_X1 U20596 ( .A1(n17877), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17773) );
  NAND4_X1 U20597 ( .A1(n17434), .A2(n17433), .A3(n17432), .A4(n17773), .ZN(
        P3_U2815) );
  INV_X1 U20598 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17783) );
  INV_X1 U20599 ( .A(n17802), .ZN(n17464) );
  NOR2_X1 U20600 ( .A1(n17783), .A2(n17464), .ZN(n17436) );
  OAI21_X1 U20601 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17436), .A(
        n17435), .ZN(n17795) );
  NOR2_X1 U20602 ( .A1(n17458), .A2(n17991), .ZN(n17490) );
  AOI21_X1 U20603 ( .B1(n17437), .B2(n17490), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17439) );
  OAI22_X1 U20604 ( .A1(n17440), .A2(n17439), .B1(n17605), .B2(n17438), .ZN(
        n17446) );
  INV_X1 U20605 ( .A(n17765), .ZN(n17781) );
  OAI221_X1 U20606 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17781), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17495), .A(n17441), .ZN(
        n17790) );
  OAI21_X1 U20607 ( .B1(n17443), .B2(n17442), .A(n17465), .ZN(n17444) );
  XNOR2_X1 U20608 ( .A(n17444), .B(n20872), .ZN(n17789) );
  OAI22_X1 U20609 ( .A1(n17494), .A2(n17790), .B1(n17470), .B2(n17789), .ZN(
        n17445) );
  AOI211_X1 U20610 ( .C1(n17940), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17446), 
        .B(n17445), .ZN(n17447) );
  OAI21_X1 U20611 ( .B1(n17626), .B2(n17795), .A(n17447), .ZN(P3_U2816) );
  INV_X1 U20612 ( .A(n17471), .ZN(n17450) );
  OAI22_X1 U20613 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17531), .B1(
        n17448), .B2(n17784), .ZN(n17449) );
  OAI21_X1 U20614 ( .B1(n17531), .B2(n17450), .A(n17449), .ZN(n17451) );
  XOR2_X1 U20615 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17451), .Z(
        n17808) );
  AOI21_X1 U20616 ( .B1(n17453), .B2(n17452), .A(n17589), .ZN(n17544) );
  OAI21_X1 U20617 ( .B1(n17454), .B2(n17581), .A(n17544), .ZN(n17455) );
  AOI21_X1 U20618 ( .B1(n17457), .B2(n17456), .A(n17455), .ZN(n17478) );
  NOR2_X1 U20619 ( .A1(n17459), .A2(n17458), .ZN(n17473) );
  OAI211_X1 U20620 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17473), .B(n17460), .ZN(n17462) );
  NAND2_X1 U20621 ( .A1(n17940), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17461) );
  OAI211_X1 U20622 ( .C1(n17478), .C2(n17463), .A(n17462), .B(n17461), .ZN(
        n17467) );
  NAND2_X1 U20623 ( .A1(n17780), .A2(n17495), .ZN(n17799) );
  AOI22_X1 U20624 ( .A1(n9632), .A2(n17464), .B1(n17529), .B2(n17799), .ZN(
        n17481) );
  INV_X1 U20625 ( .A(n17798), .ZN(n17829) );
  NAND2_X1 U20626 ( .A1(n17829), .A2(n17483), .ZN(n17482) );
  OAI22_X1 U20627 ( .A1(n17481), .A2(n17783), .B1(n17465), .B2(n17482), .ZN(
        n17466) );
  AOI211_X1 U20628 ( .C1(n17475), .C2(n17468), .A(n17467), .B(n17466), .ZN(
        n17469) );
  OAI21_X1 U20629 ( .B1(n17470), .B2(n17808), .A(n17469), .ZN(P3_U2817) );
  NAND2_X1 U20630 ( .A1(n17827), .A2(n17511), .ZN(n17484) );
  OAI21_X1 U20631 ( .B1(n17485), .B2(n17484), .A(n17471), .ZN(n17472) );
  XNOR2_X1 U20632 ( .A(n17472), .B(n17809), .ZN(n17812) );
  AOI22_X1 U20633 ( .A1(n17475), .A2(n17474), .B1(n17473), .B2(n17477), .ZN(
        n17476) );
  NAND2_X1 U20634 ( .A1(n17877), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17813) );
  OAI211_X1 U20635 ( .C1(n17478), .C2(n17477), .A(n17476), .B(n17813), .ZN(
        n17479) );
  AOI21_X1 U20636 ( .B1(n17533), .B2(n17812), .A(n17479), .ZN(n17480) );
  OAI221_X1 U20637 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17482), 
        .C1(n17809), .C2(n17481), .A(n17480), .ZN(P3_U2818) );
  INV_X1 U20638 ( .A(n17483), .ZN(n17521) );
  NAND2_X1 U20639 ( .A1(n17827), .A2(n17485), .ZN(n17833) );
  OAI21_X1 U20640 ( .B1(n17502), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17484), .ZN(n17486) );
  XNOR2_X1 U20641 ( .A(n17486), .B(n17485), .ZN(n17817) );
  NOR2_X1 U20642 ( .A1(n17950), .A2(n18510), .ZN(n17492) );
  NAND2_X1 U20643 ( .A1(n10413), .A2(n18344), .ZN(n17556) );
  NOR2_X1 U20644 ( .A1(n17555), .A2(n17556), .ZN(n17538) );
  NAND2_X1 U20645 ( .A1(n17487), .A2(n17538), .ZN(n17513) );
  NOR2_X1 U20646 ( .A1(n17499), .A2(n17513), .ZN(n17498) );
  AOI21_X1 U20647 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17551), .A(
        n17498), .ZN(n17489) );
  OAI22_X1 U20648 ( .A1(n17490), .A2(n17489), .B1(n17605), .B2(n17488), .ZN(
        n17491) );
  AOI211_X1 U20649 ( .C1(n17533), .C2(n17817), .A(n17492), .B(n17491), .ZN(
        n17497) );
  NOR2_X1 U20650 ( .A1(n17827), .A2(n17521), .ZN(n17505) );
  OAI22_X1 U20651 ( .A1(n17495), .A2(n17494), .B1(n17626), .B2(n17493), .ZN(
        n17510) );
  OAI21_X1 U20652 ( .B1(n17505), .B2(n17510), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17496) );
  OAI211_X1 U20653 ( .C1(n17521), .C2(n17833), .A(n17497), .B(n17496), .ZN(
        P3_U2819) );
  INV_X1 U20654 ( .A(n17551), .ZN(n17618) );
  AOI211_X1 U20655 ( .C1(n17513), .C2(n17499), .A(n17618), .B(n17498), .ZN(
        n17500) );
  AOI21_X1 U20656 ( .B1(n17501), .B2(n17370), .A(n17500), .ZN(n17509) );
  OAI21_X1 U20657 ( .B1(n17847), .B2(n17503), .A(n17502), .ZN(n17504) );
  XNOR2_X1 U20658 ( .A(n17504), .B(n17841), .ZN(n17838) );
  AOI22_X1 U20659 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17510), .B1(
        n17533), .B2(n17838), .ZN(n17508) );
  NAND2_X1 U20660 ( .A1(n17940), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17507) );
  OAI21_X1 U20661 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17505), .ZN(n17506) );
  NAND4_X1 U20662 ( .A1(n17509), .A2(n17508), .A3(n17507), .A4(n17506), .ZN(
        P3_U2820) );
  INV_X1 U20663 ( .A(n17510), .ZN(n17520) );
  NOR2_X1 U20664 ( .A1(n17511), .A2(n9714), .ZN(n17512) );
  XNOR2_X1 U20665 ( .A(n17512), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17844) );
  NOR2_X1 U20666 ( .A1(n17950), .A2(n18506), .ZN(n17518) );
  INV_X1 U20667 ( .A(n17513), .ZN(n17516) );
  AOI22_X1 U20668 ( .A1(n17538), .A2(n17524), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17551), .ZN(n17515) );
  OAI22_X1 U20669 ( .A1(n17516), .A2(n17515), .B1(n17605), .B2(n17514), .ZN(
        n17517) );
  AOI211_X1 U20670 ( .C1(n17533), .C2(n17844), .A(n17518), .B(n17517), .ZN(
        n17519) );
  OAI221_X1 U20671 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17521), .C1(
        n17847), .C2(n17520), .A(n17519), .ZN(P3_U2821) );
  OAI21_X1 U20672 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17523), .A(
        n17522), .ZN(n17867) );
  NAND2_X1 U20673 ( .A1(n16532), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17525) );
  AOI211_X1 U20674 ( .C1(n17526), .C2(n17525), .A(n17524), .B(n17991), .ZN(
        n17528) );
  OAI22_X1 U20675 ( .A1(n17544), .A2(n17526), .B1(n17950), .B2(n18505), .ZN(
        n17527) );
  AOI211_X1 U20676 ( .C1(n17864), .C2(n17529), .A(n17528), .B(n17527), .ZN(
        n17535) );
  OAI21_X1 U20677 ( .B1(n17531), .B2(n17864), .A(n17530), .ZN(n17861) );
  AOI22_X1 U20678 ( .A1(n17533), .A2(n17861), .B1(n17532), .B2(n17370), .ZN(
        n17534) );
  OAI211_X1 U20679 ( .C1(n17626), .C2(n17867), .A(n17535), .B(n17534), .ZN(
        P3_U2822) );
  AOI21_X1 U20680 ( .B1(n17542), .B2(n17537), .A(n17536), .ZN(n17872) );
  AOI22_X1 U20681 ( .A1(n17614), .A2(n17872), .B1(n17538), .B2(n20781), .ZN(
        n17548) );
  AOI21_X1 U20682 ( .B1(n17541), .B2(n17540), .A(n17539), .ZN(n17543) );
  XNOR2_X1 U20683 ( .A(n17543), .B(n17542), .ZN(n17873) );
  OAI22_X1 U20684 ( .A1(n17605), .A2(n17545), .B1(n17544), .B2(n20781), .ZN(
        n17546) );
  AOI21_X1 U20685 ( .B1(n9632), .B2(n17873), .A(n17546), .ZN(n17547) );
  OAI211_X1 U20686 ( .C1(n17950), .C2(n18502), .A(n17548), .B(n17547), .ZN(
        P3_U2823) );
  OAI21_X1 U20687 ( .B1(n17550), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17549), .ZN(n17884) );
  NAND2_X1 U20688 ( .A1(n17551), .A2(n17556), .ZN(n17568) );
  AOI21_X1 U20689 ( .B1(n17553), .B2(n17552), .A(n9712), .ZN(n17876) );
  AOI22_X1 U20690 ( .A1(n17614), .A2(n17876), .B1(n17940), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n17554) );
  OAI221_X1 U20691 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17556), .C1(
        n17555), .C2(n17568), .A(n17554), .ZN(n17557) );
  AOI21_X1 U20692 ( .B1(n17558), .B2(n17370), .A(n17557), .ZN(n17559) );
  OAI21_X1 U20693 ( .B1(n17626), .B2(n17884), .A(n17559), .ZN(P3_U2824) );
  OAI21_X1 U20694 ( .B1(n17562), .B2(n17561), .A(n17560), .ZN(n17891) );
  OAI21_X1 U20695 ( .B1(n17565), .B2(n17564), .A(n17563), .ZN(n17566) );
  XNOR2_X1 U20696 ( .A(n17566), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17887) );
  AOI21_X1 U20697 ( .B1(n17567), .B2(n17622), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17569) );
  OAI22_X1 U20698 ( .A1(n17605), .A2(n17570), .B1(n17569), .B2(n17568), .ZN(
        n17571) );
  AOI21_X1 U20699 ( .B1(n17614), .B2(n17887), .A(n17571), .ZN(n17572) );
  NAND2_X1 U20700 ( .A1(n17877), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n17885) );
  OAI211_X1 U20701 ( .C1(n17626), .C2(n17891), .A(n17572), .B(n17885), .ZN(
        P3_U2825) );
  OAI21_X1 U20702 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17574), .A(
        n17573), .ZN(n17903) );
  INV_X1 U20703 ( .A(n17575), .ZN(n17576) );
  OAI22_X1 U20704 ( .A1(n17626), .A2(n17903), .B1(n17991), .B2(n17576), .ZN(
        n17577) );
  AOI21_X1 U20705 ( .B1(n17940), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17577), .ZN(
        n17584) );
  AOI21_X1 U20706 ( .B1(n17580), .B2(n17579), .A(n17578), .ZN(n17892) );
  OAI21_X1 U20707 ( .B1(n17582), .B2(n17581), .A(n17622), .ZN(n17596) );
  AOI22_X1 U20708 ( .A1(n17614), .A2(n17892), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17596), .ZN(n17583) );
  OAI211_X1 U20709 ( .C1(n17605), .C2(n17585), .A(n17584), .B(n17583), .ZN(
        P3_U2826) );
  OAI21_X1 U20710 ( .B1(n17588), .B2(n17587), .A(n17586), .ZN(n17904) );
  NOR2_X1 U20711 ( .A1(n17589), .A2(n17608), .ZN(n17609) );
  OAI21_X1 U20712 ( .B1(n17592), .B2(n17591), .A(n17590), .ZN(n17593) );
  XNOR2_X1 U20713 ( .A(n17593), .B(n17905), .ZN(n17912) );
  OAI22_X1 U20714 ( .A1(n17605), .A2(n17594), .B1(n17625), .B2(n17912), .ZN(
        n17595) );
  AOI221_X1 U20715 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17596), .C1(
        n17609), .C2(n17596), .A(n17595), .ZN(n17597) );
  NAND2_X1 U20716 ( .A1(n17940), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n17910) );
  OAI211_X1 U20717 ( .C1(n17626), .C2(n17904), .A(n17597), .B(n17910), .ZN(
        P3_U2827) );
  AOI21_X1 U20718 ( .B1(n17600), .B2(n17599), .A(n17598), .ZN(n17916) );
  NOR2_X1 U20719 ( .A1(n17950), .A2(n18492), .ZN(n17915) );
  OAI21_X1 U20720 ( .B1(n17603), .B2(n17602), .A(n17601), .ZN(n17931) );
  OAI22_X1 U20721 ( .A1(n17605), .A2(n17604), .B1(n17626), .B2(n17931), .ZN(
        n17606) );
  AOI211_X1 U20722 ( .C1(n17614), .C2(n17916), .A(n17915), .B(n17606), .ZN(
        n17607) );
  OAI221_X1 U20723 ( .B1(n17609), .B2(n17608), .C1(n17609), .C2(n17991), .A(
        n17607), .ZN(P3_U2828) );
  NOR2_X1 U20724 ( .A1(n17620), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17610) );
  XNOR2_X1 U20725 ( .A(n17610), .B(n17613), .ZN(n17939) );
  AOI22_X1 U20726 ( .A1(n9632), .A2(n17939), .B1(n17940), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17616) );
  AOI21_X1 U20727 ( .B1(n17613), .B2(n17619), .A(n17612), .ZN(n17932) );
  AOI22_X1 U20728 ( .A1(n17614), .A2(n17932), .B1(n17617), .B2(n17370), .ZN(
        n17615) );
  OAI211_X1 U20729 ( .C1(n17618), .C2(n17617), .A(n17616), .B(n17615), .ZN(
        P3_U2829) );
  OAI21_X1 U20730 ( .B1(n17620), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17619), .ZN(n17946) );
  INV_X1 U20731 ( .A(n17946), .ZN(n17948) );
  INV_X1 U20732 ( .A(n17621), .ZN(n18464) );
  OAI21_X1 U20733 ( .B1(n18464), .B2(n18625), .A(n17622), .ZN(n17623) );
  AOI22_X1 U20734 ( .A1(n17877), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17623), .ZN(n17624) );
  OAI221_X1 U20735 ( .B1(n17948), .B2(n17626), .C1(n17946), .C2(n17625), .A(
        n17624), .ZN(P3_U2830) );
  AOI221_X1 U20736 ( .B1(n17634), .B2(n17627), .C1(n17684), .C2(n17627), .A(
        n17951), .ZN(n17642) );
  INV_X1 U20737 ( .A(n17628), .ZN(n17640) );
  INV_X1 U20738 ( .A(n17922), .ZN(n17850) );
  INV_X1 U20739 ( .A(n17629), .ZN(n17633) );
  INV_X1 U20740 ( .A(n18427), .ZN(n18417) );
  INV_X1 U20741 ( .A(n17689), .ZN(n17632) );
  OAI21_X1 U20742 ( .B1(n17755), .B2(n17630), .A(n18417), .ZN(n17631) );
  INV_X1 U20743 ( .A(n17631), .ZN(n17711) );
  AOI21_X1 U20744 ( .B1(n18417), .B2(n17632), .A(n17711), .ZN(n17697) );
  OAI21_X1 U20745 ( .B1(n17850), .B2(n17633), .A(n17697), .ZN(n17672) );
  AOI22_X1 U20746 ( .A1(n17952), .A2(n17635), .B1(n18417), .B2(n17634), .ZN(
        n17636) );
  OAI211_X1 U20747 ( .C1(n17638), .C2(n17690), .A(n17637), .B(n17636), .ZN(
        n17639) );
  AOI211_X1 U20748 ( .C1(n18399), .C2(n17640), .A(n17672), .B(n17639), .ZN(
        n17650) );
  OAI211_X1 U20749 ( .C1(n9629), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17650), .ZN(n17641) );
  AOI22_X1 U20750 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17896), .B1(
        n17642), .B2(n17641), .ZN(n17645) );
  INV_X1 U20751 ( .A(n17643), .ZN(n17644) );
  OAI211_X1 U20752 ( .C1(n17646), .C2(n17807), .A(n17645), .B(n17644), .ZN(
        P3_U2835) );
  INV_X1 U20753 ( .A(n17647), .ZN(n17648) );
  OAI22_X1 U20754 ( .A1(n17650), .A2(n17649), .B1(n17684), .B2(n17648), .ZN(
        n17651) );
  AOI22_X1 U20755 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17896), .B1(
        n17934), .B2(n17651), .ZN(n17654) );
  INV_X1 U20756 ( .A(n17652), .ZN(n17653) );
  OAI211_X1 U20757 ( .C1(n17655), .C2(n17807), .A(n17654), .B(n17653), .ZN(
        P3_U2836) );
  INV_X1 U20758 ( .A(n17863), .ZN(n17791) );
  NOR2_X1 U20759 ( .A1(n17950), .A2(n18539), .ZN(n17663) );
  AOI211_X1 U20760 ( .C1(n17855), .C2(n17656), .A(n17673), .B(n17672), .ZN(
        n17661) );
  NAND2_X1 U20761 ( .A1(n17658), .A2(n17657), .ZN(n17660) );
  AOI221_X1 U20762 ( .B1(n17661), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17660), .C2(n17659), .A(n17951), .ZN(n17662) );
  AOI211_X1 U20763 ( .C1(n17896), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17663), .B(n17662), .ZN(n17667) );
  AOI22_X1 U20764 ( .A1(n17947), .A2(n17665), .B1(n17862), .B2(n17664), .ZN(
        n17666) );
  OAI211_X1 U20765 ( .C1(n17791), .C2(n17668), .A(n17667), .B(n17666), .ZN(
        P3_U2837) );
  OAI22_X1 U20766 ( .A1(n17670), .A2(n17801), .B1(n17669), .B2(n17690), .ZN(
        n17671) );
  NOR3_X1 U20767 ( .A1(n17896), .A2(n17672), .A3(n17671), .ZN(n17677) );
  NOR2_X1 U20768 ( .A1(n17673), .A2(n20785), .ZN(n17674) );
  AOI21_X1 U20769 ( .B1(n17677), .B2(n17674), .A(n17940), .ZN(n17686) );
  INV_X1 U20770 ( .A(n17686), .ZN(n17675) );
  AOI211_X1 U20771 ( .C1(n17897), .C2(n17677), .A(n17676), .B(n17675), .ZN(
        n17678) );
  AOI211_X1 U20772 ( .C1(n17681), .C2(n17680), .A(n17679), .B(n17678), .ZN(
        n17682) );
  OAI21_X1 U20773 ( .B1(n17683), .B2(n17807), .A(n17682), .ZN(P3_U2838) );
  OAI21_X1 U20774 ( .B1(n17896), .B2(n17684), .A(n20785), .ZN(n17685) );
  AOI22_X1 U20775 ( .A1(n17877), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17686), 
        .B2(n17685), .ZN(n17687) );
  OAI21_X1 U20776 ( .B1(n17807), .B2(n17688), .A(n17687), .ZN(P3_U2839) );
  NAND2_X1 U20777 ( .A1(n17940), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17705) );
  OAI22_X1 U20778 ( .A1(n9629), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n17689), .B2(n17919), .ZN(n17699) );
  NOR2_X1 U20779 ( .A1(n17691), .A2(n17690), .ZN(n17769) );
  AOI21_X1 U20780 ( .B1(n18399), .B2(n17771), .A(n17769), .ZN(n17710) );
  INV_X1 U20781 ( .A(n17692), .ZN(n17741) );
  OAI21_X1 U20782 ( .B1(n17707), .B2(n17741), .A(n18438), .ZN(n17693) );
  OAI221_X1 U20783 ( .B1(n9629), .B2(n17694), .C1(n9629), .C2(n17721), .A(
        n17693), .ZN(n17719) );
  NOR2_X1 U20784 ( .A1(n18399), .A2(n17819), .ZN(n17826) );
  OAI22_X1 U20785 ( .A1(n9629), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17695), .B2(n17826), .ZN(n17696) );
  NOR2_X1 U20786 ( .A1(n17719), .A2(n17696), .ZN(n17712) );
  NAND3_X1 U20787 ( .A1(n17697), .A2(n17710), .A3(n17712), .ZN(n17698) );
  NOR3_X1 U20788 ( .A1(n17700), .A2(n17699), .A3(n17698), .ZN(n17701) );
  INV_X1 U20789 ( .A(n17896), .ZN(n17935) );
  OAI22_X1 U20790 ( .A1(n17701), .A2(n17951), .B1(n17700), .B2(n17935), .ZN(
        n17702) );
  OAI21_X1 U20791 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17703), .A(
        n17702), .ZN(n17704) );
  OAI211_X1 U20792 ( .C1(n17706), .C2(n17807), .A(n17705), .B(n17704), .ZN(
        P3_U2840) );
  NOR3_X1 U20793 ( .A1(n17708), .A2(n17951), .A3(n17707), .ZN(n17731) );
  AOI22_X1 U20794 ( .A1(n17877), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17709), 
        .B2(n17731), .ZN(n17716) );
  NOR2_X1 U20795 ( .A1(n18438), .A2(n18417), .ZN(n17779) );
  NAND2_X1 U20796 ( .A1(n17934), .A2(n17710), .ZN(n17758) );
  NOR2_X1 U20797 ( .A1(n17711), .A2(n17758), .ZN(n17724) );
  OAI211_X1 U20798 ( .C1(n17713), .C2(n17779), .A(n17724), .B(n17712), .ZN(
        n17714) );
  NAND3_X1 U20799 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17950), .A3(
        n17714), .ZN(n17715) );
  OAI211_X1 U20800 ( .C1(n17717), .C2(n17807), .A(n17716), .B(n17715), .ZN(
        P3_U2841) );
  AOI22_X1 U20801 ( .A1(n17877), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17731), 
        .B2(n17718), .ZN(n17727) );
  INV_X1 U20802 ( .A(n17719), .ZN(n17720) );
  OAI21_X1 U20803 ( .B1(n17721), .B2(n17826), .A(n17720), .ZN(n17722) );
  INV_X1 U20804 ( .A(n17722), .ZN(n17723) );
  AOI21_X1 U20805 ( .B1(n17724), .B2(n17723), .A(n17940), .ZN(n17732) );
  NOR3_X1 U20806 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17779), .A3(
        n18631), .ZN(n17725) );
  OAI21_X1 U20807 ( .B1(n17732), .B2(n17725), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17726) );
  OAI211_X1 U20808 ( .C1(n17807), .C2(n17728), .A(n17727), .B(n17726), .ZN(
        P3_U2842) );
  NOR2_X1 U20809 ( .A1(n17950), .A2(n18526), .ZN(n17729) );
  AOI221_X1 U20810 ( .B1(n17732), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), 
        .C1(n17731), .C2(n17730), .A(n17729), .ZN(n17733) );
  OAI21_X1 U20811 ( .B1(n17734), .B2(n17807), .A(n17733), .ZN(P3_U2843) );
  AOI22_X1 U20812 ( .A1(n17893), .A2(n18438), .B1(n17851), .B2(n17917), .ZN(
        n17856) );
  INV_X1 U20813 ( .A(n17856), .ZN(n17908) );
  NAND2_X1 U20814 ( .A1(n17735), .A2(n17908), .ZN(n17764) );
  AOI21_X1 U20815 ( .B1(n17736), .B2(n17764), .A(n17951), .ZN(n17834) );
  NAND2_X1 U20816 ( .A1(n10214), .A2(n17834), .ZN(n17763) );
  NOR2_X1 U20817 ( .A1(n18427), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17920) );
  NOR3_X1 U20818 ( .A1(n17920), .A2(n17737), .A3(n17762), .ZN(n17739) );
  OAI22_X1 U20819 ( .A1(n17850), .A2(n17739), .B1(n17738), .B2(n17826), .ZN(
        n17740) );
  AOI211_X1 U20820 ( .C1(n18438), .C2(n17741), .A(n17758), .B(n17740), .ZN(
        n17748) );
  AOI221_X1 U20821 ( .B1(n17850), .B2(n17748), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17748), .A(n17877), .ZN(
        n17743) );
  AOI22_X1 U20822 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17743), .B1(
        n17862), .B2(n17742), .ZN(n17745) );
  NAND2_X1 U20823 ( .A1(n17940), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17744) );
  OAI211_X1 U20824 ( .C1(n17746), .C2(n17763), .A(n17745), .B(n17744), .ZN(
        P3_U2844) );
  NOR3_X1 U20825 ( .A1(n17877), .A2(n17748), .A3(n17747), .ZN(n17749) );
  AOI21_X1 U20826 ( .B1(n17862), .B2(n17750), .A(n17749), .ZN(n17752) );
  NAND2_X1 U20827 ( .A1(n17940), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17751) );
  OAI211_X1 U20828 ( .C1(n17753), .C2(n17763), .A(n17752), .B(n17751), .ZN(
        P3_U2845) );
  AOI22_X1 U20829 ( .A1(n18438), .A2(n17754), .B1(n17952), .B2(n17821), .ZN(
        n17824) );
  OAI21_X1 U20830 ( .B1(n17774), .B2(n18417), .A(n17755), .ZN(n17756) );
  OAI211_X1 U20831 ( .C1(n17757), .C2(n17828), .A(n17824), .B(n17756), .ZN(
        n17766) );
  OAI221_X1 U20832 ( .B1(n17758), .B2(n17855), .C1(n17758), .C2(n17766), .A(
        n17835), .ZN(n17761) );
  AOI22_X1 U20833 ( .A1(n17940), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n17862), 
        .B2(n17759), .ZN(n17760) );
  OAI221_X1 U20834 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17763), 
        .C1(n17762), .C2(n17761), .A(n17760), .ZN(P3_U2846) );
  OR2_X1 U20835 ( .A1(n17765), .A2(n17764), .ZN(n17788) );
  OAI21_X1 U20836 ( .B1(n20872), .B2(n17788), .A(n17774), .ZN(n17767) );
  AOI22_X1 U20837 ( .A1(n17769), .A2(n17768), .B1(n17767), .B2(n17766), .ZN(
        n17778) );
  NAND3_X1 U20838 ( .A1(n17947), .A2(n17771), .A3(n17770), .ZN(n17772) );
  OAI211_X1 U20839 ( .C1(n17935), .C2(n17774), .A(n17773), .B(n17772), .ZN(
        n17775) );
  AOI21_X1 U20840 ( .B1(n17862), .B2(n17776), .A(n17775), .ZN(n17777) );
  OAI21_X1 U20841 ( .B1(n17778), .B2(n17951), .A(n17777), .ZN(P3_U2847) );
  INV_X1 U20842 ( .A(n17779), .ZN(n17933) );
  OAI22_X1 U20843 ( .A1(n9629), .A2(n17781), .B1(n17780), .B2(n17919), .ZN(
        n17782) );
  AOI211_X1 U20844 ( .C1(n17783), .C2(n17933), .A(n20872), .B(n17782), .ZN(
        n17785) );
  OR3_X1 U20845 ( .A1(n18595), .A2(n17784), .A3(n17821), .ZN(n17811) );
  NAND2_X1 U20846 ( .A1(n18417), .A2(n17811), .ZN(n17803) );
  NAND3_X1 U20847 ( .A1(n17824), .A2(n17785), .A3(n17803), .ZN(n17786) );
  AOI22_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17896), .B1(
        n17934), .B2(n17786), .ZN(n17787) );
  AOI21_X1 U20849 ( .B1(n20872), .B2(n17788), .A(n17787), .ZN(n17793) );
  OAI22_X1 U20850 ( .A1(n17791), .A2(n17790), .B1(n17807), .B2(n17789), .ZN(
        n17792) );
  AOI211_X1 U20851 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n17940), .A(n17793), 
        .B(n17792), .ZN(n17794) );
  OAI21_X1 U20852 ( .B1(n17930), .B2(n17795), .A(n17794), .ZN(P3_U2848) );
  INV_X1 U20853 ( .A(n17834), .ZN(n17848) );
  NOR2_X1 U20854 ( .A1(n17798), .A2(n17848), .ZN(n17797) );
  AOI22_X1 U20855 ( .A1(n17877), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n17797), 
        .B2(n17796), .ZN(n17806) );
  INV_X1 U20856 ( .A(n17828), .ZN(n17836) );
  AOI22_X1 U20857 ( .A1(n17819), .A2(n17799), .B1(n17798), .B2(n17836), .ZN(
        n17800) );
  OAI211_X1 U20858 ( .C1(n17802), .C2(n17801), .A(n17824), .B(n17800), .ZN(
        n17810) );
  OAI211_X1 U20859 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17828), .A(
        n17934), .B(n17803), .ZN(n17804) );
  OAI211_X1 U20860 ( .C1(n17810), .C2(n17804), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17950), .ZN(n17805) );
  OAI211_X1 U20861 ( .C1(n17808), .C2(n17807), .A(n17806), .B(n17805), .ZN(
        P3_U2849) );
  AOI211_X1 U20862 ( .C1(n17811), .C2(n18417), .A(n17810), .B(n17809), .ZN(
        n17816) );
  AOI22_X1 U20863 ( .A1(n17829), .A2(n17834), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17934), .ZN(n17815) );
  AOI22_X1 U20864 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17896), .B1(
        n17862), .B2(n17812), .ZN(n17814) );
  OAI211_X1 U20865 ( .C1(n17816), .C2(n17815), .A(n17814), .B(n17813), .ZN(
        P3_U2850) );
  AOI22_X1 U20866 ( .A1(n17940), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17862), 
        .B2(n17817), .ZN(n17832) );
  AOI22_X1 U20867 ( .A1(n18399), .A2(n17820), .B1(n17819), .B2(n17818), .ZN(
        n17823) );
  OAI21_X1 U20868 ( .B1(n18595), .B2(n17821), .A(n18417), .ZN(n17822) );
  NAND4_X1 U20869 ( .A1(n17824), .A2(n17934), .A3(n17823), .A4(n17822), .ZN(
        n17843) );
  AOI21_X1 U20870 ( .B1(n18417), .B2(n17847), .A(n17843), .ZN(n17825) );
  OAI21_X1 U20871 ( .B1(n17827), .B2(n17826), .A(n17825), .ZN(n17837) );
  OAI22_X1 U20872 ( .A1(n18427), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n17829), .B2(n17828), .ZN(n17830) );
  OAI211_X1 U20873 ( .C1(n17837), .C2(n17830), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17950), .ZN(n17831) );
  OAI211_X1 U20874 ( .C1(n17833), .C2(n17848), .A(n17832), .B(n17831), .ZN(
        P3_U2851) );
  NAND2_X1 U20875 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17834), .ZN(
        n17842) );
  OAI221_X1 U20876 ( .B1(n17837), .B2(n17847), .C1(n17837), .C2(n17836), .A(
        n17835), .ZN(n17840) );
  AOI22_X1 U20877 ( .A1(n17877), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17862), 
        .B2(n17838), .ZN(n17839) );
  OAI221_X1 U20878 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17842), 
        .C1(n17841), .C2(n17840), .A(n17839), .ZN(P3_U2852) );
  NAND2_X1 U20879 ( .A1(n17950), .A2(n17843), .ZN(n17846) );
  AOI22_X1 U20880 ( .A1(n17940), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n17862), 
        .B2(n17844), .ZN(n17845) );
  OAI221_X1 U20881 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17848), .C1(
        n17847), .C2(n17846), .A(n17845), .ZN(P3_U2853) );
  INV_X1 U20882 ( .A(n17849), .ZN(n17852) );
  AOI21_X1 U20883 ( .B1(n17852), .B2(n17893), .A(n17919), .ZN(n17854) );
  AOI21_X1 U20884 ( .B1(n17852), .B2(n17851), .A(n17850), .ZN(n17853) );
  NOR4_X1 U20885 ( .A1(n17854), .A2(n17920), .A3(n17853), .A4(n17951), .ZN(
        n17878) );
  NAND2_X1 U20886 ( .A1(n17855), .A2(n17857), .ZN(n17868) );
  AOI21_X1 U20887 ( .B1(n17878), .B2(n17868), .A(n17940), .ZN(n17871) );
  NOR3_X1 U20888 ( .A1(n17856), .A2(n17951), .A3(n17905), .ZN(n17899) );
  NAND3_X1 U20889 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n17899), .ZN(n17879) );
  NOR2_X1 U20890 ( .A1(n17857), .A2(n17879), .ZN(n17860) );
  NOR2_X1 U20891 ( .A1(n17950), .A2(n18505), .ZN(n17858) );
  AOI221_X1 U20892 ( .B1(n17871), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(
        n17860), .C2(n17859), .A(n17858), .ZN(n17866) );
  AOI22_X1 U20893 ( .A1(n17864), .A2(n17863), .B1(n17862), .B2(n17861), .ZN(
        n17865) );
  OAI211_X1 U20894 ( .C1(n17930), .C2(n17867), .A(n17866), .B(n17865), .ZN(
        P3_U2854) );
  NOR2_X1 U20895 ( .A1(n17950), .A2(n18502), .ZN(n17870) );
  INV_X1 U20896 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17880) );
  NOR3_X1 U20897 ( .A1(n17880), .A2(n17868), .A3(n17879), .ZN(n17869) );
  AOI211_X1 U20898 ( .C1(n17871), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17870), .B(n17869), .ZN(n17875) );
  AOI22_X1 U20899 ( .A1(n17947), .A2(n17873), .B1(n17949), .B2(n17872), .ZN(
        n17874) );
  NAND2_X1 U20900 ( .A1(n17875), .A2(n17874), .ZN(P3_U2855) );
  AOI22_X1 U20901 ( .A1(n17877), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17949), 
        .B2(n17876), .ZN(n17883) );
  NOR2_X1 U20902 ( .A1(n17940), .A2(n17878), .ZN(n17888) );
  INV_X1 U20903 ( .A(n17879), .ZN(n17881) );
  AOI22_X1 U20904 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17888), .B1(
        n17881), .B2(n17880), .ZN(n17882) );
  OAI211_X1 U20905 ( .C1(n17930), .C2(n17884), .A(n17883), .B(n17882), .ZN(
        P3_U2856) );
  INV_X1 U20906 ( .A(n17885), .ZN(n17886) );
  AOI21_X1 U20907 ( .B1(n17887), .B2(n17949), .A(n17886), .ZN(n17890) );
  OAI221_X1 U20908 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17899), .C1(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n17888), .ZN(n17889) );
  OAI211_X1 U20909 ( .C1(n17930), .C2(n17891), .A(n17890), .B(n17889), .ZN(
        P3_U2857) );
  AOI22_X1 U20910 ( .A1(n17940), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n17949), 
        .B2(n17892), .ZN(n17902) );
  NOR2_X1 U20911 ( .A1(n17919), .A2(n17893), .ZN(n17927) );
  AOI211_X1 U20912 ( .C1(n17922), .C2(n17894), .A(n17927), .B(n17920), .ZN(
        n17895) );
  AOI21_X1 U20913 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17895), .A(
        n17951), .ZN(n17909) );
  NOR2_X1 U20914 ( .A1(n17896), .A2(n17909), .ZN(n17906) );
  AOI21_X1 U20915 ( .B1(n17897), .B2(n17935), .A(n17906), .ZN(n17900) );
  INV_X1 U20916 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17898) );
  AOI22_X1 U20917 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17900), .B1(
        n17899), .B2(n17898), .ZN(n17901) );
  OAI211_X1 U20918 ( .C1(n17930), .C2(n17903), .A(n17902), .B(n17901), .ZN(
        P3_U2858) );
  INV_X1 U20919 ( .A(n17949), .ZN(n17943) );
  OAI22_X1 U20920 ( .A1(n17906), .A2(n17905), .B1(n17930), .B2(n17904), .ZN(
        n17907) );
  AOI21_X1 U20921 ( .B1(n17909), .B2(n17908), .A(n17907), .ZN(n17911) );
  OAI211_X1 U20922 ( .C1(n17912), .C2(n17943), .A(n17911), .B(n17910), .ZN(
        P3_U2859) );
  NOR2_X1 U20923 ( .A1(n17913), .A2(n17935), .ZN(n17914) );
  AOI211_X1 U20924 ( .C1(n17949), .C2(n17916), .A(n17915), .B(n17914), .ZN(
        n17929) );
  INV_X1 U20925 ( .A(n17917), .ZN(n17918) );
  NOR2_X1 U20926 ( .A1(n18576), .A2(n17918), .ZN(n17925) );
  NOR3_X1 U20927 ( .A1(n17919), .A2(n18595), .A3(n18576), .ZN(n17921) );
  AOI211_X1 U20928 ( .C1(n17922), .C2(n18576), .A(n17921), .B(n17920), .ZN(
        n17923) );
  INV_X1 U20929 ( .A(n17923), .ZN(n17924) );
  MUX2_X1 U20930 ( .A(n17925), .B(n17924), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n17926) );
  OAI21_X1 U20931 ( .B1(n17927), .B2(n17926), .A(n17934), .ZN(n17928) );
  OAI211_X1 U20932 ( .C1(n17931), .C2(n17930), .A(n17929), .B(n17928), .ZN(
        P3_U2860) );
  INV_X1 U20933 ( .A(n17932), .ZN(n17944) );
  NAND3_X1 U20934 ( .A1(n17934), .A2(n18595), .A3(n17933), .ZN(n17954) );
  AOI21_X1 U20935 ( .B1(n17935), .B2(n17954), .A(n18576), .ZN(n17938) );
  AOI211_X1 U20936 ( .C1(n9629), .C2(n18595), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n17936), .ZN(n17937) );
  AOI211_X1 U20937 ( .C1(n17947), .C2(n17939), .A(n17938), .B(n17937), .ZN(
        n17942) );
  NAND2_X1 U20938 ( .A1(n17940), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n17941) );
  OAI211_X1 U20939 ( .C1(n17944), .C2(n17943), .A(n17942), .B(n17941), .ZN(
        P3_U2861) );
  INV_X1 U20940 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18606) );
  NOR2_X1 U20941 ( .A1(n17950), .A2(n18606), .ZN(n17945) );
  AOI221_X1 U20942 ( .B1(n17949), .B2(n17948), .C1(n17947), .C2(n17946), .A(
        n17945), .ZN(n17955) );
  OAI211_X1 U20943 ( .C1(n17952), .C2(n17951), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n17950), .ZN(n17953) );
  NAND3_X1 U20944 ( .A1(n17955), .A2(n17954), .A3(n17953), .ZN(P3_U2862) );
  OAI211_X1 U20945 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n17956), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18455)
         );
  OAI21_X1 U20946 ( .B1(n17959), .B2(n17957), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17958) );
  OAI221_X1 U20947 ( .B1(n17959), .B2(n18455), .C1(n17959), .C2(n18003), .A(
        n17958), .ZN(P3_U2863) );
  INV_X1 U20948 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18445) );
  NOR2_X1 U20949 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18442), .ZN(
        n18134) );
  INV_X1 U20950 ( .A(n18134), .ZN(n18108) );
  NOR2_X1 U20951 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18445), .ZN(
        n18228) );
  NAND2_X1 U20952 ( .A1(n18303), .A2(n18228), .ZN(n18251) );
  AND2_X1 U20953 ( .A1(n18108), .A2(n18251), .ZN(n17961) );
  OAI22_X1 U20954 ( .A1(n17962), .A2(n18445), .B1(n17961), .B2(n17960), .ZN(
        P3_U2866) );
  NOR2_X1 U20955 ( .A1(n20778), .A2(n17963), .ZN(P3_U2867) );
  NAND2_X1 U20956 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17965) );
  NOR2_X1 U20957 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17965), .ZN(
        n18343) );
  NAND2_X1 U20958 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18343), .ZN(
        n18398) );
  NAND2_X1 U20959 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18344), .ZN(n18281) );
  AND2_X1 U20960 ( .A1(n18344), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18345) );
  NAND2_X1 U20961 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18249), .ZN(
        n18109) );
  NOR2_X2 U20962 ( .A1(n17965), .A2(n18109), .ZN(n18333) );
  NOR2_X2 U20963 ( .A1(n18043), .A2(n17964), .ZN(n18339) );
  NOR2_X1 U20964 ( .A1(n18445), .A2(n18133), .ZN(n18342) );
  NAND2_X1 U20965 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18342), .ZN(
        n18349) );
  NAND2_X1 U20966 ( .A1(n18423), .A2(n18249), .ZN(n18425) );
  NAND2_X1 U20967 ( .A1(n18442), .A2(n18445), .ZN(n18042) );
  NOR2_X2 U20968 ( .A1(n18425), .A2(n18042), .ZN(n18049) );
  INV_X1 U20969 ( .A(n18049), .ZN(n18064) );
  NAND2_X1 U20970 ( .A1(n18349), .A2(n18064), .ZN(n18022) );
  AND2_X1 U20971 ( .A1(n18462), .A2(n18022), .ZN(n17997) );
  AOI22_X1 U20972 ( .A1(n18345), .A2(n18333), .B1(n18339), .B2(n17997), .ZN(
        n17970) );
  INV_X1 U20973 ( .A(n18109), .ZN(n18203) );
  NOR2_X1 U20974 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18249), .ZN(
        n18179) );
  NOR2_X1 U20975 ( .A1(n18203), .A2(n18179), .ZN(n18252) );
  NOR2_X1 U20976 ( .A1(n18252), .A2(n17965), .ZN(n18304) );
  AOI21_X1 U20977 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18043), .ZN(n18301) );
  AOI22_X1 U20978 ( .A1(n18344), .A2(n18304), .B1(n18301), .B2(n18022), .ZN(
        n18000) );
  NAND2_X1 U20979 ( .A1(n17967), .A2(n17966), .ZN(n17998) );
  NOR2_X1 U20980 ( .A1(n17968), .A2(n17998), .ZN(n18278) );
  AOI22_X1 U20981 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18000), .B1(
        n18049), .B2(n18278), .ZN(n17969) );
  OAI211_X1 U20982 ( .C1(n18398), .C2(n18281), .A(n17970), .B(n17969), .ZN(
        P3_U2868) );
  INV_X1 U20983 ( .A(n18333), .ZN(n18307) );
  NAND2_X1 U20984 ( .A1(n18344), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18260) );
  INV_X1 U20985 ( .A(n18398), .ZN(n18376) );
  NAND2_X1 U20986 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18344), .ZN(n18355) );
  INV_X1 U20987 ( .A(n18355), .ZN(n18257) );
  AND2_X1 U20988 ( .A1(n18254), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U20989 ( .A1(n18376), .A2(n18257), .B1(n17997), .B2(n18350), .ZN(
        n17973) );
  NOR2_X2 U20990 ( .A1(n17971), .A2(n17998), .ZN(n18352) );
  AOI22_X1 U20991 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18000), .B1(
        n18049), .B2(n18352), .ZN(n17972) );
  OAI211_X1 U20992 ( .C1(n18307), .C2(n18260), .A(n17973), .B(n17972), .ZN(
        P3_U2869) );
  NAND2_X1 U20993 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18344), .ZN(n18313) );
  NAND2_X1 U20994 ( .A1(n18344), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18361) );
  INV_X1 U20995 ( .A(n18361), .ZN(n18310) );
  NOR2_X2 U20996 ( .A1(n18043), .A2(n17974), .ZN(n18356) );
  AOI22_X1 U20997 ( .A1(n18333), .A2(n18310), .B1(n17997), .B2(n18356), .ZN(
        n17977) );
  NOR2_X2 U20998 ( .A1(n17975), .A2(n17998), .ZN(n18358) );
  AOI22_X1 U20999 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18000), .B1(
        n18049), .B2(n18358), .ZN(n17976) );
  OAI211_X1 U21000 ( .C1(n18398), .C2(n18313), .A(n17977), .B(n17976), .ZN(
        P3_U2870) );
  NAND2_X1 U21001 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18344), .ZN(n18317) );
  NAND2_X1 U21002 ( .A1(n18344), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18367) );
  NOR2_X2 U21003 ( .A1(n18043), .A2(n17978), .ZN(n18362) );
  AOI22_X1 U21004 ( .A1(n18333), .A2(n18314), .B1(n17997), .B2(n18362), .ZN(
        n17981) );
  NOR2_X2 U21005 ( .A1(n17979), .A2(n17998), .ZN(n18364) );
  AOI22_X1 U21006 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18000), .B1(
        n18049), .B2(n18364), .ZN(n17980) );
  OAI211_X1 U21007 ( .C1(n18398), .C2(n18317), .A(n17981), .B(n17980), .ZN(
        P3_U2871) );
  NAND2_X1 U21008 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18344), .ZN(n18321) );
  NAND2_X1 U21009 ( .A1(n18344), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18373) );
  INV_X1 U21010 ( .A(n18373), .ZN(n18318) );
  NOR2_X2 U21011 ( .A1(n18043), .A2(n17982), .ZN(n18368) );
  AOI22_X1 U21012 ( .A1(n18333), .A2(n18318), .B1(n17997), .B2(n18368), .ZN(
        n17985) );
  NOR2_X2 U21013 ( .A1(n17983), .A2(n17998), .ZN(n18370) );
  AOI22_X1 U21014 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18000), .B1(
        n18049), .B2(n18370), .ZN(n17984) );
  OAI211_X1 U21015 ( .C1(n18398), .C2(n18321), .A(n17985), .B(n17984), .ZN(
        P3_U2872) );
  NAND2_X1 U21016 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18344), .ZN(n18381) );
  NOR2_X1 U21017 ( .A1(n17991), .A2(n17986), .ZN(n18375) );
  NOR2_X2 U21018 ( .A1(n18043), .A2(n17987), .ZN(n18374) );
  AOI22_X1 U21019 ( .A1(n18333), .A2(n18375), .B1(n17997), .B2(n18374), .ZN(
        n17990) );
  NOR2_X2 U21020 ( .A1(n17988), .A2(n17998), .ZN(n18377) );
  AOI22_X1 U21021 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18000), .B1(
        n18049), .B2(n18377), .ZN(n17989) );
  OAI211_X1 U21022 ( .C1(n18398), .C2(n18381), .A(n17990), .B(n17989), .ZN(
        P3_U2873) );
  NAND2_X1 U21023 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18344), .ZN(n18330) );
  NOR2_X1 U21024 ( .A1(n17991), .A2(n14953), .ZN(n18327) );
  NOR2_X2 U21025 ( .A1(n18043), .A2(n17992), .ZN(n18382) );
  AOI22_X1 U21026 ( .A1(n18333), .A2(n18327), .B1(n17997), .B2(n18382), .ZN(
        n17995) );
  NOR2_X2 U21027 ( .A1(n17993), .A2(n17998), .ZN(n18384) );
  AOI22_X1 U21028 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18000), .B1(
        n18049), .B2(n18384), .ZN(n17994) );
  OAI211_X1 U21029 ( .C1(n18398), .C2(n18330), .A(n17995), .B(n17994), .ZN(
        P3_U2874) );
  NAND2_X1 U21030 ( .A1(n18344), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18338) );
  NAND2_X1 U21031 ( .A1(n18344), .A2(BUF2_REG_23__SCAN_IN), .ZN(n18397) );
  INV_X1 U21032 ( .A(n18397), .ZN(n18332) );
  NOR2_X2 U21033 ( .A1(n18043), .A2(n17996), .ZN(n18389) );
  AOI22_X1 U21034 ( .A1(n18333), .A2(n18332), .B1(n17997), .B2(n18389), .ZN(
        n18002) );
  NOR2_X2 U21035 ( .A1(n17999), .A2(n17998), .ZN(n18392) );
  AOI22_X1 U21036 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18000), .B1(
        n18049), .B2(n18392), .ZN(n18001) );
  OAI211_X1 U21037 ( .C1(n18398), .C2(n18338), .A(n18002), .B(n18001), .ZN(
        P3_U2875) );
  INV_X1 U21038 ( .A(n18349), .ZN(n18393) );
  NAND2_X1 U21039 ( .A1(n18423), .A2(n18462), .ZN(n18180) );
  NOR2_X1 U21040 ( .A1(n18042), .A2(n18180), .ZN(n18018) );
  AOI22_X1 U21041 ( .A1(n18393), .A2(n18345), .B1(n18339), .B2(n18018), .ZN(
        n18005) );
  INV_X1 U21042 ( .A(n18042), .ZN(n18044) );
  NAND2_X1 U21043 ( .A1(n18254), .A2(n18003), .ZN(n18227) );
  NOR2_X1 U21044 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18227), .ZN(
        n18181) );
  AOI22_X1 U21045 ( .A1(n18344), .A2(n18342), .B1(n18044), .B2(n18181), .ZN(
        n18019) );
  NAND2_X1 U21046 ( .A1(n18044), .A2(n18179), .ZN(n18081) );
  INV_X1 U21047 ( .A(n18081), .ZN(n18083) );
  AOI22_X1 U21048 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18019), .B1(
        n18278), .B2(n18083), .ZN(n18004) );
  OAI211_X1 U21049 ( .C1(n18281), .C2(n18307), .A(n18005), .B(n18004), .ZN(
        P3_U2876) );
  AOI22_X1 U21050 ( .A1(n18333), .A2(n18257), .B1(n18350), .B2(n18018), .ZN(
        n18007) );
  AOI22_X1 U21051 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18019), .B1(
        n18352), .B2(n18083), .ZN(n18006) );
  OAI211_X1 U21052 ( .C1(n18349), .C2(n18260), .A(n18007), .B(n18006), .ZN(
        P3_U2877) );
  INV_X1 U21053 ( .A(n18313), .ZN(n18357) );
  AOI22_X1 U21054 ( .A1(n18333), .A2(n18357), .B1(n18356), .B2(n18018), .ZN(
        n18009) );
  AOI22_X1 U21055 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18019), .B1(
        n18358), .B2(n18083), .ZN(n18008) );
  OAI211_X1 U21056 ( .C1(n18349), .C2(n18361), .A(n18009), .B(n18008), .ZN(
        P3_U2878) );
  AOI22_X1 U21057 ( .A1(n18393), .A2(n18314), .B1(n18362), .B2(n18018), .ZN(
        n18011) );
  AOI22_X1 U21058 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18019), .B1(
        n18364), .B2(n18083), .ZN(n18010) );
  OAI211_X1 U21059 ( .C1(n18307), .C2(n18317), .A(n18011), .B(n18010), .ZN(
        P3_U2879) );
  AOI22_X1 U21060 ( .A1(n18393), .A2(n18318), .B1(n18368), .B2(n18018), .ZN(
        n18013) );
  AOI22_X1 U21061 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18019), .B1(
        n18370), .B2(n18083), .ZN(n18012) );
  OAI211_X1 U21062 ( .C1(n18307), .C2(n18321), .A(n18013), .B(n18012), .ZN(
        P3_U2880) );
  AOI22_X1 U21063 ( .A1(n18393), .A2(n18375), .B1(n18374), .B2(n18018), .ZN(
        n18015) );
  AOI22_X1 U21064 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18019), .B1(
        n18377), .B2(n18083), .ZN(n18014) );
  OAI211_X1 U21065 ( .C1(n18307), .C2(n18381), .A(n18015), .B(n18014), .ZN(
        P3_U2881) );
  INV_X1 U21066 ( .A(n18327), .ZN(n18387) );
  INV_X1 U21067 ( .A(n18330), .ZN(n18383) );
  AOI22_X1 U21068 ( .A1(n18333), .A2(n18383), .B1(n18382), .B2(n18018), .ZN(
        n18017) );
  AOI22_X1 U21069 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18019), .B1(
        n18384), .B2(n18083), .ZN(n18016) );
  OAI211_X1 U21070 ( .C1(n18349), .C2(n18387), .A(n18017), .B(n18016), .ZN(
        P3_U2882) );
  INV_X1 U21071 ( .A(n18338), .ZN(n18391) );
  AOI22_X1 U21072 ( .A1(n18333), .A2(n18391), .B1(n18389), .B2(n18018), .ZN(
        n18021) );
  AOI22_X1 U21073 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18019), .B1(
        n18392), .B2(n18083), .ZN(n18020) );
  OAI211_X1 U21074 ( .C1(n18349), .C2(n18397), .A(n18021), .B(n18020), .ZN(
        P3_U2883) );
  INV_X1 U21075 ( .A(n18278), .ZN(n18348) );
  NAND2_X1 U21076 ( .A1(n18044), .A2(n18203), .ZN(n18102) );
  INV_X1 U21077 ( .A(n18281), .ZN(n18340) );
  INV_X1 U21078 ( .A(n18462), .ZN(n18250) );
  NOR2_X1 U21079 ( .A1(n18083), .A2(n18104), .ZN(n18065) );
  NOR2_X1 U21080 ( .A1(n18250), .A2(n18065), .ZN(n18038) );
  AOI22_X1 U21081 ( .A1(n18340), .A2(n18393), .B1(n18339), .B2(n18038), .ZN(
        n18025) );
  INV_X1 U21082 ( .A(n18065), .ZN(n18023) );
  OAI221_X1 U21083 ( .B1(n18023), .B2(n18303), .C1(n18023), .C2(n18022), .A(
        n18301), .ZN(n18039) );
  AOI22_X1 U21084 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18039), .B1(
        n18049), .B2(n18345), .ZN(n18024) );
  OAI211_X1 U21085 ( .C1(n18348), .C2(n18102), .A(n18025), .B(n18024), .ZN(
        P3_U2884) );
  AOI22_X1 U21086 ( .A1(n18393), .A2(n18257), .B1(n18350), .B2(n18038), .ZN(
        n18027) );
  AOI22_X1 U21087 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18039), .B1(
        n18352), .B2(n18104), .ZN(n18026) );
  OAI211_X1 U21088 ( .C1(n18064), .C2(n18260), .A(n18027), .B(n18026), .ZN(
        P3_U2885) );
  AOI22_X1 U21089 ( .A1(n18393), .A2(n18357), .B1(n18356), .B2(n18038), .ZN(
        n18029) );
  AOI22_X1 U21090 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18039), .B1(
        n18358), .B2(n18104), .ZN(n18028) );
  OAI211_X1 U21091 ( .C1(n18064), .C2(n18361), .A(n18029), .B(n18028), .ZN(
        P3_U2886) );
  AOI22_X1 U21092 ( .A1(n18049), .A2(n18314), .B1(n18362), .B2(n18038), .ZN(
        n18031) );
  AOI22_X1 U21093 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18039), .B1(
        n18364), .B2(n18104), .ZN(n18030) );
  OAI211_X1 U21094 ( .C1(n18349), .C2(n18317), .A(n18031), .B(n18030), .ZN(
        P3_U2887) );
  AOI22_X1 U21095 ( .A1(n18049), .A2(n18318), .B1(n18368), .B2(n18038), .ZN(
        n18033) );
  AOI22_X1 U21096 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18039), .B1(
        n18370), .B2(n18104), .ZN(n18032) );
  OAI211_X1 U21097 ( .C1(n18349), .C2(n18321), .A(n18033), .B(n18032), .ZN(
        P3_U2888) );
  AOI22_X1 U21098 ( .A1(n18049), .A2(n18375), .B1(n18374), .B2(n18038), .ZN(
        n18035) );
  AOI22_X1 U21099 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18039), .B1(
        n18377), .B2(n18104), .ZN(n18034) );
  OAI211_X1 U21100 ( .C1(n18349), .C2(n18381), .A(n18035), .B(n18034), .ZN(
        P3_U2889) );
  AOI22_X1 U21101 ( .A1(n18393), .A2(n18383), .B1(n18382), .B2(n18038), .ZN(
        n18037) );
  AOI22_X1 U21102 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18039), .B1(
        n18384), .B2(n18104), .ZN(n18036) );
  OAI211_X1 U21103 ( .C1(n18064), .C2(n18387), .A(n18037), .B(n18036), .ZN(
        P3_U2890) );
  AOI22_X1 U21104 ( .A1(n18049), .A2(n18332), .B1(n18389), .B2(n18038), .ZN(
        n18041) );
  AOI22_X1 U21105 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18039), .B1(
        n18392), .B2(n18104), .ZN(n18040) );
  OAI211_X1 U21106 ( .C1(n18349), .C2(n18338), .A(n18041), .B(n18040), .ZN(
        P3_U2891) );
  NOR2_X1 U21107 ( .A1(n18423), .A2(n18042), .ZN(n18087) );
  NAND2_X1 U21108 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18087), .ZN(
        n18132) );
  INV_X1 U21109 ( .A(n18303), .ZN(n18110) );
  AOI21_X1 U21110 ( .B1(n18423), .B2(n18110), .A(n18043), .ZN(n18135) );
  OAI211_X1 U21111 ( .C1(n18125), .C2(n18566), .A(n18044), .B(n18135), .ZN(
        n18061) );
  AND2_X1 U21112 ( .A1(n18462), .A2(n18087), .ZN(n18060) );
  AOI22_X1 U21113 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18061), .B1(
        n18339), .B2(n18060), .ZN(n18046) );
  AOI22_X1 U21114 ( .A1(n18278), .A2(n18125), .B1(n18345), .B2(n18083), .ZN(
        n18045) );
  OAI211_X1 U21115 ( .C1(n18281), .C2(n18064), .A(n18046), .B(n18045), .ZN(
        P3_U2892) );
  AOI22_X1 U21116 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18061), .B1(
        n18350), .B2(n18060), .ZN(n18048) );
  AOI22_X1 U21117 ( .A1(n18049), .A2(n18257), .B1(n18352), .B2(n18125), .ZN(
        n18047) );
  OAI211_X1 U21118 ( .C1(n18260), .C2(n18081), .A(n18048), .B(n18047), .ZN(
        P3_U2893) );
  AOI22_X1 U21119 ( .A1(n18049), .A2(n18357), .B1(n18356), .B2(n18060), .ZN(
        n18051) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18061), .B1(
        n18358), .B2(n18125), .ZN(n18050) );
  OAI211_X1 U21121 ( .C1(n18361), .C2(n18081), .A(n18051), .B(n18050), .ZN(
        P3_U2894) );
  AOI22_X1 U21122 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18061), .B1(
        n18362), .B2(n18060), .ZN(n18053) );
  AOI22_X1 U21123 ( .A1(n18364), .A2(n18125), .B1(n18314), .B2(n18083), .ZN(
        n18052) );
  OAI211_X1 U21124 ( .C1(n18064), .C2(n18317), .A(n18053), .B(n18052), .ZN(
        P3_U2895) );
  AOI22_X1 U21125 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18061), .B1(
        n18368), .B2(n18060), .ZN(n18055) );
  AOI22_X1 U21126 ( .A1(n18370), .A2(n18125), .B1(n18318), .B2(n18083), .ZN(
        n18054) );
  OAI211_X1 U21127 ( .C1(n18064), .C2(n18321), .A(n18055), .B(n18054), .ZN(
        P3_U2896) );
  AOI22_X1 U21128 ( .A1(n18375), .A2(n18083), .B1(n18374), .B2(n18060), .ZN(
        n18057) );
  AOI22_X1 U21129 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18061), .B1(
        n18377), .B2(n18125), .ZN(n18056) );
  OAI211_X1 U21130 ( .C1(n18064), .C2(n18381), .A(n18057), .B(n18056), .ZN(
        P3_U2897) );
  AOI22_X1 U21131 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18061), .B1(
        n18382), .B2(n18060), .ZN(n18059) );
  AOI22_X1 U21132 ( .A1(n18384), .A2(n18125), .B1(n18327), .B2(n18083), .ZN(
        n18058) );
  OAI211_X1 U21133 ( .C1(n18064), .C2(n18330), .A(n18059), .B(n18058), .ZN(
        P3_U2898) );
  AOI22_X1 U21134 ( .A1(n18332), .A2(n18083), .B1(n18389), .B2(n18060), .ZN(
        n18063) );
  AOI22_X1 U21135 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18061), .B1(
        n18392), .B2(n18125), .ZN(n18062) );
  OAI211_X1 U21136 ( .C1(n18064), .C2(n18338), .A(n18063), .B(n18062), .ZN(
        P3_U2899) );
  INV_X1 U21137 ( .A(n18425), .ZN(n18156) );
  NAND2_X1 U21138 ( .A1(n18156), .A2(n18134), .ZN(n18150) );
  AOI21_X1 U21139 ( .B1(n18132), .B2(n18150), .A(n18250), .ZN(n18082) );
  AOI22_X1 U21140 ( .A1(n18345), .A2(n18104), .B1(n18339), .B2(n18082), .ZN(
        n18068) );
  AOI221_X1 U21141 ( .B1(n18065), .B2(n18132), .C1(n18110), .C2(n18132), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18066) );
  OAI21_X1 U21142 ( .B1(n18153), .B2(n18066), .A(n18254), .ZN(n18084) );
  AOI22_X1 U21143 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18084), .B1(
        n18278), .B2(n18153), .ZN(n18067) );
  OAI211_X1 U21144 ( .C1(n18281), .C2(n18081), .A(n18068), .B(n18067), .ZN(
        P3_U2900) );
  INV_X1 U21145 ( .A(n18260), .ZN(n18351) );
  AOI22_X1 U21146 ( .A1(n18351), .A2(n18104), .B1(n18350), .B2(n18082), .ZN(
        n18070) );
  AOI22_X1 U21147 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18084), .B1(
        n18352), .B2(n18153), .ZN(n18069) );
  OAI211_X1 U21148 ( .C1(n18355), .C2(n18081), .A(n18070), .B(n18069), .ZN(
        P3_U2901) );
  AOI22_X1 U21149 ( .A1(n18357), .A2(n18083), .B1(n18356), .B2(n18082), .ZN(
        n18072) );
  AOI22_X1 U21150 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18084), .B1(
        n18358), .B2(n18153), .ZN(n18071) );
  OAI211_X1 U21151 ( .C1(n18361), .C2(n18102), .A(n18072), .B(n18071), .ZN(
        P3_U2902) );
  AOI22_X1 U21152 ( .A1(n18314), .A2(n18104), .B1(n18362), .B2(n18082), .ZN(
        n18074) );
  AOI22_X1 U21153 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18084), .B1(
        n18364), .B2(n18153), .ZN(n18073) );
  OAI211_X1 U21154 ( .C1(n18317), .C2(n18081), .A(n18074), .B(n18073), .ZN(
        P3_U2903) );
  INV_X1 U21155 ( .A(n18321), .ZN(n18369) );
  AOI22_X1 U21156 ( .A1(n18369), .A2(n18083), .B1(n18368), .B2(n18082), .ZN(
        n18076) );
  AOI22_X1 U21157 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18084), .B1(
        n18370), .B2(n18153), .ZN(n18075) );
  OAI211_X1 U21158 ( .C1(n18373), .C2(n18102), .A(n18076), .B(n18075), .ZN(
        P3_U2904) );
  AOI22_X1 U21159 ( .A1(n18375), .A2(n18104), .B1(n18374), .B2(n18082), .ZN(
        n18078) );
  AOI22_X1 U21160 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18084), .B1(
        n18377), .B2(n18153), .ZN(n18077) );
  OAI211_X1 U21161 ( .C1(n18381), .C2(n18081), .A(n18078), .B(n18077), .ZN(
        P3_U2905) );
  AOI22_X1 U21162 ( .A1(n18327), .A2(n18104), .B1(n18382), .B2(n18082), .ZN(
        n18080) );
  AOI22_X1 U21163 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18084), .B1(
        n18384), .B2(n18153), .ZN(n18079) );
  OAI211_X1 U21164 ( .C1(n18330), .C2(n18081), .A(n18080), .B(n18079), .ZN(
        P3_U2906) );
  AOI22_X1 U21165 ( .A1(n18391), .A2(n18083), .B1(n18389), .B2(n18082), .ZN(
        n18086) );
  AOI22_X1 U21166 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18084), .B1(
        n18392), .B2(n18153), .ZN(n18085) );
  OAI211_X1 U21167 ( .C1(n18397), .C2(n18102), .A(n18086), .B(n18085), .ZN(
        P3_U2907) );
  NAND2_X1 U21168 ( .A1(n18179), .A2(n18134), .ZN(n18171) );
  NOR2_X1 U21169 ( .A1(n18180), .A2(n18108), .ZN(n18103) );
  AOI22_X1 U21170 ( .A1(n18340), .A2(n18104), .B1(n18339), .B2(n18103), .ZN(
        n18089) );
  AOI22_X1 U21171 ( .A1(n18344), .A2(n18087), .B1(n18181), .B2(n18134), .ZN(
        n18105) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18105), .B1(
        n18345), .B2(n18125), .ZN(n18088) );
  OAI211_X1 U21173 ( .C1(n18348), .C2(n18171), .A(n18089), .B(n18088), .ZN(
        P3_U2908) );
  AOI22_X1 U21174 ( .A1(n18351), .A2(n18125), .B1(n18350), .B2(n18103), .ZN(
        n18091) );
  INV_X1 U21175 ( .A(n18171), .ZN(n18176) );
  AOI22_X1 U21176 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18105), .B1(
        n18352), .B2(n18176), .ZN(n18090) );
  OAI211_X1 U21177 ( .C1(n18355), .C2(n18102), .A(n18091), .B(n18090), .ZN(
        P3_U2909) );
  AOI22_X1 U21178 ( .A1(n18310), .A2(n18125), .B1(n18356), .B2(n18103), .ZN(
        n18093) );
  AOI22_X1 U21179 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18105), .B1(
        n18358), .B2(n18176), .ZN(n18092) );
  OAI211_X1 U21180 ( .C1(n18313), .C2(n18102), .A(n18093), .B(n18092), .ZN(
        P3_U2910) );
  INV_X1 U21181 ( .A(n18317), .ZN(n18363) );
  AOI22_X1 U21182 ( .A1(n18363), .A2(n18104), .B1(n18362), .B2(n18103), .ZN(
        n18095) );
  AOI22_X1 U21183 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18105), .B1(
        n18364), .B2(n18176), .ZN(n18094) );
  OAI211_X1 U21184 ( .C1(n18367), .C2(n18132), .A(n18095), .B(n18094), .ZN(
        P3_U2911) );
  AOI22_X1 U21185 ( .A1(n18369), .A2(n18104), .B1(n18368), .B2(n18103), .ZN(
        n18097) );
  AOI22_X1 U21186 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18105), .B1(
        n18370), .B2(n18176), .ZN(n18096) );
  OAI211_X1 U21187 ( .C1(n18373), .C2(n18132), .A(n18097), .B(n18096), .ZN(
        P3_U2912) );
  AOI22_X1 U21188 ( .A1(n18375), .A2(n18125), .B1(n18374), .B2(n18103), .ZN(
        n18099) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18105), .B1(
        n18377), .B2(n18176), .ZN(n18098) );
  OAI211_X1 U21190 ( .C1(n18381), .C2(n18102), .A(n18099), .B(n18098), .ZN(
        P3_U2913) );
  AOI22_X1 U21191 ( .A1(n18327), .A2(n18125), .B1(n18382), .B2(n18103), .ZN(
        n18101) );
  AOI22_X1 U21192 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18105), .B1(
        n18384), .B2(n18176), .ZN(n18100) );
  OAI211_X1 U21193 ( .C1(n18330), .C2(n18102), .A(n18101), .B(n18100), .ZN(
        P3_U2914) );
  AOI22_X1 U21194 ( .A1(n18391), .A2(n18104), .B1(n18389), .B2(n18103), .ZN(
        n18107) );
  AOI22_X1 U21195 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18105), .B1(
        n18392), .B2(n18176), .ZN(n18106) );
  OAI211_X1 U21196 ( .C1(n18397), .C2(n18132), .A(n18107), .B(n18106), .ZN(
        P3_U2915) );
  NOR2_X1 U21197 ( .A1(n18176), .A2(n9592), .ZN(n18157) );
  NOR2_X1 U21198 ( .A1(n18250), .A2(n18157), .ZN(n18128) );
  AOI22_X1 U21199 ( .A1(n18345), .A2(n18153), .B1(n18339), .B2(n18128), .ZN(
        n18114) );
  NOR2_X1 U21200 ( .A1(n18125), .A2(n18153), .ZN(n18111) );
  OAI21_X1 U21201 ( .B1(n18111), .B2(n18110), .A(n18157), .ZN(n18112) );
  OAI211_X1 U21202 ( .C1(n9592), .C2(n18566), .A(n18254), .B(n18112), .ZN(
        n18129) );
  AOI22_X1 U21203 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18129), .B1(
        n18278), .B2(n9592), .ZN(n18113) );
  OAI211_X1 U21204 ( .C1(n18281), .C2(n18132), .A(n18114), .B(n18113), .ZN(
        P3_U2916) );
  AOI22_X1 U21205 ( .A1(n18351), .A2(n18153), .B1(n18350), .B2(n18128), .ZN(
        n18116) );
  AOI22_X1 U21206 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18129), .B1(
        n18352), .B2(n9592), .ZN(n18115) );
  OAI211_X1 U21207 ( .C1(n18355), .C2(n18132), .A(n18116), .B(n18115), .ZN(
        P3_U2917) );
  AOI22_X1 U21208 ( .A1(n18357), .A2(n18125), .B1(n18356), .B2(n18128), .ZN(
        n18118) );
  AOI22_X1 U21209 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18129), .B1(
        n18358), .B2(n9592), .ZN(n18117) );
  OAI211_X1 U21210 ( .C1(n18361), .C2(n18150), .A(n18118), .B(n18117), .ZN(
        P3_U2918) );
  AOI22_X1 U21211 ( .A1(n18363), .A2(n18125), .B1(n18362), .B2(n18128), .ZN(
        n18120) );
  AOI22_X1 U21212 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18129), .B1(
        n18364), .B2(n9592), .ZN(n18119) );
  OAI211_X1 U21213 ( .C1(n18367), .C2(n18150), .A(n18120), .B(n18119), .ZN(
        P3_U2919) );
  AOI22_X1 U21214 ( .A1(n18369), .A2(n18125), .B1(n18368), .B2(n18128), .ZN(
        n18122) );
  AOI22_X1 U21215 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18129), .B1(
        n18370), .B2(n9592), .ZN(n18121) );
  OAI211_X1 U21216 ( .C1(n18373), .C2(n18150), .A(n18122), .B(n18121), .ZN(
        P3_U2920) );
  AOI22_X1 U21217 ( .A1(n18375), .A2(n18153), .B1(n18374), .B2(n18128), .ZN(
        n18124) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18129), .B1(
        n18377), .B2(n9592), .ZN(n18123) );
  OAI211_X1 U21219 ( .C1(n18381), .C2(n18132), .A(n18124), .B(n18123), .ZN(
        P3_U2921) );
  AOI22_X1 U21220 ( .A1(n18383), .A2(n18125), .B1(n18382), .B2(n18128), .ZN(
        n18127) );
  AOI22_X1 U21221 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18129), .B1(
        n18384), .B2(n9592), .ZN(n18126) );
  OAI211_X1 U21222 ( .C1(n18387), .C2(n18150), .A(n18127), .B(n18126), .ZN(
        P3_U2922) );
  AOI22_X1 U21223 ( .A1(n18332), .A2(n18153), .B1(n18389), .B2(n18128), .ZN(
        n18131) );
  AOI22_X1 U21224 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18129), .B1(
        n18392), .B2(n9592), .ZN(n18130) );
  OAI211_X1 U21225 ( .C1(n18338), .C2(n18132), .A(n18131), .B(n18130), .ZN(
        P3_U2923) );
  INV_X1 U21226 ( .A(n18222), .ZN(n18220) );
  NOR2_X1 U21227 ( .A1(n18133), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18182) );
  AND2_X1 U21228 ( .A1(n18462), .A2(n18182), .ZN(n18151) );
  AOI22_X1 U21229 ( .A1(n18340), .A2(n18153), .B1(n18339), .B2(n18151), .ZN(
        n18137) );
  OAI211_X1 U21230 ( .C1(n18222), .C2(n18566), .A(n18135), .B(n18134), .ZN(
        n18152) );
  AOI22_X1 U21231 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18152), .B1(
        n18345), .B2(n18176), .ZN(n18136) );
  OAI211_X1 U21232 ( .C1(n18348), .C2(n18220), .A(n18137), .B(n18136), .ZN(
        P3_U2924) );
  AOI22_X1 U21233 ( .A1(n18257), .A2(n18153), .B1(n18350), .B2(n18151), .ZN(
        n18139) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18152), .B1(
        n18352), .B2(n18222), .ZN(n18138) );
  OAI211_X1 U21235 ( .C1(n18260), .C2(n18171), .A(n18139), .B(n18138), .ZN(
        P3_U2925) );
  AOI22_X1 U21236 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18152), .B1(
        n18356), .B2(n18151), .ZN(n18141) );
  AOI22_X1 U21237 ( .A1(n18358), .A2(n18222), .B1(n18310), .B2(n18176), .ZN(
        n18140) );
  OAI211_X1 U21238 ( .C1(n18313), .C2(n18150), .A(n18141), .B(n18140), .ZN(
        P3_U2926) );
  AOI22_X1 U21239 ( .A1(n18314), .A2(n18176), .B1(n18362), .B2(n18151), .ZN(
        n18143) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18152), .B1(
        n18364), .B2(n18222), .ZN(n18142) );
  OAI211_X1 U21241 ( .C1(n18317), .C2(n18150), .A(n18143), .B(n18142), .ZN(
        P3_U2927) );
  AOI22_X1 U21242 ( .A1(n18368), .A2(n18151), .B1(n18318), .B2(n18176), .ZN(
        n18145) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18152), .B1(
        n18370), .B2(n18222), .ZN(n18144) );
  OAI211_X1 U21244 ( .C1(n18321), .C2(n18150), .A(n18145), .B(n18144), .ZN(
        P3_U2928) );
  AOI22_X1 U21245 ( .A1(n18375), .A2(n18176), .B1(n18374), .B2(n18151), .ZN(
        n18147) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18152), .B1(
        n18377), .B2(n18222), .ZN(n18146) );
  OAI211_X1 U21247 ( .C1(n18381), .C2(n18150), .A(n18147), .B(n18146), .ZN(
        P3_U2929) );
  AOI22_X1 U21248 ( .A1(n18327), .A2(n18176), .B1(n18382), .B2(n18151), .ZN(
        n18149) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18152), .B1(
        n18384), .B2(n18222), .ZN(n18148) );
  OAI211_X1 U21250 ( .C1(n18330), .C2(n18150), .A(n18149), .B(n18148), .ZN(
        P3_U2930) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18152), .B1(
        n18389), .B2(n18151), .ZN(n18155) );
  AOI22_X1 U21252 ( .A1(n18391), .A2(n18153), .B1(n18392), .B2(n18222), .ZN(
        n18154) );
  OAI211_X1 U21253 ( .C1(n18397), .C2(n18171), .A(n18155), .B(n18154), .ZN(
        P3_U2931) );
  NAND2_X1 U21254 ( .A1(n18156), .A2(n18228), .ZN(n18248) );
  NAND2_X1 U21255 ( .A1(n18220), .A2(n18248), .ZN(n18204) );
  INV_X1 U21256 ( .A(n18157), .ZN(n18158) );
  OAI221_X1 U21257 ( .B1(n18204), .B2(n18303), .C1(n18204), .C2(n18158), .A(
        n18301), .ZN(n18175) );
  AND2_X1 U21258 ( .A1(n18462), .A2(n18204), .ZN(n18174) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18175), .B1(
        n18339), .B2(n18174), .ZN(n18160) );
  INV_X1 U21260 ( .A(n18248), .ZN(n18241) );
  AOI22_X1 U21261 ( .A1(n18278), .A2(n18241), .B1(n18345), .B2(n9592), .ZN(
        n18159) );
  OAI211_X1 U21262 ( .C1(n18281), .C2(n18171), .A(n18160), .B(n18159), .ZN(
        P3_U2932) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18175), .B1(
        n18350), .B2(n18174), .ZN(n18162) );
  AOI22_X1 U21264 ( .A1(n18351), .A2(n9592), .B1(n18352), .B2(n18241), .ZN(
        n18161) );
  OAI211_X1 U21265 ( .C1(n18355), .C2(n18171), .A(n18162), .B(n18161), .ZN(
        P3_U2933) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18175), .B1(
        n18356), .B2(n18174), .ZN(n18164) );
  AOI22_X1 U21267 ( .A1(n18358), .A2(n18241), .B1(n18310), .B2(n9592), .ZN(
        n18163) );
  OAI211_X1 U21268 ( .C1(n18313), .C2(n18171), .A(n18164), .B(n18163), .ZN(
        P3_U2934) );
  AOI22_X1 U21269 ( .A1(n18314), .A2(n9592), .B1(n18362), .B2(n18174), .ZN(
        n18166) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18175), .B1(
        n18364), .B2(n18241), .ZN(n18165) );
  OAI211_X1 U21271 ( .C1(n18317), .C2(n18171), .A(n18166), .B(n18165), .ZN(
        P3_U2935) );
  AOI22_X1 U21272 ( .A1(n18368), .A2(n18174), .B1(n18318), .B2(n9592), .ZN(
        n18168) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18175), .B1(
        n18370), .B2(n18241), .ZN(n18167) );
  OAI211_X1 U21274 ( .C1(n18321), .C2(n18171), .A(n18168), .B(n18167), .ZN(
        P3_U2936) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18175), .B1(
        n18374), .B2(n18174), .ZN(n18170) );
  AOI22_X1 U21276 ( .A1(n18377), .A2(n18241), .B1(n18375), .B2(n9592), .ZN(
        n18169) );
  OAI211_X1 U21277 ( .C1(n18381), .C2(n18171), .A(n18170), .B(n18169), .ZN(
        P3_U2937) );
  INV_X1 U21278 ( .A(n9592), .ZN(n18194) );
  AOI22_X1 U21279 ( .A1(n18383), .A2(n18176), .B1(n18382), .B2(n18174), .ZN(
        n18173) );
  AOI22_X1 U21280 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18175), .B1(
        n18384), .B2(n18241), .ZN(n18172) );
  OAI211_X1 U21281 ( .C1(n18387), .C2(n18194), .A(n18173), .B(n18172), .ZN(
        P3_U2938) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18175), .B1(
        n18389), .B2(n18174), .ZN(n18178) );
  AOI22_X1 U21283 ( .A1(n18391), .A2(n18176), .B1(n18392), .B2(n18241), .ZN(
        n18177) );
  OAI211_X1 U21284 ( .C1(n18397), .C2(n18194), .A(n18178), .B(n18177), .ZN(
        P3_U2939) );
  NAND2_X1 U21285 ( .A1(n18179), .A2(n18228), .ZN(n18276) );
  INV_X1 U21286 ( .A(n18228), .ZN(n18226) );
  NOR2_X1 U21287 ( .A1(n18180), .A2(n18226), .ZN(n18199) );
  AOI22_X1 U21288 ( .A1(n18345), .A2(n18222), .B1(n18339), .B2(n18199), .ZN(
        n18184) );
  AOI22_X1 U21289 ( .A1(n18344), .A2(n18182), .B1(n18181), .B2(n18228), .ZN(
        n18200) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18200), .B1(
        n18340), .B2(n9592), .ZN(n18183) );
  OAI211_X1 U21291 ( .C1(n18348), .C2(n18276), .A(n18184), .B(n18183), .ZN(
        P3_U2940) );
  AOI22_X1 U21292 ( .A1(n18351), .A2(n18222), .B1(n18350), .B2(n18199), .ZN(
        n18186) );
  INV_X1 U21293 ( .A(n18276), .ZN(n18267) );
  AOI22_X1 U21294 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18200), .B1(
        n18352), .B2(n18267), .ZN(n18185) );
  OAI211_X1 U21295 ( .C1(n18355), .C2(n18194), .A(n18186), .B(n18185), .ZN(
        P3_U2941) );
  AOI22_X1 U21296 ( .A1(n18357), .A2(n9592), .B1(n18356), .B2(n18199), .ZN(
        n18189) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18200), .B1(
        n18358), .B2(n18267), .ZN(n18188) );
  OAI211_X1 U21298 ( .C1(n18361), .C2(n18220), .A(n18189), .B(n18188), .ZN(
        P3_U2942) );
  AOI22_X1 U21299 ( .A1(n18314), .A2(n18222), .B1(n18362), .B2(n18199), .ZN(
        n18191) );
  AOI22_X1 U21300 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18200), .B1(
        n18364), .B2(n18267), .ZN(n18190) );
  OAI211_X1 U21301 ( .C1(n18317), .C2(n18194), .A(n18191), .B(n18190), .ZN(
        P3_U2943) );
  AOI22_X1 U21302 ( .A1(n18368), .A2(n18199), .B1(n18318), .B2(n18222), .ZN(
        n18193) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18200), .B1(
        n18370), .B2(n18267), .ZN(n18192) );
  OAI211_X1 U21304 ( .C1(n18321), .C2(n18194), .A(n18193), .B(n18192), .ZN(
        P3_U2944) );
  INV_X1 U21305 ( .A(n18375), .ZN(n18326) );
  INV_X1 U21306 ( .A(n18381), .ZN(n18323) );
  AOI22_X1 U21307 ( .A1(n18323), .A2(n9592), .B1(n18374), .B2(n18199), .ZN(
        n18196) );
  AOI22_X1 U21308 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18200), .B1(
        n18377), .B2(n18267), .ZN(n18195) );
  OAI211_X1 U21309 ( .C1(n18326), .C2(n18220), .A(n18196), .B(n18195), .ZN(
        P3_U2945) );
  AOI22_X1 U21310 ( .A1(n18383), .A2(n9592), .B1(n18382), .B2(n18199), .ZN(
        n18198) );
  AOI22_X1 U21311 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18200), .B1(
        n18384), .B2(n18267), .ZN(n18197) );
  OAI211_X1 U21312 ( .C1(n18387), .C2(n18220), .A(n18198), .B(n18197), .ZN(
        P3_U2946) );
  AOI22_X1 U21313 ( .A1(n18391), .A2(n9592), .B1(n18389), .B2(n18199), .ZN(
        n18202) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18200), .B1(
        n18392), .B2(n18267), .ZN(n18201) );
  OAI211_X1 U21315 ( .C1(n18397), .C2(n18220), .A(n18202), .B(n18201), .ZN(
        P3_U2947) );
  NAND2_X1 U21316 ( .A1(n18203), .A2(n18228), .ZN(n18288) );
  AOI21_X1 U21317 ( .B1(n18276), .B2(n18288), .A(n18250), .ZN(n18221) );
  AOI22_X1 U21318 ( .A1(n18340), .A2(n18222), .B1(n18339), .B2(n18221), .ZN(
        n18207) );
  NAND2_X1 U21319 ( .A1(n18276), .A2(n18288), .ZN(n18205) );
  OAI221_X1 U21320 ( .B1(n18205), .B2(n18303), .C1(n18205), .C2(n18204), .A(
        n18301), .ZN(n18223) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18223), .B1(
        n18345), .B2(n18241), .ZN(n18206) );
  OAI211_X1 U21322 ( .C1(n18348), .C2(n18288), .A(n18207), .B(n18206), .ZN(
        P3_U2948) );
  AOI22_X1 U21323 ( .A1(n18257), .A2(n18222), .B1(n18350), .B2(n18221), .ZN(
        n18209) );
  INV_X1 U21324 ( .A(n18288), .ZN(n18296) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18223), .B1(
        n18352), .B2(n18296), .ZN(n18208) );
  OAI211_X1 U21326 ( .C1(n18260), .C2(n18248), .A(n18209), .B(n18208), .ZN(
        P3_U2949) );
  AOI22_X1 U21327 ( .A1(n18310), .A2(n18241), .B1(n18356), .B2(n18221), .ZN(
        n18211) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18223), .B1(
        n18358), .B2(n18296), .ZN(n18210) );
  OAI211_X1 U21329 ( .C1(n18313), .C2(n18220), .A(n18211), .B(n18210), .ZN(
        P3_U2950) );
  AOI22_X1 U21330 ( .A1(n18314), .A2(n18241), .B1(n18362), .B2(n18221), .ZN(
        n18213) );
  AOI22_X1 U21331 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18223), .B1(
        n18364), .B2(n18296), .ZN(n18212) );
  OAI211_X1 U21332 ( .C1(n18317), .C2(n18220), .A(n18213), .B(n18212), .ZN(
        P3_U2951) );
  AOI22_X1 U21333 ( .A1(n18369), .A2(n18222), .B1(n18368), .B2(n18221), .ZN(
        n18215) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18223), .B1(
        n18370), .B2(n18296), .ZN(n18214) );
  OAI211_X1 U21335 ( .C1(n18373), .C2(n18248), .A(n18215), .B(n18214), .ZN(
        P3_U2952) );
  AOI22_X1 U21336 ( .A1(n18375), .A2(n18241), .B1(n18374), .B2(n18221), .ZN(
        n18217) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18223), .B1(
        n18377), .B2(n18296), .ZN(n18216) );
  OAI211_X1 U21338 ( .C1(n18381), .C2(n18220), .A(n18217), .B(n18216), .ZN(
        P3_U2953) );
  AOI22_X1 U21339 ( .A1(n18327), .A2(n18241), .B1(n18382), .B2(n18221), .ZN(
        n18219) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18223), .B1(
        n18384), .B2(n18296), .ZN(n18218) );
  OAI211_X1 U21341 ( .C1(n18330), .C2(n18220), .A(n18219), .B(n18218), .ZN(
        P3_U2954) );
  AOI22_X1 U21342 ( .A1(n18391), .A2(n18222), .B1(n18389), .B2(n18221), .ZN(
        n18225) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18223), .B1(
        n18392), .B2(n18296), .ZN(n18224) );
  OAI211_X1 U21344 ( .C1(n18397), .C2(n18248), .A(n18225), .B(n18224), .ZN(
        P3_U2955) );
  NOR2_X1 U21345 ( .A1(n18423), .A2(n18226), .ZN(n18277) );
  AND2_X1 U21346 ( .A1(n18462), .A2(n18277), .ZN(n18244) );
  AOI22_X1 U21347 ( .A1(n18345), .A2(n18267), .B1(n18339), .B2(n18244), .ZN(
        n18230) );
  INV_X1 U21348 ( .A(n18227), .ZN(n18341) );
  AOI22_X1 U21349 ( .A1(n18344), .A2(n18228), .B1(n18341), .B2(n18277), .ZN(
        n18245) );
  NAND2_X1 U21350 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18277), .ZN(
        n18337) );
  INV_X1 U21351 ( .A(n18337), .ZN(n18322) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18245), .B1(
        n18278), .B2(n18322), .ZN(n18229) );
  OAI211_X1 U21353 ( .C1(n18281), .C2(n18248), .A(n18230), .B(n18229), .ZN(
        P3_U2956) );
  AOI22_X1 U21354 ( .A1(n18257), .A2(n18241), .B1(n18350), .B2(n18244), .ZN(
        n18232) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18245), .B1(
        n18352), .B2(n18322), .ZN(n18231) );
  OAI211_X1 U21356 ( .C1(n18260), .C2(n18276), .A(n18232), .B(n18231), .ZN(
        P3_U2957) );
  AOI22_X1 U21357 ( .A1(n18310), .A2(n18267), .B1(n18356), .B2(n18244), .ZN(
        n18234) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18245), .B1(
        n18358), .B2(n18322), .ZN(n18233) );
  OAI211_X1 U21359 ( .C1(n18313), .C2(n18248), .A(n18234), .B(n18233), .ZN(
        P3_U2958) );
  AOI22_X1 U21360 ( .A1(n18314), .A2(n18267), .B1(n18362), .B2(n18244), .ZN(
        n18236) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18245), .B1(
        n18364), .B2(n18322), .ZN(n18235) );
  OAI211_X1 U21362 ( .C1(n18317), .C2(n18248), .A(n18236), .B(n18235), .ZN(
        P3_U2959) );
  AOI22_X1 U21363 ( .A1(n18368), .A2(n18244), .B1(n18318), .B2(n18267), .ZN(
        n18238) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18245), .B1(
        n18370), .B2(n18322), .ZN(n18237) );
  OAI211_X1 U21365 ( .C1(n18321), .C2(n18248), .A(n18238), .B(n18237), .ZN(
        P3_U2960) );
  AOI22_X1 U21366 ( .A1(n18323), .A2(n18241), .B1(n18374), .B2(n18244), .ZN(
        n18240) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18245), .B1(
        n18377), .B2(n18322), .ZN(n18239) );
  OAI211_X1 U21368 ( .C1(n18326), .C2(n18276), .A(n18240), .B(n18239), .ZN(
        P3_U2961) );
  AOI22_X1 U21369 ( .A1(n18383), .A2(n18241), .B1(n18382), .B2(n18244), .ZN(
        n18243) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18245), .B1(
        n18384), .B2(n18322), .ZN(n18242) );
  OAI211_X1 U21371 ( .C1(n18387), .C2(n18276), .A(n18243), .B(n18242), .ZN(
        P3_U2962) );
  AOI22_X1 U21372 ( .A1(n18332), .A2(n18267), .B1(n18389), .B2(n18244), .ZN(
        n18247) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18245), .B1(
        n18392), .B2(n18322), .ZN(n18246) );
  OAI211_X1 U21374 ( .C1(n18338), .C2(n18248), .A(n18247), .B(n18246), .ZN(
        P3_U2963) );
  NAND2_X1 U21375 ( .A1(n18343), .A2(n18249), .ZN(n18380) );
  NOR2_X1 U21376 ( .A1(n18322), .A2(n18390), .ZN(n18300) );
  NOR2_X1 U21377 ( .A1(n18250), .A2(n18300), .ZN(n18272) );
  AOI22_X1 U21378 ( .A1(n18345), .A2(n18296), .B1(n18339), .B2(n18272), .ZN(
        n18256) );
  OAI21_X1 U21379 ( .B1(n18252), .B2(n18251), .A(n18300), .ZN(n18253) );
  OAI211_X1 U21380 ( .C1(n18390), .C2(n18566), .A(n18254), .B(n18253), .ZN(
        n18273) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18273), .B1(
        n18340), .B2(n18267), .ZN(n18255) );
  OAI211_X1 U21382 ( .C1(n18348), .C2(n18380), .A(n18256), .B(n18255), .ZN(
        P3_U2964) );
  AOI22_X1 U21383 ( .A1(n18257), .A2(n18267), .B1(n18350), .B2(n18272), .ZN(
        n18259) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18273), .B1(
        n18352), .B2(n18390), .ZN(n18258) );
  OAI211_X1 U21385 ( .C1(n18260), .C2(n18288), .A(n18259), .B(n18258), .ZN(
        P3_U2965) );
  AOI22_X1 U21386 ( .A1(n18357), .A2(n18267), .B1(n18356), .B2(n18272), .ZN(
        n18262) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18273), .B1(
        n18358), .B2(n18390), .ZN(n18261) );
  OAI211_X1 U21388 ( .C1(n18361), .C2(n18288), .A(n18262), .B(n18261), .ZN(
        P3_U2966) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18273), .B1(
        n18362), .B2(n18272), .ZN(n18264) );
  AOI22_X1 U21390 ( .A1(n18363), .A2(n18267), .B1(n18364), .B2(n18390), .ZN(
        n18263) );
  OAI211_X1 U21391 ( .C1(n18367), .C2(n18288), .A(n18264), .B(n18263), .ZN(
        P3_U2967) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18273), .B1(
        n18368), .B2(n18272), .ZN(n18266) );
  AOI22_X1 U21393 ( .A1(n18370), .A2(n18390), .B1(n18318), .B2(n18296), .ZN(
        n18265) );
  OAI211_X1 U21394 ( .C1(n18321), .C2(n18276), .A(n18266), .B(n18265), .ZN(
        P3_U2968) );
  AOI22_X1 U21395 ( .A1(n18323), .A2(n18267), .B1(n18374), .B2(n18272), .ZN(
        n18269) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18273), .B1(
        n18377), .B2(n18390), .ZN(n18268) );
  OAI211_X1 U21397 ( .C1(n18326), .C2(n18288), .A(n18269), .B(n18268), .ZN(
        P3_U2969) );
  AOI22_X1 U21398 ( .A1(n18327), .A2(n18296), .B1(n18382), .B2(n18272), .ZN(
        n18271) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18273), .B1(
        n18384), .B2(n18390), .ZN(n18270) );
  OAI211_X1 U21400 ( .C1(n18330), .C2(n18276), .A(n18271), .B(n18270), .ZN(
        P3_U2970) );
  AOI22_X1 U21401 ( .A1(n18332), .A2(n18296), .B1(n18389), .B2(n18272), .ZN(
        n18275) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18273), .B1(
        n18392), .B2(n18390), .ZN(n18274) );
  OAI211_X1 U21403 ( .C1(n18338), .C2(n18276), .A(n18275), .B(n18274), .ZN(
        P3_U2971) );
  AND2_X1 U21404 ( .A1(n18462), .A2(n18343), .ZN(n18295) );
  AOI22_X1 U21405 ( .A1(n18345), .A2(n18322), .B1(n18339), .B2(n18295), .ZN(
        n18280) );
  AOI22_X1 U21406 ( .A1(n18344), .A2(n18277), .B1(n18343), .B2(n18341), .ZN(
        n18297) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18297), .B1(
        n18376), .B2(n18278), .ZN(n18279) );
  OAI211_X1 U21408 ( .C1(n18281), .C2(n18288), .A(n18280), .B(n18279), .ZN(
        P3_U2972) );
  AOI22_X1 U21409 ( .A1(n18351), .A2(n18322), .B1(n18350), .B2(n18295), .ZN(
        n18283) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18297), .B1(
        n18376), .B2(n18352), .ZN(n18282) );
  OAI211_X1 U21411 ( .C1(n18355), .C2(n18288), .A(n18283), .B(n18282), .ZN(
        P3_U2973) );
  AOI22_X1 U21412 ( .A1(n18357), .A2(n18296), .B1(n18356), .B2(n18295), .ZN(
        n18285) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18297), .B1(
        n18376), .B2(n18358), .ZN(n18284) );
  OAI211_X1 U21414 ( .C1(n18361), .C2(n18337), .A(n18285), .B(n18284), .ZN(
        P3_U2974) );
  AOI22_X1 U21415 ( .A1(n18314), .A2(n18322), .B1(n18362), .B2(n18295), .ZN(
        n18287) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18297), .B1(
        n18376), .B2(n18364), .ZN(n18286) );
  OAI211_X1 U21417 ( .C1(n18317), .C2(n18288), .A(n18287), .B(n18286), .ZN(
        P3_U2975) );
  AOI22_X1 U21418 ( .A1(n18369), .A2(n18296), .B1(n18368), .B2(n18295), .ZN(
        n18290) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18297), .B1(
        n18376), .B2(n18370), .ZN(n18289) );
  OAI211_X1 U21420 ( .C1(n18373), .C2(n18337), .A(n18290), .B(n18289), .ZN(
        P3_U2976) );
  AOI22_X1 U21421 ( .A1(n18323), .A2(n18296), .B1(n18374), .B2(n18295), .ZN(
        n18292) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18297), .B1(
        n18376), .B2(n18377), .ZN(n18291) );
  OAI211_X1 U21423 ( .C1(n18326), .C2(n18337), .A(n18292), .B(n18291), .ZN(
        P3_U2977) );
  AOI22_X1 U21424 ( .A1(n18383), .A2(n18296), .B1(n18382), .B2(n18295), .ZN(
        n18294) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18297), .B1(
        n18376), .B2(n18384), .ZN(n18293) );
  OAI211_X1 U21426 ( .C1(n18387), .C2(n18337), .A(n18294), .B(n18293), .ZN(
        P3_U2978) );
  AOI22_X1 U21427 ( .A1(n18391), .A2(n18296), .B1(n18389), .B2(n18295), .ZN(
        n18299) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18297), .B1(
        n18376), .B2(n18392), .ZN(n18298) );
  OAI211_X1 U21429 ( .C1(n18397), .C2(n18337), .A(n18299), .B(n18298), .ZN(
        P3_U2979) );
  AND2_X1 U21430 ( .A1(n18462), .A2(n18304), .ZN(n18331) );
  AOI22_X1 U21431 ( .A1(n18340), .A2(n18322), .B1(n18339), .B2(n18331), .ZN(
        n18306) );
  INV_X1 U21432 ( .A(n18300), .ZN(n18302) );
  OAI221_X1 U21433 ( .B1(n18304), .B2(n18303), .C1(n18304), .C2(n18302), .A(
        n18301), .ZN(n18334) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18334), .B1(
        n18345), .B2(n18390), .ZN(n18305) );
  OAI211_X1 U21435 ( .C1(n18348), .C2(n18307), .A(n18306), .B(n18305), .ZN(
        P3_U2980) );
  AOI22_X1 U21436 ( .A1(n18351), .A2(n18390), .B1(n18350), .B2(n18331), .ZN(
        n18309) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18352), .ZN(n18308) );
  OAI211_X1 U21438 ( .C1(n18355), .C2(n18337), .A(n18309), .B(n18308), .ZN(
        P3_U2981) );
  AOI22_X1 U21439 ( .A1(n18310), .A2(n18390), .B1(n18356), .B2(n18331), .ZN(
        n18312) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18358), .ZN(n18311) );
  OAI211_X1 U21441 ( .C1(n18313), .C2(n18337), .A(n18312), .B(n18311), .ZN(
        P3_U2982) );
  AOI22_X1 U21442 ( .A1(n18314), .A2(n18390), .B1(n18362), .B2(n18331), .ZN(
        n18316) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18364), .ZN(n18315) );
  OAI211_X1 U21444 ( .C1(n18317), .C2(n18337), .A(n18316), .B(n18315), .ZN(
        P3_U2983) );
  AOI22_X1 U21445 ( .A1(n18368), .A2(n18331), .B1(n18318), .B2(n18390), .ZN(
        n18320) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18370), .ZN(n18319) );
  OAI211_X1 U21447 ( .C1(n18321), .C2(n18337), .A(n18320), .B(n18319), .ZN(
        P3_U2984) );
  AOI22_X1 U21448 ( .A1(n18323), .A2(n18322), .B1(n18374), .B2(n18331), .ZN(
        n18325) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18377), .ZN(n18324) );
  OAI211_X1 U21450 ( .C1(n18326), .C2(n18380), .A(n18325), .B(n18324), .ZN(
        P3_U2985) );
  AOI22_X1 U21451 ( .A1(n18327), .A2(n18390), .B1(n18382), .B2(n18331), .ZN(
        n18329) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18384), .ZN(n18328) );
  OAI211_X1 U21453 ( .C1(n18330), .C2(n18337), .A(n18329), .B(n18328), .ZN(
        P3_U2986) );
  AOI22_X1 U21454 ( .A1(n18332), .A2(n18390), .B1(n18389), .B2(n18331), .ZN(
        n18336) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18392), .ZN(n18335) );
  OAI211_X1 U21456 ( .C1(n18338), .C2(n18337), .A(n18336), .B(n18335), .ZN(
        P3_U2987) );
  AND2_X1 U21457 ( .A1(n18462), .A2(n18342), .ZN(n18388) );
  AOI22_X1 U21458 ( .A1(n18340), .A2(n18390), .B1(n18339), .B2(n18388), .ZN(
        n18347) );
  AOI22_X1 U21459 ( .A1(n18344), .A2(n18343), .B1(n18342), .B2(n18341), .ZN(
        n18394) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18394), .B1(
        n18376), .B2(n18345), .ZN(n18346) );
  OAI211_X1 U21461 ( .C1(n18349), .C2(n18348), .A(n18347), .B(n18346), .ZN(
        P3_U2988) );
  AOI22_X1 U21462 ( .A1(n18376), .A2(n18351), .B1(n18350), .B2(n18388), .ZN(
        n18354) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18352), .ZN(n18353) );
  OAI211_X1 U21464 ( .C1(n18355), .C2(n18380), .A(n18354), .B(n18353), .ZN(
        P3_U2989) );
  AOI22_X1 U21465 ( .A1(n18357), .A2(n18390), .B1(n18356), .B2(n18388), .ZN(
        n18360) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18358), .ZN(n18359) );
  OAI211_X1 U21467 ( .C1(n18398), .C2(n18361), .A(n18360), .B(n18359), .ZN(
        P3_U2990) );
  AOI22_X1 U21468 ( .A1(n18363), .A2(n18390), .B1(n18362), .B2(n18388), .ZN(
        n18366) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18364), .ZN(n18365) );
  OAI211_X1 U21470 ( .C1(n18398), .C2(n18367), .A(n18366), .B(n18365), .ZN(
        P3_U2991) );
  AOI22_X1 U21471 ( .A1(n18369), .A2(n18390), .B1(n18368), .B2(n18388), .ZN(
        n18372) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18370), .ZN(n18371) );
  OAI211_X1 U21473 ( .C1(n18398), .C2(n18373), .A(n18372), .B(n18371), .ZN(
        P3_U2992) );
  AOI22_X1 U21474 ( .A1(n18376), .A2(n18375), .B1(n18374), .B2(n18388), .ZN(
        n18379) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18377), .ZN(n18378) );
  OAI211_X1 U21476 ( .C1(n18381), .C2(n18380), .A(n18379), .B(n18378), .ZN(
        P3_U2993) );
  AOI22_X1 U21477 ( .A1(n18383), .A2(n18390), .B1(n18382), .B2(n18388), .ZN(
        n18386) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18384), .ZN(n18385) );
  OAI211_X1 U21479 ( .C1(n18398), .C2(n18387), .A(n18386), .B(n18385), .ZN(
        P3_U2994) );
  AOI22_X1 U21480 ( .A1(n18391), .A2(n18390), .B1(n18389), .B2(n18388), .ZN(
        n18396) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18392), .ZN(n18395) );
  OAI211_X1 U21482 ( .C1(n18398), .C2(n18397), .A(n18396), .B(n18395), .ZN(
        P3_U2995) );
  NOR2_X1 U21483 ( .A1(n18438), .A2(n18399), .ZN(n18401) );
  OAI222_X1 U21484 ( .A1(n18405), .A2(n18404), .B1(n18403), .B2(n18402), .C1(
        n18401), .C2(n18400), .ZN(n18612) );
  OAI21_X1 U21485 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18406), .ZN(n18407) );
  OAI211_X1 U21486 ( .C1(n18439), .C2(n18409), .A(n18408), .B(n18407), .ZN(
        n18450) );
  NAND2_X1 U21487 ( .A1(n9629), .A2(n18598), .ZN(n18420) );
  AOI22_X1 U21488 ( .A1(n18413), .A2(n18420), .B1(n18438), .B2(n18412), .ZN(
        n18410) );
  NOR2_X1 U21489 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18410), .ZN(
        n18569) );
  INV_X1 U21490 ( .A(n18411), .ZN(n18431) );
  OAI21_X1 U21491 ( .B1(n18413), .B2(n9629), .A(n18412), .ZN(n18414) );
  AOI21_X1 U21492 ( .B1(n18431), .B2(n18415), .A(n18414), .ZN(n18570) );
  NAND2_X1 U21493 ( .A1(n18439), .A2(n18570), .ZN(n18416) );
  AOI22_X1 U21494 ( .A1(n18439), .A2(n18569), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18416), .ZN(n18448) );
  NOR2_X1 U21495 ( .A1(n18418), .A2(n18417), .ZN(n18422) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n9629), .B1(
        n18422), .B2(n18598), .ZN(n18594) );
  NOR2_X1 U21497 ( .A1(n18594), .A2(n18423), .ZN(n18426) );
  INV_X1 U21498 ( .A(n18420), .ZN(n18421) );
  OAI22_X1 U21499 ( .A1(n18422), .A2(n18585), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18421), .ZN(n18590) );
  OAI221_X1 U21500 ( .B1(n18590), .B2(n18594), .C1(n18590), .C2(n18423), .A(
        n18439), .ZN(n18424) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18426), .B1(
        n18425), .B2(n18424), .ZN(n18443) );
  INV_X1 U21502 ( .A(n18439), .ZN(n18440) );
  NOR2_X1 U21503 ( .A1(n18427), .A2(n18598), .ZN(n18428) );
  OAI21_X1 U21504 ( .B1(n18428), .B2(n18430), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18436) );
  OAI221_X1 U21505 ( .B1(n18431), .B2(n18592), .C1(n18431), .C2(n18430), .A(
        n18429), .ZN(n18435) );
  OAI211_X1 U21506 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18433), .B(n18432), .ZN(
        n18434) );
  OAI221_X1 U21507 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18436), 
        .C1(n18584), .C2(n18435), .A(n18434), .ZN(n18437) );
  AOI21_X1 U21508 ( .B1(n18438), .B2(n18578), .A(n18437), .ZN(n18581) );
  AOI22_X1 U21509 ( .A1(n18440), .A2(n18584), .B1(n18581), .B2(n18439), .ZN(
        n18444) );
  AND2_X1 U21510 ( .A1(n18443), .A2(n18444), .ZN(n18441) );
  OAI221_X1 U21511 ( .B1(n18443), .B2(n18444), .C1(n18442), .C2(n18441), .A(
        n20778), .ZN(n18447) );
  AOI21_X1 U21512 ( .B1(n20778), .B2(n18445), .A(n18444), .ZN(n18446) );
  AOI222_X1 U21513 ( .A1(n18448), .A2(n18447), .B1(n18448), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18447), .C2(n18446), .ZN(
        n18449) );
  NOR4_X1 U21514 ( .A1(n18451), .A2(n18612), .A3(n18450), .A4(n18449), .ZN(
        n18460) );
  OAI211_X1 U21515 ( .C1(n18453), .C2(n18452), .A(n18617), .B(n18460), .ZN(
        n18565) );
  INV_X1 U21516 ( .A(n18565), .ZN(n18454) );
  NOR2_X1 U21517 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18613), .ZN(n18461) );
  NOR2_X1 U21518 ( .A1(n18454), .A2(n18461), .ZN(n18463) );
  OAI211_X1 U21519 ( .C1(P3_STATE2_REG_1__SCAN_IN), .C2(n18462), .A(n18463), 
        .B(n18455), .ZN(n18457) );
  AOI22_X1 U21520 ( .A1(n18593), .A2(n18625), .B1(n18620), .B2(n18614), .ZN(
        n18456) );
  AOI22_X1 U21521 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18457), .B1(n18456), 
        .B2(n18622), .ZN(n18458) );
  OAI21_X1 U21522 ( .B1(n18460), .B2(n18459), .A(n18458), .ZN(P3_U2996) );
  NAND2_X1 U21523 ( .A1(n18620), .A2(n18614), .ZN(n18466) );
  NAND3_X1 U21524 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n18461), .ZN(n18469) );
  NAND3_X1 U21525 ( .A1(n18464), .A2(n18463), .A3(n18462), .ZN(n18465) );
  NAND4_X1 U21526 ( .A1(n18467), .A2(n18466), .A3(n18469), .A4(n18465), .ZN(
        P3_U2997) );
  OAI21_X1 U21527 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18468), .ZN(n18471) );
  INV_X1 U21528 ( .A(n18469), .ZN(n18470) );
  AOI21_X1 U21529 ( .B1(n18472), .B2(n18471), .A(n18470), .ZN(P3_U2998) );
  AND2_X1 U21530 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n9595), .ZN(P3_U2999) );
  AND2_X1 U21531 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n9594), .ZN(P3_U3000) );
  AND2_X1 U21532 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n9595), .ZN(P3_U3001) );
  AND2_X1 U21533 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n9594), .ZN(P3_U3002) );
  AND2_X1 U21534 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n9595), .ZN(P3_U3003) );
  AND2_X1 U21535 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n9594), .ZN(P3_U3004) );
  AND2_X1 U21536 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n9595), .ZN(P3_U3005) );
  AND2_X1 U21537 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n9594), .ZN(P3_U3006) );
  AND2_X1 U21538 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n9594), .ZN(P3_U3007) );
  AND2_X1 U21539 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n9595), .ZN(P3_U3008) );
  AND2_X1 U21540 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n9594), .ZN(P3_U3009) );
  AND2_X1 U21541 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n9595), .ZN(P3_U3010) );
  AND2_X1 U21542 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n9594), .ZN(P3_U3011) );
  AND2_X1 U21543 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n9595), .ZN(P3_U3012) );
  AND2_X1 U21544 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n9594), .ZN(P3_U3013) );
  AND2_X1 U21545 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n9595), .ZN(P3_U3014) );
  AND2_X1 U21546 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n9594), .ZN(P3_U3015) );
  AND2_X1 U21547 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n9595), .ZN(P3_U3016) );
  AND2_X1 U21548 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n9595), .ZN(P3_U3017) );
  AND2_X1 U21549 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n9594), .ZN(P3_U3018) );
  AND2_X1 U21550 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n9595), .ZN(P3_U3019) );
  AND2_X1 U21551 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n9594), .ZN(P3_U3020) );
  AND2_X1 U21552 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n9594), .ZN(P3_U3021)
         );
  AND2_X1 U21553 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n9595), .ZN(P3_U3022)
         );
  AND2_X1 U21554 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n9594), .ZN(P3_U3023)
         );
  AND2_X1 U21555 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n9595), .ZN(P3_U3024)
         );
  AND2_X1 U21556 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n9594), .ZN(P3_U3025)
         );
  AND2_X1 U21557 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n9595), .ZN(P3_U3026)
         );
  AND2_X1 U21558 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n9594), .ZN(P3_U3027)
         );
  AND2_X1 U21559 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n9595), .ZN(P3_U3028)
         );
  INV_X1 U21560 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18627) );
  AOI21_X1 U21561 ( .B1(HOLD), .B2(n18474), .A(n18627), .ZN(n18476) );
  NOR2_X1 U21562 ( .A1(n18613), .A2(n18483), .ZN(n18482) );
  OAI21_X1 U21563 ( .B1(n18482), .B2(n18488), .A(n18490), .ZN(n18475) );
  NAND3_X1 U21564 ( .A1(NA), .A2(n18488), .A3(n18483), .ZN(n18481) );
  OAI211_X1 U21565 ( .C1(n18610), .C2(n18476), .A(n18475), .B(n18481), .ZN(
        P3_U3029) );
  NOR2_X1 U21566 ( .A1(n18490), .A2(n20585), .ZN(n18486) );
  NOR3_X1 U21567 ( .A1(n18486), .A2(n18627), .A3(n18488), .ZN(n18477) );
  NOR2_X1 U21568 ( .A1(n18477), .A2(n18482), .ZN(n18479) );
  OAI211_X1 U21569 ( .C1(n20585), .C2(n18480), .A(n18479), .B(n18478), .ZN(
        P3_U3030) );
  AOI21_X1 U21570 ( .B1(n18488), .B2(n18481), .A(n18482), .ZN(n18489) );
  INV_X1 U21571 ( .A(NA), .ZN(n20592) );
  AOI22_X1 U21572 ( .A1(n18483), .A2(n18627), .B1(n20592), .B2(n18482), .ZN(
        n18484) );
  INV_X1 U21573 ( .A(n18484), .ZN(n18485) );
  OAI22_X1 U21574 ( .A1(n18486), .A2(n18485), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18487) );
  OAI22_X1 U21575 ( .A1(n18489), .A2(n18490), .B1(n18488), .B2(n18487), .ZN(
        P3_U3031) );
  OAI222_X1 U21576 ( .A1(n18600), .A2(n18552), .B1(n18491), .B2(n18610), .C1(
        n18492), .C2(n18538), .ZN(P3_U3032) );
  OAI222_X1 U21577 ( .A1(n18538), .A2(n18494), .B1(n18493), .B2(n18610), .C1(
        n18492), .C2(n18552), .ZN(P3_U3033) );
  OAI222_X1 U21578 ( .A1(n18538), .A2(n18496), .B1(n18495), .B2(n18610), .C1(
        n18494), .C2(n18552), .ZN(P3_U3034) );
  OAI222_X1 U21579 ( .A1(n18538), .A2(n18498), .B1(n18497), .B2(n18610), .C1(
        n18496), .C2(n18552), .ZN(P3_U3035) );
  OAI222_X1 U21580 ( .A1(n18538), .A2(n18500), .B1(n18499), .B2(n18610), .C1(
        n18498), .C2(n18552), .ZN(P3_U3036) );
  OAI222_X1 U21581 ( .A1(n18538), .A2(n18502), .B1(n18501), .B2(n18610), .C1(
        n18500), .C2(n18552), .ZN(P3_U3037) );
  OAI222_X1 U21582 ( .A1(n18538), .A2(n18505), .B1(n18503), .B2(n18610), .C1(
        n18502), .C2(n18552), .ZN(P3_U3038) );
  OAI222_X1 U21583 ( .A1(n18505), .A2(n18552), .B1(n18504), .B2(n18610), .C1(
        n18506), .C2(n18538), .ZN(P3_U3039) );
  INV_X1 U21584 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18508) );
  OAI222_X1 U21585 ( .A1(n18538), .A2(n18508), .B1(n18507), .B2(n18610), .C1(
        n18506), .C2(n18552), .ZN(P3_U3040) );
  OAI222_X1 U21586 ( .A1(n18538), .A2(n18510), .B1(n18509), .B2(n18610), .C1(
        n18508), .C2(n18552), .ZN(P3_U3041) );
  OAI222_X1 U21587 ( .A1(n18538), .A2(n18513), .B1(n18511), .B2(n18610), .C1(
        n18510), .C2(n18552), .ZN(P3_U3042) );
  INV_X1 U21588 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18514) );
  OAI222_X1 U21589 ( .A1(n18513), .A2(n18552), .B1(n18512), .B2(n18610), .C1(
        n18514), .C2(n18538), .ZN(P3_U3043) );
  INV_X1 U21590 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18517) );
  OAI222_X1 U21591 ( .A1(n18538), .A2(n18517), .B1(n18515), .B2(n18610), .C1(
        n18514), .C2(n18552), .ZN(P3_U3044) );
  INV_X1 U21592 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18518) );
  OAI222_X1 U21593 ( .A1(n18517), .A2(n18552), .B1(n18516), .B2(n18610), .C1(
        n18518), .C2(n18538), .ZN(P3_U3045) );
  INV_X1 U21594 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18520) );
  OAI222_X1 U21595 ( .A1(n18538), .A2(n18520), .B1(n18519), .B2(n18610), .C1(
        n18518), .C2(n18552), .ZN(P3_U3046) );
  INV_X1 U21596 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18522) );
  OAI222_X1 U21597 ( .A1(n18538), .A2(n18522), .B1(n18521), .B2(n18610), .C1(
        n18520), .C2(n18552), .ZN(P3_U3047) );
  OAI222_X1 U21598 ( .A1(n18538), .A2(n18524), .B1(n18523), .B2(n18610), .C1(
        n18522), .C2(n18552), .ZN(P3_U3048) );
  OAI222_X1 U21599 ( .A1(n18538), .A2(n18526), .B1(n18525), .B2(n18610), .C1(
        n18524), .C2(n18552), .ZN(P3_U3049) );
  OAI222_X1 U21600 ( .A1(n18538), .A2(n18528), .B1(n18527), .B2(n18610), .C1(
        n18526), .C2(n18552), .ZN(P3_U3050) );
  OAI222_X1 U21601 ( .A1(n18538), .A2(n18530), .B1(n18529), .B2(n18610), .C1(
        n18528), .C2(n18552), .ZN(P3_U3051) );
  OAI222_X1 U21602 ( .A1(n18538), .A2(n18532), .B1(n18531), .B2(n18610), .C1(
        n18530), .C2(n18552), .ZN(P3_U3052) );
  OAI222_X1 U21603 ( .A1(n18538), .A2(n18535), .B1(n18533), .B2(n18610), .C1(
        n18532), .C2(n18552), .ZN(P3_U3053) );
  OAI222_X1 U21604 ( .A1(n18535), .A2(n18552), .B1(n18534), .B2(n18610), .C1(
        n18536), .C2(n18538), .ZN(P3_U3054) );
  OAI222_X1 U21605 ( .A1(n18538), .A2(n18539), .B1(n18537), .B2(n18610), .C1(
        n18536), .C2(n18552), .ZN(P3_U3055) );
  OAI222_X1 U21606 ( .A1(n18538), .A2(n18541), .B1(n18540), .B2(n18610), .C1(
        n18539), .C2(n18552), .ZN(P3_U3056) );
  OAI222_X1 U21607 ( .A1(n18538), .A2(n18543), .B1(n18542), .B2(n18610), .C1(
        n18541), .C2(n18552), .ZN(P3_U3057) );
  INV_X1 U21608 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18546) );
  OAI222_X1 U21609 ( .A1(n18538), .A2(n18546), .B1(n18544), .B2(n18610), .C1(
        n18543), .C2(n18552), .ZN(P3_U3058) );
  INV_X1 U21610 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18547) );
  OAI222_X1 U21611 ( .A1(n18546), .A2(n18552), .B1(n18545), .B2(n18610), .C1(
        n18547), .C2(n18538), .ZN(P3_U3059) );
  OAI222_X1 U21612 ( .A1(n18538), .A2(n18551), .B1(n18548), .B2(n18610), .C1(
        n18547), .C2(n18552), .ZN(P3_U3060) );
  OAI222_X1 U21613 ( .A1(n18552), .A2(n18551), .B1(n18550), .B2(n18610), .C1(
        n18549), .C2(n18538), .ZN(P3_U3061) );
  INV_X1 U21614 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18553) );
  AOI22_X1 U21615 ( .A1(n18610), .A2(n18554), .B1(n18553), .B2(n18629), .ZN(
        P3_U3274) );
  INV_X1 U21616 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18602) );
  INV_X1 U21617 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18555) );
  AOI22_X1 U21618 ( .A1(n18610), .A2(n18602), .B1(n18555), .B2(n18629), .ZN(
        P3_U3275) );
  INV_X1 U21619 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18556) );
  AOI22_X1 U21620 ( .A1(n18610), .A2(n18557), .B1(n18556), .B2(n18629), .ZN(
        P3_U3276) );
  INV_X1 U21621 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18608) );
  INV_X1 U21622 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18558) );
  AOI22_X1 U21623 ( .A1(n18610), .A2(n18608), .B1(n18558), .B2(n18629), .ZN(
        P3_U3277) );
  INV_X1 U21624 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18560) );
  AOI21_X1 U21625 ( .B1(n9595), .B2(n18560), .A(n18559), .ZN(P3_U3280) );
  OAI21_X1 U21626 ( .B1(n18563), .B2(n18562), .A(n18561), .ZN(P3_U3281) );
  OAI221_X1 U21627 ( .B1(n18566), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18566), 
        .C2(n18565), .A(n18564), .ZN(P3_U3282) );
  INV_X1 U21628 ( .A(n18567), .ZN(n18568) );
  AOI22_X1 U21629 ( .A1(n18632), .A2(n18569), .B1(n18593), .B2(n18568), .ZN(
        n18574) );
  INV_X1 U21630 ( .A(n18570), .ZN(n18571) );
  AOI21_X1 U21631 ( .B1(n18632), .B2(n18571), .A(n18599), .ZN(n18573) );
  OAI22_X1 U21632 ( .A1(n18599), .A2(n18574), .B1(n18573), .B2(n18572), .ZN(
        P3_U3285) );
  AOI22_X1 U21633 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18576), .B2(n18575), .ZN(
        n18586) );
  NOR2_X1 U21634 ( .A1(n18577), .A2(n18595), .ZN(n18587) );
  INV_X1 U21635 ( .A(n18593), .ZN(n18579) );
  OAI22_X1 U21636 ( .A1(n18581), .A2(n18580), .B1(n18579), .B2(n18578), .ZN(
        n18582) );
  AOI21_X1 U21637 ( .B1(n18586), .B2(n18587), .A(n18582), .ZN(n18583) );
  AOI22_X1 U21638 ( .A1(n18599), .A2(n18584), .B1(n18583), .B2(n18596), .ZN(
        P3_U3288) );
  INV_X1 U21639 ( .A(n18585), .ZN(n18589) );
  INV_X1 U21640 ( .A(n18586), .ZN(n18588) );
  AOI222_X1 U21641 ( .A1(n18590), .A2(n18632), .B1(n18593), .B2(n18589), .C1(
        n18588), .C2(n18587), .ZN(n18591) );
  AOI22_X1 U21642 ( .A1(n18599), .A2(n18592), .B1(n18591), .B2(n18596), .ZN(
        P3_U3289) );
  AOI222_X1 U21643 ( .A1(n18595), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18632), 
        .B2(n18594), .C1(n18598), .C2(n18593), .ZN(n18597) );
  AOI22_X1 U21644 ( .A1(n18599), .A2(n18598), .B1(n18597), .B2(n18596), .ZN(
        P3_U3290) );
  AOI21_X1 U21645 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18601) );
  AOI22_X1 U21646 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18601), .B2(n18600), .ZN(n18603) );
  AOI22_X1 U21647 ( .A1(n18604), .A2(n18603), .B1(n18602), .B2(n18607), .ZN(
        P3_U3292) );
  NOR2_X1 U21648 ( .A1(n18607), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18605) );
  AOI22_X1 U21649 ( .A1(n18608), .A2(n18607), .B1(n18606), .B2(n18605), .ZN(
        P3_U3293) );
  INV_X1 U21650 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18609) );
  AOI22_X1 U21651 ( .A1(n18610), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18609), 
        .B2(n18629), .ZN(P3_U3294) );
  MUX2_X1 U21652 ( .A(P3_MORE_REG_SCAN_IN), .B(n18612), .S(n18611), .Z(
        P3_U3295) );
  AOI21_X1 U21653 ( .B1(n18614), .B2(n18613), .A(n18634), .ZN(n18615) );
  OAI21_X1 U21654 ( .B1(n18617), .B2(n18616), .A(n18615), .ZN(n18628) );
  OAI21_X1 U21655 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18619), .A(n18618), 
        .ZN(n18621) );
  AOI211_X1 U21656 ( .C1(n18633), .C2(n18621), .A(n18620), .B(n18631), .ZN(
        n18623) );
  NOR2_X1 U21657 ( .A1(n18623), .A2(n18622), .ZN(n18624) );
  OAI21_X1 U21658 ( .B1(n18625), .B2(n18624), .A(n18628), .ZN(n18626) );
  OAI21_X1 U21659 ( .B1(n18628), .B2(n18627), .A(n18626), .ZN(P3_U3296) );
  OAI22_X1 U21660 ( .A1(n18629), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18610), .ZN(n18630) );
  INV_X1 U21661 ( .A(n18630), .ZN(P3_U3297) );
  AOI21_X1 U21662 ( .B1(n18632), .B2(n18631), .A(n18634), .ZN(n18636) );
  INV_X1 U21663 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18635) );
  AOI22_X1 U21664 ( .A1(n18636), .A2(n18635), .B1(n18634), .B2(n18633), .ZN(
        P3_U3298) );
  INV_X1 U21665 ( .A(n18636), .ZN(n18638) );
  OAI21_X1 U21666 ( .B1(n18638), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18637), 
        .ZN(n18639) );
  INV_X1 U21667 ( .A(n18639), .ZN(P3_U3299) );
  INV_X1 U21668 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18640) );
  NAND2_X1 U21669 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19634), .ZN(n19624) );
  NAND2_X1 U21670 ( .A1(n19622), .A2(n20756), .ZN(n19623) );
  OAI21_X1 U21671 ( .B1(n19622), .B2(n19624), .A(n19623), .ZN(n19689) );
  OAI21_X1 U21672 ( .B1(n19622), .B2(n18640), .A(n9597), .ZN(P2_U2815) );
  INV_X1 U21673 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18642) );
  OAI22_X1 U21674 ( .A1(n18643), .A2(n18642), .B1(n19751), .B2(n18641), .ZN(
        P2_U2816) );
  AOI21_X1 U21675 ( .B1(n19622), .B2(n19634), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18644) );
  AOI22_X1 U21676 ( .A1(n19761), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18644), 
        .B2(n19758), .ZN(P2_U2817) );
  AOI21_X1 U21677 ( .B1(n19628), .B2(n18645), .A(n9597), .ZN(n19685) );
  INV_X1 U21678 ( .A(n19685), .ZN(n19687) );
  OAI21_X1 U21679 ( .B1(n19689), .B2(n19692), .A(n19687), .ZN(P2_U2818) );
  NOR4_X1 U21680 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18649) );
  NOR4_X1 U21681 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18648) );
  NOR4_X1 U21682 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18647) );
  NOR4_X1 U21683 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18646) );
  NAND4_X1 U21684 ( .A1(n18649), .A2(n18648), .A3(n18647), .A4(n18646), .ZN(
        n18655) );
  NOR4_X1 U21685 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18653) );
  AOI211_X1 U21686 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_7__SCAN_IN), .B(
        P2_DATAWIDTH_REG_25__SCAN_IN), .ZN(n18652) );
  NOR4_X1 U21687 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18651) );
  NOR4_X1 U21688 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18650) );
  NAND4_X1 U21689 ( .A1(n18653), .A2(n18652), .A3(n18651), .A4(n18650), .ZN(
        n18654) );
  NOR2_X1 U21690 ( .A1(n18655), .A2(n18654), .ZN(n18663) );
  INV_X1 U21691 ( .A(n18663), .ZN(n18662) );
  NOR2_X1 U21692 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18662), .ZN(n18656) );
  INV_X1 U21693 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19684) );
  AOI22_X1 U21694 ( .A1(n18656), .A2(n18657), .B1(n18662), .B2(n19684), .ZN(
        P2_U2820) );
  INV_X1 U21695 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19688) );
  INV_X1 U21696 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19686) );
  NAND3_X1 U21697 ( .A1(n18657), .A2(n19688), .A3(n19686), .ZN(n18661) );
  INV_X1 U21698 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19682) );
  AOI22_X1 U21699 ( .A1(n18656), .A2(n18661), .B1(n18662), .B2(n19682), .ZN(
        P2_U2821) );
  NAND2_X1 U21700 ( .A1(n18656), .A2(n19688), .ZN(n18660) );
  OAI21_X1 U21701 ( .B1(n18657), .B2(n19636), .A(n18663), .ZN(n18658) );
  OAI21_X1 U21702 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18663), .A(n18658), 
        .ZN(n18659) );
  OAI221_X1 U21703 ( .B1(n18660), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18660), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18659), .ZN(P2_U2822) );
  INV_X1 U21704 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19680) );
  OAI221_X1 U21705 ( .B1(n18663), .B2(n19680), .C1(n18662), .C2(n18661), .A(
        n18660), .ZN(P2_U2823) );
  INV_X1 U21706 ( .A(n18664), .ZN(n18666) );
  AOI21_X1 U21707 ( .B1(n18669), .B2(n18666), .A(n18665), .ZN(n18667) );
  AOI21_X1 U21708 ( .B1(n18865), .B2(n18668), .A(n18667), .ZN(n18676) );
  AOI22_X1 U21709 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n18867), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n18866), .ZN(n18675) );
  AOI22_X1 U21710 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18874), .B1(
        n18669), .B2(n18857), .ZN(n18674) );
  OAI22_X1 U21711 ( .A1(n18671), .A2(n18870), .B1(n18836), .B2(n18670), .ZN(
        n18672) );
  INV_X1 U21712 ( .A(n18672), .ZN(n18673) );
  NAND4_X1 U21713 ( .A1(n18676), .A2(n18675), .A3(n18674), .A4(n18673), .ZN(
        P2_U2835) );
  NAND2_X1 U21714 ( .A1(n13945), .A2(n18677), .ZN(n18678) );
  XOR2_X1 U21715 ( .A(n18679), .B(n18678), .Z(n18688) );
  OAI21_X1 U21716 ( .B1(n20834), .B2(n18774), .A(n18772), .ZN(n18682) );
  OAI22_X1 U21717 ( .A1(n18680), .A2(n18852), .B1(n20750), .B2(n18832), .ZN(
        n18681) );
  AOI211_X1 U21718 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18866), .A(n18682), .B(
        n18681), .ZN(n18687) );
  OAI22_X1 U21719 ( .A1(n18684), .A2(n18870), .B1(n18683), .B2(n18836), .ZN(
        n18685) );
  INV_X1 U21720 ( .A(n18685), .ZN(n18686) );
  OAI211_X1 U21721 ( .C1(n18877), .C2(n18688), .A(n18687), .B(n18686), .ZN(
        P2_U2836) );
  NOR2_X1 U21722 ( .A1(n10466), .A2(n18689), .ZN(n18691) );
  XOR2_X1 U21723 ( .A(n18691), .B(n18690), .Z(n18699) );
  AOI22_X1 U21724 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n18866), .ZN(n18692) );
  OAI21_X1 U21725 ( .B1(n18693), .B2(n18852), .A(n18692), .ZN(n18694) );
  AOI211_X1 U21726 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18867), .A(n18822), 
        .B(n18694), .ZN(n18698) );
  AOI22_X1 U21727 ( .A1(n18696), .A2(n18863), .B1(n18695), .B2(n18840), .ZN(
        n18697) );
  OAI211_X1 U21728 ( .C1(n18877), .C2(n18699), .A(n18698), .B(n18697), .ZN(
        P2_U2837) );
  NAND2_X1 U21729 ( .A1(n13945), .A2(n18700), .ZN(n18701) );
  XOR2_X1 U21730 ( .A(n18702), .B(n18701), .Z(n18713) );
  OAI21_X1 U21731 ( .B1(n19656), .B2(n18774), .A(n18772), .ZN(n18706) );
  OAI22_X1 U21732 ( .A1(n18704), .A2(n18852), .B1(n18703), .B2(n18832), .ZN(
        n18705) );
  AOI211_X1 U21733 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18866), .A(n18706), .B(
        n18705), .ZN(n18712) );
  INV_X1 U21734 ( .A(n18707), .ZN(n18710) );
  INV_X1 U21735 ( .A(n18708), .ZN(n18709) );
  AOI22_X1 U21736 ( .A1(n18710), .A2(n18863), .B1(n18840), .B2(n18709), .ZN(
        n18711) );
  OAI211_X1 U21737 ( .C1(n18877), .C2(n18713), .A(n18712), .B(n18711), .ZN(
        P2_U2838) );
  NOR2_X1 U21738 ( .A1(n10466), .A2(n18714), .ZN(n18716) );
  XOR2_X1 U21739 ( .A(n18716), .B(n18715), .Z(n18723) );
  AOI22_X1 U21740 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_16__SCAN_IN), .B2(n18866), .ZN(n18717) );
  OAI21_X1 U21741 ( .B1(n18718), .B2(n18852), .A(n18717), .ZN(n18719) );
  AOI211_X1 U21742 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18867), .A(n18822), 
        .B(n18719), .ZN(n18722) );
  NOR2_X1 U21743 ( .A1(n18880), .A2(n18870), .ZN(n18720) );
  AOI21_X1 U21744 ( .B1(n18913), .B2(n18863), .A(n18720), .ZN(n18721) );
  OAI211_X1 U21745 ( .C1(n18877), .C2(n18723), .A(n18722), .B(n18721), .ZN(
        P2_U2839) );
  OAI22_X1 U21746 ( .A1(n18725), .A2(n18852), .B1(n18724), .B2(n18837), .ZN(
        n18726) );
  AOI211_X1 U21747 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18867), .A(n18822), 
        .B(n18726), .ZN(n18735) );
  NAND2_X1 U21748 ( .A1(n13945), .A2(n18727), .ZN(n18728) );
  XNOR2_X1 U21749 ( .A(n18729), .B(n18728), .ZN(n18733) );
  OAI22_X1 U21750 ( .A1(n18731), .A2(n18836), .B1(n18730), .B2(n18870), .ZN(
        n18732) );
  AOI21_X1 U21751 ( .B1(n18827), .B2(n18733), .A(n18732), .ZN(n18734) );
  OAI211_X1 U21752 ( .C1(n18736), .C2(n18832), .A(n18735), .B(n18734), .ZN(
        P2_U2840) );
  OR2_X1 U21753 ( .A1(n10466), .A2(n18737), .ZN(n18746) );
  XNOR2_X1 U21754 ( .A(n18746), .B(n18738), .ZN(n18745) );
  AOI22_X1 U21755 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n18866), .ZN(n18739) );
  OAI21_X1 U21756 ( .B1(n18740), .B2(n18852), .A(n18739), .ZN(n18741) );
  AOI211_X1 U21757 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18867), .A(n18822), 
        .B(n18741), .ZN(n18744) );
  AOI22_X1 U21758 ( .A1(n18917), .A2(n18863), .B1(n18840), .B2(n18742), .ZN(
        n18743) );
  OAI211_X1 U21759 ( .C1(n18877), .C2(n18745), .A(n18744), .B(n18743), .ZN(
        P2_U2841) );
  AOI211_X1 U21760 ( .C1(n18755), .C2(n18747), .A(n18877), .B(n18746), .ZN(
        n18753) );
  NAND2_X1 U21761 ( .A1(n18748), .A2(n18865), .ZN(n18751) );
  AOI22_X1 U21762 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18874), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n18867), .ZN(n18750) );
  NAND2_X1 U21763 ( .A1(n18866), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n18749) );
  NAND4_X1 U21764 ( .A1(n18751), .A2(n18750), .A3(n18772), .A4(n18749), .ZN(
        n18752) );
  NOR2_X1 U21765 ( .A1(n18753), .A2(n18752), .ZN(n18757) );
  AOI22_X1 U21766 ( .A1(n18857), .A2(n18755), .B1(n18840), .B2(n18754), .ZN(
        n18756) );
  OAI211_X1 U21767 ( .C1(n18758), .C2(n18836), .A(n18757), .B(n18756), .ZN(
        P2_U2842) );
  AOI22_X1 U21768 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n18866), .ZN(n18759) );
  OAI21_X1 U21769 ( .B1(n18760), .B2(n18852), .A(n18759), .ZN(n18761) );
  AOI211_X1 U21770 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n18867), .A(n18822), 
        .B(n18761), .ZN(n18769) );
  NAND2_X1 U21771 ( .A1(n13945), .A2(n18762), .ZN(n18763) );
  XNOR2_X1 U21772 ( .A(n18764), .B(n18763), .ZN(n18767) );
  INV_X1 U21773 ( .A(n18765), .ZN(n18766) );
  AOI22_X1 U21774 ( .A1(n18767), .A2(n18827), .B1(n18840), .B2(n18766), .ZN(
        n18768) );
  OAI211_X1 U21775 ( .C1(n18770), .C2(n18836), .A(n18769), .B(n18768), .ZN(
        P2_U2844) );
  AOI22_X1 U21776 ( .A1(n18771), .A2(n18865), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n18866), .ZN(n18773) );
  OAI211_X1 U21777 ( .C1(n11030), .C2(n18774), .A(n18773), .B(n18772), .ZN(
        n18775) );
  AOI21_X1 U21778 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18874), .A(
        n18775), .ZN(n18781) );
  NOR2_X1 U21779 ( .A1(n10466), .A2(n18776), .ZN(n18778) );
  XNOR2_X1 U21780 ( .A(n18778), .B(n18777), .ZN(n18779) );
  AOI22_X1 U21781 ( .A1(n18779), .A2(n18827), .B1(n18840), .B2(n18897), .ZN(
        n18780) );
  OAI211_X1 U21782 ( .C1(n18925), .C2(n18836), .A(n18781), .B(n18780), .ZN(
        P2_U2845) );
  INV_X1 U21783 ( .A(n18782), .ZN(n18783) );
  OAI22_X1 U21784 ( .A1(n18783), .A2(n18852), .B1(n12324), .B2(n18837), .ZN(
        n18784) );
  AOI211_X1 U21785 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18867), .A(n18822), .B(
        n18784), .ZN(n18793) );
  NAND2_X1 U21786 ( .A1(n13945), .A2(n18785), .ZN(n18786) );
  XNOR2_X1 U21787 ( .A(n18787), .B(n18786), .ZN(n18791) );
  OAI22_X1 U21788 ( .A1(n18789), .A2(n18836), .B1(n18870), .B2(n18788), .ZN(
        n18790) );
  AOI21_X1 U21789 ( .B1(n18827), .B2(n18791), .A(n18790), .ZN(n18792) );
  OAI211_X1 U21790 ( .C1(n18794), .C2(n18832), .A(n18793), .B(n18792), .ZN(
        P2_U2846) );
  NOR2_X1 U21791 ( .A1(n10466), .A2(n18795), .ZN(n18797) );
  XOR2_X1 U21792 ( .A(n18797), .B(n18796), .Z(n18807) );
  INV_X1 U21793 ( .A(n18798), .ZN(n18800) );
  AOI22_X1 U21794 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n18866), .ZN(n18799) );
  OAI21_X1 U21795 ( .B1(n18800), .B2(n18852), .A(n18799), .ZN(n18801) );
  AOI211_X1 U21796 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n18867), .A(n18822), .B(
        n18801), .ZN(n18806) );
  OAI22_X1 U21797 ( .A1(n18803), .A2(n18870), .B1(n18802), .B2(n18836), .ZN(
        n18804) );
  INV_X1 U21798 ( .A(n18804), .ZN(n18805) );
  OAI211_X1 U21799 ( .C1(n18877), .C2(n18807), .A(n18806), .B(n18805), .ZN(
        P2_U2847) );
  AOI22_X1 U21800 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_6__SCAN_IN), .B2(n18866), .ZN(n18808) );
  OAI21_X1 U21801 ( .B1(n18809), .B2(n18852), .A(n18808), .ZN(n18810) );
  AOI211_X1 U21802 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n18867), .A(n18822), .B(
        n18810), .ZN(n18817) );
  NOR2_X1 U21803 ( .A1(n10466), .A2(n18811), .ZN(n18813) );
  XNOR2_X1 U21804 ( .A(n18813), .B(n18812), .ZN(n18815) );
  AOI22_X1 U21805 ( .A1(n18815), .A2(n18827), .B1(n18840), .B2(n18814), .ZN(
        n18816) );
  OAI211_X1 U21806 ( .C1(n18836), .C2(n18818), .A(n18817), .B(n18816), .ZN(
        P2_U2849) );
  AOI22_X1 U21807 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n18874), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n18866), .ZN(n18819) );
  OAI21_X1 U21808 ( .B1(n18820), .B2(n18852), .A(n18819), .ZN(n18821) );
  AOI211_X1 U21809 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18867), .A(n18822), .B(
        n18821), .ZN(n18830) );
  NAND2_X1 U21810 ( .A1(n13945), .A2(n18823), .ZN(n18824) );
  XNOR2_X1 U21811 ( .A(n18825), .B(n18824), .ZN(n18828) );
  AOI22_X1 U21812 ( .A1(n18828), .A2(n18827), .B1(n18840), .B2(n18826), .ZN(
        n18829) );
  OAI211_X1 U21813 ( .C1(n18836), .C2(n18935), .A(n18830), .B(n18829), .ZN(
        P2_U2850) );
  INV_X1 U21814 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18831) );
  OAI22_X1 U21815 ( .A1(n18833), .A2(n18852), .B1(n18832), .B2(n18831), .ZN(
        n18834) );
  INV_X1 U21816 ( .A(n18834), .ZN(n18848) );
  INV_X1 U21817 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18902) );
  OAI22_X1 U21818 ( .A1(n18837), .A2(n18902), .B1(n18836), .B2(n18835), .ZN(
        n18838) );
  AOI211_X1 U21819 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n18867), .A(n18839), .B(
        n18838), .ZN(n18847) );
  INV_X1 U21820 ( .A(n18931), .ZN(n18900) );
  AOI22_X1 U21821 ( .A1(n18900), .A2(n18873), .B1(n18840), .B2(n18984), .ZN(
        n18846) );
  INV_X1 U21822 ( .A(n18988), .ZN(n18844) );
  NOR2_X1 U21823 ( .A1(n10466), .A2(n18841), .ZN(n18843) );
  AOI21_X1 U21824 ( .B1(n18844), .B2(n18843), .A(n18877), .ZN(n18842) );
  OAI21_X1 U21825 ( .B1(n18844), .B2(n18843), .A(n18842), .ZN(n18845) );
  NAND4_X1 U21826 ( .A1(n18848), .A2(n18847), .A3(n18846), .A4(n18845), .ZN(
        P2_U2851) );
  NAND2_X1 U21827 ( .A1(n18866), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n18850) );
  AOI22_X1 U21828 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18867), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18874), .ZN(n18849) );
  OAI211_X1 U21829 ( .C1(n18852), .C2(n18851), .A(n18850), .B(n18849), .ZN(
        n18855) );
  NOR2_X1 U21830 ( .A1(n18853), .A2(n18870), .ZN(n18854) );
  AOI211_X1 U21831 ( .C1(n18863), .C2(n19717), .A(n18855), .B(n18854), .ZN(
        n18859) );
  AOI22_X1 U21832 ( .A1(n18857), .A2(n18856), .B1(n19715), .B2(n18873), .ZN(
        n18858) );
  OAI211_X1 U21833 ( .C1(n18877), .C2(n18860), .A(n18859), .B(n18858), .ZN(
        P2_U2854) );
  AOI22_X1 U21834 ( .A1(n18865), .A2(n18864), .B1(n18863), .B2(n18862), .ZN(
        n18869) );
  AOI22_X1 U21835 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(n18867), .B1(n18866), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n18868) );
  OAI211_X1 U21836 ( .C1(n18871), .C2(n18870), .A(n18869), .B(n18868), .ZN(
        n18872) );
  AOI21_X1 U21837 ( .B1(n19287), .B2(n18873), .A(n18872), .ZN(n18876) );
  NAND2_X1 U21838 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18874), .ZN(
        n18875) );
  OAI211_X1 U21839 ( .C1(n14020), .C2(n18877), .A(n18876), .B(n18875), .ZN(
        P2_U2855) );
  NOR2_X1 U21840 ( .A1(n9648), .A2(n18878), .ZN(n18879) );
  OR2_X1 U21841 ( .A1(n13991), .A2(n18879), .ZN(n18910) );
  OAI22_X1 U21842 ( .A1(n18910), .A2(n18893), .B1(n18888), .B2(n18880), .ZN(
        n18881) );
  INV_X1 U21843 ( .A(n18881), .ZN(n18882) );
  OAI21_X1 U21844 ( .B1(n18903), .B2(n12358), .A(n18882), .ZN(P2_U2871) );
  AOI21_X1 U21845 ( .B1(n18895), .B2(n18884), .A(n18883), .ZN(n18885) );
  NOR3_X1 U21846 ( .A1(n9704), .A2(n18885), .A3(n18893), .ZN(n18886) );
  AOI21_X1 U21847 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n18888), .A(n18886), .ZN(
        n18887) );
  OAI21_X1 U21848 ( .B1(n18889), .B2(n18888), .A(n18887), .ZN(P2_U2875) );
  AOI21_X1 U21849 ( .B1(n18892), .B2(n18891), .A(n18890), .ZN(n18894) );
  NOR3_X1 U21850 ( .A1(n18895), .A2(n18894), .A3(n18893), .ZN(n18896) );
  AOI21_X1 U21851 ( .B1(n18897), .B2(n18903), .A(n18896), .ZN(n18898) );
  OAI21_X1 U21852 ( .B1(n18903), .B2(n9959), .A(n18898), .ZN(P2_U2877) );
  AOI22_X1 U21853 ( .A1(n18900), .A2(n18899), .B1(n18903), .B2(n18984), .ZN(
        n18901) );
  OAI21_X1 U21854 ( .B1(n18903), .B2(n18902), .A(n18901), .ZN(P2_U2883) );
  AOI22_X1 U21855 ( .A1(n18908), .A2(BUF2_REG_31__SCAN_IN), .B1(n18912), .B2(
        n18904), .ZN(n18906) );
  AOI22_X1 U21856 ( .A1(n18909), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n18921), .ZN(n18905) );
  NAND2_X1 U21857 ( .A1(n18906), .A2(n18905), .ZN(P2_U2888) );
  AOI22_X1 U21858 ( .A1(n18907), .A2(n19030), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n18921), .ZN(n18916) );
  AOI22_X1 U21859 ( .A1(n18909), .A2(BUF1_REG_16__SCAN_IN), .B1(n18908), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n18915) );
  NOR2_X1 U21860 ( .A1(n18910), .A2(n18930), .ZN(n18911) );
  AOI21_X1 U21861 ( .B1(n18913), .B2(n18912), .A(n18911), .ZN(n18914) );
  NAND3_X1 U21862 ( .A1(n18916), .A2(n18915), .A3(n18914), .ZN(P2_U2903) );
  INV_X1 U21863 ( .A(n18917), .ZN(n18920) );
  INV_X1 U21864 ( .A(n18918), .ZN(n18971) );
  AOI22_X1 U21865 ( .A1(n18923), .A2(n18971), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n18921), .ZN(n18919) );
  OAI21_X1 U21866 ( .B1(n18936), .B2(n18920), .A(n18919), .ZN(P2_U2905) );
  AOI22_X1 U21867 ( .A1(n18923), .A2(n18922), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n18921), .ZN(n18924) );
  OAI21_X1 U21868 ( .B1(n18936), .B2(n18925), .A(n18924), .ZN(P2_U2909) );
  INV_X1 U21869 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18960) );
  OAI22_X1 U21870 ( .A1(n18928), .A2(n18927), .B1(n18926), .B2(n18960), .ZN(
        n18929) );
  INV_X1 U21871 ( .A(n18929), .ZN(n18934) );
  OR3_X1 U21872 ( .A1(n18932), .A2(n18931), .A3(n18930), .ZN(n18933) );
  OAI211_X1 U21873 ( .C1(n18936), .C2(n18935), .A(n18934), .B(n18933), .ZN(
        P2_U2914) );
  INV_X1 U21874 ( .A(n18967), .ZN(n18941) );
  NOR2_X1 U21875 ( .A1(n18941), .A2(n18937), .ZN(P2_U2920) );
  INV_X1 U21876 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n18940) );
  INV_X1 U21877 ( .A(n20720), .ZN(n18938) );
  AOI22_X1 U21878 ( .A1(n18938), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n20716), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n18939) );
  OAI21_X1 U21879 ( .B1(n18941), .B2(n18940), .A(n18939), .ZN(P2_U2921) );
  AOI22_X1 U21880 ( .A1(n20716), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18942) );
  OAI21_X1 U21881 ( .B1(n13237), .B2(n18969), .A(n18942), .ZN(P2_U2936) );
  INV_X1 U21882 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18944) );
  AOI22_X1 U21883 ( .A1(n20716), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18943) );
  OAI21_X1 U21884 ( .B1(n18944), .B2(n18969), .A(n18943), .ZN(P2_U2937) );
  AOI22_X1 U21885 ( .A1(n20716), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18945) );
  OAI21_X1 U21886 ( .B1(n18946), .B2(n18969), .A(n18945), .ZN(P2_U2938) );
  AOI22_X1 U21887 ( .A1(n20716), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18947) );
  OAI21_X1 U21888 ( .B1(n18948), .B2(n18969), .A(n18947), .ZN(P2_U2939) );
  AOI22_X1 U21889 ( .A1(n20716), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18949) );
  OAI21_X1 U21890 ( .B1(n18950), .B2(n18969), .A(n18949), .ZN(P2_U2940) );
  AOI22_X1 U21891 ( .A1(n20716), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18951) );
  OAI21_X1 U21892 ( .B1(n11031), .B2(n18969), .A(n18951), .ZN(P2_U2941) );
  AOI22_X1 U21893 ( .A1(n20716), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18952) );
  OAI21_X1 U21894 ( .B1(n18953), .B2(n18969), .A(n18952), .ZN(P2_U2942) );
  AOI22_X1 U21895 ( .A1(n20716), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18954) );
  OAI21_X1 U21896 ( .B1(n10999), .B2(n18969), .A(n18954), .ZN(P2_U2943) );
  AOI22_X1 U21897 ( .A1(n20716), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18955) );
  OAI21_X1 U21898 ( .B1(n18956), .B2(n18969), .A(n18955), .ZN(P2_U2944) );
  AOI22_X1 U21899 ( .A1(n20716), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18957) );
  OAI21_X1 U21900 ( .B1(n18958), .B2(n18969), .A(n18957), .ZN(P2_U2945) );
  AOI22_X1 U21901 ( .A1(n20716), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18959) );
  OAI21_X1 U21902 ( .B1(n18960), .B2(n18969), .A(n18959), .ZN(P2_U2946) );
  AOI22_X1 U21903 ( .A1(n20716), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18961) );
  OAI21_X1 U21904 ( .B1(n13783), .B2(n18969), .A(n18961), .ZN(P2_U2947) );
  AOI22_X1 U21905 ( .A1(n20716), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n18962) );
  OAI21_X1 U21906 ( .B1(n10894), .B2(n18969), .A(n18962), .ZN(P2_U2948) );
  AOI22_X1 U21907 ( .A1(n20716), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18963) );
  OAI21_X1 U21908 ( .B1(n18964), .B2(n18969), .A(n18963), .ZN(P2_U2949) );
  AOI22_X1 U21909 ( .A1(n20716), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18965) );
  OAI21_X1 U21910 ( .B1(n18966), .B2(n18969), .A(n18965), .ZN(P2_U2950) );
  AOI22_X1 U21911 ( .A1(n20716), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18967), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18968) );
  OAI21_X1 U21912 ( .B1(n10842), .B2(n18969), .A(n18968), .ZN(P2_U2951) );
  AOI22_X1 U21913 ( .A1(P2_UWORD_REG_14__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n18973) );
  NAND2_X1 U21914 ( .A1(n18972), .A2(n18971), .ZN(n18975) );
  NAND2_X1 U21915 ( .A1(n18973), .A2(n18975), .ZN(P2_U2966) );
  AOI22_X1 U21916 ( .A1(P2_LWORD_REG_14__SCAN_IN), .A2(n18970), .B1(n18974), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n18976) );
  NAND2_X1 U21917 ( .A1(n18976), .A2(n18975), .ZN(P2_U2981) );
  AOI22_X1 U21918 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18977), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n18839), .ZN(n18987) );
  INV_X1 U21919 ( .A(n18978), .ZN(n18982) );
  OAI22_X1 U21920 ( .A1(n18982), .A2(n18981), .B1(n18980), .B2(n18979), .ZN(
        n18983) );
  AOI21_X1 U21921 ( .B1(n18985), .B2(n18984), .A(n18983), .ZN(n18986) );
  OAI211_X1 U21922 ( .C1(n18989), .C2(n18988), .A(n18987), .B(n18986), .ZN(
        P2_U3010) );
  NAND3_X1 U21923 ( .A1(n18992), .A2(n18991), .A3(n18990), .ZN(n18995) );
  NAND2_X1 U21924 ( .A1(n18993), .A2(n19708), .ZN(n18994) );
  OAI211_X1 U21925 ( .C1(n18997), .C2(n18996), .A(n18995), .B(n18994), .ZN(
        n18998) );
  INV_X1 U21926 ( .A(n18998), .ZN(n19016) );
  INV_X1 U21927 ( .A(n18999), .ZN(n19014) );
  NAND2_X1 U21928 ( .A1(n19000), .A2(n19009), .ZN(n19005) );
  NAND2_X1 U21929 ( .A1(n19002), .A2(n19001), .ZN(n19003) );
  NAND3_X1 U21930 ( .A1(n19005), .A2(n19004), .A3(n19003), .ZN(n19006) );
  NAND2_X1 U21931 ( .A1(n19006), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19013) );
  NAND2_X1 U21932 ( .A1(n19008), .A2(n19007), .ZN(n19012) );
  NAND2_X1 U21933 ( .A1(n19010), .A2(n19009), .ZN(n19011) );
  AND4_X1 U21934 ( .A1(n19014), .A2(n19013), .A3(n19012), .A4(n19011), .ZN(
        n19015) );
  OAI211_X1 U21935 ( .C1(n14224), .C2(n19017), .A(n19016), .B(n19015), .ZN(
        P2_U3044) );
  INV_X1 U21936 ( .A(n19105), .ZN(n19018) );
  NAND3_X1 U21937 ( .A1(n19609), .A2(n19690), .A3(n19018), .ZN(n19019) );
  NAND2_X1 U21938 ( .A1(n19690), .A2(n19692), .ZN(n19505) );
  NAND2_X1 U21939 ( .A1(n19019), .A2(n19505), .ZN(n19031) );
  NOR3_X1 U21940 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19109), .ZN(n19032) );
  INV_X1 U21941 ( .A(n19020), .ZN(n19021) );
  AND2_X1 U21942 ( .A1(n19021), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19600) );
  NOR2_X1 U21943 ( .A1(n19032), .A2(n19600), .ZN(n19035) );
  AOI21_X1 U21944 ( .B1(n19022), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19023) );
  OAI21_X1 U21945 ( .B1(n19023), .B2(n19032), .A(n19554), .ZN(n19024) );
  AOI22_X1 U21946 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19076), .ZN(n19455) );
  OR2_X1 U21947 ( .A1(n19072), .A2(n19028), .ZN(n19443) );
  INV_X1 U21948 ( .A(n19032), .ZN(n19073) );
  OAI22_X1 U21949 ( .A1(n19609), .A2(n19455), .B1(n19443), .B2(n19073), .ZN(
        n19029) );
  INV_X1 U21950 ( .A(n19029), .ZN(n19038) );
  INV_X1 U21951 ( .A(n19031), .ZN(n19036) );
  OAI21_X1 U21952 ( .B1(n19033), .B2(n19032), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19034) );
  AOI22_X1 U21953 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19076), .ZN(n19563) );
  AOI22_X1 U21954 ( .A1(n19553), .A2(n19078), .B1(n19105), .B2(n19510), .ZN(
        n19037) );
  OAI211_X1 U21955 ( .C1(n19082), .C2(n19039), .A(n19038), .B(n19037), .ZN(
        P2_U3048) );
  AOI22_X1 U21956 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19076), .ZN(n19461) );
  OR2_X1 U21957 ( .A1(n19072), .A2(n12750), .ZN(n19456) );
  OAI22_X1 U21958 ( .A1(n19609), .A2(n19461), .B1(n19456), .B2(n19073), .ZN(
        n19040) );
  INV_X1 U21959 ( .A(n19040), .ZN(n19043) );
  AND2_X1 U21960 ( .A1(n19554), .A2(n19041), .ZN(n19565) );
  AOI22_X1 U21961 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19076), .ZN(n19569) );
  AOI22_X1 U21962 ( .A1(n19565), .A2(n19078), .B1(n19105), .B2(n19518), .ZN(
        n19042) );
  OAI211_X1 U21963 ( .C1(n19082), .C2(n19044), .A(n19043), .B(n19042), .ZN(
        P2_U3049) );
  AOI22_X1 U21964 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19076), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19077), .ZN(n19467) );
  OR2_X1 U21965 ( .A1(n19072), .A2(n19045), .ZN(n19462) );
  OAI22_X1 U21966 ( .A1(n19609), .A2(n19467), .B1(n19462), .B2(n19073), .ZN(
        n19046) );
  INV_X1 U21967 ( .A(n19046), .ZN(n19049) );
  AND2_X1 U21968 ( .A1(n19554), .A2(n19047), .ZN(n19571) );
  AOI22_X1 U21969 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19076), .ZN(n19575) );
  AOI22_X1 U21970 ( .A1(n19571), .A2(n19078), .B1(n19105), .B2(n19522), .ZN(
        n19048) );
  OAI211_X1 U21971 ( .C1(n19082), .C2(n10878), .A(n19049), .B(n19048), .ZN(
        P2_U3050) );
  INV_X1 U21972 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19054) );
  AOI22_X1 U21973 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19076), .ZN(n19473) );
  OR2_X1 U21974 ( .A1(n19072), .A2(n10623), .ZN(n19468) );
  OAI22_X1 U21975 ( .A1(n19609), .A2(n19473), .B1(n19468), .B2(n19073), .ZN(
        n19050) );
  INV_X1 U21976 ( .A(n19050), .ZN(n19053) );
  AND2_X1 U21977 ( .A1(n19554), .A2(n19051), .ZN(n19577) );
  AOI22_X1 U21978 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19076), .ZN(n19581) );
  AOI22_X1 U21979 ( .A1(n19577), .A2(n19078), .B1(n19105), .B2(n19526), .ZN(
        n19052) );
  OAI211_X1 U21980 ( .C1(n19082), .C2(n19054), .A(n19053), .B(n19052), .ZN(
        P2_U3051) );
  INV_X1 U21981 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19060) );
  AOI22_X1 U21982 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19076), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19077), .ZN(n19479) );
  OR2_X1 U21983 ( .A1(n19072), .A2(n19055), .ZN(n19474) );
  OAI22_X1 U21984 ( .A1(n19609), .A2(n19479), .B1(n19474), .B2(n19073), .ZN(
        n19056) );
  INV_X1 U21985 ( .A(n19056), .ZN(n19059) );
  AND2_X1 U21986 ( .A1(n19554), .A2(n19057), .ZN(n19583) );
  AOI22_X1 U21987 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19076), .ZN(n19587) );
  AOI22_X1 U21988 ( .A1(n19583), .A2(n19078), .B1(n19105), .B2(n19530), .ZN(
        n19058) );
  OAI211_X1 U21989 ( .C1(n19082), .C2(n19060), .A(n19059), .B(n19058), .ZN(
        P2_U3052) );
  AOI22_X1 U21990 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19076), .ZN(n19485) );
  OR2_X1 U21991 ( .A1(n19072), .A2(n19061), .ZN(n19480) );
  OAI22_X1 U21992 ( .A1(n19609), .A2(n19485), .B1(n19480), .B2(n19073), .ZN(
        n19062) );
  INV_X1 U21993 ( .A(n19062), .ZN(n19065) );
  AND2_X1 U21994 ( .A1(n19554), .A2(n19063), .ZN(n19589) );
  AOI22_X1 U21995 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19076), .ZN(n19593) );
  AOI22_X1 U21996 ( .A1(n19589), .A2(n19078), .B1(n19105), .B2(n19534), .ZN(
        n19064) );
  OAI211_X1 U21997 ( .C1(n19082), .C2(n13527), .A(n19065), .B(n19064), .ZN(
        P2_U3053) );
  AOI22_X1 U21998 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19076), .ZN(n19491) );
  OR2_X1 U21999 ( .A1(n19072), .A2(n12795), .ZN(n19486) );
  OAI22_X1 U22000 ( .A1(n19609), .A2(n19491), .B1(n19486), .B2(n19073), .ZN(
        n19066) );
  INV_X1 U22001 ( .A(n19066), .ZN(n19069) );
  AND2_X1 U22002 ( .A1(n19554), .A2(n19067), .ZN(n19595) );
  AOI22_X1 U22003 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19076), .ZN(n19599) );
  AOI22_X1 U22004 ( .A1(n19595), .A2(n19078), .B1(n19105), .B2(n19538), .ZN(
        n19068) );
  OAI211_X1 U22005 ( .C1(n19082), .C2(n19070), .A(n19069), .B(n19068), .ZN(
        P2_U3054) );
  AOI22_X1 U22006 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19076), .ZN(n19501) );
  OR2_X1 U22007 ( .A1(n19072), .A2(n19071), .ZN(n19493) );
  OAI22_X1 U22008 ( .A1(n19609), .A2(n19501), .B1(n19493), .B2(n19073), .ZN(
        n19074) );
  INV_X1 U22009 ( .A(n19074), .ZN(n19080) );
  AND2_X1 U22010 ( .A1(n19554), .A2(n19075), .ZN(n19602) );
  AOI22_X1 U22011 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19077), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19076), .ZN(n19610) );
  AOI22_X1 U22012 ( .A1(n19602), .A2(n19078), .B1(n19105), .B2(n19543), .ZN(
        n19079) );
  OAI211_X1 U22013 ( .C1(n19082), .C2(n19081), .A(n19080), .B(n19079), .ZN(
        P2_U3055) );
  OR2_X1 U22014 ( .A1(n19109), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19086) );
  INV_X1 U22015 ( .A(n19083), .ZN(n19613) );
  NOR2_X1 U22016 ( .A1(n19729), .A2(n19086), .ZN(n19103) );
  NOR3_X1 U22017 ( .A1(n19084), .A2(n19103), .A3(n19549), .ZN(n19085) );
  AOI211_X2 U22018 ( .C1(n19086), .C2(n19549), .A(n19613), .B(n19085), .ZN(
        n19104) );
  INV_X1 U22019 ( .A(n19443), .ZN(n19552) );
  AOI22_X1 U22020 ( .A1(n19104), .A2(n19553), .B1(n19552), .B2(n19103), .ZN(
        n19090) );
  AND2_X1 U22021 ( .A1(n19320), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19261) );
  NAND2_X1 U22022 ( .A1(n19261), .A2(n19321), .ZN(n19087) );
  AOI21_X1 U22023 ( .B1(n19087), .B2(n19086), .A(n19085), .ZN(n19088) );
  OAI211_X1 U22024 ( .C1(n19103), .C2(n19700), .A(n19088), .B(n19554), .ZN(
        n19106) );
  INV_X1 U22025 ( .A(n19455), .ZN(n19560) );
  AOI22_X1 U22026 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19106), .B1(
        n19105), .B2(n19560), .ZN(n19089) );
  OAI211_X1 U22027 ( .C1(n19563), .C2(n19140), .A(n19090), .B(n19089), .ZN(
        P2_U3056) );
  INV_X1 U22028 ( .A(n19456), .ZN(n19564) );
  AOI22_X1 U22029 ( .A1(n19104), .A2(n19565), .B1(n19564), .B2(n19103), .ZN(
        n19092) );
  INV_X1 U22030 ( .A(n19461), .ZN(n19566) );
  AOI22_X1 U22031 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19106), .B1(
        n19105), .B2(n19566), .ZN(n19091) );
  OAI211_X1 U22032 ( .C1(n19569), .C2(n19140), .A(n19092), .B(n19091), .ZN(
        P2_U3057) );
  INV_X1 U22033 ( .A(n19462), .ZN(n19570) );
  AOI22_X1 U22034 ( .A1(n19104), .A2(n19571), .B1(n19570), .B2(n19103), .ZN(
        n19094) );
  INV_X1 U22035 ( .A(n19467), .ZN(n19572) );
  AOI22_X1 U22036 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19106), .B1(
        n19105), .B2(n19572), .ZN(n19093) );
  OAI211_X1 U22037 ( .C1(n19575), .C2(n19140), .A(n19094), .B(n19093), .ZN(
        P2_U3058) );
  INV_X1 U22038 ( .A(n19468), .ZN(n19576) );
  AOI22_X1 U22039 ( .A1(n19104), .A2(n19577), .B1(n19576), .B2(n19103), .ZN(
        n19096) );
  INV_X1 U22040 ( .A(n19473), .ZN(n19578) );
  AOI22_X1 U22041 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19106), .B1(
        n19105), .B2(n19578), .ZN(n19095) );
  OAI211_X1 U22042 ( .C1(n19581), .C2(n19140), .A(n19096), .B(n19095), .ZN(
        P2_U3059) );
  AOI22_X1 U22043 ( .A1(n19104), .A2(n19583), .B1(n19582), .B2(n19103), .ZN(
        n19098) );
  INV_X1 U22044 ( .A(n19479), .ZN(n19584) );
  AOI22_X1 U22045 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19106), .B1(
        n19105), .B2(n19584), .ZN(n19097) );
  OAI211_X1 U22046 ( .C1(n19587), .C2(n19140), .A(n19098), .B(n19097), .ZN(
        P2_U3060) );
  INV_X1 U22047 ( .A(n19480), .ZN(n19588) );
  AOI22_X1 U22048 ( .A1(n19104), .A2(n19589), .B1(n19588), .B2(n19103), .ZN(
        n19100) );
  INV_X1 U22049 ( .A(n19485), .ZN(n19590) );
  AOI22_X1 U22050 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19106), .B1(
        n19105), .B2(n19590), .ZN(n19099) );
  OAI211_X1 U22051 ( .C1(n19593), .C2(n19140), .A(n19100), .B(n19099), .ZN(
        P2_U3061) );
  INV_X1 U22052 ( .A(n19486), .ZN(n19594) );
  AOI22_X1 U22053 ( .A1(n19104), .A2(n19595), .B1(n19594), .B2(n19103), .ZN(
        n19102) );
  INV_X1 U22054 ( .A(n19491), .ZN(n19596) );
  AOI22_X1 U22055 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19106), .B1(
        n19105), .B2(n19596), .ZN(n19101) );
  OAI211_X1 U22056 ( .C1(n19599), .C2(n19140), .A(n19102), .B(n19101), .ZN(
        P2_U3062) );
  AOI22_X1 U22057 ( .A1(n19104), .A2(n19602), .B1(n19601), .B2(n19103), .ZN(
        n19108) );
  INV_X1 U22058 ( .A(n19501), .ZN(n19604) );
  AOI22_X1 U22059 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19106), .B1(
        n19105), .B2(n19604), .ZN(n19107) );
  OAI211_X1 U22060 ( .C1(n19610), .C2(n19140), .A(n19108), .B(n19107), .ZN(
        P2_U3063) );
  NOR2_X1 U22061 ( .A1(n19719), .A2(n19109), .ZN(n19149) );
  AND2_X1 U22062 ( .A1(n19149), .A2(n19729), .ZN(n19135) );
  OAI21_X1 U22063 ( .B1(n19110), .B2(n19135), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19112) );
  NAND2_X1 U22064 ( .A1(n19111), .A2(n19142), .ZN(n19116) );
  NAND2_X1 U22065 ( .A1(n19112), .A2(n19116), .ZN(n19136) );
  AOI22_X1 U22066 ( .A1(n19136), .A2(n19553), .B1(n19552), .B2(n19135), .ZN(
        n19122) );
  INV_X1 U22067 ( .A(n19135), .ZN(n19113) );
  OAI21_X1 U22068 ( .B1(n19114), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19113), 
        .ZN(n19119) );
  INV_X1 U22069 ( .A(n19140), .ZN(n19115) );
  OAI21_X1 U22070 ( .B1(n19166), .B2(n19115), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19117) );
  NAND2_X1 U22071 ( .A1(n19117), .A2(n19116), .ZN(n19118) );
  MUX2_X1 U22072 ( .A(n19119), .B(n19118), .S(n19690), .Z(n19120) );
  NAND2_X1 U22073 ( .A1(n19120), .A2(n19554), .ZN(n19137) );
  AOI22_X1 U22074 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19137), .B1(
        n19166), .B2(n19510), .ZN(n19121) );
  OAI211_X1 U22075 ( .C1(n19455), .C2(n19140), .A(n19122), .B(n19121), .ZN(
        P2_U3064) );
  AOI22_X1 U22076 ( .A1(n19136), .A2(n19565), .B1(n19564), .B2(n19135), .ZN(
        n19124) );
  AOI22_X1 U22077 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19137), .B1(
        n19166), .B2(n19518), .ZN(n19123) );
  OAI211_X1 U22078 ( .C1(n19461), .C2(n19140), .A(n19124), .B(n19123), .ZN(
        P2_U3065) );
  AOI22_X1 U22079 ( .A1(n19136), .A2(n19571), .B1(n19570), .B2(n19135), .ZN(
        n19126) );
  AOI22_X1 U22080 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19137), .B1(
        n19166), .B2(n19522), .ZN(n19125) );
  OAI211_X1 U22081 ( .C1(n19467), .C2(n19140), .A(n19126), .B(n19125), .ZN(
        P2_U3066) );
  AOI22_X1 U22082 ( .A1(n19136), .A2(n19577), .B1(n19576), .B2(n19135), .ZN(
        n19128) );
  AOI22_X1 U22083 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19137), .B1(
        n19166), .B2(n19526), .ZN(n19127) );
  OAI211_X1 U22084 ( .C1(n19473), .C2(n19140), .A(n19128), .B(n19127), .ZN(
        P2_U3067) );
  AOI22_X1 U22085 ( .A1(n19136), .A2(n19583), .B1(n19582), .B2(n19135), .ZN(
        n19130) );
  AOI22_X1 U22086 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19137), .B1(
        n19166), .B2(n19530), .ZN(n19129) );
  OAI211_X1 U22087 ( .C1(n19479), .C2(n19140), .A(n19130), .B(n19129), .ZN(
        P2_U3068) );
  AOI22_X1 U22088 ( .A1(n19136), .A2(n19589), .B1(n19588), .B2(n19135), .ZN(
        n19132) );
  AOI22_X1 U22089 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19137), .B1(
        n19166), .B2(n19534), .ZN(n19131) );
  OAI211_X1 U22090 ( .C1(n19485), .C2(n19140), .A(n19132), .B(n19131), .ZN(
        P2_U3069) );
  AOI22_X1 U22091 ( .A1(n19136), .A2(n19595), .B1(n19594), .B2(n19135), .ZN(
        n19134) );
  AOI22_X1 U22092 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19137), .B1(
        n19166), .B2(n19538), .ZN(n19133) );
  OAI211_X1 U22093 ( .C1(n19491), .C2(n19140), .A(n19134), .B(n19133), .ZN(
        P2_U3070) );
  AOI22_X1 U22094 ( .A1(n19136), .A2(n19602), .B1(n19601), .B2(n19135), .ZN(
        n19139) );
  AOI22_X1 U22095 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19137), .B1(
        n19166), .B2(n19543), .ZN(n19138) );
  OAI211_X1 U22096 ( .C1(n19501), .C2(n19140), .A(n19139), .B(n19138), .ZN(
        P2_U3071) );
  AOI21_X1 U22097 ( .B1(n19261), .B2(n19375), .A(n19416), .ZN(n19145) );
  INV_X1 U22098 ( .A(n19141), .ZN(n19147) );
  INV_X1 U22099 ( .A(n19378), .ZN(n19143) );
  NAND2_X1 U22100 ( .A1(n19143), .A2(n19142), .ZN(n19146) );
  AOI21_X1 U22101 ( .B1(n19147), .B2(n19146), .A(n19549), .ZN(n19144) );
  INV_X1 U22102 ( .A(n19553), .ZN(n19444) );
  INV_X1 U22103 ( .A(n19146), .ZN(n19165) );
  AOI22_X1 U22104 ( .A1(n19166), .A2(n19560), .B1(n19165), .B2(n19552), .ZN(
        n19152) );
  INV_X1 U22105 ( .A(n19145), .ZN(n19150) );
  OAI211_X1 U22106 ( .C1(n19147), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19146), 
        .B(n19416), .ZN(n19148) );
  OAI211_X1 U22107 ( .C1(n19150), .C2(n19149), .A(n19554), .B(n19148), .ZN(
        n19167) );
  AOI22_X1 U22108 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19167), .B1(
        n19178), .B2(n19510), .ZN(n19151) );
  OAI211_X1 U22109 ( .C1(n19170), .C2(n19444), .A(n19152), .B(n19151), .ZN(
        P2_U3072) );
  INV_X1 U22110 ( .A(n19565), .ZN(n19457) );
  AOI22_X1 U22111 ( .A1(n19178), .A2(n19518), .B1(n19165), .B2(n19564), .ZN(
        n19154) );
  AOI22_X1 U22112 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19566), .ZN(n19153) );
  OAI211_X1 U22113 ( .C1(n19170), .C2(n19457), .A(n19154), .B(n19153), .ZN(
        P2_U3073) );
  INV_X1 U22114 ( .A(n19571), .ZN(n19463) );
  AOI22_X1 U22115 ( .A1(n19178), .A2(n19522), .B1(n19165), .B2(n19570), .ZN(
        n19156) );
  AOI22_X1 U22116 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19572), .ZN(n19155) );
  OAI211_X1 U22117 ( .C1(n19170), .C2(n19463), .A(n19156), .B(n19155), .ZN(
        P2_U3074) );
  INV_X1 U22118 ( .A(n19577), .ZN(n19469) );
  AOI22_X1 U22119 ( .A1(n19178), .A2(n19526), .B1(n19165), .B2(n19576), .ZN(
        n19158) );
  AOI22_X1 U22120 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19578), .ZN(n19157) );
  OAI211_X1 U22121 ( .C1(n19170), .C2(n19469), .A(n19158), .B(n19157), .ZN(
        P2_U3075) );
  INV_X1 U22122 ( .A(n19583), .ZN(n19475) );
  AOI22_X1 U22123 ( .A1(n19166), .A2(n19584), .B1(n19165), .B2(n19582), .ZN(
        n19160) );
  AOI22_X1 U22124 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19167), .B1(
        n19178), .B2(n19530), .ZN(n19159) );
  OAI211_X1 U22125 ( .C1(n19170), .C2(n19475), .A(n19160), .B(n19159), .ZN(
        P2_U3076) );
  INV_X1 U22126 ( .A(n19589), .ZN(n19481) );
  AOI22_X1 U22127 ( .A1(n19166), .A2(n19590), .B1(n19165), .B2(n19588), .ZN(
        n19162) );
  AOI22_X1 U22128 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19167), .B1(
        n19178), .B2(n19534), .ZN(n19161) );
  OAI211_X1 U22129 ( .C1(n19170), .C2(n19481), .A(n19162), .B(n19161), .ZN(
        P2_U3077) );
  INV_X1 U22130 ( .A(n19595), .ZN(n19487) );
  AOI22_X1 U22131 ( .A1(n19178), .A2(n19538), .B1(n19165), .B2(n19594), .ZN(
        n19164) );
  AOI22_X1 U22132 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19596), .ZN(n19163) );
  OAI211_X1 U22133 ( .C1(n19170), .C2(n19487), .A(n19164), .B(n19163), .ZN(
        P2_U3078) );
  INV_X1 U22134 ( .A(n19602), .ZN(n19494) );
  AOI22_X1 U22135 ( .A1(n19178), .A2(n19543), .B1(n19165), .B2(n19601), .ZN(
        n19169) );
  AOI22_X1 U22136 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19604), .ZN(n19168) );
  OAI211_X1 U22137 ( .C1(n19170), .C2(n19494), .A(n19169), .B(n19168), .ZN(
        P2_U3079) );
  NAND3_X1 U22138 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19704), .A3(
        n19719), .ZN(n19208) );
  NOR2_X1 U22139 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19208), .ZN(
        n19196) );
  OAI21_X1 U22140 ( .B1(n12201), .B2(n19196), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19172) );
  NAND3_X1 U22141 ( .A1(n19409), .A2(n19704), .A3(n19408), .ZN(n19171) );
  NAND2_X1 U22142 ( .A1(n19172), .A2(n19171), .ZN(n19197) );
  AOI22_X1 U22143 ( .A1(n19197), .A2(n19553), .B1(n19552), .B2(n19196), .ZN(
        n19183) );
  INV_X1 U22144 ( .A(n19196), .ZN(n19173) );
  OAI211_X1 U22145 ( .C1(n19174), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19416), 
        .B(n19173), .ZN(n19181) );
  INV_X1 U22146 ( .A(n19175), .ZN(n19176) );
  NAND2_X1 U22147 ( .A1(n19176), .A2(n19408), .ZN(n19414) );
  NOR2_X2 U22148 ( .A1(n19232), .A2(n19451), .ZN(n19222) );
  OAI21_X1 U22149 ( .B1(n19178), .B2(n19222), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19179) );
  OAI21_X1 U22150 ( .B1(n19414), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19179), .ZN(n19180) );
  NAND3_X1 U22151 ( .A1(n19181), .A2(n19554), .A3(n19180), .ZN(n19198) );
  AOI22_X1 U22152 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19198), .B1(
        n19222), .B2(n19510), .ZN(n19182) );
  OAI211_X1 U22153 ( .C1(n19455), .C2(n19201), .A(n19183), .B(n19182), .ZN(
        P2_U3080) );
  AOI22_X1 U22154 ( .A1(n19197), .A2(n19565), .B1(n19564), .B2(n19196), .ZN(
        n19185) );
  AOI22_X1 U22155 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19198), .B1(
        n19222), .B2(n19518), .ZN(n19184) );
  OAI211_X1 U22156 ( .C1(n19461), .C2(n19201), .A(n19185), .B(n19184), .ZN(
        P2_U3081) );
  AOI22_X1 U22157 ( .A1(n19197), .A2(n19571), .B1(n19570), .B2(n19196), .ZN(
        n19187) );
  AOI22_X1 U22158 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19198), .B1(
        n19222), .B2(n19522), .ZN(n19186) );
  OAI211_X1 U22159 ( .C1(n19467), .C2(n19201), .A(n19187), .B(n19186), .ZN(
        P2_U3082) );
  AOI22_X1 U22160 ( .A1(n19197), .A2(n19577), .B1(n19576), .B2(n19196), .ZN(
        n19189) );
  AOI22_X1 U22161 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19198), .B1(
        n19222), .B2(n19526), .ZN(n19188) );
  OAI211_X1 U22162 ( .C1(n19473), .C2(n19201), .A(n19189), .B(n19188), .ZN(
        P2_U3083) );
  AOI22_X1 U22163 ( .A1(n19197), .A2(n19583), .B1(n19582), .B2(n19196), .ZN(
        n19191) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19198), .B1(
        n19222), .B2(n19530), .ZN(n19190) );
  OAI211_X1 U22165 ( .C1(n19479), .C2(n19201), .A(n19191), .B(n19190), .ZN(
        P2_U3084) );
  AOI22_X1 U22166 ( .A1(n19197), .A2(n19589), .B1(n19588), .B2(n19196), .ZN(
        n19193) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19198), .B1(
        n19222), .B2(n19534), .ZN(n19192) );
  OAI211_X1 U22168 ( .C1(n19485), .C2(n19201), .A(n19193), .B(n19192), .ZN(
        P2_U3085) );
  AOI22_X1 U22169 ( .A1(n19197), .A2(n19595), .B1(n19594), .B2(n19196), .ZN(
        n19195) );
  AOI22_X1 U22170 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19198), .B1(
        n19222), .B2(n19538), .ZN(n19194) );
  OAI211_X1 U22171 ( .C1(n19491), .C2(n19201), .A(n19195), .B(n19194), .ZN(
        P2_U3086) );
  AOI22_X1 U22172 ( .A1(n19197), .A2(n19602), .B1(n19601), .B2(n19196), .ZN(
        n19200) );
  AOI22_X1 U22173 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19198), .B1(
        n19222), .B2(n19543), .ZN(n19199) );
  OAI211_X1 U22174 ( .C1(n19501), .C2(n19201), .A(n19200), .B(n19199), .ZN(
        P2_U3087) );
  INV_X1 U22175 ( .A(n19222), .ZN(n19229) );
  NOR2_X1 U22176 ( .A1(n19729), .A2(n19208), .ZN(n19230) );
  AOI22_X1 U22177 ( .A1(n19249), .A2(n19510), .B1(n19230), .B2(n19552), .ZN(
        n19211) );
  AOI21_X1 U22178 ( .B1(n19261), .B2(n19446), .A(n19416), .ZN(n19205) );
  INV_X1 U22179 ( .A(n19230), .ZN(n19203) );
  OAI21_X1 U22180 ( .B1(n19206), .B2(n19549), .A(n19700), .ZN(n19202) );
  AOI22_X1 U22181 ( .A1(n19205), .A2(n19208), .B1(n19203), .B2(n19202), .ZN(
        n19204) );
  NAND2_X1 U22182 ( .A1(n19204), .A2(n19554), .ZN(n19226) );
  INV_X1 U22183 ( .A(n19205), .ZN(n19209) );
  OAI21_X1 U22184 ( .B1(n19206), .B2(n19230), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19207) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19226), .B1(
        n19553), .B2(n19225), .ZN(n19210) );
  OAI211_X1 U22186 ( .C1(n19455), .C2(n19229), .A(n19211), .B(n19210), .ZN(
        P2_U3088) );
  AOI22_X1 U22187 ( .A1(n19249), .A2(n19518), .B1(n19230), .B2(n19564), .ZN(
        n19213) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19226), .B1(
        n19565), .B2(n19225), .ZN(n19212) );
  OAI211_X1 U22189 ( .C1(n19461), .C2(n19229), .A(n19213), .B(n19212), .ZN(
        P2_U3089) );
  AOI22_X1 U22190 ( .A1(n19222), .A2(n19572), .B1(n19570), .B2(n19230), .ZN(
        n19215) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19226), .B1(
        n19571), .B2(n19225), .ZN(n19214) );
  OAI211_X1 U22192 ( .C1(n19575), .C2(n19257), .A(n19215), .B(n19214), .ZN(
        P2_U3090) );
  AOI22_X1 U22193 ( .A1(n19222), .A2(n19578), .B1(n19230), .B2(n19576), .ZN(
        n19217) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19226), .B1(
        n19577), .B2(n19225), .ZN(n19216) );
  OAI211_X1 U22195 ( .C1(n19581), .C2(n19257), .A(n19217), .B(n19216), .ZN(
        P2_U3091) );
  AOI22_X1 U22196 ( .A1(n19249), .A2(n19530), .B1(n19230), .B2(n19582), .ZN(
        n19219) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19226), .B1(
        n19583), .B2(n19225), .ZN(n19218) );
  OAI211_X1 U22198 ( .C1(n19479), .C2(n19229), .A(n19219), .B(n19218), .ZN(
        P2_U3092) );
  AOI22_X1 U22199 ( .A1(n19249), .A2(n19534), .B1(n19230), .B2(n19588), .ZN(
        n19221) );
  AOI22_X1 U22200 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19226), .B1(
        n19589), .B2(n19225), .ZN(n19220) );
  OAI211_X1 U22201 ( .C1(n19485), .C2(n19229), .A(n19221), .B(n19220), .ZN(
        P2_U3093) );
  AOI22_X1 U22202 ( .A1(n19222), .A2(n19596), .B1(n19230), .B2(n19594), .ZN(
        n19224) );
  AOI22_X1 U22203 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19226), .B1(
        n19595), .B2(n19225), .ZN(n19223) );
  OAI211_X1 U22204 ( .C1(n19599), .C2(n19257), .A(n19224), .B(n19223), .ZN(
        P2_U3094) );
  AOI22_X1 U22205 ( .A1(n19249), .A2(n19543), .B1(n19230), .B2(n19601), .ZN(
        n19228) );
  AOI22_X1 U22206 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19226), .B1(
        n19602), .B2(n19225), .ZN(n19227) );
  OAI211_X1 U22207 ( .C1(n19501), .C2(n19229), .A(n19228), .B(n19227), .ZN(
        P2_U3095) );
  INV_X1 U22208 ( .A(n19265), .ZN(n19260) );
  NOR2_X1 U22209 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19260), .ZN(
        n19252) );
  NOR2_X1 U22210 ( .A1(n19230), .A2(n19252), .ZN(n19234) );
  OAI21_X1 U22211 ( .B1(n12205), .B2(n19252), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19231) );
  AOI22_X1 U22212 ( .A1(n19253), .A2(n19553), .B1(n19552), .B2(n19252), .ZN(
        n19238) );
  OAI21_X1 U22213 ( .B1(n19249), .B2(n19283), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19235) );
  AOI211_X1 U22214 ( .C1(n12205), .C2(n19700), .A(n19690), .B(n19252), .ZN(
        n19233) );
  AOI211_X1 U22215 ( .C1(n19235), .C2(n19234), .A(n19509), .B(n19233), .ZN(
        n19236) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19254), .B1(
        n19283), .B2(n19510), .ZN(n19237) );
  OAI211_X1 U22217 ( .C1(n19455), .C2(n19257), .A(n19238), .B(n19237), .ZN(
        P2_U3096) );
  AOI22_X1 U22218 ( .A1(n19253), .A2(n19565), .B1(n19564), .B2(n19252), .ZN(
        n19240) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19254), .B1(
        n19283), .B2(n19518), .ZN(n19239) );
  OAI211_X1 U22220 ( .C1(n19461), .C2(n19257), .A(n19240), .B(n19239), .ZN(
        P2_U3097) );
  AOI22_X1 U22221 ( .A1(n19253), .A2(n19571), .B1(n19570), .B2(n19252), .ZN(
        n19242) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19254), .B1(
        n19283), .B2(n19522), .ZN(n19241) );
  OAI211_X1 U22223 ( .C1(n19467), .C2(n19257), .A(n19242), .B(n19241), .ZN(
        P2_U3098) );
  AOI22_X1 U22224 ( .A1(n19253), .A2(n19577), .B1(n19576), .B2(n19252), .ZN(
        n19244) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19254), .B1(
        n19283), .B2(n19526), .ZN(n19243) );
  OAI211_X1 U22226 ( .C1(n19473), .C2(n19257), .A(n19244), .B(n19243), .ZN(
        P2_U3099) );
  AOI22_X1 U22227 ( .A1(n19253), .A2(n19583), .B1(n19582), .B2(n19252), .ZN(
        n19246) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19254), .B1(
        n19283), .B2(n19530), .ZN(n19245) );
  OAI211_X1 U22229 ( .C1(n19479), .C2(n19257), .A(n19246), .B(n19245), .ZN(
        P2_U3100) );
  AOI22_X1 U22230 ( .A1(n19253), .A2(n19589), .B1(n19588), .B2(n19252), .ZN(
        n19248) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19254), .B1(
        n19283), .B2(n19534), .ZN(n19247) );
  OAI211_X1 U22232 ( .C1(n19485), .C2(n19257), .A(n19248), .B(n19247), .ZN(
        P2_U3101) );
  INV_X1 U22233 ( .A(n19283), .ZN(n19273) );
  AOI22_X1 U22234 ( .A1(n19253), .A2(n19595), .B1(n19594), .B2(n19252), .ZN(
        n19251) );
  AOI22_X1 U22235 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19254), .B1(
        n19249), .B2(n19596), .ZN(n19250) );
  OAI211_X1 U22236 ( .C1(n19599), .C2(n19273), .A(n19251), .B(n19250), .ZN(
        P2_U3102) );
  AOI22_X1 U22237 ( .A1(n19253), .A2(n19602), .B1(n19601), .B2(n19252), .ZN(
        n19256) );
  AOI22_X1 U22238 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19254), .B1(
        n19283), .B2(n19543), .ZN(n19255) );
  OAI211_X1 U22239 ( .C1(n19501), .C2(n19257), .A(n19256), .B(n19255), .ZN(
        P2_U3103) );
  INV_X1 U22240 ( .A(n19290), .ZN(n19293) );
  INV_X1 U22241 ( .A(n19262), .ZN(n19259) );
  AOI211_X2 U22242 ( .C1(n19260), .C2(n19549), .A(n19613), .B(n19259), .ZN(
        n19282) );
  AOI22_X1 U22243 ( .A1(n19282), .A2(n19553), .B1(n19293), .B2(n19552), .ZN(
        n19267) );
  AND2_X1 U22244 ( .A1(n19261), .A2(n19696), .ZN(n19691) );
  OAI211_X1 U22245 ( .C1(n19293), .C2(n19700), .A(n19262), .B(n19554), .ZN(
        n19263) );
  INV_X1 U22246 ( .A(n19263), .ZN(n19264) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19560), .ZN(n19266) );
  OAI211_X1 U22248 ( .C1(n19563), .C2(n19315), .A(n19267), .B(n19266), .ZN(
        P2_U3104) );
  AOI22_X1 U22249 ( .A1(n19282), .A2(n19565), .B1(n19293), .B2(n19564), .ZN(
        n19269) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19566), .ZN(n19268) );
  OAI211_X1 U22251 ( .C1(n19569), .C2(n19315), .A(n19269), .B(n19268), .ZN(
        P2_U3105) );
  AOI22_X1 U22252 ( .A1(n19282), .A2(n19571), .B1(n19293), .B2(n19570), .ZN(
        n19272) );
  INV_X1 U22253 ( .A(n19315), .ZN(n19270) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19284), .B1(
        n19270), .B2(n19522), .ZN(n19271) );
  OAI211_X1 U22255 ( .C1(n19467), .C2(n19273), .A(n19272), .B(n19271), .ZN(
        P2_U3106) );
  AOI22_X1 U22256 ( .A1(n19282), .A2(n19577), .B1(n19293), .B2(n19576), .ZN(
        n19275) );
  AOI22_X1 U22257 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19578), .ZN(n19274) );
  OAI211_X1 U22258 ( .C1(n19581), .C2(n19315), .A(n19275), .B(n19274), .ZN(
        P2_U3107) );
  AOI22_X1 U22259 ( .A1(n19282), .A2(n19583), .B1(n19293), .B2(n19582), .ZN(
        n19277) );
  AOI22_X1 U22260 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19584), .ZN(n19276) );
  OAI211_X1 U22261 ( .C1(n19587), .C2(n19315), .A(n19277), .B(n19276), .ZN(
        P2_U3108) );
  AOI22_X1 U22262 ( .A1(n19282), .A2(n19589), .B1(n19293), .B2(n19588), .ZN(
        n19279) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19590), .ZN(n19278) );
  OAI211_X1 U22264 ( .C1(n19593), .C2(n19315), .A(n19279), .B(n19278), .ZN(
        P2_U3109) );
  AOI22_X1 U22265 ( .A1(n19282), .A2(n19595), .B1(n19293), .B2(n19594), .ZN(
        n19281) );
  AOI22_X1 U22266 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19596), .ZN(n19280) );
  OAI211_X1 U22267 ( .C1(n19599), .C2(n19315), .A(n19281), .B(n19280), .ZN(
        P2_U3110) );
  AOI22_X1 U22268 ( .A1(n19282), .A2(n19602), .B1(n19293), .B2(n19601), .ZN(
        n19286) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19604), .ZN(n19285) );
  OAI211_X1 U22270 ( .C1(n19610), .C2(n19315), .A(n19286), .B(n19285), .ZN(
        P2_U3111) );
  NAND2_X1 U22271 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19710), .ZN(
        n19383) );
  NOR3_X2 U22272 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19383), .ZN(n19310) );
  AOI22_X1 U22273 ( .A1(n19342), .A2(n19510), .B1(n19552), .B2(n19310), .ZN(
        n19297) );
  NAND2_X1 U22274 ( .A1(n19690), .A2(n19315), .ZN(n19288) );
  OAI21_X1 U22275 ( .B1(n19342), .B2(n19288), .A(n19505), .ZN(n19292) );
  OAI21_X1 U22276 ( .B1(n12232), .B2(n19549), .A(n19700), .ZN(n19289) );
  AOI21_X1 U22277 ( .B1(n19292), .B2(n19290), .A(n19289), .ZN(n19291) );
  OAI21_X1 U22278 ( .B1(n19293), .B2(n19310), .A(n19292), .ZN(n19295) );
  OAI21_X1 U22279 ( .B1(n12232), .B2(n19310), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19294) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19312), .B1(
        n19553), .B2(n19311), .ZN(n19296) );
  OAI211_X1 U22281 ( .C1(n19455), .C2(n19315), .A(n19297), .B(n19296), .ZN(
        P2_U3112) );
  AOI22_X1 U22282 ( .A1(n19342), .A2(n19518), .B1(n19564), .B2(n19310), .ZN(
        n19299) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19565), .ZN(n19298) );
  OAI211_X1 U22284 ( .C1(n19461), .C2(n19315), .A(n19299), .B(n19298), .ZN(
        P2_U3113) );
  AOI22_X1 U22285 ( .A1(n19342), .A2(n19522), .B1(n19570), .B2(n19310), .ZN(
        n19301) );
  AOI22_X1 U22286 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19571), .ZN(n19300) );
  OAI211_X1 U22287 ( .C1(n19467), .C2(n19315), .A(n19301), .B(n19300), .ZN(
        P2_U3114) );
  AOI22_X1 U22288 ( .A1(n19342), .A2(n19526), .B1(n19576), .B2(n19310), .ZN(
        n19303) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19577), .ZN(n19302) );
  OAI211_X1 U22290 ( .C1(n19473), .C2(n19315), .A(n19303), .B(n19302), .ZN(
        P2_U3115) );
  AOI22_X1 U22291 ( .A1(n19342), .A2(n19530), .B1(n19582), .B2(n19310), .ZN(
        n19305) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19583), .ZN(n19304) );
  OAI211_X1 U22293 ( .C1(n19479), .C2(n19315), .A(n19305), .B(n19304), .ZN(
        P2_U3116) );
  AOI22_X1 U22294 ( .A1(n19342), .A2(n19534), .B1(n19588), .B2(n19310), .ZN(
        n19307) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19589), .ZN(n19306) );
  OAI211_X1 U22296 ( .C1(n19485), .C2(n19315), .A(n19307), .B(n19306), .ZN(
        P2_U3117) );
  AOI22_X1 U22297 ( .A1(n19342), .A2(n19538), .B1(n19594), .B2(n19310), .ZN(
        n19309) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19595), .ZN(n19308) );
  OAI211_X1 U22299 ( .C1(n19491), .C2(n19315), .A(n19309), .B(n19308), .ZN(
        P2_U3118) );
  AOI22_X1 U22300 ( .A1(n19342), .A2(n19543), .B1(n19601), .B2(n19310), .ZN(
        n19314) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19602), .ZN(n19313) );
  OAI211_X1 U22302 ( .C1(n19501), .C2(n19315), .A(n19314), .B(n19313), .ZN(
        P2_U3119) );
  OR2_X1 U22303 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19383), .ZN(
        n19322) );
  NOR2_X1 U22304 ( .A1(n19416), .A2(n19322), .ZN(n19317) );
  NOR3_X2 U22305 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19729), .A3(
        n19383), .ZN(n19349) );
  INV_X1 U22306 ( .A(n19349), .ZN(n19318) );
  AOI21_X1 U22307 ( .B1(n19319), .B2(n19318), .A(n19549), .ZN(n19316) );
  NOR2_X1 U22308 ( .A1(n19317), .A2(n19316), .ZN(n19346) );
  AOI22_X1 U22309 ( .A1(n19342), .A2(n19560), .B1(n19552), .B2(n19349), .ZN(
        n19329) );
  OAI21_X1 U22310 ( .B1(n19319), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19318), 
        .ZN(n19325) );
  NOR2_X1 U22311 ( .A1(n19320), .A2(n19692), .ZN(n19558) );
  NAND2_X1 U22312 ( .A1(n19558), .A2(n19321), .ZN(n19323) );
  NAND2_X1 U22313 ( .A1(n19323), .A2(n19322), .ZN(n19324) );
  MUX2_X1 U22314 ( .A(n19325), .B(n19324), .S(n19690), .Z(n19326) );
  NAND2_X1 U22315 ( .A1(n19326), .A2(n19554), .ZN(n19343) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19343), .B1(
        n19350), .B2(n19510), .ZN(n19328) );
  OAI211_X1 U22317 ( .C1(n19346), .C2(n19444), .A(n19329), .B(n19328), .ZN(
        P2_U3120) );
  AOI22_X1 U22318 ( .A1(n19350), .A2(n19518), .B1(n19564), .B2(n19349), .ZN(
        n19331) );
  AOI22_X1 U22319 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19343), .B1(
        n19342), .B2(n19566), .ZN(n19330) );
  OAI211_X1 U22320 ( .C1(n19346), .C2(n19457), .A(n19331), .B(n19330), .ZN(
        P2_U3121) );
  AOI22_X1 U22321 ( .A1(n19342), .A2(n19572), .B1(n19570), .B2(n19349), .ZN(
        n19333) );
  AOI22_X1 U22322 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19343), .B1(
        n19350), .B2(n19522), .ZN(n19332) );
  OAI211_X1 U22323 ( .C1(n19346), .C2(n19463), .A(n19333), .B(n19332), .ZN(
        P2_U3122) );
  AOI22_X1 U22324 ( .A1(n19342), .A2(n19578), .B1(n19576), .B2(n19349), .ZN(
        n19335) );
  AOI22_X1 U22325 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19343), .B1(
        n19350), .B2(n19526), .ZN(n19334) );
  OAI211_X1 U22326 ( .C1(n19346), .C2(n19469), .A(n19335), .B(n19334), .ZN(
        P2_U3123) );
  AOI22_X1 U22327 ( .A1(n19350), .A2(n19530), .B1(n19582), .B2(n19349), .ZN(
        n19337) );
  AOI22_X1 U22328 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19343), .B1(
        n19342), .B2(n19584), .ZN(n19336) );
  OAI211_X1 U22329 ( .C1(n19346), .C2(n19475), .A(n19337), .B(n19336), .ZN(
        P2_U3124) );
  AOI22_X1 U22330 ( .A1(n19350), .A2(n19534), .B1(n19588), .B2(n19349), .ZN(
        n19339) );
  AOI22_X1 U22331 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19343), .B1(
        n19342), .B2(n19590), .ZN(n19338) );
  OAI211_X1 U22332 ( .C1(n19346), .C2(n19481), .A(n19339), .B(n19338), .ZN(
        P2_U3125) );
  AOI22_X1 U22333 ( .A1(n19342), .A2(n19596), .B1(n19594), .B2(n19349), .ZN(
        n19341) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19343), .B1(
        n19350), .B2(n19538), .ZN(n19340) );
  OAI211_X1 U22335 ( .C1(n19346), .C2(n19487), .A(n19341), .B(n19340), .ZN(
        P2_U3126) );
  AOI22_X1 U22336 ( .A1(n19350), .A2(n19543), .B1(n19601), .B2(n19349), .ZN(
        n19345) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19343), .B1(
        n19342), .B2(n19604), .ZN(n19344) );
  OAI211_X1 U22338 ( .C1(n19346), .C2(n19494), .A(n19345), .B(n19344), .ZN(
        P2_U3127) );
  NOR3_X2 U22339 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19719), .A3(
        n19383), .ZN(n19369) );
  OAI21_X1 U22340 ( .B1(n12231), .B2(n19369), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19347) );
  AOI22_X1 U22341 ( .A1(n19370), .A2(n19553), .B1(n19552), .B2(n19369), .ZN(
        n19356) );
  AOI221_X1 U22342 ( .B1(n19350), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19404), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19349), .ZN(n19351) );
  MUX2_X1 U22343 ( .A(n19352), .B(n19351), .S(n19549), .Z(n19353) );
  NOR2_X1 U22344 ( .A1(n19353), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19354) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19371), .B1(
        n19404), .B2(n19510), .ZN(n19355) );
  OAI211_X1 U22346 ( .C1(n19455), .C2(n19374), .A(n19356), .B(n19355), .ZN(
        P2_U3128) );
  AOI22_X1 U22347 ( .A1(n19370), .A2(n19565), .B1(n19564), .B2(n19369), .ZN(
        n19358) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19371), .B1(
        n19404), .B2(n19518), .ZN(n19357) );
  OAI211_X1 U22349 ( .C1(n19461), .C2(n19374), .A(n19358), .B(n19357), .ZN(
        P2_U3129) );
  AOI22_X1 U22350 ( .A1(n19370), .A2(n19571), .B1(n19570), .B2(n19369), .ZN(
        n19360) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19371), .B1(
        n19404), .B2(n19522), .ZN(n19359) );
  OAI211_X1 U22352 ( .C1(n19467), .C2(n19374), .A(n19360), .B(n19359), .ZN(
        P2_U3130) );
  AOI22_X1 U22353 ( .A1(n19370), .A2(n19577), .B1(n19576), .B2(n19369), .ZN(
        n19362) );
  AOI22_X1 U22354 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19371), .B1(
        n19404), .B2(n19526), .ZN(n19361) );
  OAI211_X1 U22355 ( .C1(n19473), .C2(n19374), .A(n19362), .B(n19361), .ZN(
        P2_U3131) );
  AOI22_X1 U22356 ( .A1(n19370), .A2(n19583), .B1(n19582), .B2(n19369), .ZN(
        n19364) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19371), .B1(
        n19404), .B2(n19530), .ZN(n19363) );
  OAI211_X1 U22358 ( .C1(n19479), .C2(n19374), .A(n19364), .B(n19363), .ZN(
        P2_U3132) );
  AOI22_X1 U22359 ( .A1(n19370), .A2(n19589), .B1(n19588), .B2(n19369), .ZN(
        n19366) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19371), .B1(
        n19404), .B2(n19534), .ZN(n19365) );
  OAI211_X1 U22361 ( .C1(n19485), .C2(n19374), .A(n19366), .B(n19365), .ZN(
        P2_U3133) );
  AOI22_X1 U22362 ( .A1(n19370), .A2(n19595), .B1(n19594), .B2(n19369), .ZN(
        n19368) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19371), .B1(
        n19404), .B2(n19538), .ZN(n19367) );
  OAI211_X1 U22364 ( .C1(n19491), .C2(n19374), .A(n19368), .B(n19367), .ZN(
        P2_U3134) );
  AOI22_X1 U22365 ( .A1(n19370), .A2(n19602), .B1(n19601), .B2(n19369), .ZN(
        n19373) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19371), .B1(
        n19404), .B2(n19543), .ZN(n19372) );
  OAI211_X1 U22367 ( .C1(n19501), .C2(n19374), .A(n19373), .B(n19372), .ZN(
        P2_U3135) );
  INV_X1 U22368 ( .A(n19383), .ZN(n19377) );
  NAND2_X1 U22369 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19377), .ZN(
        n19381) );
  NOR2_X1 U22370 ( .A1(n19378), .A2(n19383), .ZN(n19402) );
  OAI21_X1 U22371 ( .B1(n19379), .B2(n19402), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19380) );
  OAI21_X1 U22372 ( .B1(n19381), .B2(n19416), .A(n19380), .ZN(n19403) );
  AOI22_X1 U22373 ( .A1(n19403), .A2(n19553), .B1(n19552), .B2(n19402), .ZN(
        n19389) );
  AOI21_X1 U22374 ( .B1(n19382), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19387) );
  INV_X1 U22375 ( .A(n19558), .ZN(n19385) );
  OAI22_X1 U22376 ( .A1(n19385), .A2(n19384), .B1(n19719), .B2(n19383), .ZN(
        n19386) );
  OAI211_X1 U22377 ( .C1(n19402), .C2(n19387), .A(n19386), .B(n19554), .ZN(
        n19405) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19405), .B1(
        n19404), .B2(n19560), .ZN(n19388) );
  OAI211_X1 U22379 ( .C1(n19563), .C2(n19438), .A(n19389), .B(n19388), .ZN(
        P2_U3136) );
  AOI22_X1 U22380 ( .A1(n19403), .A2(n19565), .B1(n19564), .B2(n19402), .ZN(
        n19391) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19405), .B1(
        n19404), .B2(n19566), .ZN(n19390) );
  OAI211_X1 U22382 ( .C1(n19569), .C2(n19438), .A(n19391), .B(n19390), .ZN(
        P2_U3137) );
  AOI22_X1 U22383 ( .A1(n19403), .A2(n19571), .B1(n19570), .B2(n19402), .ZN(
        n19393) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19405), .B1(
        n19404), .B2(n19572), .ZN(n19392) );
  OAI211_X1 U22385 ( .C1(n19575), .C2(n19438), .A(n19393), .B(n19392), .ZN(
        P2_U3138) );
  AOI22_X1 U22386 ( .A1(n19403), .A2(n19577), .B1(n19576), .B2(n19402), .ZN(
        n19395) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19405), .B1(
        n19404), .B2(n19578), .ZN(n19394) );
  OAI211_X1 U22388 ( .C1(n19581), .C2(n19438), .A(n19395), .B(n19394), .ZN(
        P2_U3139) );
  AOI22_X1 U22389 ( .A1(n19403), .A2(n19583), .B1(n19582), .B2(n19402), .ZN(
        n19397) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19405), .B1(
        n19404), .B2(n19584), .ZN(n19396) );
  OAI211_X1 U22391 ( .C1(n19587), .C2(n19438), .A(n19397), .B(n19396), .ZN(
        P2_U3140) );
  AOI22_X1 U22392 ( .A1(n19403), .A2(n19589), .B1(n19588), .B2(n19402), .ZN(
        n19399) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19405), .B1(
        n19404), .B2(n19590), .ZN(n19398) );
  OAI211_X1 U22394 ( .C1(n19593), .C2(n19438), .A(n19399), .B(n19398), .ZN(
        P2_U3141) );
  AOI22_X1 U22395 ( .A1(n19403), .A2(n19595), .B1(n19594), .B2(n19402), .ZN(
        n19401) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19405), .B1(
        n19404), .B2(n19596), .ZN(n19400) );
  OAI211_X1 U22397 ( .C1(n19599), .C2(n19438), .A(n19401), .B(n19400), .ZN(
        P2_U3142) );
  AOI22_X1 U22398 ( .A1(n19403), .A2(n19602), .B1(n19601), .B2(n19402), .ZN(
        n19407) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19405), .B1(
        n19404), .B2(n19604), .ZN(n19406) );
  OAI211_X1 U22400 ( .C1(n19610), .C2(n19438), .A(n19407), .B(n19406), .ZN(
        P2_U3143) );
  NAND3_X1 U22401 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19719), .ZN(n19448) );
  NOR2_X1 U22402 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19448), .ZN(
        n19433) );
  OAI21_X1 U22403 ( .B1(n12249), .B2(n19433), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19411) );
  NAND3_X1 U22404 ( .A1(n19409), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n19408), .ZN(n19410) );
  NAND2_X1 U22405 ( .A1(n19411), .A2(n19410), .ZN(n19434) );
  AOI22_X1 U22406 ( .A1(n19434), .A2(n19553), .B1(n19552), .B2(n19433), .ZN(
        n19420) );
  INV_X1 U22407 ( .A(n19438), .ZN(n19412) );
  OAI21_X1 U22408 ( .B1(n19412), .B2(n19439), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19413) );
  OAI21_X1 U22409 ( .B1(n19704), .B2(n19414), .A(n19413), .ZN(n19418) );
  INV_X1 U22410 ( .A(n19433), .ZN(n19415) );
  OAI211_X1 U22411 ( .C1(n12250), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19416), 
        .B(n19415), .ZN(n19417) );
  NAND3_X1 U22412 ( .A1(n19418), .A2(n19554), .A3(n19417), .ZN(n19435) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19435), .B1(
        n19439), .B2(n19510), .ZN(n19419) );
  OAI211_X1 U22414 ( .C1(n19455), .C2(n19438), .A(n19420), .B(n19419), .ZN(
        P2_U3144) );
  AOI22_X1 U22415 ( .A1(n19434), .A2(n19565), .B1(n19564), .B2(n19433), .ZN(
        n19422) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19435), .B1(
        n19439), .B2(n19518), .ZN(n19421) );
  OAI211_X1 U22417 ( .C1(n19461), .C2(n19438), .A(n19422), .B(n19421), .ZN(
        P2_U3145) );
  AOI22_X1 U22418 ( .A1(n19434), .A2(n19571), .B1(n19570), .B2(n19433), .ZN(
        n19424) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19435), .B1(
        n19439), .B2(n19522), .ZN(n19423) );
  OAI211_X1 U22420 ( .C1(n19467), .C2(n19438), .A(n19424), .B(n19423), .ZN(
        P2_U3146) );
  AOI22_X1 U22421 ( .A1(n19434), .A2(n19577), .B1(n19576), .B2(n19433), .ZN(
        n19426) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19435), .B1(
        n19439), .B2(n19526), .ZN(n19425) );
  OAI211_X1 U22423 ( .C1(n19473), .C2(n19438), .A(n19426), .B(n19425), .ZN(
        P2_U3147) );
  AOI22_X1 U22424 ( .A1(n19434), .A2(n19583), .B1(n19582), .B2(n19433), .ZN(
        n19428) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19435), .B1(
        n19439), .B2(n19530), .ZN(n19427) );
  OAI211_X1 U22426 ( .C1(n19479), .C2(n19438), .A(n19428), .B(n19427), .ZN(
        P2_U3148) );
  AOI22_X1 U22427 ( .A1(n19434), .A2(n19589), .B1(n19588), .B2(n19433), .ZN(
        n19430) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19435), .B1(
        n19439), .B2(n19534), .ZN(n19429) );
  OAI211_X1 U22429 ( .C1(n19485), .C2(n19438), .A(n19430), .B(n19429), .ZN(
        P2_U3149) );
  AOI22_X1 U22430 ( .A1(n19434), .A2(n19595), .B1(n19594), .B2(n19433), .ZN(
        n19432) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19435), .B1(
        n19439), .B2(n19538), .ZN(n19431) );
  OAI211_X1 U22432 ( .C1(n19491), .C2(n19438), .A(n19432), .B(n19431), .ZN(
        P2_U3150) );
  AOI22_X1 U22433 ( .A1(n19434), .A2(n19602), .B1(n19601), .B2(n19433), .ZN(
        n19437) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19435), .B1(
        n19439), .B2(n19543), .ZN(n19436) );
  OAI211_X1 U22435 ( .C1(n19501), .C2(n19438), .A(n19437), .B(n19436), .ZN(
        P2_U3151) );
  NOR2_X1 U22436 ( .A1(n19729), .A2(n19448), .ZN(n19507) );
  INV_X1 U22437 ( .A(n19507), .ZN(n19492) );
  AND2_X1 U22438 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19492), .ZN(n19440) );
  INV_X1 U22439 ( .A(n19448), .ZN(n19441) );
  AOI21_X1 U22440 ( .B1(n19700), .B2(n19441), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19442) );
  OAI22_X1 U22441 ( .A1(n19495), .A2(n19444), .B1(n19443), .B2(n19492), .ZN(
        n19445) );
  INV_X1 U22442 ( .A(n19445), .ZN(n19454) );
  NAND2_X1 U22443 ( .A1(n19558), .A2(n19446), .ZN(n19449) );
  AOI21_X1 U22444 ( .B1(n19449), .B2(n19448), .A(n19447), .ZN(n19450) );
  OAI211_X1 U22445 ( .C1(n19507), .C2(n19700), .A(n19450), .B(n19554), .ZN(
        n19497) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19497), .B1(
        n19542), .B2(n19510), .ZN(n19453) );
  OAI211_X1 U22447 ( .C1(n19455), .C2(n19500), .A(n19454), .B(n19453), .ZN(
        P2_U3152) );
  OAI22_X1 U22448 ( .A1(n19495), .A2(n19457), .B1(n19456), .B2(n19492), .ZN(
        n19458) );
  INV_X1 U22449 ( .A(n19458), .ZN(n19460) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19497), .B1(
        n19542), .B2(n19518), .ZN(n19459) );
  OAI211_X1 U22451 ( .C1(n19461), .C2(n19500), .A(n19460), .B(n19459), .ZN(
        P2_U3153) );
  OAI22_X1 U22452 ( .A1(n19495), .A2(n19463), .B1(n19462), .B2(n19492), .ZN(
        n19464) );
  INV_X1 U22453 ( .A(n19464), .ZN(n19466) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19497), .B1(
        n19542), .B2(n19522), .ZN(n19465) );
  OAI211_X1 U22455 ( .C1(n19467), .C2(n19500), .A(n19466), .B(n19465), .ZN(
        P2_U3154) );
  OAI22_X1 U22456 ( .A1(n19495), .A2(n19469), .B1(n19468), .B2(n19492), .ZN(
        n19470) );
  INV_X1 U22457 ( .A(n19470), .ZN(n19472) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19497), .B1(
        n19542), .B2(n19526), .ZN(n19471) );
  OAI211_X1 U22459 ( .C1(n19473), .C2(n19500), .A(n19472), .B(n19471), .ZN(
        P2_U3155) );
  OAI22_X1 U22460 ( .A1(n19495), .A2(n19475), .B1(n19474), .B2(n19492), .ZN(
        n19476) );
  INV_X1 U22461 ( .A(n19476), .ZN(n19478) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19497), .B1(
        n19542), .B2(n19530), .ZN(n19477) );
  OAI211_X1 U22463 ( .C1(n19479), .C2(n19500), .A(n19478), .B(n19477), .ZN(
        P2_U3156) );
  OAI22_X1 U22464 ( .A1(n19495), .A2(n19481), .B1(n19480), .B2(n19492), .ZN(
        n19482) );
  INV_X1 U22465 ( .A(n19482), .ZN(n19484) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19497), .B1(
        n19542), .B2(n19534), .ZN(n19483) );
  OAI211_X1 U22467 ( .C1(n19485), .C2(n19500), .A(n19484), .B(n19483), .ZN(
        P2_U3157) );
  OAI22_X1 U22468 ( .A1(n19495), .A2(n19487), .B1(n19486), .B2(n19492), .ZN(
        n19488) );
  INV_X1 U22469 ( .A(n19488), .ZN(n19490) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19497), .B1(
        n19542), .B2(n19538), .ZN(n19489) );
  OAI211_X1 U22471 ( .C1(n19491), .C2(n19500), .A(n19490), .B(n19489), .ZN(
        P2_U3158) );
  OAI22_X1 U22472 ( .A1(n19495), .A2(n19494), .B1(n19493), .B2(n19492), .ZN(
        n19496) );
  INV_X1 U22473 ( .A(n19496), .ZN(n19499) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19497), .B1(
        n19542), .B2(n19543), .ZN(n19498) );
  OAI211_X1 U22475 ( .C1(n19501), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        P2_U3159) );
  INV_X1 U22476 ( .A(n19542), .ZN(n19502) );
  NAND2_X1 U22477 ( .A1(n19502), .A2(n19690), .ZN(n19506) );
  OAI21_X1 U22478 ( .B1(n19506), .B2(n19605), .A(n19505), .ZN(n19511) );
  NOR3_X2 U22479 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19704), .A3(
        n19548), .ZN(n19541) );
  NOR2_X1 U22480 ( .A1(n19541), .A2(n19507), .ZN(n19513) );
  AOI211_X1 U22481 ( .C1(n12248), .C2(n19700), .A(n19690), .B(n19541), .ZN(
        n19508) );
  AOI22_X1 U22482 ( .A1(n19605), .A2(n19510), .B1(n19552), .B2(n19541), .ZN(
        n19516) );
  INV_X1 U22483 ( .A(n19511), .ZN(n19514) );
  OAI21_X1 U22484 ( .B1(n12248), .B2(n19541), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19512) );
  AOI22_X1 U22485 ( .A1(n19553), .A2(n19544), .B1(n19542), .B2(n19560), .ZN(
        n19515) );
  OAI211_X1 U22486 ( .C1(n19547), .C2(n19517), .A(n19516), .B(n19515), .ZN(
        P2_U3160) );
  INV_X1 U22487 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n19521) );
  AOI22_X1 U22488 ( .A1(n19542), .A2(n19566), .B1(n19564), .B2(n19541), .ZN(
        n19520) );
  AOI22_X1 U22489 ( .A1(n19565), .A2(n19544), .B1(n19605), .B2(n19518), .ZN(
        n19519) );
  OAI211_X1 U22490 ( .C1(n19547), .C2(n19521), .A(n19520), .B(n19519), .ZN(
        P2_U3161) );
  INV_X1 U22491 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19525) );
  AOI22_X1 U22492 ( .A1(n19542), .A2(n19572), .B1(n19570), .B2(n19541), .ZN(
        n19524) );
  AOI22_X1 U22493 ( .A1(n19571), .A2(n19544), .B1(n19605), .B2(n19522), .ZN(
        n19523) );
  OAI211_X1 U22494 ( .C1(n19547), .C2(n19525), .A(n19524), .B(n19523), .ZN(
        P2_U3162) );
  INV_X1 U22495 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n19529) );
  AOI22_X1 U22496 ( .A1(n19542), .A2(n19578), .B1(n19576), .B2(n19541), .ZN(
        n19528) );
  AOI22_X1 U22497 ( .A1(n19577), .A2(n19544), .B1(n19605), .B2(n19526), .ZN(
        n19527) );
  OAI211_X1 U22498 ( .C1(n19547), .C2(n19529), .A(n19528), .B(n19527), .ZN(
        P2_U3163) );
  INV_X1 U22499 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19533) );
  AOI22_X1 U22500 ( .A1(n19605), .A2(n19530), .B1(n19582), .B2(n19541), .ZN(
        n19532) );
  AOI22_X1 U22501 ( .A1(n19583), .A2(n19544), .B1(n19542), .B2(n19584), .ZN(
        n19531) );
  OAI211_X1 U22502 ( .C1(n19547), .C2(n19533), .A(n19532), .B(n19531), .ZN(
        P2_U3164) );
  INV_X1 U22503 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n19537) );
  AOI22_X1 U22504 ( .A1(n19542), .A2(n19590), .B1(n19588), .B2(n19541), .ZN(
        n19536) );
  AOI22_X1 U22505 ( .A1(n19589), .A2(n19544), .B1(n19605), .B2(n19534), .ZN(
        n19535) );
  OAI211_X1 U22506 ( .C1(n19547), .C2(n19537), .A(n19536), .B(n19535), .ZN(
        P2_U3165) );
  AOI22_X1 U22507 ( .A1(n19542), .A2(n19596), .B1(n19594), .B2(n19541), .ZN(
        n19540) );
  AOI22_X1 U22508 ( .A1(n19595), .A2(n19544), .B1(n19605), .B2(n19538), .ZN(
        n19539) );
  OAI211_X1 U22509 ( .C1(n19547), .C2(n12970), .A(n19540), .B(n19539), .ZN(
        P2_U3166) );
  INV_X1 U22510 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20818) );
  AOI22_X1 U22511 ( .A1(n19542), .A2(n19604), .B1(n19601), .B2(n19541), .ZN(
        n19546) );
  AOI22_X1 U22512 ( .A1(n19602), .A2(n19544), .B1(n19605), .B2(n19543), .ZN(
        n19545) );
  OAI211_X1 U22513 ( .C1(n19547), .C2(n20818), .A(n19546), .B(n19545), .ZN(
        P2_U3167) );
  NOR2_X1 U22514 ( .A1(n19704), .A2(n19548), .ZN(n19559) );
  INV_X1 U22515 ( .A(n19559), .ZN(n19550) );
  OAI21_X1 U22516 ( .B1(n19550), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19549), 
        .ZN(n19551) );
  AOI22_X1 U22517 ( .A1(n19603), .A2(n19553), .B1(n19552), .B2(n19600), .ZN(
        n19562) );
  OAI211_X1 U22518 ( .C1(n19600), .C2(n19700), .A(n19555), .B(n19554), .ZN(
        n19556) );
  INV_X1 U22519 ( .A(n19556), .ZN(n19557) );
  OAI221_X1 U22520 ( .B1(n19559), .B2(n19696), .C1(n19559), .C2(n19558), .A(
        n19557), .ZN(n19606) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19560), .ZN(n19561) );
  OAI211_X1 U22522 ( .C1(n19563), .C2(n19609), .A(n19562), .B(n19561), .ZN(
        P2_U3168) );
  AOI22_X1 U22523 ( .A1(n19603), .A2(n19565), .B1(n19564), .B2(n19600), .ZN(
        n19568) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19566), .ZN(n19567) );
  OAI211_X1 U22525 ( .C1(n19569), .C2(n19609), .A(n19568), .B(n19567), .ZN(
        P2_U3169) );
  AOI22_X1 U22526 ( .A1(n19603), .A2(n19571), .B1(n19570), .B2(n19600), .ZN(
        n19574) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19572), .ZN(n19573) );
  OAI211_X1 U22528 ( .C1(n19575), .C2(n19609), .A(n19574), .B(n19573), .ZN(
        P2_U3170) );
  AOI22_X1 U22529 ( .A1(n19603), .A2(n19577), .B1(n19576), .B2(n19600), .ZN(
        n19580) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19578), .ZN(n19579) );
  OAI211_X1 U22531 ( .C1(n19581), .C2(n19609), .A(n19580), .B(n19579), .ZN(
        P2_U3171) );
  AOI22_X1 U22532 ( .A1(n19603), .A2(n19583), .B1(n19582), .B2(n19600), .ZN(
        n19586) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19584), .ZN(n19585) );
  OAI211_X1 U22534 ( .C1(n19587), .C2(n19609), .A(n19586), .B(n19585), .ZN(
        P2_U3172) );
  AOI22_X1 U22535 ( .A1(n19603), .A2(n19589), .B1(n19588), .B2(n19600), .ZN(
        n19592) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19590), .ZN(n19591) );
  OAI211_X1 U22537 ( .C1(n19593), .C2(n19609), .A(n19592), .B(n19591), .ZN(
        P2_U3173) );
  AOI22_X1 U22538 ( .A1(n19603), .A2(n19595), .B1(n19594), .B2(n19600), .ZN(
        n19598) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19596), .ZN(n19597) );
  OAI211_X1 U22540 ( .C1(n19599), .C2(n19609), .A(n19598), .B(n19597), .ZN(
        P2_U3174) );
  AOI22_X1 U22541 ( .A1(n19603), .A2(n19602), .B1(n19601), .B2(n19600), .ZN(
        n19608) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19604), .ZN(n19607) );
  OAI211_X1 U22543 ( .C1(n19610), .C2(n19609), .A(n19608), .B(n19607), .ZN(
        P2_U3175) );
  OR3_X1 U22544 ( .A1(n19613), .A2(n19612), .A3(n19611), .ZN(n19614) );
  OAI221_X1 U22545 ( .B1(n14021), .B2(n19616), .C1(n14021), .C2(n19615), .A(
        n19614), .ZN(P2_U3177) );
  AND2_X1 U22546 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n9598), .ZN(P2_U3179) );
  AND2_X1 U22547 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n9597), .ZN(P2_U3180) );
  AND2_X1 U22548 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n9598), .ZN(P2_U3181) );
  AND2_X1 U22549 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n9597), .ZN(P2_U3182) );
  AND2_X1 U22550 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n9598), .ZN(P2_U3183) );
  AND2_X1 U22551 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n9597), .ZN(P2_U3184) );
  AND2_X1 U22552 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n9598), .ZN(P2_U3185) );
  AND2_X1 U22553 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n9597), .ZN(P2_U3186) );
  AND2_X1 U22554 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n9597), .ZN(P2_U3187) );
  AND2_X1 U22555 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n9598), .ZN(P2_U3188) );
  AND2_X1 U22556 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n9597), .ZN(P2_U3189) );
  AND2_X1 U22557 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n9598), .ZN(P2_U3190) );
  AND2_X1 U22558 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n9597), .ZN(P2_U3191) );
  AND2_X1 U22559 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n9598), .ZN(P2_U3192) );
  AND2_X1 U22560 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n9597), .ZN(P2_U3193) );
  AND2_X1 U22561 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n9598), .ZN(P2_U3194) );
  AND2_X1 U22562 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n9597), .ZN(P2_U3195) );
  AND2_X1 U22563 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n9598), .ZN(P2_U3196) );
  AND2_X1 U22564 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n9598), .ZN(P2_U3197) );
  AND2_X1 U22565 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n9597), .ZN(P2_U3198) );
  AND2_X1 U22566 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n9598), .ZN(P2_U3199) );
  AND2_X1 U22567 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n9597), .ZN(P2_U3200) );
  AND2_X1 U22568 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n9597), .ZN(P2_U3201)
         );
  AND2_X1 U22569 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n9598), .ZN(P2_U3202)
         );
  AND2_X1 U22570 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n9597), .ZN(P2_U3203)
         );
  AND2_X1 U22571 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n9598), .ZN(P2_U3204)
         );
  AND2_X1 U22572 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n9597), .ZN(P2_U3205)
         );
  AND2_X1 U22573 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n9598), .ZN(P2_U3206)
         );
  AND2_X1 U22574 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n9597), .ZN(P2_U3207)
         );
  AND2_X1 U22575 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n9598), .ZN(P2_U3208)
         );
  OAI21_X1 U22576 ( .B1(n20592), .B2(n19623), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19633) );
  INV_X1 U22577 ( .A(n19633), .ZN(n19621) );
  NAND2_X1 U22578 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19618), .ZN(n19631) );
  INV_X1 U22579 ( .A(n19631), .ZN(n19627) );
  INV_X1 U22580 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19757) );
  NOR3_X1 U22581 ( .A1(n19627), .A2(n19757), .A3(n19622), .ZN(n19620) );
  OAI211_X1 U22582 ( .C1(HOLD), .C2(n19757), .A(n19758), .B(n19628), .ZN(
        n19619) );
  OAI21_X1 U22583 ( .B1(n19621), .B2(n19620), .A(n19619), .ZN(P2_U3209) );
  NOR2_X1 U22584 ( .A1(HOLD), .A2(n19622), .ZN(n19632) );
  AOI21_X1 U22585 ( .B1(n19634), .B2(n19623), .A(n19632), .ZN(n19625) );
  OAI22_X1 U22586 ( .A1(n19625), .A2(n19757), .B1(n20585), .B2(n19624), .ZN(
        n19626) );
  OR3_X1 U22587 ( .A1(n19752), .A2(n19627), .A3(n19626), .ZN(P2_U3210) );
  OAI22_X1 U22588 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19628), .B1(NA), 
        .B2(n19631), .ZN(n19629) );
  OAI211_X1 U22589 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19629), .ZN(n19630) );
  OAI221_X1 U22590 ( .B1(n19633), .B2(n19632), .C1(n19633), .C2(n19631), .A(
        n19630), .ZN(P2_U3211) );
  OAI222_X1 U22591 ( .A1(n19675), .A2(n19636), .B1(n19635), .B2(n19761), .C1(
        n14224), .C2(n19678), .ZN(P2_U3212) );
  OAI222_X1 U22592 ( .A1(n19675), .A2(n14224), .B1(n19637), .B2(n19761), .C1(
        n10913), .C2(n19678), .ZN(P2_U3213) );
  OAI222_X1 U22593 ( .A1(n19675), .A2(n10913), .B1(n19638), .B2(n19761), .C1(
        n10927), .C2(n19678), .ZN(P2_U3214) );
  OAI222_X1 U22594 ( .A1(n19678), .A2(n10606), .B1(n19639), .B2(n19761), .C1(
        n10927), .C2(n19675), .ZN(P2_U3215) );
  OAI222_X1 U22595 ( .A1(n19678), .A2(n19641), .B1(n19640), .B2(n19761), .C1(
        n10606), .C2(n19675), .ZN(P2_U3216) );
  OAI222_X1 U22596 ( .A1(n19678), .A2(n19643), .B1(n19642), .B2(n19761), .C1(
        n19641), .C2(n19675), .ZN(P2_U3217) );
  OAI222_X1 U22597 ( .A1(n19678), .A2(n10998), .B1(n19644), .B2(n19761), .C1(
        n19643), .C2(n19675), .ZN(P2_U3218) );
  OAI222_X1 U22598 ( .A1(n19678), .A2(n19646), .B1(n19645), .B2(n19761), .C1(
        n10998), .C2(n19675), .ZN(P2_U3219) );
  OAI222_X1 U22599 ( .A1(n19678), .A2(n11030), .B1(n19647), .B2(n19761), .C1(
        n19646), .C2(n19675), .ZN(P2_U3220) );
  OAI222_X1 U22600 ( .A1(n19678), .A2(n15369), .B1(n19648), .B2(n19761), .C1(
        n11030), .C2(n19675), .ZN(P2_U3221) );
  OAI222_X1 U22601 ( .A1(n19678), .A2(n13908), .B1(n19649), .B2(n19761), .C1(
        n15369), .C2(n19675), .ZN(P2_U3222) );
  OAI222_X1 U22602 ( .A1(n19678), .A2(n19651), .B1(n19650), .B2(n19761), .C1(
        n13908), .C2(n19675), .ZN(P2_U3223) );
  OAI222_X1 U22603 ( .A1(n19678), .A2(n11095), .B1(n19652), .B2(n19761), .C1(
        n19651), .C2(n19675), .ZN(P2_U3224) );
  OAI222_X1 U22604 ( .A1(n19678), .A2(n10711), .B1(n19653), .B2(n19761), .C1(
        n11095), .C2(n19675), .ZN(P2_U3225) );
  OAI222_X1 U22605 ( .A1(n19678), .A2(n11111), .B1(n19654), .B2(n19761), .C1(
        n10711), .C2(n19675), .ZN(P2_U3226) );
  OAI222_X1 U22606 ( .A1(n19678), .A2(n19656), .B1(n19655), .B2(n19761), .C1(
        n11111), .C2(n19675), .ZN(P2_U3227) );
  OAI222_X1 U22607 ( .A1(n19678), .A2(n10807), .B1(n19657), .B2(n19761), .C1(
        n19656), .C2(n19675), .ZN(P2_U3228) );
  OAI222_X1 U22608 ( .A1(n19678), .A2(n20834), .B1(n19658), .B2(n19761), .C1(
        n10807), .C2(n19675), .ZN(P2_U3229) );
  OAI222_X1 U22609 ( .A1(n19678), .A2(n11119), .B1(n19659), .B2(n19761), .C1(
        n20834), .C2(n19675), .ZN(P2_U3230) );
  OAI222_X1 U22610 ( .A1(n19678), .A2(n19661), .B1(n19660), .B2(n19761), .C1(
        n11119), .C2(n19675), .ZN(P2_U3231) );
  OAI222_X1 U22611 ( .A1(n19678), .A2(n19663), .B1(n19662), .B2(n19761), .C1(
        n19661), .C2(n19675), .ZN(P2_U3232) );
  OAI222_X1 U22612 ( .A1(n19678), .A2(n11125), .B1(n19664), .B2(n19761), .C1(
        n19663), .C2(n19675), .ZN(P2_U3233) );
  OAI222_X1 U22613 ( .A1(n19678), .A2(n11127), .B1(n19665), .B2(n19761), .C1(
        n11125), .C2(n19675), .ZN(P2_U3234) );
  OAI222_X1 U22614 ( .A1(n19678), .A2(n14792), .B1(n19666), .B2(n19761), .C1(
        n11127), .C2(n19675), .ZN(P2_U3235) );
  OAI222_X1 U22615 ( .A1(n19678), .A2(n15016), .B1(n19667), .B2(n19761), .C1(
        n14792), .C2(n19675), .ZN(P2_U3236) );
  OAI222_X1 U22616 ( .A1(n19678), .A2(n19670), .B1(n19668), .B2(n19761), .C1(
        n15016), .C2(n19675), .ZN(P2_U3237) );
  OAI222_X1 U22617 ( .A1(n19675), .A2(n19670), .B1(n19669), .B2(n19761), .C1(
        n19671), .C2(n19678), .ZN(P2_U3238) );
  OAI222_X1 U22618 ( .A1(n19678), .A2(n19673), .B1(n19672), .B2(n19761), .C1(
        n19671), .C2(n19675), .ZN(P2_U3239) );
  OAI222_X1 U22619 ( .A1(n19678), .A2(n19676), .B1(n19674), .B2(n19761), .C1(
        n19673), .C2(n19675), .ZN(P2_U3240) );
  INV_X1 U22620 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19677) );
  OAI222_X1 U22621 ( .A1(n19678), .A2(n19677), .B1(n20840), .B2(n19761), .C1(
        n19676), .C2(n19675), .ZN(P2_U3241) );
  INV_X1 U22622 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19679) );
  AOI22_X1 U22623 ( .A1(n19761), .A2(n19680), .B1(n19679), .B2(n19758), .ZN(
        P2_U3585) );
  MUX2_X1 U22624 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19761), .Z(P2_U3586) );
  INV_X1 U22625 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19681) );
  AOI22_X1 U22626 ( .A1(n19761), .A2(n19682), .B1(n19681), .B2(n19758), .ZN(
        P2_U3587) );
  INV_X1 U22627 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19683) );
  AOI22_X1 U22628 ( .A1(n19761), .A2(n19684), .B1(n19683), .B2(n19758), .ZN(
        P2_U3588) );
  AOI21_X1 U22629 ( .B1(n9598), .B2(n19686), .A(n19685), .ZN(P2_U3591) );
  OAI21_X1 U22630 ( .B1(n19689), .B2(n19688), .A(n19687), .ZN(P2_U3592) );
  NAND2_X1 U22631 ( .A1(n19691), .A2(n19690), .ZN(n19699) );
  NOR2_X1 U22632 ( .A1(n19693), .A2(n19692), .ZN(n19695) );
  INV_X1 U22633 ( .A(n19694), .ZN(n19723) );
  AOI21_X1 U22634 ( .B1(n19696), .B2(n19695), .A(n19723), .ZN(n19707) );
  NAND2_X1 U22635 ( .A1(n19707), .A2(n19697), .ZN(n19698) );
  OAI211_X1 U22636 ( .C1(n19701), .C2(n19700), .A(n19699), .B(n19698), .ZN(
        n19702) );
  INV_X1 U22637 ( .A(n19702), .ZN(n19703) );
  AOI22_X1 U22638 ( .A1(n19727), .A2(n19704), .B1(n19703), .B2(n19728), .ZN(
        P2_U3602) );
  OAI21_X1 U22639 ( .B1(n19712), .B2(n19714), .A(n19705), .ZN(n19706) );
  AOI22_X1 U22640 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19708), .B1(n19707), 
        .B2(n19706), .ZN(n19709) );
  AOI22_X1 U22641 ( .A1(n19727), .A2(n19710), .B1(n19709), .B2(n19728), .ZN(
        P2_U3603) );
  AND2_X1 U22642 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19711) );
  OR3_X1 U22643 ( .A1(n19712), .A2(n19723), .A3(n19711), .ZN(n19713) );
  OAI21_X1 U22644 ( .B1(n19715), .B2(n19714), .A(n19713), .ZN(n19716) );
  AOI21_X1 U22645 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19717), .A(n19716), 
        .ZN(n19718) );
  AOI22_X1 U22646 ( .A1(n19727), .A2(n19719), .B1(n19718), .B2(n19728), .ZN(
        P2_U3604) );
  INV_X1 U22647 ( .A(n19720), .ZN(n19722) );
  OAI22_X1 U22648 ( .A1(n19724), .A2(n19723), .B1(n19722), .B2(n19721), .ZN(
        n19725) );
  AOI21_X1 U22649 ( .B1(n19729), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19725), 
        .ZN(n19726) );
  OAI22_X1 U22650 ( .A1(n19729), .A2(n19728), .B1(n19727), .B2(n19726), .ZN(
        P2_U3605) );
  INV_X1 U22651 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19730) );
  AOI22_X1 U22652 ( .A1(n19761), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19730), 
        .B2(n19758), .ZN(P2_U3608) );
  INV_X1 U22653 ( .A(n19731), .ZN(n19733) );
  AOI22_X1 U22654 ( .A1(n19735), .A2(n19734), .B1(n19733), .B2(n19732), .ZN(
        n19738) );
  OAI21_X1 U22655 ( .B1(n19738), .B2(n19737), .A(n19736), .ZN(n19740) );
  MUX2_X1 U22656 ( .A(P2_MORE_REG_SCAN_IN), .B(n19740), .S(n19739), .Z(
        P2_U3609) );
  OAI21_X1 U22657 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19742), .A(n19741), 
        .ZN(n19743) );
  AOI21_X1 U22658 ( .B1(n20716), .B2(n19747), .A(n19743), .ZN(n19756) );
  INV_X1 U22659 ( .A(n19744), .ZN(n19745) );
  NOR3_X1 U22660 ( .A1(n19745), .A2(n19752), .A3(n12750), .ZN(n19749) );
  AOI21_X1 U22661 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19747), .A(n19746), 
        .ZN(n19748) );
  NOR2_X1 U22662 ( .A1(n19749), .A2(n19748), .ZN(n19755) );
  AOI211_X1 U22663 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19752), .A(n19751), 
        .B(n19750), .ZN(n19753) );
  NOR2_X1 U22664 ( .A1(n19756), .A2(n19753), .ZN(n19754) );
  AOI22_X1 U22665 ( .A1(n19757), .A2(n19756), .B1(n19755), .B2(n19754), .ZN(
        P2_U3610) );
  INV_X1 U22666 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19759) );
  AOI22_X1 U22667 ( .A1(n19761), .A2(n19760), .B1(n19759), .B2(n19758), .ZN(
        P2_U3611) );
  AOI21_X1 U22668 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20599), .A(n20598), 
        .ZN(n19768) );
  INV_X1 U22669 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19762) );
  NAND2_X1 U22670 ( .A1(n20598), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20636) );
  AOI21_X1 U22671 ( .B1(n19768), .B2(n19762), .A(n20715), .ZN(P1_U2802) );
  OAI21_X1 U22672 ( .B1(n19764), .B2(n19763), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19765) );
  OAI21_X1 U22673 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19766), .A(n19765), 
        .ZN(P1_U2803) );
  NOR2_X1 U22674 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19769) );
  OAI21_X1 U22675 ( .B1(n19769), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20712), .ZN(
        n19767) );
  OAI21_X1 U22676 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20712), .A(n19767), 
        .ZN(P1_U2804) );
  NOR2_X1 U22677 ( .A1(n20715), .A2(n19768), .ZN(n20663) );
  OAI21_X1 U22678 ( .B1(BS16), .B2(n19769), .A(n20663), .ZN(n20661) );
  OAI21_X1 U22679 ( .B1(n20663), .B2(n20771), .A(n20661), .ZN(P1_U2805) );
  OAI21_X1 U22680 ( .B1(n19771), .B2(n19770), .A(n19943), .ZN(P1_U2806) );
  NOR4_X1 U22681 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19775) );
  NOR4_X1 U22682 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19774) );
  NOR4_X1 U22683 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19773) );
  NOR4_X1 U22684 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19772) );
  NAND4_X1 U22685 ( .A1(n19775), .A2(n19774), .A3(n19773), .A4(n19772), .ZN(
        n19781) );
  NOR4_X1 U22686 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19779) );
  AOI211_X1 U22687 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19778) );
  NOR4_X1 U22688 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19777) );
  NOR4_X1 U22689 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19776) );
  NAND4_X1 U22690 ( .A1(n19779), .A2(n19778), .A3(n19777), .A4(n19776), .ZN(
        n19780) );
  NOR2_X1 U22691 ( .A1(n19781), .A2(n19780), .ZN(n20698) );
  INV_X1 U22692 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20656) );
  NOR3_X1 U22693 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19783) );
  OAI21_X1 U22694 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19783), .A(n20698), .ZN(
        n19782) );
  OAI21_X1 U22695 ( .B1(n20698), .B2(n20656), .A(n19782), .ZN(P1_U2807) );
  INV_X1 U22696 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20662) );
  AOI21_X1 U22697 ( .B1(n20600), .B2(n20662), .A(n19783), .ZN(n19784) );
  INV_X1 U22698 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20653) );
  INV_X1 U22699 ( .A(n20698), .ZN(n20695) );
  AOI22_X1 U22700 ( .A1(n20698), .A2(n19784), .B1(n20653), .B2(n20695), .ZN(
        P1_U2808) );
  NAND2_X1 U22701 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19789) );
  NOR2_X1 U22702 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19789), .ZN(n19788) );
  AOI22_X1 U22703 ( .A1(n19785), .A2(n19833), .B1(n19832), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n19786) );
  OAI211_X1 U22704 ( .C1(n19813), .C2(n11729), .A(n19786), .B(n19964), .ZN(
        n19787) );
  AOI21_X1 U22705 ( .B1(n19788), .B2(n19807), .A(n19787), .ZN(n19796) );
  INV_X1 U22706 ( .A(n19789), .ZN(n19792) );
  OAI21_X1 U22707 ( .B1(n19830), .B2(n19791), .A(n19790), .ZN(n19825) );
  OAI21_X1 U22708 ( .B1(n19793), .B2(n19792), .A(n19825), .ZN(n19801) );
  AOI22_X1 U22709 ( .A1(n19794), .A2(n19802), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n19801), .ZN(n19795) );
  OAI211_X1 U22710 ( .C1(n19797), .C2(n19818), .A(n19796), .B(n19795), .ZN(
        P1_U2833) );
  NAND2_X1 U22711 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19807), .ZN(n19799) );
  AOI22_X1 U22712 ( .A1(n19848), .A2(n19833), .B1(n19832), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n19798) );
  OAI21_X1 U22713 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n19799), .A(n19798), .ZN(
        n19800) );
  AOI211_X1 U22714 ( .C1(n19838), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19977), .B(n19800), .ZN(n19804) );
  AOI22_X1 U22715 ( .A1(n19851), .A2(n19802), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n19801), .ZN(n19803) );
  OAI211_X1 U22716 ( .C1(n19805), .C2(n19818), .A(n19804), .B(n19803), .ZN(
        P1_U2834) );
  INV_X1 U22717 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20607) );
  NOR2_X1 U22718 ( .A1(n19825), .A2(n20607), .ZN(n19815) );
  NAND2_X1 U22719 ( .A1(n19806), .A2(n19833), .ZN(n19811) );
  INV_X1 U22720 ( .A(n19807), .ZN(n19808) );
  NOR2_X1 U22721 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19808), .ZN(n19809) );
  AOI211_X1 U22722 ( .C1(n19832), .C2(P1_EBX_REG_5__SCAN_IN), .A(n19977), .B(
        n19809), .ZN(n19810) );
  OAI211_X1 U22723 ( .C1(n19813), .C2(n19812), .A(n19811), .B(n19810), .ZN(
        n19814) );
  AOI211_X1 U22724 ( .C1(n19816), .C2(n19843), .A(n19815), .B(n19814), .ZN(
        n19817) );
  OAI21_X1 U22725 ( .B1(n19819), .B2(n19818), .A(n19817), .ZN(P1_U2835) );
  AOI22_X1 U22726 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19838), .B1(
        n19833), .B2(n19949), .ZN(n19829) );
  INV_X1 U22727 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20604) );
  NAND2_X1 U22728 ( .A1(n19821), .A2(n19820), .ZN(n19824) );
  INV_X1 U22729 ( .A(n19938), .ZN(n19822) );
  AOI22_X1 U22730 ( .A1(n19837), .A2(n19822), .B1(n19832), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n19823) );
  OAI211_X1 U22731 ( .C1(n20604), .C2(n19825), .A(n19824), .B(n19823), .ZN(
        n19826) );
  AOI21_X1 U22732 ( .B1(n19933), .B2(n19843), .A(n19826), .ZN(n19828) );
  NAND4_X1 U22733 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(n19835), .A4(n20604), .ZN(n19827) );
  NAND4_X1 U22734 ( .A1(n19829), .A2(n19828), .A3(n19964), .A4(n19827), .ZN(
        P1_U2836) );
  AOI21_X1 U22735 ( .B1(n19831), .B2(n20600), .A(n19830), .ZN(n19847) );
  INV_X1 U22736 ( .A(n19965), .ZN(n19834) );
  AOI22_X1 U22737 ( .A1(n19834), .A2(n19833), .B1(n19832), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n19846) );
  AOI22_X1 U22738 ( .A1(n19837), .A2(n19836), .B1(n19835), .B2(n13514), .ZN(
        n19840) );
  NAND2_X1 U22739 ( .A1(n19838), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19839) );
  OAI211_X1 U22740 ( .C1(n20678), .C2(n19841), .A(n19840), .B(n19839), .ZN(
        n19842) );
  AOI21_X1 U22741 ( .B1(n19844), .B2(n19843), .A(n19842), .ZN(n19845) );
  OAI211_X1 U22742 ( .C1(n19847), .C2(n13514), .A(n19846), .B(n19845), .ZN(
        P1_U2838) );
  AOI22_X1 U22743 ( .A1(n19851), .A2(n19850), .B1(n19849), .B2(n19848), .ZN(
        n19852) );
  OAI21_X1 U22744 ( .B1(n19854), .B2(n19853), .A(n19852), .ZN(P1_U2866) );
  AOI22_X1 U22745 ( .A1(n20709), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19856) );
  OAI21_X1 U22746 ( .B1(n19857), .B2(n19886), .A(n19856), .ZN(P1_U2921) );
  INV_X1 U22747 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U22748 ( .A1(n20709), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19858) );
  OAI21_X1 U22749 ( .B1(n19859), .B2(n19886), .A(n19858), .ZN(P1_U2922) );
  INV_X1 U22750 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19861) );
  AOI22_X1 U22751 ( .A1(n20709), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19860) );
  OAI21_X1 U22752 ( .B1(n19861), .B2(n19886), .A(n19860), .ZN(P1_U2923) );
  AOI22_X1 U22753 ( .A1(n20709), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19862) );
  OAI21_X1 U22754 ( .B1(n14081), .B2(n19886), .A(n19862), .ZN(P1_U2924) );
  INV_X1 U22755 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U22756 ( .A1(n20709), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19863) );
  OAI21_X1 U22757 ( .B1(n19864), .B2(n19886), .A(n19863), .ZN(P1_U2925) );
  INV_X1 U22758 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U22759 ( .A1(n20709), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19865) );
  OAI21_X1 U22760 ( .B1(n19866), .B2(n19886), .A(n19865), .ZN(P1_U2926) );
  INV_X1 U22761 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U22762 ( .A1(n20709), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19867) );
  OAI21_X1 U22763 ( .B1(n19868), .B2(n19886), .A(n19867), .ZN(P1_U2927) );
  AOI22_X1 U22764 ( .A1(n20709), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19869) );
  OAI21_X1 U22765 ( .B1(n19870), .B2(n19886), .A(n19869), .ZN(P1_U2928) );
  AOI22_X1 U22766 ( .A1(n19884), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19871) );
  OAI21_X1 U22767 ( .B1(n19872), .B2(n19886), .A(n19871), .ZN(P1_U2929) );
  AOI22_X1 U22768 ( .A1(n19884), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19873) );
  OAI21_X1 U22769 ( .B1(n13847), .B2(n19886), .A(n19873), .ZN(P1_U2930) );
  AOI22_X1 U22770 ( .A1(n19884), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19874) );
  OAI21_X1 U22771 ( .B1(n11704), .B2(n19886), .A(n19874), .ZN(P1_U2931) );
  AOI22_X1 U22772 ( .A1(n19884), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19875), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19876) );
  OAI21_X1 U22773 ( .B1(n19877), .B2(n19886), .A(n19876), .ZN(P1_U2932) );
  AOI22_X1 U22774 ( .A1(n19884), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19878) );
  OAI21_X1 U22775 ( .B1(n19879), .B2(n19886), .A(n19878), .ZN(P1_U2933) );
  AOI22_X1 U22776 ( .A1(n19884), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19880) );
  OAI21_X1 U22777 ( .B1(n20850), .B2(n19886), .A(n19880), .ZN(P1_U2934) );
  AOI22_X1 U22778 ( .A1(n19884), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19881) );
  OAI21_X1 U22779 ( .B1(n19882), .B2(n19886), .A(n19881), .ZN(P1_U2935) );
  AOI22_X1 U22780 ( .A1(n19884), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19883), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19885) );
  OAI21_X1 U22781 ( .B1(n19887), .B2(n19886), .A(n19885), .ZN(P1_U2936) );
  AOI22_X1 U22782 ( .A1(n19925), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n19920), .ZN(n19889) );
  OAI21_X1 U22783 ( .B1(n20018), .B2(n19927), .A(n19889), .ZN(P1_U2937) );
  AOI22_X1 U22784 ( .A1(n19925), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n19920), .ZN(n19890) );
  OAI21_X1 U22785 ( .B1(n20026), .B2(n19927), .A(n19890), .ZN(P1_U2938) );
  AOI22_X1 U22786 ( .A1(n19925), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n19920), .ZN(n19891) );
  OAI21_X1 U22787 ( .B1(n20030), .B2(n19927), .A(n19891), .ZN(P1_U2939) );
  AOI22_X1 U22788 ( .A1(n19925), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n19920), .ZN(n19892) );
  OAI21_X1 U22789 ( .B1(n20033), .B2(n19927), .A(n19892), .ZN(P1_U2940) );
  AOI22_X1 U22790 ( .A1(n19925), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n19920), .ZN(n19893) );
  OAI21_X1 U22791 ( .B1(n20037), .B2(n19927), .A(n19893), .ZN(P1_U2941) );
  AOI22_X1 U22792 ( .A1(n19925), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n19920), .ZN(n19894) );
  OAI21_X1 U22793 ( .B1(n20041), .B2(n19927), .A(n19894), .ZN(P1_U2942) );
  AOI22_X1 U22794 ( .A1(n19925), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n19920), .ZN(n19895) );
  OAI21_X1 U22795 ( .B1(n20045), .B2(n19927), .A(n19895), .ZN(P1_U2943) );
  AOI22_X1 U22796 ( .A1(n19925), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n19920), .ZN(n19896) );
  OAI21_X1 U22797 ( .B1(n20051), .B2(n19927), .A(n19896), .ZN(P1_U2944) );
  AOI22_X1 U22798 ( .A1(n19925), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n19920), .ZN(n19897) );
  OAI21_X1 U22799 ( .B1(n20018), .B2(n19927), .A(n19897), .ZN(P1_U2952) );
  AOI22_X1 U22800 ( .A1(n19925), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n19920), .ZN(n19898) );
  OAI21_X1 U22801 ( .B1(n20026), .B2(n19927), .A(n19898), .ZN(P1_U2953) );
  AOI22_X1 U22802 ( .A1(n19925), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n19920), .ZN(n19899) );
  OAI21_X1 U22803 ( .B1(n20030), .B2(n19927), .A(n19899), .ZN(P1_U2954) );
  AOI22_X1 U22804 ( .A1(n19925), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n19920), .ZN(n19900) );
  OAI21_X1 U22805 ( .B1(n20033), .B2(n19927), .A(n19900), .ZN(P1_U2955) );
  AOI22_X1 U22806 ( .A1(n19925), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n19920), .ZN(n19901) );
  OAI21_X1 U22807 ( .B1(n20037), .B2(n19927), .A(n19901), .ZN(P1_U2956) );
  AOI22_X1 U22808 ( .A1(n19925), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n19920), .ZN(n19902) );
  OAI21_X1 U22809 ( .B1(n20041), .B2(n19927), .A(n19902), .ZN(P1_U2957) );
  AOI22_X1 U22810 ( .A1(n19925), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n19920), .ZN(n19903) );
  OAI21_X1 U22811 ( .B1(n20045), .B2(n19927), .A(n19903), .ZN(P1_U2958) );
  AOI22_X1 U22812 ( .A1(n19925), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19920), .ZN(n19904) );
  OAI21_X1 U22813 ( .B1(n20051), .B2(n19927), .A(n19904), .ZN(P1_U2959) );
  AOI22_X1 U22814 ( .A1(n19925), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n19920), .ZN(n19907) );
  NAND2_X1 U22815 ( .A1(n19922), .A2(n19905), .ZN(n19906) );
  NAND2_X1 U22816 ( .A1(n19907), .A2(n19906), .ZN(P1_U2961) );
  AOI22_X1 U22817 ( .A1(n19925), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19920), .ZN(n19910) );
  NAND2_X1 U22818 ( .A1(n19922), .A2(n19908), .ZN(n19909) );
  NAND2_X1 U22819 ( .A1(n19910), .A2(n19909), .ZN(P1_U2962) );
  AOI22_X1 U22820 ( .A1(n19925), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19920), .ZN(n19913) );
  NAND2_X1 U22821 ( .A1(n19922), .A2(n19911), .ZN(n19912) );
  NAND2_X1 U22822 ( .A1(n19913), .A2(n19912), .ZN(P1_U2963) );
  AOI22_X1 U22823 ( .A1(n19925), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19920), .ZN(n19916) );
  NAND2_X1 U22824 ( .A1(n19922), .A2(n19914), .ZN(n19915) );
  NAND2_X1 U22825 ( .A1(n19916), .A2(n19915), .ZN(P1_U2964) );
  AOI22_X1 U22826 ( .A1(n19925), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n19920), .ZN(n19919) );
  NAND2_X1 U22827 ( .A1(n19922), .A2(n19917), .ZN(n19918) );
  NAND2_X1 U22828 ( .A1(n19919), .A2(n19918), .ZN(P1_U2965) );
  AOI22_X1 U22829 ( .A1(n19925), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19920), .ZN(n19924) );
  NAND2_X1 U22830 ( .A1(n19922), .A2(n19921), .ZN(n19923) );
  NAND2_X1 U22831 ( .A1(n19924), .A2(n19923), .ZN(P1_U2966) );
  AOI22_X1 U22832 ( .A1(n19925), .A2(P1_EAX_REG_15__SCAN_IN), .B1(
        P1_LWORD_REG_15__SCAN_IN), .B2(n19920), .ZN(n19926) );
  OAI21_X1 U22833 ( .B1(n19928), .B2(n19927), .A(n19926), .ZN(P1_U2967) );
  AOI22_X1 U22834 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19937) );
  OAI21_X1 U22835 ( .B1(n19931), .B2(n19930), .A(n19929), .ZN(n19932) );
  INV_X1 U22836 ( .A(n19932), .ZN(n19950) );
  AOI22_X1 U22837 ( .A1(n19950), .A2(n19935), .B1(n19934), .B2(n19933), .ZN(
        n19936) );
  OAI211_X1 U22838 ( .C1(n19942), .C2(n19938), .A(n19937), .B(n19936), .ZN(
        P1_U2995) );
  AOI22_X1 U22839 ( .A1(n19939), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19977), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n19946) );
  OAI21_X1 U22840 ( .B1(n19941), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19940), .ZN(n19983) );
  OAI22_X1 U22841 ( .A1(n19983), .A2(n19943), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19942), .ZN(n19944) );
  INV_X1 U22842 ( .A(n19944), .ZN(n19945) );
  OAI211_X1 U22843 ( .C1(n20006), .C2(n19947), .A(n19946), .B(n19945), .ZN(
        P1_U2998) );
  OAI21_X1 U22844 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n19948), .ZN(n19953) );
  AOI22_X1 U22845 ( .A1(n19979), .A2(n19949), .B1(n19977), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n19952) );
  AOI22_X1 U22846 ( .A1(n19950), .A2(n19957), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19958), .ZN(n19951) );
  OAI211_X1 U22847 ( .C1(n19961), .C2(n19953), .A(n19952), .B(n19951), .ZN(
        P1_U3027) );
  AOI21_X1 U22848 ( .B1(n19979), .B2(n19955), .A(n19954), .ZN(n19960) );
  AOI22_X1 U22849 ( .A1(n19958), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n19957), .B2(n19956), .ZN(n19959) );
  OAI211_X1 U22850 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n19961), .A(
        n19960), .B(n19959), .ZN(P1_U3028) );
  NAND2_X1 U22851 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19963) );
  OAI21_X1 U22852 ( .B1(n19963), .B2(n9764), .A(n19962), .ZN(n19967) );
  OAI22_X1 U22853 ( .A1(n19995), .A2(n19965), .B1(n13514), .B2(n19964), .ZN(
        n19966) );
  AOI21_X1 U22854 ( .B1(n19968), .B2(n19967), .A(n19966), .ZN(n19974) );
  NOR2_X1 U22855 ( .A1(n19969), .A2(n19996), .ZN(n19972) );
  NOR3_X1 U22856 ( .A1(n19970), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        n19987), .ZN(n19971) );
  AOI21_X1 U22857 ( .B1(n19972), .B2(n13511), .A(n19971), .ZN(n19973) );
  OAI211_X1 U22858 ( .C1(n19975), .C2(n9764), .A(n19974), .B(n19973), .ZN(
        P1_U3029) );
  INV_X1 U22859 ( .A(n19976), .ZN(n19978) );
  AOI22_X1 U22860 ( .A1(n19979), .A2(n19978), .B1(n19977), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n19990) );
  NOR2_X1 U22861 ( .A1(n19992), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19980) );
  OR2_X1 U22862 ( .A1(n19981), .A2(n19980), .ZN(n19999) );
  INV_X1 U22863 ( .A(n19999), .ZN(n19982) );
  OAI22_X1 U22864 ( .A1(n19983), .A2(n19996), .B1(n19982), .B2(n19987), .ZN(
        n19984) );
  INV_X1 U22865 ( .A(n19984), .ZN(n19989) );
  NAND3_X1 U22866 ( .A1(n19987), .A2(n19986), .A3(n19985), .ZN(n19988) );
  NAND3_X1 U22867 ( .A1(n19990), .A2(n19989), .A3(n19988), .ZN(P1_U3030) );
  INV_X1 U22868 ( .A(n19991), .ZN(n19993) );
  NAND3_X1 U22869 ( .A1(n19993), .A2(n20798), .A3(n19992), .ZN(n20000) );
  OAI22_X1 U22870 ( .A1(n19997), .A2(n19996), .B1(n19995), .B2(n19994), .ZN(
        n19998) );
  AOI221_X1 U22871 ( .B1(n20001), .B2(n20000), .C1(n19999), .C2(n20000), .A(
        n19998), .ZN(n20003) );
  NAND2_X1 U22872 ( .A1(n20003), .A2(n20002), .ZN(P1_U3031) );
  NOR2_X1 U22873 ( .A1(n20004), .A2(n20688), .ZN(P1_U3032) );
  INV_X1 U22874 ( .A(n20383), .ZN(n20011) );
  AOI22_X1 U22875 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20048), .B1(DATAI_24_), 
        .B2(n20008), .ZN(n20533) );
  INV_X1 U22876 ( .A(n20533), .ZN(n20481) );
  OR2_X1 U22877 ( .A1(n20012), .A2(n20024), .ZN(n20215) );
  NAND3_X1 U22878 ( .A1(n20673), .A2(n20681), .A3(n20690), .ZN(n20058) );
  NOR2_X1 U22879 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20058), .ZN(
        n20050) );
  AOI22_X1 U22880 ( .A1(n20575), .A2(n20481), .B1(n20523), .B2(n20050), .ZN(
        n20023) );
  INV_X1 U22881 ( .A(n20019), .ZN(n20013) );
  NOR2_X1 U22882 ( .A1(n20013), .A2(n20700), .ZN(n20408) );
  NOR2_X1 U22883 ( .A1(n20059), .A2(n20408), .ZN(n20350) );
  NOR3_X1 U22884 ( .A1(n20075), .A2(n20377), .A3(n20575), .ZN(n20014) );
  NAND2_X1 U22885 ( .A1(n20771), .A2(n20519), .ZN(n20668) );
  INV_X1 U22886 ( .A(n20668), .ZN(n20683) );
  NOR2_X1 U22887 ( .A1(n20014), .A2(n20683), .ZN(n20021) );
  INV_X1 U22888 ( .A(n20021), .ZN(n20016) );
  INV_X1 U22889 ( .A(n20678), .ZN(n20015) );
  OR2_X1 U22890 ( .A1(n20666), .A2(n20015), .ZN(n20056) );
  OR2_X1 U22891 ( .A1(n20056), .A2(n20687), .ZN(n20020) );
  NAND2_X1 U22892 ( .A1(n20348), .A2(n20290), .ZN(n20160) );
  AOI22_X1 U22893 ( .A1(n20016), .A2(n20020), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20160), .ZN(n20017) );
  NOR2_X2 U22894 ( .A1(n20018), .A2(n20059), .ZN(n20524) );
  OR2_X1 U22895 ( .A1(n20019), .A2(n20700), .ZN(n20352) );
  AOI22_X1 U22896 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20053), .B1(
        n20524), .B2(n20052), .ZN(n20022) );
  OAI211_X1 U22897 ( .C1(n20484), .C2(n20084), .A(n20023), .B(n20022), .ZN(
        P1_U3033) );
  AOI22_X1 U22898 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20048), .B1(DATAI_17_), 
        .B2(n20008), .ZN(n20488) );
  AOI22_X1 U22899 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20048), .B1(DATAI_25_), 
        .B2(n20008), .ZN(n20539) );
  INV_X1 U22900 ( .A(n20539), .ZN(n20485) );
  AOI22_X1 U22901 ( .A1(n20575), .A2(n20485), .B1(n20534), .B2(n20050), .ZN(
        n20028) );
  NOR2_X2 U22902 ( .A1(n20026), .A2(n20059), .ZN(n20535) );
  AOI22_X1 U22903 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20053), .B1(
        n20535), .B2(n20052), .ZN(n20027) );
  OAI211_X1 U22904 ( .C1(n20488), .C2(n20084), .A(n20028), .B(n20027), .ZN(
        P1_U3034) );
  AOI22_X1 U22905 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20048), .B1(DATAI_26_), 
        .B2(n20008), .ZN(n20545) );
  INV_X1 U22906 ( .A(n20545), .ZN(n20489) );
  AOI22_X1 U22907 ( .A1(n20575), .A2(n20489), .B1(n20540), .B2(n20050), .ZN(
        n20032) );
  NOR2_X2 U22908 ( .A1(n20030), .A2(n20059), .ZN(n20541) );
  AOI22_X1 U22909 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20053), .B1(
        n20541), .B2(n20052), .ZN(n20031) );
  OAI211_X1 U22910 ( .C1(n20492), .C2(n20084), .A(n20032), .B(n20031), .ZN(
        P1_U3035) );
  AOI22_X1 U22911 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20048), .B1(DATAI_19_), 
        .B2(n20008), .ZN(n20496) );
  AOI22_X1 U22912 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20048), .B1(DATAI_27_), 
        .B2(n20008), .ZN(n20551) );
  INV_X1 U22913 ( .A(n20551), .ZN(n20493) );
  AOI22_X1 U22914 ( .A1(n20575), .A2(n20493), .B1(n20546), .B2(n20050), .ZN(
        n20035) );
  NOR2_X2 U22915 ( .A1(n20033), .A2(n20059), .ZN(n20547) );
  AOI22_X1 U22916 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20053), .B1(
        n20547), .B2(n20052), .ZN(n20034) );
  OAI211_X1 U22917 ( .C1(n20496), .C2(n20084), .A(n20035), .B(n20034), .ZN(
        P1_U3036) );
  AOI22_X1 U22918 ( .A1(DATAI_20_), .A2(n20008), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20048), .ZN(n20500) );
  AOI22_X1 U22919 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20048), .B1(DATAI_28_), 
        .B2(n20008), .ZN(n20557) );
  INV_X1 U22920 ( .A(n20557), .ZN(n20497) );
  AOI22_X1 U22921 ( .A1(n20575), .A2(n20497), .B1(n20552), .B2(n20050), .ZN(
        n20039) );
  NOR2_X2 U22922 ( .A1(n20037), .A2(n20059), .ZN(n20553) );
  AOI22_X1 U22923 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20053), .B1(
        n20553), .B2(n20052), .ZN(n20038) );
  OAI211_X1 U22924 ( .C1(n20500), .C2(n20084), .A(n20039), .B(n20038), .ZN(
        P1_U3037) );
  AOI22_X1 U22925 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20048), .B1(DATAI_29_), 
        .B2(n20008), .ZN(n20563) );
  INV_X1 U22926 ( .A(n20563), .ZN(n20501) );
  AOI22_X1 U22927 ( .A1(n20575), .A2(n20501), .B1(n20558), .B2(n20050), .ZN(
        n20043) );
  NOR2_X2 U22928 ( .A1(n20041), .A2(n20059), .ZN(n20559) );
  AOI22_X1 U22929 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20053), .B1(
        n20559), .B2(n20052), .ZN(n20042) );
  OAI211_X1 U22930 ( .C1(n20504), .C2(n20084), .A(n20043), .B(n20042), .ZN(
        P1_U3038) );
  AOI22_X1 U22931 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20048), .B1(DATAI_30_), 
        .B2(n20008), .ZN(n20569) );
  INV_X1 U22932 ( .A(n20569), .ZN(n20505) );
  AOI22_X1 U22933 ( .A1(n20575), .A2(n20505), .B1(n20564), .B2(n20050), .ZN(
        n20047) );
  NOR2_X2 U22934 ( .A1(n20045), .A2(n20059), .ZN(n20565) );
  AOI22_X1 U22935 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20053), .B1(
        n20565), .B2(n20052), .ZN(n20046) );
  OAI211_X1 U22936 ( .C1(n20508), .C2(n20084), .A(n20047), .B(n20046), .ZN(
        P1_U3039) );
  AOI22_X1 U22937 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20048), .B1(DATAI_23_), 
        .B2(n20008), .ZN(n20516) );
  AOI22_X1 U22938 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20048), .B1(DATAI_31_), 
        .B2(n20008), .ZN(n20580) );
  INV_X1 U22939 ( .A(n20580), .ZN(n20511) );
  AOI22_X1 U22940 ( .A1(n20575), .A2(n20511), .B1(n20571), .B2(n20050), .ZN(
        n20055) );
  NOR2_X2 U22941 ( .A1(n20051), .A2(n20059), .ZN(n20573) );
  AOI22_X1 U22942 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20053), .B1(
        n20573), .B2(n20052), .ZN(n20054) );
  OAI211_X1 U22943 ( .C1(n20516), .C2(n20084), .A(n20055), .B(n20054), .ZN(
        P1_U3040) );
  INV_X1 U22944 ( .A(n20056), .ZN(n20123) );
  INV_X1 U22945 ( .A(n20057), .ZN(n20187) );
  NOR2_X1 U22946 ( .A1(n20446), .A2(n20058), .ZN(n20078) );
  AOI21_X1 U22947 ( .B1(n20123), .B2(n20187), .A(n20078), .ZN(n20060) );
  OAI22_X1 U22948 ( .A1(n20060), .A2(n20377), .B1(n20058), .B2(n20700), .ZN(
        n20079) );
  AOI22_X1 U22949 ( .A1(n20524), .A2(n20079), .B1(n20523), .B2(n20078), .ZN(
        n20064) );
  INV_X1 U22950 ( .A(n20058), .ZN(n20062) );
  INV_X1 U22951 ( .A(n20118), .ZN(n20125) );
  OAI211_X1 U22952 ( .C1(n20125), .C2(n20771), .A(n20060), .B(n20519), .ZN(
        n20061) );
  OAI211_X1 U22953 ( .C1(n20519), .C2(n20062), .A(n20527), .B(n20061), .ZN(
        n20081) );
  AOI22_X1 U22954 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20081), .B1(
        n20075), .B2(n20481), .ZN(n20063) );
  OAI211_X1 U22955 ( .C1(n20484), .C2(n20117), .A(n20064), .B(n20063), .ZN(
        P1_U3041) );
  AOI22_X1 U22956 ( .A1(n20535), .A2(n20079), .B1(n20534), .B2(n20078), .ZN(
        n20066) );
  INV_X1 U22957 ( .A(n20117), .ZN(n20080) );
  INV_X1 U22958 ( .A(n20488), .ZN(n20536) );
  AOI22_X1 U22959 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20081), .B1(
        n20080), .B2(n20536), .ZN(n20065) );
  OAI211_X1 U22960 ( .C1(n20539), .C2(n20084), .A(n20066), .B(n20065), .ZN(
        P1_U3042) );
  AOI22_X1 U22961 ( .A1(n20541), .A2(n20079), .B1(n20540), .B2(n20078), .ZN(
        n20068) );
  AOI22_X1 U22962 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20081), .B1(
        n20075), .B2(n20489), .ZN(n20067) );
  OAI211_X1 U22963 ( .C1(n20492), .C2(n20117), .A(n20068), .B(n20067), .ZN(
        P1_U3043) );
  AOI22_X1 U22964 ( .A1(n20547), .A2(n20079), .B1(n20546), .B2(n20078), .ZN(
        n20070) );
  AOI22_X1 U22965 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20081), .B1(
        n20075), .B2(n20493), .ZN(n20069) );
  OAI211_X1 U22966 ( .C1(n20496), .C2(n20117), .A(n20070), .B(n20069), .ZN(
        P1_U3044) );
  AOI22_X1 U22967 ( .A1(n20553), .A2(n20079), .B1(n20552), .B2(n20078), .ZN(
        n20072) );
  AOI22_X1 U22968 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20081), .B1(
        n20075), .B2(n20497), .ZN(n20071) );
  OAI211_X1 U22969 ( .C1(n20500), .C2(n20117), .A(n20072), .B(n20071), .ZN(
        P1_U3045) );
  AOI22_X1 U22970 ( .A1(n20559), .A2(n20079), .B1(n20558), .B2(n20078), .ZN(
        n20074) );
  AOI22_X1 U22971 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20081), .B1(
        n20075), .B2(n20501), .ZN(n20073) );
  OAI211_X1 U22972 ( .C1(n20504), .C2(n20117), .A(n20074), .B(n20073), .ZN(
        P1_U3046) );
  AOI22_X1 U22973 ( .A1(n20565), .A2(n20079), .B1(n20564), .B2(n20078), .ZN(
        n20077) );
  AOI22_X1 U22974 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20081), .B1(
        n20075), .B2(n20505), .ZN(n20076) );
  OAI211_X1 U22975 ( .C1(n20508), .C2(n20117), .A(n20077), .B(n20076), .ZN(
        P1_U3047) );
  AOI22_X1 U22976 ( .A1(n20573), .A2(n20079), .B1(n20571), .B2(n20078), .ZN(
        n20083) );
  INV_X1 U22977 ( .A(n20516), .ZN(n20574) );
  AOI22_X1 U22978 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20081), .B1(
        n20080), .B2(n20574), .ZN(n20082) );
  OAI211_X1 U22979 ( .C1(n20580), .C2(n20084), .A(n20083), .B(n20082), .ZN(
        P1_U3048) );
  NAND3_X1 U22980 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20673), .A3(
        n20681), .ZN(n20128) );
  OR2_X1 U22981 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20128), .ZN(
        n20111) );
  OAI22_X1 U22982 ( .A1(n20117), .A2(n20533), .B1(n20111), .B2(n20215), .ZN(
        n20085) );
  INV_X1 U22983 ( .A(n20085), .ZN(n20092) );
  NAND2_X1 U22984 ( .A1(n20152), .A2(n20117), .ZN(n20086) );
  AOI21_X1 U22985 ( .B1(n20086), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20377), 
        .ZN(n20088) );
  NAND2_X1 U22986 ( .A1(n20123), .A2(n20687), .ZN(n20089) );
  AOI22_X1 U22987 ( .A1(n20088), .A2(n20089), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20111), .ZN(n20087) );
  OAI21_X1 U22988 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20348), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20219) );
  NAND3_X1 U22989 ( .A1(n20350), .A2(n20087), .A3(n20219), .ZN(n20114) );
  INV_X1 U22990 ( .A(n20088), .ZN(n20090) );
  INV_X1 U22991 ( .A(n20348), .ZN(n20291) );
  NAND2_X1 U22992 ( .A1(n20291), .A2(n20673), .ZN(n20222) );
  OAI22_X1 U22993 ( .A1(n20090), .A2(n20089), .B1(n20222), .B2(n20352), .ZN(
        n20113) );
  AOI22_X1 U22994 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20114), .B1(
        n20524), .B2(n20113), .ZN(n20091) );
  OAI211_X1 U22995 ( .C1(n20484), .C2(n20152), .A(n20092), .B(n20091), .ZN(
        P1_U3049) );
  INV_X1 U22996 ( .A(n20534), .ZN(n20227) );
  OAI22_X1 U22997 ( .A1(n20152), .A2(n20488), .B1(n20227), .B2(n20111), .ZN(
        n20093) );
  INV_X1 U22998 ( .A(n20093), .ZN(n20095) );
  AOI22_X1 U22999 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20114), .B1(
        n20535), .B2(n20113), .ZN(n20094) );
  OAI211_X1 U23000 ( .C1(n20539), .C2(n20117), .A(n20095), .B(n20094), .ZN(
        P1_U3050) );
  INV_X1 U23001 ( .A(n20540), .ZN(n20231) );
  OAI22_X1 U23002 ( .A1(n20117), .A2(n20545), .B1(n20111), .B2(n20231), .ZN(
        n20096) );
  INV_X1 U23003 ( .A(n20096), .ZN(n20098) );
  AOI22_X1 U23004 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20114), .B1(
        n20541), .B2(n20113), .ZN(n20097) );
  OAI211_X1 U23005 ( .C1(n20492), .C2(n20152), .A(n20098), .B(n20097), .ZN(
        P1_U3051) );
  INV_X1 U23006 ( .A(n20546), .ZN(n20235) );
  OAI22_X1 U23007 ( .A1(n20152), .A2(n20496), .B1(n20111), .B2(n20235), .ZN(
        n20099) );
  INV_X1 U23008 ( .A(n20099), .ZN(n20101) );
  AOI22_X1 U23009 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20114), .B1(
        n20547), .B2(n20113), .ZN(n20100) );
  OAI211_X1 U23010 ( .C1(n20551), .C2(n20117), .A(n20101), .B(n20100), .ZN(
        P1_U3052) );
  INV_X1 U23011 ( .A(n20552), .ZN(n20239) );
  OAI22_X1 U23012 ( .A1(n20152), .A2(n20500), .B1(n20111), .B2(n20239), .ZN(
        n20102) );
  INV_X1 U23013 ( .A(n20102), .ZN(n20104) );
  AOI22_X1 U23014 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20114), .B1(
        n20553), .B2(n20113), .ZN(n20103) );
  OAI211_X1 U23015 ( .C1(n20557), .C2(n20117), .A(n20104), .B(n20103), .ZN(
        P1_U3053) );
  INV_X1 U23016 ( .A(n20558), .ZN(n20243) );
  OAI22_X1 U23017 ( .A1(n20152), .A2(n20504), .B1(n20111), .B2(n20243), .ZN(
        n20105) );
  INV_X1 U23018 ( .A(n20105), .ZN(n20107) );
  AOI22_X1 U23019 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20114), .B1(
        n20559), .B2(n20113), .ZN(n20106) );
  OAI211_X1 U23020 ( .C1(n20563), .C2(n20117), .A(n20107), .B(n20106), .ZN(
        P1_U3054) );
  INV_X1 U23021 ( .A(n20564), .ZN(n20247) );
  OAI22_X1 U23022 ( .A1(n20117), .A2(n20569), .B1(n20111), .B2(n20247), .ZN(
        n20108) );
  INV_X1 U23023 ( .A(n20108), .ZN(n20110) );
  AOI22_X1 U23024 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20114), .B1(
        n20565), .B2(n20113), .ZN(n20109) );
  OAI211_X1 U23025 ( .C1(n20508), .C2(n20152), .A(n20110), .B(n20109), .ZN(
        P1_U3055) );
  INV_X1 U23026 ( .A(n20571), .ZN(n20252) );
  OAI22_X1 U23027 ( .A1(n20152), .A2(n20516), .B1(n20111), .B2(n20252), .ZN(
        n20112) );
  INV_X1 U23028 ( .A(n20112), .ZN(n20116) );
  AOI22_X1 U23029 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20114), .B1(
        n20573), .B2(n20113), .ZN(n20115) );
  OAI211_X1 U23030 ( .C1(n20580), .C2(n20117), .A(n20116), .B(n20115), .ZN(
        P1_U3056) );
  OR2_X1 U23031 ( .A1(n20375), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20151) );
  OAI22_X1 U23032 ( .A1(n20152), .A2(n20533), .B1(n20215), .B2(n20151), .ZN(
        n20119) );
  INV_X1 U23033 ( .A(n20119), .ZN(n20132) );
  NOR2_X1 U23034 ( .A1(n20121), .A2(n20120), .ZN(n20517) );
  INV_X1 U23035 ( .A(n20151), .ZN(n20122) );
  AOI21_X1 U23036 ( .B1(n20123), .B2(n20517), .A(n20122), .ZN(n20129) );
  NAND2_X1 U23037 ( .A1(n20010), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20124) );
  AND2_X1 U23038 ( .A1(n20124), .A2(n20519), .ZN(n20675) );
  AOI21_X1 U23039 ( .B1(n20125), .B2(n20519), .A(n20675), .ZN(n20130) );
  INV_X1 U23040 ( .A(n20130), .ZN(n20126) );
  AOI22_X1 U23041 ( .A1(n20129), .A2(n20126), .B1(n20377), .B2(n20128), .ZN(
        n20127) );
  NAND2_X1 U23042 ( .A1(n20527), .A2(n20127), .ZN(n20155) );
  OAI22_X1 U23043 ( .A1(n20130), .A2(n20129), .B1(n20700), .B2(n20128), .ZN(
        n20154) );
  AOI22_X1 U23044 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20155), .B1(
        n20524), .B2(n20154), .ZN(n20131) );
  OAI211_X1 U23045 ( .C1(n20484), .C2(n20186), .A(n20132), .B(n20131), .ZN(
        P1_U3057) );
  OAI22_X1 U23046 ( .A1(n20186), .A2(n20488), .B1(n20227), .B2(n20151), .ZN(
        n20133) );
  INV_X1 U23047 ( .A(n20133), .ZN(n20135) );
  AOI22_X1 U23048 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20155), .B1(
        n20535), .B2(n20154), .ZN(n20134) );
  OAI211_X1 U23049 ( .C1(n20539), .C2(n20152), .A(n20135), .B(n20134), .ZN(
        P1_U3058) );
  OAI22_X1 U23050 ( .A1(n20152), .A2(n20545), .B1(n20151), .B2(n20231), .ZN(
        n20136) );
  INV_X1 U23051 ( .A(n20136), .ZN(n20138) );
  AOI22_X1 U23052 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20155), .B1(
        n20541), .B2(n20154), .ZN(n20137) );
  OAI211_X1 U23053 ( .C1(n20492), .C2(n20186), .A(n20138), .B(n20137), .ZN(
        P1_U3059) );
  OAI22_X1 U23054 ( .A1(n20152), .A2(n20551), .B1(n20235), .B2(n20151), .ZN(
        n20139) );
  INV_X1 U23055 ( .A(n20139), .ZN(n20141) );
  AOI22_X1 U23056 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20155), .B1(
        n20547), .B2(n20154), .ZN(n20140) );
  OAI211_X1 U23057 ( .C1(n20496), .C2(n20186), .A(n20141), .B(n20140), .ZN(
        P1_U3060) );
  OAI22_X1 U23058 ( .A1(n20186), .A2(n20500), .B1(n20239), .B2(n20151), .ZN(
        n20142) );
  INV_X1 U23059 ( .A(n20142), .ZN(n20144) );
  AOI22_X1 U23060 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20155), .B1(
        n20553), .B2(n20154), .ZN(n20143) );
  OAI211_X1 U23061 ( .C1(n20557), .C2(n20152), .A(n20144), .B(n20143), .ZN(
        P1_U3061) );
  OAI22_X1 U23062 ( .A1(n20186), .A2(n20504), .B1(n20243), .B2(n20151), .ZN(
        n20145) );
  INV_X1 U23063 ( .A(n20145), .ZN(n20147) );
  AOI22_X1 U23064 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20155), .B1(
        n20559), .B2(n20154), .ZN(n20146) );
  OAI211_X1 U23065 ( .C1(n20563), .C2(n20152), .A(n20147), .B(n20146), .ZN(
        P1_U3062) );
  OAI22_X1 U23066 ( .A1(n20152), .A2(n20569), .B1(n20151), .B2(n20247), .ZN(
        n20148) );
  INV_X1 U23067 ( .A(n20148), .ZN(n20150) );
  AOI22_X1 U23068 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20155), .B1(
        n20565), .B2(n20154), .ZN(n20149) );
  OAI211_X1 U23069 ( .C1(n20508), .C2(n20186), .A(n20150), .B(n20149), .ZN(
        P1_U3063) );
  OAI22_X1 U23070 ( .A1(n20152), .A2(n20580), .B1(n20252), .B2(n20151), .ZN(
        n20153) );
  INV_X1 U23071 ( .A(n20153), .ZN(n20157) );
  AOI22_X1 U23072 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20155), .B1(
        n20573), .B2(n20154), .ZN(n20156) );
  OAI211_X1 U23073 ( .C1(n20516), .C2(n20186), .A(n20157), .B(n20156), .ZN(
        P1_U3064) );
  OR2_X1 U23074 ( .A1(n20678), .A2(n20159), .ZN(n20218) );
  NAND2_X1 U23075 ( .A1(n13829), .A2(n20519), .ZN(n20161) );
  INV_X1 U23076 ( .A(n20408), .ZN(n20471) );
  OAI22_X1 U23077 ( .A1(n20218), .A2(n20161), .B1(n20471), .B2(n20160), .ZN(
        n20182) );
  NAND3_X1 U23078 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20673), .A3(
        n20690), .ZN(n20188) );
  NOR2_X1 U23079 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20188), .ZN(
        n20181) );
  AOI22_X1 U23080 ( .A1(n20524), .A2(n20182), .B1(n20523), .B2(n20181), .ZN(
        n20167) );
  INV_X1 U23081 ( .A(n20218), .ZN(n20260) );
  AOI21_X1 U23082 ( .B1(n20186), .B2(n20203), .A(n20771), .ZN(n20162) );
  AOI21_X1 U23083 ( .B1(n20260), .B2(n13829), .A(n20162), .ZN(n20163) );
  NOR2_X1 U23084 ( .A1(n20163), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20165) );
  INV_X1 U23085 ( .A(n20186), .ZN(n20178) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20183), .B1(
        n20178), .B2(n20481), .ZN(n20166) );
  OAI211_X1 U23087 ( .C1(n20484), .C2(n20203), .A(n20167), .B(n20166), .ZN(
        P1_U3065) );
  AOI22_X1 U23088 ( .A1(n20535), .A2(n20182), .B1(n20534), .B2(n20181), .ZN(
        n20169) );
  AOI22_X1 U23089 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20183), .B1(
        n20210), .B2(n20536), .ZN(n20168) );
  OAI211_X1 U23090 ( .C1(n20539), .C2(n20186), .A(n20169), .B(n20168), .ZN(
        P1_U3066) );
  AOI22_X1 U23091 ( .A1(n20541), .A2(n20182), .B1(n20540), .B2(n20181), .ZN(
        n20171) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20183), .B1(
        n20178), .B2(n20489), .ZN(n20170) );
  OAI211_X1 U23093 ( .C1(n20492), .C2(n20203), .A(n20171), .B(n20170), .ZN(
        P1_U3067) );
  AOI22_X1 U23094 ( .A1(n20547), .A2(n20182), .B1(n20546), .B2(n20181), .ZN(
        n20173) );
  INV_X1 U23095 ( .A(n20496), .ZN(n20548) );
  AOI22_X1 U23096 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20183), .B1(
        n20210), .B2(n20548), .ZN(n20172) );
  OAI211_X1 U23097 ( .C1(n20551), .C2(n20186), .A(n20173), .B(n20172), .ZN(
        P1_U3068) );
  AOI22_X1 U23098 ( .A1(n20553), .A2(n20182), .B1(n20552), .B2(n20181), .ZN(
        n20175) );
  INV_X1 U23099 ( .A(n20500), .ZN(n20554) );
  AOI22_X1 U23100 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20183), .B1(
        n20210), .B2(n20554), .ZN(n20174) );
  OAI211_X1 U23101 ( .C1(n20557), .C2(n20186), .A(n20175), .B(n20174), .ZN(
        P1_U3069) );
  AOI22_X1 U23102 ( .A1(n20559), .A2(n20182), .B1(n20558), .B2(n20181), .ZN(
        n20177) );
  INV_X1 U23103 ( .A(n20504), .ZN(n20560) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20183), .B1(
        n20210), .B2(n20560), .ZN(n20176) );
  OAI211_X1 U23105 ( .C1(n20563), .C2(n20186), .A(n20177), .B(n20176), .ZN(
        P1_U3070) );
  AOI22_X1 U23106 ( .A1(n20565), .A2(n20182), .B1(n20564), .B2(n20181), .ZN(
        n20180) );
  AOI22_X1 U23107 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20183), .B1(
        n20178), .B2(n20505), .ZN(n20179) );
  OAI211_X1 U23108 ( .C1(n20508), .C2(n20203), .A(n20180), .B(n20179), .ZN(
        P1_U3071) );
  AOI22_X1 U23109 ( .A1(n20573), .A2(n20182), .B1(n20571), .B2(n20181), .ZN(
        n20185) );
  AOI22_X1 U23110 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20183), .B1(
        n20210), .B2(n20574), .ZN(n20184) );
  OAI211_X1 U23111 ( .C1(n20580), .C2(n20186), .A(n20185), .B(n20184), .ZN(
        P1_U3072) );
  NOR2_X1 U23112 ( .A1(n20446), .A2(n20188), .ZN(n20208) );
  AOI21_X1 U23113 ( .B1(n20260), .B2(n20187), .A(n20208), .ZN(n20189) );
  OAI22_X1 U23114 ( .A1(n20189), .A2(n20377), .B1(n20188), .B2(n20700), .ZN(
        n20209) );
  AOI22_X1 U23115 ( .A1(n20524), .A2(n20209), .B1(n20523), .B2(n20208), .ZN(
        n20193) );
  INV_X1 U23116 ( .A(n20188), .ZN(n20191) );
  OAI211_X1 U23117 ( .C1(n20214), .C2(n20771), .A(n20189), .B(n20519), .ZN(
        n20190) );
  OAI211_X1 U23118 ( .C1(n20519), .C2(n20191), .A(n20527), .B(n20190), .ZN(
        n20211) );
  AOI22_X1 U23119 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20211), .B1(
        n20210), .B2(n20481), .ZN(n20192) );
  OAI211_X1 U23120 ( .C1(n20484), .C2(n20253), .A(n20193), .B(n20192), .ZN(
        P1_U3073) );
  AOI22_X1 U23121 ( .A1(n20535), .A2(n20209), .B1(n20534), .B2(n20208), .ZN(
        n20195) );
  AOI22_X1 U23122 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20211), .B1(
        n20210), .B2(n20485), .ZN(n20194) );
  OAI211_X1 U23123 ( .C1(n20488), .C2(n20253), .A(n20195), .B(n20194), .ZN(
        P1_U3074) );
  AOI22_X1 U23124 ( .A1(n20541), .A2(n20209), .B1(n20540), .B2(n20208), .ZN(
        n20197) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20211), .B1(
        n20210), .B2(n20489), .ZN(n20196) );
  OAI211_X1 U23126 ( .C1(n20492), .C2(n20253), .A(n20197), .B(n20196), .ZN(
        P1_U3075) );
  AOI22_X1 U23127 ( .A1(n20547), .A2(n20209), .B1(n20546), .B2(n20208), .ZN(
        n20199) );
  INV_X1 U23128 ( .A(n20253), .ZN(n20200) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20211), .B1(
        n20200), .B2(n20548), .ZN(n20198) );
  OAI211_X1 U23130 ( .C1(n20551), .C2(n20203), .A(n20199), .B(n20198), .ZN(
        P1_U3076) );
  AOI22_X1 U23131 ( .A1(n20553), .A2(n20209), .B1(n20552), .B2(n20208), .ZN(
        n20202) );
  AOI22_X1 U23132 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20211), .B1(
        n20200), .B2(n20554), .ZN(n20201) );
  OAI211_X1 U23133 ( .C1(n20557), .C2(n20203), .A(n20202), .B(n20201), .ZN(
        P1_U3077) );
  AOI22_X1 U23134 ( .A1(n20559), .A2(n20209), .B1(n20558), .B2(n20208), .ZN(
        n20205) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20211), .B1(
        n20210), .B2(n20501), .ZN(n20204) );
  OAI211_X1 U23136 ( .C1(n20504), .C2(n20253), .A(n20205), .B(n20204), .ZN(
        P1_U3078) );
  AOI22_X1 U23137 ( .A1(n20565), .A2(n20209), .B1(n20564), .B2(n20208), .ZN(
        n20207) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20211), .B1(
        n20210), .B2(n20505), .ZN(n20206) );
  OAI211_X1 U23139 ( .C1(n20508), .C2(n20253), .A(n20207), .B(n20206), .ZN(
        P1_U3079) );
  AOI22_X1 U23140 ( .A1(n20573), .A2(n20209), .B1(n20571), .B2(n20208), .ZN(
        n20213) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20211), .B1(
        n20210), .B2(n20511), .ZN(n20212) );
  OAI211_X1 U23142 ( .C1(n20516), .C2(n20253), .A(n20213), .B(n20212), .ZN(
        P1_U3080) );
  INV_X1 U23143 ( .A(n20010), .ZN(n20525) );
  OR2_X1 U23144 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20261), .ZN(
        n20251) );
  OAI22_X1 U23145 ( .A1(n20253), .A2(n20533), .B1(n20215), .B2(n20251), .ZN(
        n20216) );
  INV_X1 U23146 ( .A(n20216), .ZN(n20226) );
  NAND3_X1 U23147 ( .A1(n20288), .A2(n20519), .A3(n20253), .ZN(n20217) );
  NAND2_X1 U23148 ( .A1(n20217), .A2(n20668), .ZN(n20221) );
  OR2_X1 U23149 ( .A1(n20218), .A2(n13829), .ZN(n20223) );
  AOI22_X1 U23150 ( .A1(n20221), .A2(n20223), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20251), .ZN(n20220) );
  NAND3_X1 U23151 ( .A1(n20478), .A2(n20220), .A3(n20219), .ZN(n20256) );
  INV_X1 U23152 ( .A(n20221), .ZN(n20224) );
  OAI22_X1 U23153 ( .A1(n20224), .A2(n20223), .B1(n20222), .B2(n20471), .ZN(
        n20255) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20256), .B1(
        n20524), .B2(n20255), .ZN(n20225) );
  OAI211_X1 U23155 ( .C1(n20484), .C2(n20288), .A(n20226), .B(n20225), .ZN(
        P1_U3081) );
  OAI22_X1 U23156 ( .A1(n20253), .A2(n20539), .B1(n20227), .B2(n20251), .ZN(
        n20228) );
  INV_X1 U23157 ( .A(n20228), .ZN(n20230) );
  AOI22_X1 U23158 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20256), .B1(
        n20535), .B2(n20255), .ZN(n20229) );
  OAI211_X1 U23159 ( .C1(n20488), .C2(n20288), .A(n20230), .B(n20229), .ZN(
        P1_U3082) );
  OAI22_X1 U23160 ( .A1(n20253), .A2(n20545), .B1(n20231), .B2(n20251), .ZN(
        n20232) );
  INV_X1 U23161 ( .A(n20232), .ZN(n20234) );
  AOI22_X1 U23162 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20256), .B1(
        n20541), .B2(n20255), .ZN(n20233) );
  OAI211_X1 U23163 ( .C1(n20492), .C2(n20288), .A(n20234), .B(n20233), .ZN(
        P1_U3083) );
  OAI22_X1 U23164 ( .A1(n20288), .A2(n20496), .B1(n20235), .B2(n20251), .ZN(
        n20236) );
  INV_X1 U23165 ( .A(n20236), .ZN(n20238) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20256), .B1(
        n20547), .B2(n20255), .ZN(n20237) );
  OAI211_X1 U23167 ( .C1(n20551), .C2(n20253), .A(n20238), .B(n20237), .ZN(
        P1_U3084) );
  OAI22_X1 U23168 ( .A1(n20253), .A2(n20557), .B1(n20239), .B2(n20251), .ZN(
        n20240) );
  INV_X1 U23169 ( .A(n20240), .ZN(n20242) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20256), .B1(
        n20553), .B2(n20255), .ZN(n20241) );
  OAI211_X1 U23171 ( .C1(n20500), .C2(n20288), .A(n20242), .B(n20241), .ZN(
        P1_U3085) );
  OAI22_X1 U23172 ( .A1(n20288), .A2(n20504), .B1(n20243), .B2(n20251), .ZN(
        n20244) );
  INV_X1 U23173 ( .A(n20244), .ZN(n20246) );
  AOI22_X1 U23174 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20256), .B1(
        n20559), .B2(n20255), .ZN(n20245) );
  OAI211_X1 U23175 ( .C1(n20563), .C2(n20253), .A(n20246), .B(n20245), .ZN(
        P1_U3086) );
  OAI22_X1 U23176 ( .A1(n20253), .A2(n20569), .B1(n20247), .B2(n20251), .ZN(
        n20248) );
  INV_X1 U23177 ( .A(n20248), .ZN(n20250) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20256), .B1(
        n20565), .B2(n20255), .ZN(n20249) );
  OAI211_X1 U23179 ( .C1(n20508), .C2(n20288), .A(n20250), .B(n20249), .ZN(
        P1_U3087) );
  OAI22_X1 U23180 ( .A1(n20253), .A2(n20580), .B1(n20252), .B2(n20251), .ZN(
        n20254) );
  INV_X1 U23181 ( .A(n20254), .ZN(n20258) );
  AOI22_X1 U23182 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20256), .B1(
        n20573), .B2(n20255), .ZN(n20257) );
  OAI211_X1 U23183 ( .C1(n20516), .C2(n20288), .A(n20258), .B(n20257), .ZN(
        P1_U3088) );
  NAND2_X1 U23184 ( .A1(n20664), .A2(n20259), .ZN(n20282) );
  AOI21_X1 U23185 ( .B1(n20260), .B2(n20517), .A(n20283), .ZN(n20263) );
  OAI22_X1 U23186 ( .A1(n20263), .A2(n20377), .B1(n20261), .B2(n20700), .ZN(
        n20284) );
  AOI22_X1 U23187 ( .A1(n20524), .A2(n20284), .B1(n20523), .B2(n20283), .ZN(
        n20268) );
  NOR2_X1 U23188 ( .A1(n20262), .A2(n20377), .ZN(n20264) );
  OAI21_X1 U23189 ( .B1(n20264), .B2(n20675), .A(n20263), .ZN(n20265) );
  OAI211_X1 U23190 ( .C1(n20266), .C2(n20519), .A(n20527), .B(n20265), .ZN(
        n20285) );
  INV_X1 U23191 ( .A(n20288), .ZN(n20279) );
  AOI22_X1 U23192 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20285), .B1(
        n20279), .B2(n20481), .ZN(n20267) );
  OAI211_X1 U23193 ( .C1(n20484), .C2(n20282), .A(n20268), .B(n20267), .ZN(
        P1_U3089) );
  AOI22_X1 U23194 ( .A1(n20535), .A2(n20284), .B1(n20534), .B2(n20283), .ZN(
        n20270) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20285), .B1(
        n20279), .B2(n20485), .ZN(n20269) );
  OAI211_X1 U23196 ( .C1(n20488), .C2(n20282), .A(n20270), .B(n20269), .ZN(
        P1_U3090) );
  AOI22_X1 U23197 ( .A1(n20541), .A2(n20284), .B1(n20540), .B2(n20283), .ZN(
        n20272) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20285), .B1(
        n20279), .B2(n20489), .ZN(n20271) );
  OAI211_X1 U23199 ( .C1(n20492), .C2(n20282), .A(n20272), .B(n20271), .ZN(
        P1_U3091) );
  AOI22_X1 U23200 ( .A1(n20547), .A2(n20284), .B1(n20546), .B2(n20283), .ZN(
        n20274) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20285), .B1(
        n20313), .B2(n20548), .ZN(n20273) );
  OAI211_X1 U23202 ( .C1(n20551), .C2(n20288), .A(n20274), .B(n20273), .ZN(
        P1_U3092) );
  AOI22_X1 U23203 ( .A1(n20553), .A2(n20284), .B1(n20552), .B2(n20283), .ZN(
        n20276) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20285), .B1(
        n20313), .B2(n20554), .ZN(n20275) );
  OAI211_X1 U23205 ( .C1(n20557), .C2(n20288), .A(n20276), .B(n20275), .ZN(
        P1_U3093) );
  AOI22_X1 U23206 ( .A1(n20559), .A2(n20284), .B1(n20558), .B2(n20283), .ZN(
        n20278) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20285), .B1(
        n20279), .B2(n20501), .ZN(n20277) );
  OAI211_X1 U23208 ( .C1(n20504), .C2(n20282), .A(n20278), .B(n20277), .ZN(
        P1_U3094) );
  AOI22_X1 U23209 ( .A1(n20565), .A2(n20284), .B1(n20564), .B2(n20283), .ZN(
        n20281) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20285), .B1(
        n20279), .B2(n20505), .ZN(n20280) );
  OAI211_X1 U23211 ( .C1(n20508), .C2(n20282), .A(n20281), .B(n20280), .ZN(
        P1_U3095) );
  AOI22_X1 U23212 ( .A1(n20573), .A2(n20284), .B1(n20571), .B2(n20283), .ZN(
        n20287) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20285), .B1(
        n20313), .B2(n20574), .ZN(n20286) );
  OAI211_X1 U23214 ( .C1(n20580), .C2(n20288), .A(n20287), .B(n20286), .ZN(
        P1_U3096) );
  NAND2_X1 U23215 ( .A1(n20666), .A2(n20678), .ZN(n20346) );
  INV_X1 U23216 ( .A(n20346), .ZN(n20376) );
  NAND3_X1 U23217 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20681), .A3(
        n20690), .ZN(n20319) );
  NOR2_X1 U23218 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20319), .ZN(
        n20311) );
  AOI21_X1 U23219 ( .B1(n20376), .B2(n13829), .A(n20311), .ZN(n20294) );
  NOR2_X1 U23220 ( .A1(n20291), .A2(n20290), .ZN(n20414) );
  INV_X1 U23221 ( .A(n20414), .ZN(n20292) );
  OAI22_X1 U23222 ( .A1(n20294), .A2(n20377), .B1(n20292), .B2(n20352), .ZN(
        n20312) );
  AOI22_X1 U23223 ( .A1(n20524), .A2(n20312), .B1(n20523), .B2(n20311), .ZN(
        n20298) );
  INV_X1 U23224 ( .A(n20343), .ZN(n20293) );
  OAI21_X1 U23225 ( .B1(n20293), .B2(n20313), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20295) );
  NAND2_X1 U23226 ( .A1(n20295), .A2(n20294), .ZN(n20296) );
  OAI211_X1 U23227 ( .C1(n20311), .C2(n20780), .A(n20350), .B(n20296), .ZN(
        n20314) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20314), .B1(
        n20313), .B2(n20481), .ZN(n20297) );
  OAI211_X1 U23229 ( .C1(n20484), .C2(n20343), .A(n20298), .B(n20297), .ZN(
        P1_U3097) );
  AOI22_X1 U23230 ( .A1(n20535), .A2(n20312), .B1(n20534), .B2(n20311), .ZN(
        n20300) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20314), .B1(
        n20313), .B2(n20485), .ZN(n20299) );
  OAI211_X1 U23232 ( .C1(n20488), .C2(n20343), .A(n20300), .B(n20299), .ZN(
        P1_U3098) );
  AOI22_X1 U23233 ( .A1(n20541), .A2(n20312), .B1(n20540), .B2(n20311), .ZN(
        n20302) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20314), .B1(
        n20313), .B2(n20489), .ZN(n20301) );
  OAI211_X1 U23235 ( .C1(n20492), .C2(n20343), .A(n20302), .B(n20301), .ZN(
        P1_U3099) );
  AOI22_X1 U23236 ( .A1(n20547), .A2(n20312), .B1(n20546), .B2(n20311), .ZN(
        n20304) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20314), .B1(
        n20313), .B2(n20493), .ZN(n20303) );
  OAI211_X1 U23238 ( .C1(n20496), .C2(n20343), .A(n20304), .B(n20303), .ZN(
        P1_U3100) );
  AOI22_X1 U23239 ( .A1(n20553), .A2(n20312), .B1(n20552), .B2(n20311), .ZN(
        n20306) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20314), .B1(
        n20313), .B2(n20497), .ZN(n20305) );
  OAI211_X1 U23241 ( .C1(n20500), .C2(n20343), .A(n20306), .B(n20305), .ZN(
        P1_U3101) );
  AOI22_X1 U23242 ( .A1(n20559), .A2(n20312), .B1(n20558), .B2(n20311), .ZN(
        n20308) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20314), .B1(
        n20313), .B2(n20501), .ZN(n20307) );
  OAI211_X1 U23244 ( .C1(n20504), .C2(n20343), .A(n20308), .B(n20307), .ZN(
        P1_U3102) );
  AOI22_X1 U23245 ( .A1(n20565), .A2(n20312), .B1(n20564), .B2(n20311), .ZN(
        n20310) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20314), .B1(
        n20313), .B2(n20505), .ZN(n20309) );
  OAI211_X1 U23247 ( .C1(n20508), .C2(n20343), .A(n20310), .B(n20309), .ZN(
        P1_U3103) );
  AOI22_X1 U23248 ( .A1(n20573), .A2(n20312), .B1(n20571), .B2(n20311), .ZN(
        n20316) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20314), .B1(
        n20313), .B2(n20511), .ZN(n20315) );
  OAI211_X1 U23250 ( .C1(n20516), .C2(n20343), .A(n20316), .B(n20315), .ZN(
        P1_U3104) );
  OR2_X1 U23251 ( .A1(n20346), .A2(n20057), .ZN(n20318) );
  NOR2_X1 U23252 ( .A1(n20446), .A2(n20319), .ZN(n20338) );
  INV_X1 U23253 ( .A(n20338), .ZN(n20317) );
  AND2_X1 U23254 ( .A1(n20318), .A2(n20317), .ZN(n20320) );
  OAI22_X1 U23255 ( .A1(n20320), .A2(n20377), .B1(n20319), .B2(n20700), .ZN(
        n20339) );
  AOI22_X1 U23256 ( .A1(n20524), .A2(n20339), .B1(n20523), .B2(n20338), .ZN(
        n20325) );
  INV_X1 U23257 ( .A(n20319), .ZN(n20323) );
  OAI21_X1 U23258 ( .B1(n20377), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20665), 
        .ZN(n20321) );
  NAND2_X1 U23259 ( .A1(n20321), .A2(n20320), .ZN(n20322) );
  OAI211_X1 U23260 ( .C1(n20519), .C2(n20323), .A(n20527), .B(n20322), .ZN(
        n20340) );
  INV_X1 U23261 ( .A(n20484), .ZN(n20530) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20340), .B1(
        n20370), .B2(n20530), .ZN(n20324) );
  OAI211_X1 U23263 ( .C1(n20533), .C2(n20343), .A(n20325), .B(n20324), .ZN(
        P1_U3105) );
  AOI22_X1 U23264 ( .A1(n20535), .A2(n20339), .B1(n20534), .B2(n20338), .ZN(
        n20327) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20340), .B1(
        n20370), .B2(n20536), .ZN(n20326) );
  OAI211_X1 U23266 ( .C1(n20539), .C2(n20343), .A(n20327), .B(n20326), .ZN(
        P1_U3106) );
  AOI22_X1 U23267 ( .A1(n20541), .A2(n20339), .B1(n20540), .B2(n20338), .ZN(
        n20329) );
  INV_X1 U23268 ( .A(n20492), .ZN(n20542) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20340), .B1(
        n20370), .B2(n20542), .ZN(n20328) );
  OAI211_X1 U23270 ( .C1(n20545), .C2(n20343), .A(n20329), .B(n20328), .ZN(
        P1_U3107) );
  AOI22_X1 U23271 ( .A1(n20547), .A2(n20339), .B1(n20546), .B2(n20338), .ZN(
        n20331) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20340), .B1(
        n20370), .B2(n20548), .ZN(n20330) );
  OAI211_X1 U23273 ( .C1(n20551), .C2(n20343), .A(n20331), .B(n20330), .ZN(
        P1_U3108) );
  AOI22_X1 U23274 ( .A1(n20553), .A2(n20339), .B1(n20552), .B2(n20338), .ZN(
        n20333) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20340), .B1(
        n20370), .B2(n20554), .ZN(n20332) );
  OAI211_X1 U23276 ( .C1(n20557), .C2(n20343), .A(n20333), .B(n20332), .ZN(
        P1_U3109) );
  AOI22_X1 U23277 ( .A1(n20559), .A2(n20339), .B1(n20558), .B2(n20338), .ZN(
        n20335) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20340), .B1(
        n20370), .B2(n20560), .ZN(n20334) );
  OAI211_X1 U23279 ( .C1(n20563), .C2(n20343), .A(n20335), .B(n20334), .ZN(
        P1_U3110) );
  AOI22_X1 U23280 ( .A1(n20565), .A2(n20339), .B1(n20564), .B2(n20338), .ZN(
        n20337) );
  INV_X1 U23281 ( .A(n20508), .ZN(n20566) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20340), .B1(
        n20370), .B2(n20566), .ZN(n20336) );
  OAI211_X1 U23283 ( .C1(n20569), .C2(n20343), .A(n20337), .B(n20336), .ZN(
        P1_U3111) );
  AOI22_X1 U23284 ( .A1(n20573), .A2(n20339), .B1(n20571), .B2(n20338), .ZN(
        n20342) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20340), .B1(
        n20370), .B2(n20574), .ZN(n20341) );
  OAI211_X1 U23286 ( .C1(n20580), .C2(n20343), .A(n20342), .B(n20341), .ZN(
        P1_U3112) );
  NAND3_X1 U23287 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20681), .ZN(n20379) );
  NOR2_X1 U23288 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20379), .ZN(
        n20369) );
  AOI22_X1 U23289 ( .A1(n20370), .A2(n20481), .B1(n20523), .B2(n20369), .ZN(
        n20356) );
  INV_X1 U23290 ( .A(n20370), .ZN(n20344) );
  NAND3_X1 U23291 ( .A1(n20344), .A2(n20519), .A3(n20403), .ZN(n20345) );
  NAND2_X1 U23292 ( .A1(n20345), .A2(n20668), .ZN(n20351) );
  OR2_X1 U23293 ( .A1(n20346), .A2(n13829), .ZN(n20353) );
  INV_X1 U23294 ( .A(n20369), .ZN(n20347) );
  AOI22_X1 U23295 ( .A1(n20351), .A2(n20353), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20347), .ZN(n20349) );
  OR2_X1 U23296 ( .A1(n20348), .A2(n20673), .ZN(n20472) );
  NAND2_X1 U23297 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20472), .ZN(n20477) );
  NAND3_X1 U23298 ( .A1(n20350), .A2(n20349), .A3(n20477), .ZN(n20372) );
  INV_X1 U23299 ( .A(n20351), .ZN(n20354) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20372), .B1(
        n20524), .B2(n20371), .ZN(n20355) );
  OAI211_X1 U23301 ( .C1(n20484), .C2(n20403), .A(n20356), .B(n20355), .ZN(
        P1_U3113) );
  AOI22_X1 U23302 ( .A1(n20370), .A2(n20485), .B1(n20534), .B2(n20369), .ZN(
        n20358) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20372), .B1(
        n20535), .B2(n20371), .ZN(n20357) );
  OAI211_X1 U23304 ( .C1(n20488), .C2(n20403), .A(n20358), .B(n20357), .ZN(
        P1_U3114) );
  AOI22_X1 U23305 ( .A1(n20370), .A2(n20489), .B1(n20540), .B2(n20369), .ZN(
        n20360) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20372), .B1(
        n20541), .B2(n20371), .ZN(n20359) );
  OAI211_X1 U23307 ( .C1(n20492), .C2(n20403), .A(n20360), .B(n20359), .ZN(
        P1_U3115) );
  AOI22_X1 U23308 ( .A1(n20370), .A2(n20493), .B1(n20546), .B2(n20369), .ZN(
        n20362) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20372), .B1(
        n20547), .B2(n20371), .ZN(n20361) );
  OAI211_X1 U23310 ( .C1(n20496), .C2(n20403), .A(n20362), .B(n20361), .ZN(
        P1_U3116) );
  AOI22_X1 U23311 ( .A1(n20370), .A2(n20497), .B1(n20552), .B2(n20369), .ZN(
        n20364) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20372), .B1(
        n20553), .B2(n20371), .ZN(n20363) );
  OAI211_X1 U23313 ( .C1(n20500), .C2(n20403), .A(n20364), .B(n20363), .ZN(
        P1_U3117) );
  AOI22_X1 U23314 ( .A1(n20370), .A2(n20501), .B1(n20558), .B2(n20369), .ZN(
        n20366) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20372), .B1(
        n20559), .B2(n20371), .ZN(n20365) );
  OAI211_X1 U23316 ( .C1(n20504), .C2(n20403), .A(n20366), .B(n20365), .ZN(
        P1_U3118) );
  AOI22_X1 U23317 ( .A1(n20370), .A2(n20505), .B1(n20564), .B2(n20369), .ZN(
        n20368) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20372), .B1(
        n20565), .B2(n20371), .ZN(n20367) );
  OAI211_X1 U23319 ( .C1(n20508), .C2(n20403), .A(n20368), .B(n20367), .ZN(
        P1_U3119) );
  AOI22_X1 U23320 ( .A1(n20370), .A2(n20511), .B1(n20571), .B2(n20369), .ZN(
        n20374) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20372), .B1(
        n20573), .B2(n20371), .ZN(n20373) );
  OAI211_X1 U23322 ( .C1(n20516), .C2(n20403), .A(n20374), .B(n20373), .ZN(
        P1_U3120) );
  NOR2_X1 U23323 ( .A1(n20375), .A2(n20673), .ZN(n20398) );
  AOI21_X1 U23324 ( .B1(n20376), .B2(n20517), .A(n20398), .ZN(n20378) );
  OAI22_X1 U23325 ( .A1(n20378), .A2(n20377), .B1(n20379), .B2(n20700), .ZN(
        n20399) );
  AOI22_X1 U23326 ( .A1(n20524), .A2(n20399), .B1(n20523), .B2(n20398), .ZN(
        n20385) );
  INV_X1 U23327 ( .A(n20379), .ZN(n20382) );
  INV_X1 U23328 ( .A(n20380), .ZN(n20684) );
  NAND3_X1 U23329 ( .A1(n9617), .A2(n20684), .A3(n20010), .ZN(n20676) );
  NOR2_X1 U23330 ( .A1(n20676), .A2(n11701), .ZN(n20381) );
  OAI21_X1 U23331 ( .B1(n20382), .B2(n20381), .A(n20527), .ZN(n20400) );
  AOI22_X1 U23332 ( .A1(n20400), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n20437), .B2(n20530), .ZN(n20384) );
  OAI211_X1 U23333 ( .C1(n20533), .C2(n20403), .A(n20385), .B(n20384), .ZN(
        P1_U3121) );
  AOI22_X1 U23334 ( .A1(n20535), .A2(n20399), .B1(n20534), .B2(n20398), .ZN(
        n20387) );
  AOI22_X1 U23335 ( .A1(n20400), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n20437), .B2(n20536), .ZN(n20386) );
  OAI211_X1 U23336 ( .C1(n20539), .C2(n20403), .A(n20387), .B(n20386), .ZN(
        P1_U3122) );
  AOI22_X1 U23337 ( .A1(n20541), .A2(n20399), .B1(n20540), .B2(n20398), .ZN(
        n20389) );
  AOI22_X1 U23338 ( .A1(n20400), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n20437), .B2(n20542), .ZN(n20388) );
  OAI211_X1 U23339 ( .C1(n20545), .C2(n20403), .A(n20389), .B(n20388), .ZN(
        P1_U3123) );
  AOI22_X1 U23340 ( .A1(n20547), .A2(n20399), .B1(n20546), .B2(n20398), .ZN(
        n20391) );
  AOI22_X1 U23341 ( .A1(n20400), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n20437), .B2(n20548), .ZN(n20390) );
  OAI211_X1 U23342 ( .C1(n20551), .C2(n20403), .A(n20391), .B(n20390), .ZN(
        P1_U3124) );
  AOI22_X1 U23343 ( .A1(n20553), .A2(n20399), .B1(n20552), .B2(n20398), .ZN(
        n20393) );
  AOI22_X1 U23344 ( .A1(n20400), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n20437), .B2(n20554), .ZN(n20392) );
  OAI211_X1 U23345 ( .C1(n20557), .C2(n20403), .A(n20393), .B(n20392), .ZN(
        P1_U3125) );
  AOI22_X1 U23346 ( .A1(n20559), .A2(n20399), .B1(n20558), .B2(n20398), .ZN(
        n20395) );
  AOI22_X1 U23347 ( .A1(n20400), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n20437), .B2(n20560), .ZN(n20394) );
  OAI211_X1 U23348 ( .C1(n20563), .C2(n20403), .A(n20395), .B(n20394), .ZN(
        P1_U3126) );
  AOI22_X1 U23349 ( .A1(n20565), .A2(n20399), .B1(n20564), .B2(n20398), .ZN(
        n20397) );
  AOI22_X1 U23350 ( .A1(n20400), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n20437), .B2(n20566), .ZN(n20396) );
  OAI211_X1 U23351 ( .C1(n20569), .C2(n20403), .A(n20397), .B(n20396), .ZN(
        P1_U3127) );
  AOI22_X1 U23352 ( .A1(n20573), .A2(n20399), .B1(n20571), .B2(n20398), .ZN(
        n20402) );
  AOI22_X1 U23353 ( .A1(n20400), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n20437), .B2(n20574), .ZN(n20401) );
  OAI211_X1 U23354 ( .C1(n20580), .C2(n20403), .A(n20402), .B(n20401), .ZN(
        P1_U3128) );
  INV_X1 U23355 ( .A(n20465), .ZN(n20405) );
  NAND2_X1 U23356 ( .A1(n20405), .A2(n20519), .ZN(n20406) );
  OAI21_X1 U23357 ( .B1(n20406), .B2(n20437), .A(n20668), .ZN(n20412) );
  OR2_X1 U23358 ( .A1(n20678), .A2(n20407), .ZN(n20444) );
  NOR2_X1 U23359 ( .A1(n20444), .A2(n20687), .ZN(n20409) );
  INV_X1 U23360 ( .A(n20524), .ZN(n20417) );
  NAND3_X1 U23361 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20690), .ZN(n20445) );
  NOR2_X1 U23362 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20445), .ZN(
        n20436) );
  AOI22_X1 U23363 ( .A1(n20465), .A2(n20530), .B1(n20523), .B2(n20436), .ZN(
        n20416) );
  INV_X1 U23364 ( .A(n20409), .ZN(n20411) );
  INV_X1 U23365 ( .A(n20436), .ZN(n20410) );
  AOI22_X1 U23366 ( .A1(n20412), .A2(n20411), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20410), .ZN(n20413) );
  OAI211_X1 U23367 ( .C1(n20414), .C2(n20700), .A(n20478), .B(n20413), .ZN(
        n20438) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20481), .ZN(n20415) );
  OAI211_X1 U23369 ( .C1(n20442), .C2(n20417), .A(n20416), .B(n20415), .ZN(
        P1_U3129) );
  INV_X1 U23370 ( .A(n20535), .ZN(n20420) );
  AOI22_X1 U23371 ( .A1(n20465), .A2(n20536), .B1(n20534), .B2(n20436), .ZN(
        n20419) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20485), .ZN(n20418) );
  OAI211_X1 U23373 ( .C1(n20442), .C2(n20420), .A(n20419), .B(n20418), .ZN(
        P1_U3130) );
  INV_X1 U23374 ( .A(n20541), .ZN(n20423) );
  AOI22_X1 U23375 ( .A1(n20465), .A2(n20542), .B1(n20540), .B2(n20436), .ZN(
        n20422) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20489), .ZN(n20421) );
  OAI211_X1 U23377 ( .C1(n20442), .C2(n20423), .A(n20422), .B(n20421), .ZN(
        P1_U3131) );
  INV_X1 U23378 ( .A(n20547), .ZN(n20426) );
  AOI22_X1 U23379 ( .A1(n20465), .A2(n20548), .B1(n20546), .B2(n20436), .ZN(
        n20425) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20493), .ZN(n20424) );
  OAI211_X1 U23381 ( .C1(n20442), .C2(n20426), .A(n20425), .B(n20424), .ZN(
        P1_U3132) );
  INV_X1 U23382 ( .A(n20553), .ZN(n20429) );
  AOI22_X1 U23383 ( .A1(n20465), .A2(n20554), .B1(n20552), .B2(n20436), .ZN(
        n20428) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20497), .ZN(n20427) );
  OAI211_X1 U23385 ( .C1(n20442), .C2(n20429), .A(n20428), .B(n20427), .ZN(
        P1_U3133) );
  INV_X1 U23386 ( .A(n20559), .ZN(n20432) );
  AOI22_X1 U23387 ( .A1(n20465), .A2(n20560), .B1(n20558), .B2(n20436), .ZN(
        n20431) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20501), .ZN(n20430) );
  OAI211_X1 U23389 ( .C1(n20442), .C2(n20432), .A(n20431), .B(n20430), .ZN(
        P1_U3134) );
  INV_X1 U23390 ( .A(n20565), .ZN(n20435) );
  AOI22_X1 U23391 ( .A1(n20465), .A2(n20566), .B1(n20564), .B2(n20436), .ZN(
        n20434) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20505), .ZN(n20433) );
  OAI211_X1 U23393 ( .C1(n20442), .C2(n20435), .A(n20434), .B(n20433), .ZN(
        P1_U3135) );
  INV_X1 U23394 ( .A(n20573), .ZN(n20441) );
  AOI22_X1 U23395 ( .A1(n20465), .A2(n20574), .B1(n20571), .B2(n20436), .ZN(
        n20440) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20511), .ZN(n20439) );
  OAI211_X1 U23397 ( .C1(n20442), .C2(n20441), .A(n20440), .B(n20439), .ZN(
        P1_U3136) );
  INV_X1 U23398 ( .A(n20444), .ZN(n20475) );
  NAND2_X1 U23399 ( .A1(n20475), .A2(n20519), .ZN(n20522) );
  INV_X1 U23400 ( .A(n20445), .ZN(n20448) );
  NOR2_X1 U23401 ( .A1(n20446), .A2(n20445), .ZN(n20463) );
  AOI22_X1 U23402 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20448), .B1(n20463), 
        .B2(n20519), .ZN(n20447) );
  OAI21_X1 U23403 ( .B1(n20522), .B2(n20057), .A(n20447), .ZN(n20464) );
  AOI22_X1 U23404 ( .A1(n20524), .A2(n20464), .B1(n20523), .B2(n20463), .ZN(
        n20450) );
  NAND2_X1 U23405 ( .A1(n20470), .A2(n20684), .ZN(n20526) );
  NOR2_X1 U23406 ( .A1(n20526), .A2(n20010), .ZN(n20669) );
  OAI21_X1 U23407 ( .B1(n20448), .B2(n20669), .A(n20527), .ZN(n20466) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20481), .ZN(n20449) );
  OAI211_X1 U23409 ( .C1(n20484), .C2(n20480), .A(n20450), .B(n20449), .ZN(
        P1_U3137) );
  AOI22_X1 U23410 ( .A1(n20535), .A2(n20464), .B1(n20534), .B2(n20463), .ZN(
        n20452) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20485), .ZN(n20451) );
  OAI211_X1 U23412 ( .C1(n20488), .C2(n20480), .A(n20452), .B(n20451), .ZN(
        P1_U3138) );
  AOI22_X1 U23413 ( .A1(n20541), .A2(n20464), .B1(n20540), .B2(n20463), .ZN(
        n20454) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20489), .ZN(n20453) );
  OAI211_X1 U23415 ( .C1(n20492), .C2(n20480), .A(n20454), .B(n20453), .ZN(
        P1_U3139) );
  AOI22_X1 U23416 ( .A1(n20547), .A2(n20464), .B1(n20546), .B2(n20463), .ZN(
        n20456) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20493), .ZN(n20455) );
  OAI211_X1 U23418 ( .C1(n20496), .C2(n20480), .A(n20456), .B(n20455), .ZN(
        P1_U3140) );
  AOI22_X1 U23419 ( .A1(n20553), .A2(n20464), .B1(n20552), .B2(n20463), .ZN(
        n20458) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20497), .ZN(n20457) );
  OAI211_X1 U23421 ( .C1(n20500), .C2(n20480), .A(n20458), .B(n20457), .ZN(
        P1_U3141) );
  AOI22_X1 U23422 ( .A1(n20559), .A2(n20464), .B1(n20558), .B2(n20463), .ZN(
        n20460) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20501), .ZN(n20459) );
  OAI211_X1 U23424 ( .C1(n20504), .C2(n20480), .A(n20460), .B(n20459), .ZN(
        P1_U3142) );
  AOI22_X1 U23425 ( .A1(n20565), .A2(n20464), .B1(n20564), .B2(n20463), .ZN(
        n20462) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20505), .ZN(n20461) );
  OAI211_X1 U23427 ( .C1(n20508), .C2(n20480), .A(n20462), .B(n20461), .ZN(
        P1_U3143) );
  AOI22_X1 U23428 ( .A1(n20573), .A2(n20464), .B1(n20571), .B2(n20463), .ZN(
        n20468) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20511), .ZN(n20467) );
  OAI211_X1 U23430 ( .C1(n20516), .C2(n20480), .A(n20468), .B(n20467), .ZN(
        P1_U3144) );
  OAI22_X1 U23431 ( .A1(n20522), .A2(n13829), .B1(n20472), .B2(n20471), .ZN(
        n20510) );
  NOR2_X1 U23432 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20473), .ZN(
        n20509) );
  AOI22_X1 U23433 ( .A1(n20524), .A2(n20510), .B1(n20523), .B2(n20509), .ZN(
        n20483) );
  AOI21_X1 U23434 ( .B1(n20480), .B2(n20579), .A(n20771), .ZN(n20474) );
  AOI21_X1 U23435 ( .B1(n20475), .B2(n20687), .A(n20474), .ZN(n20476) );
  NOR2_X1 U23436 ( .A1(n20476), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20479) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20481), .ZN(n20482) );
  OAI211_X1 U23438 ( .C1(n20484), .C2(n20579), .A(n20483), .B(n20482), .ZN(
        P1_U3145) );
  AOI22_X1 U23439 ( .A1(n20535), .A2(n20510), .B1(n20534), .B2(n20509), .ZN(
        n20487) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20485), .ZN(n20486) );
  OAI211_X1 U23441 ( .C1(n20488), .C2(n20579), .A(n20487), .B(n20486), .ZN(
        P1_U3146) );
  AOI22_X1 U23442 ( .A1(n20541), .A2(n20510), .B1(n20540), .B2(n20509), .ZN(
        n20491) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20489), .ZN(n20490) );
  OAI211_X1 U23444 ( .C1(n20492), .C2(n20579), .A(n20491), .B(n20490), .ZN(
        P1_U3147) );
  AOI22_X1 U23445 ( .A1(n20547), .A2(n20510), .B1(n20546), .B2(n20509), .ZN(
        n20495) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20493), .ZN(n20494) );
  OAI211_X1 U23447 ( .C1(n20496), .C2(n20579), .A(n20495), .B(n20494), .ZN(
        P1_U3148) );
  AOI22_X1 U23448 ( .A1(n20553), .A2(n20510), .B1(n20552), .B2(n20509), .ZN(
        n20499) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20497), .ZN(n20498) );
  OAI211_X1 U23450 ( .C1(n20500), .C2(n20579), .A(n20499), .B(n20498), .ZN(
        P1_U3149) );
  AOI22_X1 U23451 ( .A1(n20559), .A2(n20510), .B1(n20558), .B2(n20509), .ZN(
        n20503) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20501), .ZN(n20502) );
  OAI211_X1 U23453 ( .C1(n20504), .C2(n20579), .A(n20503), .B(n20502), .ZN(
        P1_U3150) );
  AOI22_X1 U23454 ( .A1(n20565), .A2(n20510), .B1(n20564), .B2(n20509), .ZN(
        n20507) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20505), .ZN(n20506) );
  OAI211_X1 U23456 ( .C1(n20508), .C2(n20579), .A(n20507), .B(n20506), .ZN(
        P1_U3151) );
  AOI22_X1 U23457 ( .A1(n20573), .A2(n20510), .B1(n20571), .B2(n20509), .ZN(
        n20515) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20511), .ZN(n20514) );
  OAI211_X1 U23459 ( .C1(n20516), .C2(n20579), .A(n20515), .B(n20514), .ZN(
        P1_U3152) );
  INV_X1 U23460 ( .A(n20517), .ZN(n20521) );
  INV_X1 U23461 ( .A(n20518), .ZN(n20570) );
  AOI22_X1 U23462 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20529), .B1(n20570), 
        .B2(n20519), .ZN(n20520) );
  OAI21_X1 U23463 ( .B1(n20522), .B2(n20521), .A(n20520), .ZN(n20572) );
  AOI22_X1 U23464 ( .A1(n20524), .A2(n20572), .B1(n20523), .B2(n20570), .ZN(
        n20532) );
  NOR2_X1 U23465 ( .A1(n20526), .A2(n20525), .ZN(n20528) );
  OAI21_X1 U23466 ( .B1(n20529), .B2(n20528), .A(n20527), .ZN(n20576) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20530), .ZN(n20531) );
  OAI211_X1 U23468 ( .C1(n20533), .C2(n20579), .A(n20532), .B(n20531), .ZN(
        P1_U3153) );
  AOI22_X1 U23469 ( .A1(n20535), .A2(n20572), .B1(n20534), .B2(n20570), .ZN(
        n20538) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20536), .ZN(n20537) );
  OAI211_X1 U23471 ( .C1(n20539), .C2(n20579), .A(n20538), .B(n20537), .ZN(
        P1_U3154) );
  AOI22_X1 U23472 ( .A1(n20541), .A2(n20572), .B1(n20540), .B2(n20570), .ZN(
        n20544) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20542), .ZN(n20543) );
  OAI211_X1 U23474 ( .C1(n20545), .C2(n20579), .A(n20544), .B(n20543), .ZN(
        P1_U3155) );
  AOI22_X1 U23475 ( .A1(n20547), .A2(n20572), .B1(n20546), .B2(n20570), .ZN(
        n20550) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20548), .ZN(n20549) );
  OAI211_X1 U23477 ( .C1(n20551), .C2(n20579), .A(n20550), .B(n20549), .ZN(
        P1_U3156) );
  AOI22_X1 U23478 ( .A1(n20553), .A2(n20572), .B1(n20552), .B2(n20570), .ZN(
        n20556) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20554), .ZN(n20555) );
  OAI211_X1 U23480 ( .C1(n20557), .C2(n20579), .A(n20556), .B(n20555), .ZN(
        P1_U3157) );
  AOI22_X1 U23481 ( .A1(n20559), .A2(n20572), .B1(n20558), .B2(n20570), .ZN(
        n20562) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20560), .ZN(n20561) );
  OAI211_X1 U23483 ( .C1(n20563), .C2(n20579), .A(n20562), .B(n20561), .ZN(
        P1_U3158) );
  AOI22_X1 U23484 ( .A1(n20565), .A2(n20572), .B1(n20564), .B2(n20570), .ZN(
        n20568) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20566), .ZN(n20567) );
  OAI211_X1 U23486 ( .C1(n20569), .C2(n20579), .A(n20568), .B(n20567), .ZN(
        P1_U3159) );
  AOI22_X1 U23487 ( .A1(n20573), .A2(n20572), .B1(n20571), .B2(n20570), .ZN(
        n20578) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20574), .ZN(n20577) );
  OAI211_X1 U23489 ( .C1(n20580), .C2(n20579), .A(n20578), .B(n20577), .ZN(
        P1_U3160) );
  INV_X1 U23490 ( .A(n20581), .ZN(n20583) );
  OAI211_X1 U23491 ( .C1(n20584), .C2(n20700), .A(n20583), .B(n20582), .ZN(
        P1_U3163) );
  AND2_X1 U23492 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20659), .ZN(
        P1_U3164) );
  AND2_X1 U23493 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20659), .ZN(
        P1_U3165) );
  AND2_X1 U23494 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20659), .ZN(
        P1_U3166) );
  AND2_X1 U23495 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20659), .ZN(
        P1_U3167) );
  AND2_X1 U23496 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20659), .ZN(
        P1_U3168) );
  AND2_X1 U23497 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20659), .ZN(
        P1_U3169) );
  AND2_X1 U23498 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20659), .ZN(
        P1_U3170) );
  AND2_X1 U23499 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20659), .ZN(
        P1_U3171) );
  AND2_X1 U23500 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20659), .ZN(
        P1_U3172) );
  AND2_X1 U23501 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20659), .ZN(
        P1_U3173) );
  AND2_X1 U23502 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20659), .ZN(
        P1_U3174) );
  AND2_X1 U23503 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20659), .ZN(
        P1_U3175) );
  AND2_X1 U23504 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20659), .ZN(
        P1_U3176) );
  AND2_X1 U23505 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20659), .ZN(
        P1_U3177) );
  AND2_X1 U23506 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20659), .ZN(
        P1_U3178) );
  AND2_X1 U23507 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20659), .ZN(
        P1_U3179) );
  AND2_X1 U23508 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20659), .ZN(
        P1_U3180) );
  AND2_X1 U23509 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20659), .ZN(
        P1_U3181) );
  AND2_X1 U23510 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20659), .ZN(
        P1_U3182) );
  AND2_X1 U23511 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20659), .ZN(
        P1_U3183) );
  AND2_X1 U23512 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20659), .ZN(
        P1_U3184) );
  AND2_X1 U23513 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20659), .ZN(
        P1_U3185) );
  AND2_X1 U23514 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20659), .ZN(P1_U3186) );
  AND2_X1 U23515 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20659), .ZN(P1_U3187) );
  AND2_X1 U23516 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20659), .ZN(P1_U3188) );
  AND2_X1 U23517 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20659), .ZN(P1_U3189) );
  AND2_X1 U23518 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20659), .ZN(P1_U3190) );
  AND2_X1 U23519 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20659), .ZN(P1_U3191) );
  AND2_X1 U23520 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20659), .ZN(P1_U3192) );
  AND2_X1 U23521 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20659), .ZN(P1_U3193) );
  NAND2_X1 U23522 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20593), .ZN(n20591) );
  INV_X1 U23523 ( .A(n20591), .ZN(n20589) );
  INV_X1 U23524 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20594) );
  NOR2_X1 U23525 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20586) );
  OAI22_X1 U23526 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20592), .B1(n20586), 
        .B2(n20585), .ZN(n20587) );
  NOR2_X1 U23527 ( .A1(n20594), .A2(n20587), .ZN(n20588) );
  OAI22_X1 U23528 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20589), .B1(n20715), 
        .B2(n20588), .ZN(P1_U3194) );
  OAI211_X1 U23529 ( .C1(NA), .C2(n20708), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20599), .ZN(n20590) );
  OAI211_X1 U23530 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20594), .A(HOLD), .B(
        n20590), .ZN(n20597) );
  OAI211_X1 U23531 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20592), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20591), .ZN(n20596) );
  OR4_X1 U23532 ( .A1(n20594), .A2(n20598), .A3(n20593), .A4(NA), .ZN(n20595)
         );
  OAI211_X1 U23533 ( .C1(n20598), .C2(n20597), .A(n20596), .B(n20595), .ZN(
        P1_U3196) );
  NAND2_X1 U23534 ( .A1(n20715), .A2(n20599), .ZN(n20646) );
  INV_X1 U23535 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20601) );
  NAND2_X1 U23536 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20715), .ZN(n20643) );
  OAI222_X1 U23537 ( .A1(n20646), .A2(n13514), .B1(n20601), .B2(n20715), .C1(
        n20600), .C2(n20643), .ZN(P1_U3197) );
  AOI22_X1 U23538 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20649), .ZN(n20602) );
  OAI21_X1 U23539 ( .B1(n13514), .B2(n20643), .A(n20602), .ZN(P1_U3198) );
  OAI222_X1 U23540 ( .A1(n20643), .A2(n13771), .B1(n20603), .B2(n20715), .C1(
        n20604), .C2(n20646), .ZN(P1_U3199) );
  INV_X1 U23541 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20605) );
  OAI222_X1 U23542 ( .A1(n20646), .A2(n20607), .B1(n20605), .B2(n20715), .C1(
        n20604), .C2(n20643), .ZN(P1_U3200) );
  AOI22_X1 U23543 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20649), .ZN(n20606) );
  OAI21_X1 U23544 ( .B1(n20607), .B2(n20643), .A(n20606), .ZN(P1_U3201) );
  INV_X1 U23545 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20609) );
  AOI22_X1 U23546 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20649), .ZN(n20608) );
  OAI21_X1 U23547 ( .B1(n20609), .B2(n20643), .A(n20608), .ZN(P1_U3202) );
  INV_X1 U23548 ( .A(n20643), .ZN(n20650) );
  AOI22_X1 U23549 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20650), .ZN(n20610) );
  OAI21_X1 U23550 ( .B1(n20612), .B2(n20646), .A(n20610), .ZN(P1_U3203) );
  AOI22_X1 U23551 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20649), .ZN(n20611) );
  OAI21_X1 U23552 ( .B1(n20612), .B2(n20643), .A(n20611), .ZN(P1_U3204) );
  AOI22_X1 U23553 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20649), .ZN(n20613) );
  OAI21_X1 U23554 ( .B1(n14036), .B2(n20643), .A(n20613), .ZN(P1_U3205) );
  AOI22_X1 U23555 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20650), .ZN(n20614) );
  OAI21_X1 U23556 ( .B1(n20616), .B2(n20646), .A(n20614), .ZN(P1_U3206) );
  INV_X1 U23557 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20615) );
  OAI222_X1 U23558 ( .A1(n20643), .A2(n20616), .B1(n20615), .B2(n20715), .C1(
        n20619), .C2(n20646), .ZN(P1_U3207) );
  INV_X1 U23559 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20618) );
  OAI222_X1 U23560 ( .A1(n20643), .A2(n20619), .B1(n20618), .B2(n20715), .C1(
        n20617), .C2(n20646), .ZN(P1_U3208) );
  AOI222_X1 U23561 ( .A1(n20650), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20636), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20649), .ZN(n20620) );
  INV_X1 U23562 ( .A(n20620), .ZN(P1_U3209) );
  AOI222_X1 U23563 ( .A1(n20650), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20636), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20649), .ZN(n20621) );
  INV_X1 U23564 ( .A(n20621), .ZN(P1_U3210) );
  INV_X1 U23565 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20622) );
  OAI222_X1 U23566 ( .A1(n20643), .A2(n20623), .B1(n20622), .B2(n20715), .C1(
        n20625), .C2(n20646), .ZN(P1_U3211) );
  AOI22_X1 U23567 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20649), .ZN(n20624) );
  OAI21_X1 U23568 ( .B1(n20625), .B2(n20643), .A(n20624), .ZN(P1_U3212) );
  AOI22_X1 U23569 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20650), .ZN(n20626) );
  OAI21_X1 U23570 ( .B1(n20628), .B2(n20646), .A(n20626), .ZN(P1_U3213) );
  INV_X1 U23571 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20627) );
  OAI222_X1 U23572 ( .A1(n20643), .A2(n20628), .B1(n20627), .B2(n20715), .C1(
        n20630), .C2(n20646), .ZN(P1_U3214) );
  AOI22_X1 U23573 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20649), .ZN(n20629) );
  OAI21_X1 U23574 ( .B1(n20630), .B2(n20643), .A(n20629), .ZN(P1_U3215) );
  AOI22_X1 U23575 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20712), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20650), .ZN(n20631) );
  OAI21_X1 U23576 ( .B1(n20839), .B2(n20646), .A(n20631), .ZN(P1_U3216) );
  INV_X1 U23577 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20632) );
  OAI222_X1 U23578 ( .A1(n20643), .A2(n20839), .B1(n20632), .B2(n20715), .C1(
        n20635), .C2(n20646), .ZN(P1_U3217) );
  INV_X1 U23579 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20634) );
  OAI222_X1 U23580 ( .A1(n20643), .A2(n20635), .B1(n20634), .B2(n20715), .C1(
        n20633), .C2(n20646), .ZN(P1_U3218) );
  AOI222_X1 U23581 ( .A1(n20650), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20636), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20649), .ZN(n20637) );
  INV_X1 U23582 ( .A(n20637), .ZN(P1_U3219) );
  AOI222_X1 U23583 ( .A1(n20650), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20712), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20649), .ZN(n20638) );
  INV_X1 U23584 ( .A(n20638), .ZN(P1_U3220) );
  INV_X1 U23585 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20639) );
  OAI222_X1 U23586 ( .A1(n20643), .A2(n20640), .B1(n20639), .B2(n20715), .C1(
        n14497), .C2(n20646), .ZN(P1_U3221) );
  INV_X1 U23587 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20641) );
  OAI222_X1 U23588 ( .A1(n20643), .A2(n14497), .B1(n20641), .B2(n20715), .C1(
        n20644), .C2(n20646), .ZN(P1_U3222) );
  AOI22_X1 U23589 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20649), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20712), .ZN(n20642) );
  OAI21_X1 U23590 ( .B1(n20644), .B2(n20643), .A(n20642), .ZN(P1_U3223) );
  AOI22_X1 U23591 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20650), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20712), .ZN(n20645) );
  OAI21_X1 U23592 ( .B1(n20647), .B2(n20646), .A(n20645), .ZN(P1_U3224) );
  AOI222_X1 U23593 ( .A1(n20649), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20712), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20650), .ZN(n20648) );
  INV_X1 U23594 ( .A(n20648), .ZN(P1_U3225) );
  AOI222_X1 U23595 ( .A1(n20650), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20712), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20649), .ZN(n20651) );
  INV_X1 U23596 ( .A(n20651), .ZN(P1_U3226) );
  INV_X1 U23597 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20652) );
  AOI22_X1 U23598 ( .A1(n20715), .A2(n20653), .B1(n20652), .B2(n20712), .ZN(
        P1_U3458) );
  INV_X1 U23599 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20693) );
  INV_X1 U23600 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20654) );
  AOI22_X1 U23601 ( .A1(n20715), .A2(n20693), .B1(n20654), .B2(n20712), .ZN(
        P1_U3459) );
  INV_X1 U23602 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20655) );
  AOI22_X1 U23603 ( .A1(n20715), .A2(n20656), .B1(n20655), .B2(n20712), .ZN(
        P1_U3460) );
  INV_X1 U23604 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20696) );
  INV_X1 U23605 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20657) );
  AOI22_X1 U23606 ( .A1(n20715), .A2(n20696), .B1(n20657), .B2(n20712), .ZN(
        P1_U3461) );
  INV_X1 U23607 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20660) );
  INV_X1 U23608 ( .A(n20661), .ZN(n20658) );
  AOI21_X1 U23609 ( .B1(n20660), .B2(n20659), .A(n20658), .ZN(P1_U3464) );
  OAI21_X1 U23610 ( .B1(n20663), .B2(n20662), .A(n20661), .ZN(P1_U3465) );
  INV_X1 U23611 ( .A(n20688), .ZN(n20691) );
  OR2_X1 U23612 ( .A1(n20665), .A2(n20664), .ZN(n20671) );
  INV_X1 U23613 ( .A(n20666), .ZN(n20667) );
  OAI22_X1 U23614 ( .A1(n11701), .A2(n20668), .B1(n20667), .B2(n20682), .ZN(
        n20670) );
  AOI211_X1 U23615 ( .C1(n20684), .C2(n20671), .A(n20670), .B(n20669), .ZN(
        n20672) );
  AOI22_X1 U23616 ( .A1(n20691), .A2(n20673), .B1(n20672), .B2(n20688), .ZN(
        P1_U3475) );
  NAND2_X1 U23617 ( .A1(n20675), .A2(n20674), .ZN(n20677) );
  OAI211_X1 U23618 ( .C1(n20682), .C2(n20678), .A(n20677), .B(n20676), .ZN(
        n20679) );
  INV_X1 U23619 ( .A(n20679), .ZN(n20680) );
  AOI22_X1 U23620 ( .A1(n20691), .A2(n20681), .B1(n20680), .B2(n20688), .ZN(
        P1_U3476) );
  INV_X1 U23621 ( .A(n20682), .ZN(n20686) );
  MUX2_X1 U23622 ( .A(n20684), .B(n20683), .S(n20010), .Z(n20685) );
  AOI21_X1 U23623 ( .B1(n20687), .B2(n20686), .A(n20685), .ZN(n20689) );
  AOI22_X1 U23624 ( .A1(n20691), .A2(n20690), .B1(n20689), .B2(n20688), .ZN(
        P1_U3477) );
  AOI211_X1 U23625 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20692) );
  AOI21_X1 U23626 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20692), .ZN(n20694) );
  AOI22_X1 U23627 ( .A1(n20698), .A2(n20694), .B1(n20693), .B2(n20695), .ZN(
        P1_U3481) );
  NOR2_X1 U23628 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20697) );
  AOI22_X1 U23629 ( .A1(n20698), .A2(n20697), .B1(n20696), .B2(n20695), .ZN(
        P1_U3482) );
  INV_X1 U23630 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20699) );
  AOI22_X1 U23631 ( .A1(n20715), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20699), 
        .B2(n20712), .ZN(P1_U3483) );
  AOI21_X1 U23632 ( .B1(n20701), .B2(n20771), .A(n20700), .ZN(n20704) );
  AOI22_X1 U23633 ( .A1(n20705), .A2(n20704), .B1(n20703), .B2(n20702), .ZN(
        n20711) );
  AOI211_X1 U23634 ( .C1(n20709), .C2(n20708), .A(n20707), .B(n20706), .ZN(
        n20710) );
  MUX2_X1 U23635 ( .A(n20711), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20710), 
        .Z(P1_U3485) );
  INV_X1 U23636 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20714) );
  AOI22_X1 U23637 ( .A1(n20715), .A2(n20714), .B1(n20713), .B2(n20712), .ZN(
        P1_U3486) );
  NAND2_X1 U23638 ( .A1(n18967), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n20718) );
  NAND2_X1 U23639 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n20716), .ZN(n20717) );
  OAI211_X1 U23640 ( .C1(n20720), .C2(n20719), .A(n20718), .B(n20717), .ZN(
        n20721) );
  INV_X1 U23641 ( .A(n20721), .ZN(n20886) );
  NAND4_X1 U23642 ( .A1(keyinput0), .A2(keyinput42), .A3(keyinput27), .A4(
        keyinput33), .ZN(n20725) );
  NAND4_X1 U23643 ( .A1(keyinput32), .A2(keyinput41), .A3(keyinput40), .A4(
        keyinput30), .ZN(n20724) );
  NAND4_X1 U23644 ( .A1(keyinput23), .A2(keyinput62), .A3(keyinput6), .A4(
        keyinput11), .ZN(n20723) );
  NAND4_X1 U23645 ( .A1(keyinput19), .A2(keyinput39), .A3(keyinput50), .A4(
        keyinput5), .ZN(n20722) );
  NOR4_X1 U23646 ( .A1(n20725), .A2(n20724), .A3(n20723), .A4(n20722), .ZN(
        n20884) );
  NAND3_X1 U23647 ( .A1(keyinput54), .A2(keyinput51), .A3(keyinput2), .ZN(
        n20745) );
  NOR2_X1 U23648 ( .A1(keyinput10), .A2(keyinput63), .ZN(n20729) );
  NAND4_X1 U23649 ( .A1(keyinput49), .A2(keyinput17), .A3(keyinput12), .A4(
        keyinput24), .ZN(n20727) );
  NAND2_X1 U23650 ( .A1(keyinput20), .A2(keyinput8), .ZN(n20726) );
  NOR4_X1 U23651 ( .A1(keyinput34), .A2(keyinput45), .A3(n20727), .A4(n20726), 
        .ZN(n20728) );
  NAND4_X1 U23652 ( .A1(keyinput35), .A2(keyinput56), .A3(n20729), .A4(n20728), 
        .ZN(n20744) );
  NOR3_X1 U23653 ( .A1(keyinput58), .A2(keyinput14), .A3(keyinput37), .ZN(
        n20742) );
  NAND2_X1 U23654 ( .A1(keyinput44), .A2(keyinput21), .ZN(n20733) );
  NOR3_X1 U23655 ( .A1(keyinput13), .A2(keyinput9), .A3(keyinput59), .ZN(
        n20731) );
  NOR3_X1 U23656 ( .A1(keyinput3), .A2(keyinput52), .A3(keyinput38), .ZN(
        n20730) );
  NAND4_X1 U23657 ( .A1(keyinput7), .A2(n20731), .A3(keyinput36), .A4(n20730), 
        .ZN(n20732) );
  NOR4_X1 U23658 ( .A1(keyinput26), .A2(keyinput48), .A3(n20733), .A4(n20732), 
        .ZN(n20741) );
  NAND3_X1 U23659 ( .A1(keyinput25), .A2(keyinput29), .A3(keyinput61), .ZN(
        n20739) );
  INV_X1 U23660 ( .A(keyinput60), .ZN(n20734) );
  NAND4_X1 U23661 ( .A1(keyinput31), .A2(keyinput18), .A3(keyinput28), .A4(
        n20734), .ZN(n20738) );
  NOR3_X1 U23662 ( .A1(keyinput47), .A2(keyinput15), .A3(keyinput22), .ZN(
        n20736) );
  INV_X1 U23663 ( .A(keyinput53), .ZN(n20846) );
  NOR3_X1 U23664 ( .A1(keyinput4), .A2(keyinput1), .A3(n20846), .ZN(n20735) );
  NAND4_X1 U23665 ( .A1(keyinput16), .A2(n20736), .A3(keyinput57), .A4(n20735), 
        .ZN(n20737) );
  NOR4_X1 U23666 ( .A1(keyinput46), .A2(n20739), .A3(n20738), .A4(n20737), 
        .ZN(n20740) );
  NAND4_X1 U23667 ( .A1(keyinput55), .A2(n20742), .A3(n20741), .A4(n20740), 
        .ZN(n20743) );
  NOR4_X1 U23668 ( .A1(keyinput43), .A2(n20745), .A3(n20744), .A4(n20743), 
        .ZN(n20883) );
  INV_X1 U23669 ( .A(keyinput0), .ZN(n20748) );
  INV_X1 U23670 ( .A(keyinput42), .ZN(n20747) );
  AOI22_X1 U23671 ( .A1(n20748), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20747), .ZN(n20746) );
  OAI221_X1 U23672 ( .B1(n20748), .B2(P3_ADDRESS_REG_4__SCAN_IN), .C1(n20747), 
        .C2(P3_UWORD_REG_12__SCAN_IN), .A(n20746), .ZN(n20760) );
  INV_X1 U23673 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n20751) );
  AOI22_X1 U23674 ( .A1(n20751), .A2(keyinput27), .B1(n20750), .B2(keyinput33), 
        .ZN(n20749) );
  OAI221_X1 U23675 ( .B1(n20751), .B2(keyinput27), .C1(n20750), .C2(keyinput33), .A(n20749), .ZN(n20759) );
  INV_X1 U23676 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n20753) );
  AOI22_X1 U23677 ( .A1(n11119), .A2(keyinput32), .B1(keyinput41), .B2(n20753), 
        .ZN(n20752) );
  OAI221_X1 U23678 ( .B1(n11119), .B2(keyinput32), .C1(n20753), .C2(keyinput41), .A(n20752), .ZN(n20758) );
  INV_X1 U23679 ( .A(keyinput30), .ZN(n20755) );
  AOI22_X1 U23680 ( .A1(n20756), .A2(keyinput40), .B1(
        P2_READREQUEST_REG_SCAN_IN), .B2(n20755), .ZN(n20754) );
  OAI221_X1 U23681 ( .B1(n20756), .B2(keyinput40), .C1(n20755), .C2(
        P2_READREQUEST_REG_SCAN_IN), .A(n20754), .ZN(n20757) );
  NOR4_X1 U23682 ( .A1(n20760), .A2(n20759), .A3(n20758), .A4(n20757), .ZN(
        n20813) );
  AOI22_X1 U23683 ( .A1(n20763), .A2(keyinput23), .B1(n20762), .B2(keyinput62), 
        .ZN(n20761) );
  OAI221_X1 U23684 ( .B1(n20763), .B2(keyinput23), .C1(n20762), .C2(keyinput62), .A(n20761), .ZN(n20775) );
  INV_X1 U23685 ( .A(keyinput11), .ZN(n20765) );
  AOI22_X1 U23686 ( .A1(n20766), .A2(keyinput6), .B1(P3_UWORD_REG_7__SCAN_IN), 
        .B2(n20765), .ZN(n20764) );
  OAI221_X1 U23687 ( .B1(n20766), .B2(keyinput6), .C1(n20765), .C2(
        P3_UWORD_REG_7__SCAN_IN), .A(n20764), .ZN(n20774) );
  AOI22_X1 U23688 ( .A1(n20768), .A2(keyinput19), .B1(n12979), .B2(keyinput39), 
        .ZN(n20767) );
  OAI221_X1 U23689 ( .B1(n20768), .B2(keyinput19), .C1(n12979), .C2(keyinput39), .A(n20767), .ZN(n20773) );
  INV_X1 U23690 ( .A(DATAI_3_), .ZN(n20770) );
  AOI22_X1 U23691 ( .A1(n20771), .A2(keyinput50), .B1(keyinput5), .B2(n20770), 
        .ZN(n20769) );
  OAI221_X1 U23692 ( .B1(n20771), .B2(keyinput50), .C1(n20770), .C2(keyinput5), 
        .A(n20769), .ZN(n20772) );
  NOR4_X1 U23693 ( .A1(n20775), .A2(n20774), .A3(n20773), .A4(n20772), .ZN(
        n20812) );
  INV_X1 U23694 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n20777) );
  AOI22_X1 U23695 ( .A1(n20778), .A2(keyinput7), .B1(n20777), .B2(keyinput13), 
        .ZN(n20776) );
  OAI221_X1 U23696 ( .B1(n20778), .B2(keyinput7), .C1(n20777), .C2(keyinput13), 
        .A(n20776), .ZN(n20783) );
  AOI22_X1 U23697 ( .A1(n20781), .A2(keyinput37), .B1(n20780), .B2(keyinput55), 
        .ZN(n20779) );
  OAI221_X1 U23698 ( .B1(n20781), .B2(keyinput37), .C1(n20780), .C2(keyinput55), .A(n20779), .ZN(n20782) );
  NOR2_X1 U23699 ( .A1(n20783), .A2(n20782), .ZN(n20793) );
  INV_X1 U23700 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20786) );
  AOI22_X1 U23701 ( .A1(n20786), .A2(keyinput58), .B1(keyinput14), .B2(n20785), 
        .ZN(n20784) );
  OAI221_X1 U23702 ( .B1(n20786), .B2(keyinput58), .C1(n20785), .C2(keyinput14), .A(n20784), .ZN(n20787) );
  INV_X1 U23703 ( .A(n20787), .ZN(n20792) );
  INV_X1 U23704 ( .A(keyinput59), .ZN(n20789) );
  INV_X1 U23705 ( .A(P3_LWORD_REG_7__SCAN_IN), .ZN(n20788) );
  XNOR2_X1 U23706 ( .A(n20789), .B(n20788), .ZN(n20791) );
  XNOR2_X1 U23707 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B(keyinput9), .ZN(
        n20790) );
  AND4_X1 U23708 ( .A1(n20793), .A2(n20792), .A3(n20791), .A4(n20790), .ZN(
        n20811) );
  INV_X1 U23709 ( .A(keyinput44), .ZN(n20795) );
  AOI22_X1 U23710 ( .A1(n20796), .A2(keyinput21), .B1(P3_LWORD_REG_10__SCAN_IN), .B2(n20795), .ZN(n20794) );
  OAI221_X1 U23711 ( .B1(n20796), .B2(keyinput21), .C1(n20795), .C2(
        P3_LWORD_REG_10__SCAN_IN), .A(n20794), .ZN(n20809) );
  INV_X1 U23712 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n20799) );
  AOI22_X1 U23713 ( .A1(n20799), .A2(keyinput26), .B1(n20798), .B2(keyinput48), 
        .ZN(n20797) );
  OAI221_X1 U23714 ( .B1(n20799), .B2(keyinput26), .C1(n20798), .C2(keyinput48), .A(n20797), .ZN(n20808) );
  INV_X1 U23715 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n20801) );
  AOI22_X1 U23716 ( .A1(n20802), .A2(keyinput3), .B1(keyinput52), .B2(n20801), 
        .ZN(n20800) );
  OAI221_X1 U23717 ( .B1(n20802), .B2(keyinput3), .C1(n20801), .C2(keyinput52), 
        .A(n20800), .ZN(n20807) );
  INV_X1 U23718 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n20805) );
  AOI22_X1 U23719 ( .A1(n20805), .A2(keyinput36), .B1(keyinput38), .B2(n20804), 
        .ZN(n20803) );
  OAI221_X1 U23720 ( .B1(n20805), .B2(keyinput36), .C1(n20804), .C2(keyinput38), .A(n20803), .ZN(n20806) );
  NOR4_X1 U23721 ( .A1(n20809), .A2(n20808), .A3(n20807), .A4(n20806), .ZN(
        n20810) );
  NAND4_X1 U23722 ( .A1(n20813), .A2(n20812), .A3(n20811), .A4(n20810), .ZN(
        n20882) );
  AOI22_X1 U23723 ( .A1(n20816), .A2(keyinput12), .B1(keyinput24), .B2(n20815), 
        .ZN(n20814) );
  OAI221_X1 U23724 ( .B1(n20816), .B2(keyinput12), .C1(n20815), .C2(keyinput24), .A(n20814), .ZN(n20829) );
  INV_X1 U23725 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n20819) );
  AOI22_X1 U23726 ( .A1(n20819), .A2(keyinput49), .B1(n20818), .B2(keyinput17), 
        .ZN(n20817) );
  OAI221_X1 U23727 ( .B1(n20819), .B2(keyinput49), .C1(n20818), .C2(keyinput17), .A(n20817), .ZN(n20828) );
  INV_X1 U23728 ( .A(keyinput8), .ZN(n20821) );
  AOI22_X1 U23729 ( .A1(n20822), .A2(keyinput34), .B1(
        P2_DATAWIDTH_REG_7__SCAN_IN), .B2(n20821), .ZN(n20820) );
  OAI221_X1 U23730 ( .B1(n20822), .B2(keyinput34), .C1(n20821), .C2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A(n20820), .ZN(n20827) );
  INV_X1 U23731 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n20824) );
  AOI22_X1 U23732 ( .A1(n20825), .A2(keyinput20), .B1(keyinput45), .B2(n20824), 
        .ZN(n20823) );
  OAI221_X1 U23733 ( .B1(n20825), .B2(keyinput20), .C1(n20824), .C2(keyinput45), .A(n20823), .ZN(n20826) );
  NOR4_X1 U23734 ( .A1(n20829), .A2(n20828), .A3(n20827), .A4(n20826), .ZN(
        n20880) );
  INV_X1 U23735 ( .A(keyinput51), .ZN(n20831) );
  AOI22_X1 U23736 ( .A1(n14792), .A2(keyinput2), .B1(P1_M_IO_N_REG_SCAN_IN), 
        .B2(n20831), .ZN(n20830) );
  OAI221_X1 U23737 ( .B1(n14792), .B2(keyinput2), .C1(n20831), .C2(
        P1_M_IO_N_REG_SCAN_IN), .A(n20830), .ZN(n20844) );
  INV_X1 U23738 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n20833) );
  AOI22_X1 U23739 ( .A1(n20834), .A2(keyinput43), .B1(n20833), .B2(keyinput54), 
        .ZN(n20832) );
  OAI221_X1 U23740 ( .B1(n20834), .B2(keyinput43), .C1(n20833), .C2(keyinput54), .A(n20832), .ZN(n20843) );
  INV_X1 U23741 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20837) );
  INV_X1 U23742 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20836) );
  AOI22_X1 U23743 ( .A1(n20837), .A2(keyinput10), .B1(n20836), .B2(keyinput63), 
        .ZN(n20835) );
  OAI221_X1 U23744 ( .B1(n20837), .B2(keyinput10), .C1(n20836), .C2(keyinput63), .A(n20835), .ZN(n20842) );
  AOI22_X1 U23745 ( .A1(n20840), .A2(keyinput35), .B1(keyinput56), .B2(n20839), 
        .ZN(n20838) );
  OAI221_X1 U23746 ( .B1(n20840), .B2(keyinput35), .C1(n20839), .C2(keyinput56), .A(n20838), .ZN(n20841) );
  NOR4_X1 U23747 ( .A1(n20844), .A2(n20843), .A3(n20842), .A4(n20841), .ZN(
        n20879) );
  INV_X1 U23748 ( .A(keyinput57), .ZN(n20847) );
  AOI22_X1 U23749 ( .A1(n20847), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20846), .ZN(n20845) );
  OAI221_X1 U23750 ( .B1(n20847), .B2(P2_DATAO_REG_6__SCAN_IN), .C1(n20846), 
        .C2(P3_LWORD_REG_1__SCAN_IN), .A(n20845), .ZN(n20860) );
  AOI22_X1 U23751 ( .A1(n20850), .A2(keyinput4), .B1(n20849), .B2(keyinput1), 
        .ZN(n20848) );
  OAI221_X1 U23752 ( .B1(n20850), .B2(keyinput4), .C1(n20849), .C2(keyinput1), 
        .A(n20848), .ZN(n20859) );
  INV_X1 U23753 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n20853) );
  AOI22_X1 U23754 ( .A1(n20853), .A2(keyinput18), .B1(n20852), .B2(keyinput28), 
        .ZN(n20851) );
  OAI221_X1 U23755 ( .B1(n20853), .B2(keyinput18), .C1(n20852), .C2(keyinput28), .A(n20851), .ZN(n20858) );
  INV_X1 U23756 ( .A(keyinput31), .ZN(n20855) );
  AOI22_X1 U23757 ( .A1(n20856), .A2(keyinput60), .B1(
        P2_DATAWIDTH_REG_25__SCAN_IN), .B2(n20855), .ZN(n20854) );
  OAI221_X1 U23758 ( .B1(n20856), .B2(keyinput60), .C1(n20855), .C2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A(n20854), .ZN(n20857) );
  NOR4_X1 U23759 ( .A1(n20860), .A2(n20859), .A3(n20858), .A4(n20857), .ZN(
        n20878) );
  INV_X1 U23760 ( .A(keyinput22), .ZN(n20862) );
  AOI22_X1 U23761 ( .A1(n20863), .A2(keyinput16), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n20862), .ZN(n20861) );
  OAI221_X1 U23762 ( .B1(n20863), .B2(keyinput16), .C1(n20862), .C2(
        P3_ADDRESS_REG_10__SCAN_IN), .A(n20861), .ZN(n20876) );
  INV_X1 U23763 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20865) );
  AOI22_X1 U23764 ( .A1(n20866), .A2(keyinput47), .B1(n20865), .B2(keyinput15), 
        .ZN(n20864) );
  OAI221_X1 U23765 ( .B1(n20866), .B2(keyinput47), .C1(n20865), .C2(keyinput15), .A(n20864), .ZN(n20875) );
  AOI22_X1 U23766 ( .A1(n20869), .A2(keyinput61), .B1(n20868), .B2(keyinput46), 
        .ZN(n20867) );
  OAI221_X1 U23767 ( .B1(n20869), .B2(keyinput61), .C1(n20868), .C2(keyinput46), .A(n20867), .ZN(n20874) );
  INV_X1 U23768 ( .A(keyinput29), .ZN(n20871) );
  AOI22_X1 U23769 ( .A1(n20872), .A2(keyinput25), .B1(P3_LWORD_REG_3__SCAN_IN), 
        .B2(n20871), .ZN(n20870) );
  OAI221_X1 U23770 ( .B1(n20872), .B2(keyinput25), .C1(n20871), .C2(
        P3_LWORD_REG_3__SCAN_IN), .A(n20870), .ZN(n20873) );
  NOR4_X1 U23771 ( .A1(n20876), .A2(n20875), .A3(n20874), .A4(n20873), .ZN(
        n20877) );
  NAND4_X1 U23772 ( .A1(n20880), .A2(n20879), .A3(n20878), .A4(n20877), .ZN(
        n20881) );
  AOI211_X1 U23773 ( .C1(n20884), .C2(n20883), .A(n20882), .B(n20881), .ZN(
        n20885) );
  XNOR2_X1 U23774 ( .A(n20886), .B(n20885), .ZN(P2_U2931) );
  INV_X1 U11131 ( .A(n17032), .ZN(n17999) );
  CLKBUF_X1 U11097 ( .A(n11496), .Z(n11371) );
  CLKBUF_X1 U11112 ( .A(n11419), .Z(n9610) );
  CLKBUF_X1 U11151 ( .A(n11309), .Z(n13409) );
  CLKBUF_X1 U11156 ( .A(n12623), .Z(n12693) );
  NAND2_X1 U11309 ( .A1(n10051), .A2(n10054), .ZN(n15007) );
  CLKBUF_X1 U11318 ( .A(n10270), .Z(n16940) );
  CLKBUF_X3 U11367 ( .A(n16754), .Z(n16871) );
  CLKBUF_X2 U11371 ( .A(n10611), .Z(n13188) );
  CLKBUF_X1 U11375 ( .A(n18419), .Z(n9629) );
  CLKBUF_X1 U11403 ( .A(n10577), .Z(n19028) );
  CLKBUF_X1 U11534 ( .A(n15049), .Z(n9612) );
  CLKBUF_X1 U12054 ( .A(n17611), .Z(n9632) );
  CLKBUF_X1 U12285 ( .A(n18614), .Z(n17194) );
endmodule

