

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040;

  INV_X4 U5095 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5096 ( .A(n6915), .ZN(n6901) );
  NAND2_X1 U5097 ( .A1(n6503), .A2(n5034), .ZN(n9819) );
  INV_X2 U5098 ( .A(n6831), .ZN(n6645) );
  INV_X1 U5100 ( .A(n6308), .ZN(n6274) );
  AND2_X1 U5102 ( .A1(n9746), .A2(n6770), .ZN(n6788) );
  AND2_X1 U5103 ( .A1(n6405), .A2(n8726), .ZN(n6508) );
  INV_X1 U5104 ( .A(n9819), .ZN(n9807) );
  NAND2_X1 U5105 ( .A1(n7950), .A2(n8198), .ZN(n10871) );
  AND2_X1 U5106 ( .A1(n6470), .A2(n6430), .ZN(n6915) );
  NAND3_X1 U5107 ( .A1(n5347), .A2(n5346), .A3(n10861), .ZN(n8006) );
  INV_X1 U5108 ( .A(n10781), .ZN(n10764) );
  OAI211_X1 U5109 ( .C1(n7286), .C2(n7446), .A(n5679), .B(n5678), .ZN(n10806)
         );
  NAND2_X1 U5110 ( .A1(n9698), .A2(n5031), .ZN(n5638) );
  NAND2_X1 U5111 ( .A1(n9095), .A2(n9100), .ZN(n9094) );
  OAI211_X1 U5112 ( .C1(n6503), .C2(n7259), .A(n6452), .B(n6451), .ZN(n7980)
         );
  CLKBUF_X1 U5114 ( .A(n6508), .Z(n5032) );
  BUF_X4 U5115 ( .A(n6508), .Z(n5033) );
  OAI22_X2 U5116 ( .A1(n6312), .A2(n6311), .B1(n6310), .B2(n6309), .ZN(n6338)
         );
  XNOR2_X2 U5117 ( .A(n5158), .B(n9669), .ZN(n6952) );
  XNOR2_X2 U5118 ( .A(n5591), .B(n5590), .ZN(n6363) );
  INV_X2 U5119 ( .A(n6918), .ZN(n6850) );
  NAND2_X2 U5120 ( .A1(n5797), .A2(n5796), .ZN(n10905) );
  AND2_X1 U5121 ( .A1(n5215), .A2(n5216), .ZN(n7149) );
  OAI21_X1 U5122 ( .B1(n5520), .B2(n5044), .A(n5519), .ZN(n9755) );
  NAND2_X1 U5123 ( .A1(n5520), .A2(n5517), .ZN(n5516) );
  NAND2_X1 U5124 ( .A1(n9187), .A2(n5054), .ZN(n9027) );
  NAND2_X1 U5125 ( .A1(n6788), .A2(n6789), .ZN(n9786) );
  NAND2_X1 U5126 ( .A1(n9079), .A2(n8655), .ZN(n9062) );
  NAND2_X1 U5127 ( .A1(n9094), .A2(n5058), .ZN(n9079) );
  INV_X1 U5128 ( .A(n5494), .ZN(n5489) );
  NAND2_X1 U5129 ( .A1(n7813), .A2(n7814), .ZN(n7812) );
  NAND2_X1 U5130 ( .A1(n8322), .A2(n8321), .ZN(n10968) );
  NAND2_X1 U5131 ( .A1(n7643), .A2(n6569), .ZN(n7813) );
  NAND2_X1 U5132 ( .A1(n7644), .A2(n7645), .ZN(n7643) );
  AND2_X1 U5133 ( .A1(n6525), .A2(n7569), .ZN(n6526) );
  NAND2_X1 U5134 ( .A1(n5813), .A2(n5812), .ZN(n8257) );
  NAND2_X2 U5135 ( .A1(n7841), .A2(n11014), .ZN(n11019) );
  NOR2_X1 U5136 ( .A1(n8903), .A2(n7513), .ZN(n7584) );
  OAI21_X1 U5137 ( .B1(n5855), .B2(n5457), .A(n5455), .ZN(n5890) );
  NAND2_X1 U5138 ( .A1(n5765), .A2(n5764), .ZN(n10879) );
  NAND4_X1 U5139 ( .A1(n5665), .A2(n5664), .A3(n5663), .A4(n5662), .ZN(n8898)
         );
  NAND2_X1 U5140 ( .A1(n5313), .A2(n5314), .ZN(n8903) );
  AND2_X2 U5141 ( .A1(n7857), .A2(n7858), .ZN(n6918) );
  NAND4_X2 U5142 ( .A1(n5600), .A2(n5599), .A3(n5598), .A4(n5597), .ZN(n8901)
         );
  NAND2_X1 U5143 ( .A1(n5431), .A2(n5430), .ZN(n10781) );
  INV_X1 U5144 ( .A(n8641), .ZN(n7609) );
  INV_X1 U5145 ( .A(n5207), .ZN(n10743) );
  OAI211_X1 U5146 ( .C1(n7189), .C2(n9819), .A(n6517), .B(n6516), .ZN(n5207)
         );
  INV_X1 U5147 ( .A(n10104), .ZN(n8625) );
  NAND2_X1 U5148 ( .A1(n8124), .A2(n10785), .ZN(n10024) );
  INV_X1 U5149 ( .A(n8124), .ZN(n10086) );
  NAND2_X2 U5150 ( .A1(n5578), .A2(n5579), .ZN(n6090) );
  OR2_X1 U5151 ( .A1(n5695), .A2(n7195), .ZN(n5323) );
  AND4_X1 U5152 ( .A1(n6501), .A2(n6500), .A3(n6499), .A4(n6498), .ZN(n6507)
         );
  NAND2_X1 U5153 ( .A1(n6976), .A2(n7433), .ZN(n7109) );
  OAI211_X1 U5154 ( .C1(n6503), .C2(n7244), .A(n6490), .B(n6489), .ZN(n7994)
         );
  CLKBUF_X3 U5155 ( .A(n6497), .Z(n9815) );
  NAND2_X1 U5156 ( .A1(n9916), .A2(n7822), .ZN(n7858) );
  XNOR2_X1 U5157 ( .A(n6422), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U5158 ( .A1(n6413), .A2(n8726), .ZN(n6497) );
  CLKBUF_X2 U5159 ( .A(n6831), .Z(n9813) );
  NAND2_X1 U5160 ( .A1(n6406), .A2(n6405), .ZN(n6831) );
  NAND2_X1 U5161 ( .A1(n6399), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6422) );
  INV_X1 U5162 ( .A(n6406), .ZN(n8726) );
  INV_X1 U5163 ( .A(n6405), .ZN(n6413) );
  XNOR2_X1 U5164 ( .A(n6403), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U5165 ( .A1(n6398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U5166 ( .A1(n7182), .A2(P1_U3084), .ZN(n8813) );
  BUF_X8 U5167 ( .A(n5650), .Z(n5034) );
  NOR2_X1 U5168 ( .A1(n6515), .A2(n6372), .ZN(n6559) );
  NOR2_X1 U5169 ( .A1(n6376), .A2(n6375), .ZN(n6377) );
  AND3_X1 U5170 ( .A1(n7288), .A2(n5357), .A3(n5614), .ZN(n5627) );
  INV_X2 U5171 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9620) );
  INV_X1 U5172 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6370) );
  INV_X1 U5173 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9640) );
  INV_X1 U5174 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5841) );
  NOR2_X1 U5175 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5561) );
  NOR2_X1 U5176 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5562) );
  NOR2_X1 U5177 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5563) );
  NOR2_X1 U5178 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5130) );
  NOR2_X1 U5179 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5129) );
  NOR2_X1 U5180 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5128) );
  NOR2_X1 U5181 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5127) );
  INV_X1 U5182 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9653) );
  INV_X2 U5183 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5184 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U5185 ( .A1(n5777), .A2(n9489), .ZN(n5836) );
  INV_X1 U5186 ( .A(n5031), .ZN(n5579) );
  AND2_X1 U5187 ( .A1(n5571), .A2(n5572), .ZN(n5495) );
  NOR2_X1 U5188 ( .A1(n10476), .A2(n10284), .ZN(n9918) );
  AND2_X1 U5189 ( .A1(n10476), .A2(n10284), .ZN(n9910) );
  AND2_X1 U5190 ( .A1(n5397), .A2(n6424), .ZN(n6385) );
  NOR2_X1 U5191 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5397) );
  AND2_X1 U5192 ( .A1(n6377), .A2(n5543), .ZN(n5544) );
  AND2_X1 U5193 ( .A1(n5545), .A2(n5547), .ZN(n5543) );
  INV_X1 U5194 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5545) );
  INV_X1 U5195 ( .A(n11030), .ZN(n10275) );
  AND2_X1 U5196 ( .A1(n11030), .A2(n10272), .ZN(n10273) );
  INV_X1 U5197 ( .A(n5650), .ZN(n7182) );
  INV_X1 U5198 ( .A(n5136), .ZN(n5135) );
  NAND2_X1 U5199 ( .A1(n5279), .A2(n5277), .ZN(n7087) );
  AOI21_X1 U5200 ( .B1(n5280), .B2(n5283), .A(n5278), .ZN(n5277) );
  INV_X1 U5201 ( .A(n7083), .ZN(n5278) );
  OR2_X1 U5202 ( .A1(n7035), .A2(n5321), .ZN(n7039) );
  AND2_X1 U5203 ( .A1(n5292), .A2(n5443), .ZN(n5290) );
  AND2_X1 U5204 ( .A1(n7025), .A2(n7020), .ZN(n5443) );
  OAI21_X1 U5205 ( .B1(n9148), .B2(n8598), .A(n6303), .ZN(n6333) );
  OR2_X1 U5206 ( .A1(n9167), .A2(n8879), .ZN(n6295) );
  NAND2_X1 U5207 ( .A1(n5245), .A2(n5045), .ZN(n5244) );
  NAND2_X1 U5208 ( .A1(n5248), .A2(n5249), .ZN(n5245) );
  OR2_X1 U5209 ( .A1(n9199), .A2(n9102), .ZN(n8655) );
  NOR2_X1 U5210 ( .A1(n5826), .A2(n5378), .ZN(n5374) );
  INV_X1 U5211 ( .A(n5739), .ZN(n5378) );
  NAND2_X1 U5212 ( .A1(n8250), .A2(n5334), .ZN(n8416) );
  AND2_X1 U5213 ( .A1(n5040), .A2(n10964), .ZN(n5334) );
  INV_X1 U5214 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5589) );
  AND2_X1 U5215 ( .A1(n5221), .A2(n5220), .ZN(n5219) );
  INV_X1 U5216 ( .A(n9795), .ZN(n5220) );
  OR2_X1 U5217 ( .A1(n5512), .A2(n5036), .ZN(n5221) );
  OR2_X1 U5218 ( .A1(n10493), .A2(n10344), .ZN(n9921) );
  NAND2_X1 U5219 ( .A1(n10493), .A2(n10344), .ZN(n10296) );
  NOR2_X1 U5220 ( .A1(n8786), .A2(n5420), .ZN(n5419) );
  INV_X1 U5221 ( .A(n8783), .ZN(n5420) );
  OR2_X1 U5222 ( .A1(n10557), .A2(n10453), .ZN(n9972) );
  OR2_X1 U5223 ( .A1(n10543), .A2(n10556), .ZN(n9976) );
  OR2_X1 U5224 ( .A1(n5559), .A2(n8486), .ZN(n5406) );
  OR2_X1 U5225 ( .A1(n5559), .A2(n5408), .ZN(n5407) );
  NAND2_X1 U5226 ( .A1(n7899), .A2(n10770), .ZN(n9894) );
  NAND2_X1 U5227 ( .A1(n9886), .A2(n9885), .ZN(n5199) );
  AOI21_X1 U5228 ( .B1(n8086), .B2(n7855), .A(n5558), .ZN(n7904) );
  NOR2_X1 U5229 ( .A1(n7854), .A2(n10035), .ZN(n5558) );
  NAND2_X1 U5230 ( .A1(n6030), .A2(n6029), .ZN(n6050) );
  NAND2_X1 U5231 ( .A1(n6028), .A2(n6027), .ZN(n6030) );
  NAND2_X1 U5232 ( .A1(n5984), .A2(n5983), .ZN(n5993) );
  NAND2_X1 U5233 ( .A1(n5982), .A2(n5981), .ZN(n5984) );
  OAI21_X1 U5234 ( .B1(n5966), .B2(n5965), .A(n5967), .ZN(n5982) );
  NAND2_X1 U5235 ( .A1(n5893), .A2(n5892), .ZN(n5911) );
  NAND2_X1 U5236 ( .A1(n5890), .A2(n5889), .ZN(n5893) );
  NAND2_X1 U5237 ( .A1(n5874), .A2(n5856), .ZN(n5289) );
  NAND2_X1 U5238 ( .A1(n5837), .A2(n5836), .ZN(n5855) );
  AND2_X1 U5239 ( .A1(n5759), .A2(n5758), .ZN(n5768) );
  NAND2_X1 U5240 ( .A1(n7039), .A2(n5319), .ZN(n8730) );
  OR2_X1 U5241 ( .A1(n5321), .A2(n5320), .ZN(n5319) );
  INV_X1 U5242 ( .A(n8699), .ZN(n5320) );
  XNOR2_X1 U5243 ( .A(n7087), .B(n7085), .ZN(n8719) );
  INV_X1 U5244 ( .A(n5314), .ZN(n5310) );
  OR2_X1 U5245 ( .A1(n7091), .A2(n7090), .ZN(n8831) );
  OAI21_X1 U5246 ( .B1(n7961), .B2(n5297), .A(n5294), .ZN(n8096) );
  XNOR2_X1 U5247 ( .A(n7606), .B(n7109), .ZN(n8636) );
  AND2_X1 U5248 ( .A1(n5583), .A2(n5582), .ZN(n5313) );
  OR2_X1 U5249 ( .A1(n6090), .A2(n7779), .ZN(n5582) );
  NAND2_X1 U5250 ( .A1(n9000), .A2(n9137), .ZN(n5380) );
  NAND2_X1 U5251 ( .A1(n5359), .A2(n5362), .ZN(n5267) );
  NAND2_X1 U5252 ( .A1(n5359), .A2(n5269), .ZN(n5268) );
  NAND2_X1 U5253 ( .A1(n5363), .A2(n6314), .ZN(n5362) );
  OR2_X1 U5254 ( .A1(n9178), .A2(n9040), .ZN(n5109) );
  NAND2_X1 U5255 ( .A1(n9009), .A2(n9019), .ZN(n5110) );
  NAND2_X1 U5256 ( .A1(n5266), .A2(n5265), .ZN(n9136) );
  OR2_X1 U5257 ( .A1(n9223), .A2(n6247), .ZN(n5265) );
  NAND2_X1 U5258 ( .A1(n5256), .A2(n5254), .ZN(n5266) );
  AND2_X1 U5259 ( .A1(n5257), .A2(n5255), .ZN(n5254) );
  NOR2_X1 U5260 ( .A1(n9223), .A2(n5327), .ZN(n5326) );
  INV_X1 U5261 ( .A(n5328), .ZN(n5327) );
  OR2_X1 U5262 ( .A1(n8387), .A2(n5259), .ZN(n5256) );
  NAND2_X1 U5263 ( .A1(n6243), .A2(n5262), .ZN(n5259) );
  NAND2_X1 U5264 ( .A1(n9690), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5574) );
  NOR2_X1 U5265 ( .A1(n5318), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U5266 ( .A1(n5570), .A2(n5507), .ZN(n5506) );
  INV_X1 U5267 ( .A(n5509), .ZN(n5507) );
  OR2_X1 U5268 ( .A1(n10493), .A2(n10298), .ZN(n8788) );
  OR2_X1 U5269 ( .A1(n10500), .A2(n10358), .ZN(n8787) );
  NOR2_X1 U5270 ( .A1(n10341), .A2(n5417), .ZN(n5416) );
  INV_X1 U5271 ( .A(n8785), .ZN(n5417) );
  NAND2_X1 U5272 ( .A1(n10352), .A2(n10001), .ZN(n8803) );
  OR2_X1 U5273 ( .A1(n10508), .A2(n10387), .ZN(n10351) );
  NAND2_X1 U5274 ( .A1(n8157), .A2(n8156), .ZN(n8427) );
  INV_X1 U5275 ( .A(n6503), .ZN(n7243) );
  NAND2_X1 U5276 ( .A1(n8794), .A2(n8793), .ZN(n10476) );
  OR2_X1 U5277 ( .A1(n6381), .A2(n5385), .ZN(n6402) );
  INV_X1 U5278 ( .A(n5386), .ZN(n5385) );
  AND2_X1 U5279 ( .A1(n6385), .A2(n6378), .ZN(n6391) );
  AND2_X1 U5280 ( .A1(n5676), .A2(n5691), .ZN(n5466) );
  INV_X1 U5281 ( .A(n8790), .ZN(n10297) );
  AND2_X1 U5282 ( .A1(n9824), .A2(n9823), .ZN(n11030) );
  OR2_X1 U5283 ( .A1(n9820), .A2(n9819), .ZN(n9824) );
  NAND2_X1 U5284 ( .A1(n9931), .A2(n9930), .ZN(n9934) );
  AOI21_X1 U5285 ( .B1(n5141), .B2(n5078), .A(n5138), .ZN(n5137) );
  INV_X1 U5286 ( .A(n9971), .ZN(n5138) );
  OAI21_X1 U5287 ( .B1(n5148), .B2(n5147), .A(n5050), .ZN(n9951) );
  AOI21_X1 U5288 ( .B1(n5137), .B2(n5139), .A(n10549), .ZN(n5136) );
  INV_X1 U5289 ( .A(n5141), .ZN(n5139) );
  INV_X1 U5290 ( .A(n5137), .ZN(n5133) );
  NAND2_X1 U5291 ( .A1(n5134), .A2(n5131), .ZN(n5140) );
  INV_X1 U5292 ( .A(n5758), .ZN(n5476) );
  AND2_X1 U5293 ( .A1(n5748), .A2(n5755), .ZN(n5752) );
  OAI21_X1 U5294 ( .B1(n5153), .B2(n5152), .A(n5063), .ZN(n10013) );
  NAND2_X1 U5295 ( .A1(n10009), .A2(n10010), .ZN(n5152) );
  NOR2_X1 U5296 ( .A1(n5928), .A2(n5454), .ZN(n5453) );
  INV_X1 U5297 ( .A(n5913), .ZN(n5454) );
  INV_X1 U5298 ( .A(n8148), .ZN(n5297) );
  AND2_X1 U5299 ( .A1(n7016), .A2(n5295), .ZN(n5294) );
  NAND2_X1 U5300 ( .A1(n8148), .A2(n5296), .ZN(n5295) );
  INV_X1 U5301 ( .A(n7010), .ZN(n5296) );
  NAND2_X1 U5302 ( .A1(n5973), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5987) );
  INV_X1 U5303 ( .A(n5974), .ZN(n5973) );
  NAND2_X1 U5304 ( .A1(n8214), .A2(n5102), .ZN(n8400) );
  NAND2_X1 U5305 ( .A1(n8221), .A2(n8383), .ZN(n5102) );
  AND2_X1 U5306 ( .A1(n6301), .A2(n6302), .ZN(n8660) );
  OR2_X1 U5307 ( .A1(n9162), .A2(n8817), .ZN(n6176) );
  NAND2_X1 U5308 ( .A1(n8987), .A2(n5342), .ZN(n5341) );
  OR2_X1 U5309 ( .A1(n9054), .A2(n9034), .ZN(n6280) );
  OR2_X1 U5310 ( .A1(n5987), .A2(n9318), .ZN(n6004) );
  NAND2_X1 U5311 ( .A1(n5252), .A2(n6263), .ZN(n5250) );
  NAND2_X1 U5312 ( .A1(n6329), .A2(n5253), .ZN(n5252) );
  NAND2_X1 U5313 ( .A1(n9112), .A2(n6258), .ZN(n5253) );
  NAND2_X1 U5314 ( .A1(n6263), .A2(n6258), .ZN(n5251) );
  OR2_X1 U5315 ( .A1(n9199), .A2(n9204), .ZN(n5333) );
  OR2_X1 U5316 ( .A1(n9223), .A2(n9138), .ZN(n8649) );
  INV_X1 U5317 ( .A(n8517), .ZN(n5500) );
  NOR2_X1 U5318 ( .A1(n9229), .A2(n8760), .ZN(n5328) );
  OR2_X1 U5319 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  NAND2_X1 U5320 ( .A1(n7787), .A2(n5698), .ZN(n5369) );
  OR2_X1 U5321 ( .A1(n8898), .A2(n10820), .ZN(n5681) );
  OR2_X1 U5322 ( .A1(n8900), .A2(n7739), .ZN(n7716) );
  OR2_X1 U5323 ( .A1(n7949), .A2(n10868), .ZN(n8198) );
  OAI21_X1 U5324 ( .B1(n6167), .B2(n5317), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6355) );
  OAI22_X1 U5325 ( .A1(n7831), .A2(n6920), .B1(n7850), .B2(n6854), .ZN(n6491)
         );
  NAND4_X1 U5326 ( .A1(n6370), .A2(n9620), .A3(n5511), .A4(n6461), .ZN(n6515)
         );
  INV_X1 U5327 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5511) );
  OR2_X1 U5328 ( .A1(n10481), .A2(n8790), .ZN(n9825) );
  OR2_X1 U5329 ( .A1(n10500), .A2(n10321), .ZN(n10008) );
  NOR2_X1 U5330 ( .A1(n10419), .A2(n5192), .ZN(n5191) );
  INV_X1 U5331 ( .A(n9984), .ZN(n5192) );
  NOR2_X1 U5332 ( .A1(n10399), .A2(n5189), .ZN(n5188) );
  INV_X1 U5333 ( .A(n9862), .ZN(n5189) );
  NAND2_X1 U5334 ( .A1(n10443), .A2(n5191), .ZN(n5190) );
  OR2_X1 U5335 ( .A1(n10518), .A2(n10385), .ZN(n9863) );
  AOI21_X1 U5336 ( .B1(n5424), .B2(n10457), .A(n5059), .ZN(n5423) );
  OR2_X1 U5337 ( .A1(n8485), .A2(n5078), .ZN(n8489) );
  OR2_X1 U5338 ( .A1(n8569), .A2(n10555), .ZN(n9969) );
  NAND2_X1 U5339 ( .A1(n10922), .A2(n8431), .ZN(n5396) );
  OR2_X1 U5340 ( .A1(n10917), .A2(n8428), .ZN(n9952) );
  INV_X1 U5341 ( .A(n9942), .ZN(n5183) );
  INV_X1 U5342 ( .A(n9944), .ZN(n5182) );
  NAND2_X1 U5343 ( .A1(n5199), .A2(n5197), .ZN(n8062) );
  NOR2_X1 U5344 ( .A1(n5198), .A2(n9844), .ZN(n5197) );
  OAI21_X1 U5345 ( .B1(n10916), .B2(n5404), .A(n5403), .ZN(n10550) );
  AOI21_X1 U5346 ( .B1(n5407), .B2(n5406), .A(n5085), .ZN(n5403) );
  NAND2_X1 U5347 ( .A1(n6733), .A2(n6732), .ZN(n10557) );
  NOR2_X1 U5348 ( .A1(n8473), .A2(n9831), .ZN(n8500) );
  INV_X1 U5349 ( .A(n5474), .ZN(n6119) );
  OAI21_X1 U5350 ( .B1(n6084), .B2(n5470), .A(n5468), .ZN(n5474) );
  INV_X1 U5351 ( .A(n5469), .ZN(n5468) );
  OAI21_X1 U5352 ( .B1(n5472), .B2(n5470), .A(n6117), .ZN(n5469) );
  NAND2_X1 U5353 ( .A1(n5463), .A2(n5460), .ZN(n6082) );
  INV_X1 U5354 ( .A(n5461), .ZN(n5460) );
  OAI21_X1 U5355 ( .B1(n6066), .B2(n5462), .A(n6067), .ZN(n5461) );
  NAND2_X1 U5356 ( .A1(n5998), .A2(n5997), .ZN(n6014) );
  AND2_X1 U5357 ( .A1(n5983), .A2(n5970), .ZN(n5981) );
  NAND2_X1 U5358 ( .A1(n5945), .A2(n5944), .ZN(n5966) );
  NAND2_X1 U5359 ( .A1(n5942), .A2(n5941), .ZN(n5945) );
  XNOR2_X1 U5360 ( .A(n5891), .B(SI_15_), .ZN(n5888) );
  INV_X1 U5361 ( .A(n5458), .ZN(n5457) );
  AOI21_X1 U5362 ( .B1(n5458), .B2(n5456), .A(n5060), .ZN(n5455) );
  NOR2_X1 U5363 ( .A1(n5874), .A2(n5459), .ZN(n5458) );
  XNOR2_X1 U5364 ( .A(n5774), .B(n5773), .ZN(n5792) );
  NAND2_X1 U5365 ( .A1(n6056), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U5366 ( .A1(n8725), .A2(n7088), .ZN(n7091) );
  NAND2_X1 U5367 ( .A1(n8685), .A2(n5440), .ZN(n7961) );
  AND2_X1 U5368 ( .A1(n7009), .A2(n7004), .ZN(n5440) );
  NAND2_X1 U5369 ( .A1(n6996), .A2(n10728), .ZN(n5307) );
  AND2_X1 U5370 ( .A1(n7042), .A2(n8730), .ZN(n7043) );
  XNOR2_X1 U5371 ( .A(n8744), .B(n7103), .ZN(n8754) );
  AOI21_X1 U5372 ( .B1(n6164), .B2(n6169), .A(n6170), .ZN(n6342) );
  INV_X1 U5373 ( .A(n6333), .ZN(n6169) );
  AND2_X1 U5374 ( .A1(n5584), .A2(n5581), .ZN(n5314) );
  XNOR2_X1 U5375 ( .A(n8400), .B(n8394), .ZN(n8216) );
  NAND2_X1 U5376 ( .A1(n8216), .A2(n8418), .ZN(n8402) );
  INV_X1 U5377 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5569) );
  OR2_X1 U5378 ( .A1(n9820), .A2(n6137), .ZN(n6139) );
  AOI21_X1 U5379 ( .B1(n5490), .B2(n5488), .A(n8969), .ZN(n5487) );
  INV_X1 U5380 ( .A(n5492), .ZN(n5488) );
  INV_X1 U5381 ( .A(n8992), .ZN(n8817) );
  NAND2_X1 U5382 ( .A1(n8988), .A2(n6295), .ZN(n8975) );
  NOR2_X1 U5383 ( .A1(n8989), .A2(n5493), .ZN(n5492) );
  NAND2_X1 U5384 ( .A1(n8990), .A2(n8989), .ZN(n8988) );
  NOR2_X1 U5385 ( .A1(n9011), .A2(n9173), .ZN(n9002) );
  AND2_X1 U5386 ( .A1(n6295), .A2(n6296), .ZN(n8989) );
  NAND2_X1 U5387 ( .A1(n8999), .A2(n8658), .ZN(n5494) );
  INV_X1 U5388 ( .A(n5364), .ZN(n5363) );
  OAI21_X1 U5389 ( .B1(n9019), .B2(n6288), .A(n6178), .ZN(n5364) );
  INV_X1 U5390 ( .A(n9019), .ZN(n5365) );
  NOR2_X1 U5391 ( .A1(n9051), .A2(n9182), .ZN(n9010) );
  NAND2_X1 U5392 ( .A1(n9027), .A2(n8657), .ZN(n9009) );
  AOI21_X1 U5393 ( .B1(n5035), .B2(n9072), .A(n5372), .ZN(n5371) );
  INV_X1 U5394 ( .A(n6281), .ZN(n5372) );
  NOR2_X1 U5395 ( .A1(n9194), .A2(n9089), .ZN(n8656) );
  NAND2_X1 U5396 ( .A1(n5243), .A2(n9061), .ZN(n5373) );
  INV_X1 U5397 ( .A(n5373), .ZN(n9069) );
  INV_X1 U5398 ( .A(n5250), .ZN(n5249) );
  INV_X1 U5399 ( .A(n5251), .ZN(n5247) );
  OR2_X1 U5400 ( .A1(n9099), .A2(n8653), .ZN(n5554) );
  OR2_X1 U5401 ( .A1(n9211), .A2(n8652), .ZN(n6258) );
  NAND2_X1 U5402 ( .A1(n9209), .A2(n5108), .ZN(n9095) );
  NAND2_X1 U5403 ( .A1(n9140), .A2(n9211), .ZN(n5108) );
  AOI21_X1 U5404 ( .B1(n9136), .B2(n9125), .A(n5939), .ZN(n9108) );
  AND2_X1 U5405 ( .A1(n8417), .A2(n5091), .ZN(n9127) );
  OAI21_X1 U5406 ( .B1(n8412), .B2(n5497), .A(n5496), .ZN(n8537) );
  NAND2_X1 U5407 ( .A1(n8510), .A2(n5505), .ZN(n5497) );
  NAND2_X1 U5408 ( .A1(n5499), .A2(n5505), .ZN(n5496) );
  NAND2_X1 U5409 ( .A1(n9229), .A2(n8887), .ZN(n5505) );
  NAND2_X1 U5410 ( .A1(n5258), .A2(n6243), .ZN(n5257) );
  INV_X1 U5411 ( .A(n5260), .ZN(n5258) );
  AOI21_X1 U5412 ( .B1(n5261), .B2(n5262), .A(n5066), .ZN(n5260) );
  INV_X1 U5413 ( .A(n5504), .ZN(n5503) );
  OAI22_X1 U5414 ( .A1(n8514), .A2(n8411), .B1(n8760), .B2(n8888), .ZN(n5504)
         );
  OR2_X1 U5415 ( .A1(n8760), .A2(n8687), .ZN(n8509) );
  AND2_X1 U5416 ( .A1(n6243), .A2(n6242), .ZN(n8517) );
  NOR2_X1 U5417 ( .A1(n8416), .A2(n8744), .ZN(n8417) );
  NAND2_X1 U5418 ( .A1(n5846), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5862) );
  INV_X1 U5419 ( .A(n5847), .ZN(n5846) );
  AND2_X1 U5420 ( .A1(n6237), .A2(n6236), .ZN(n8382) );
  NAND2_X1 U5421 ( .A1(n10968), .A2(n5084), .ZN(n8381) );
  INV_X1 U5422 ( .A(n8889), .ZN(n8747) );
  NAND2_X1 U5423 ( .A1(n5376), .A2(n5375), .ZN(n8387) );
  NOR2_X1 U5424 ( .A1(n5377), .A2(n5062), .ZN(n5375) );
  NAND2_X1 U5425 ( .A1(n10905), .A2(n8892), .ZN(n5483) );
  NOR2_X1 U5426 ( .A1(n8614), .A2(n5481), .ZN(n5480) );
  INV_X1 U5427 ( .A(n5483), .ZN(n5481) );
  AND2_X1 U5428 ( .A1(n6225), .A2(n6222), .ZN(n8614) );
  NAND2_X1 U5429 ( .A1(n8270), .A2(n8269), .ZN(n8319) );
  NAND2_X1 U5430 ( .A1(n7940), .A2(n5739), .ZN(n8191) );
  INV_X1 U5431 ( .A(n5695), .ZN(n5953) );
  INV_X1 U5432 ( .A(n7286), .ZN(n5952) );
  INV_X1 U5433 ( .A(n9070), .ZN(n10798) );
  NAND2_X1 U5434 ( .A1(n5495), .A2(n5055), .ZN(n5318) );
  INV_X1 U5435 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U5436 ( .A1(n6355), .A2(n5589), .ZN(n6357) );
  INV_X1 U5437 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6147) );
  XNOR2_X1 U5438 ( .A(n5444), .B(P2_IR_REG_20__SCAN_IN), .ZN(n7588) );
  NAND2_X1 U5439 ( .A1(n5445), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U5440 ( .A1(n6166), .A2(n6165), .ZN(n5445) );
  NOR2_X1 U5441 ( .A1(n5568), .A2(n5567), .ZN(n5324) );
  INV_X1 U5442 ( .A(n5205), .ZN(n5203) );
  AOI21_X1 U5443 ( .B1(n5219), .B2(n5036), .A(n5089), .ZN(n5218) );
  AND2_X1 U5444 ( .A1(n6663), .A2(n6408), .ZN(n6682) );
  INV_X1 U5445 ( .A(n5514), .ZN(n5513) );
  OAI21_X1 U5446 ( .B1(n9754), .B2(n5515), .A(n5522), .ZN(n5514) );
  NAND2_X1 U5447 ( .A1(n5044), .A2(n5519), .ZN(n5515) );
  AND2_X1 U5448 ( .A1(n5224), .A2(n5538), .ZN(n5223) );
  INV_X1 U5449 ( .A(n5539), .ZN(n5538) );
  AOI22_X1 U5450 ( .A1(n7834), .A2(n6915), .B1(n5207), .B2(n6434), .ZN(n6528)
         );
  XNOR2_X1 U5451 ( .A(n6506), .B(n6918), .ZN(n6522) );
  OAI22_X1 U5452 ( .A1(n6507), .A2(n6920), .B1(n10719), .B2(n6854), .ZN(n6506)
         );
  OAI22_X1 U5453 ( .A1(n6507), .A2(n6901), .B1(n10719), .B2(n6920), .ZN(n6520)
         );
  NAND2_X1 U5454 ( .A1(n7812), .A2(n6593), .ZN(n8029) );
  NOR2_X1 U5455 ( .A1(n5525), .A2(n5524), .ZN(n5523) );
  INV_X1 U5456 ( .A(n6620), .ZN(n5525) );
  INV_X1 U5457 ( .A(n8018), .ZN(n5524) );
  NOR2_X1 U5458 ( .A1(n6468), .A2(n5548), .ZN(n7497) );
  AOI21_X1 U5459 ( .B1(n8014), .B2(n6434), .A(n6462), .ZN(n6463) );
  NOR2_X1 U5460 ( .A1(n6639), .A2(n8231), .ZN(n5204) );
  INV_X1 U5461 ( .A(n6623), .ZN(n5202) );
  NOR2_X1 U5462 ( .A1(n6552), .A2(n6551), .ZN(n6570) );
  NOR2_X1 U5463 ( .A1(n9754), .A2(n5518), .ZN(n5517) );
  INV_X1 U5464 ( .A(n5519), .ZN(n5518) );
  NOR2_X1 U5465 ( .A1(n10647), .A2(n10646), .ZN(n10645) );
  NOR2_X1 U5466 ( .A1(n7687), .A2(n7686), .ZN(n7868) );
  NOR2_X1 U5467 ( .A1(n7868), .A2(n5177), .ZN(n7872) );
  AND2_X1 U5468 ( .A1(n7869), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5177) );
  OR2_X1 U5469 ( .A1(n7872), .A2(n7871), .ZN(n5176) );
  NOR2_X1 U5470 ( .A1(n10188), .A2(n5174), .ZN(n10195) );
  AND2_X1 U5471 ( .A1(n10189), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5174) );
  OR2_X1 U5472 ( .A1(n10190), .A2(n8499), .ZN(n5173) );
  AOI21_X1 U5473 ( .B1(n8803), .B2(n5390), .A(n5387), .ZN(n10283) );
  AND2_X1 U5474 ( .A1(n8805), .A2(n9872), .ZN(n5390) );
  NAND2_X1 U5475 ( .A1(n5388), .A2(n9919), .ZN(n5387) );
  NAND2_X1 U5476 ( .A1(n8805), .A2(n5389), .ZN(n5388) );
  NAND2_X1 U5477 ( .A1(n5409), .A2(n5413), .ZN(n10313) );
  INV_X1 U5478 ( .A(n5414), .ZN(n5413) );
  OAI21_X1 U5479 ( .B1(n5416), .B2(n5415), .A(n10316), .ZN(n5414) );
  NAND2_X1 U5480 ( .A1(n9921), .A2(n10296), .ZN(n10316) );
  AND4_X1 U5481 ( .A1(n6882), .A2(n6881), .A3(n6880), .A4(n6879), .ZN(n10344)
         );
  AND2_X1 U5482 ( .A1(n10008), .A2(n10007), .ZN(n10341) );
  OR2_X1 U5483 ( .A1(n10376), .A2(n8802), .ZN(n10352) );
  NAND2_X1 U5484 ( .A1(n5427), .A2(n5426), .ZN(n10382) );
  AOI21_X1 U5485 ( .B1(n5428), .B2(n9986), .A(n5056), .ZN(n5426) );
  NOR2_X1 U5486 ( .A1(n10427), .A2(n10518), .ZN(n10409) );
  NAND2_X1 U5487 ( .A1(n9863), .A2(n9988), .ZN(n10399) );
  AND2_X1 U5488 ( .A1(n10399), .A2(n5074), .ZN(n5428) );
  AND2_X1 U5489 ( .A1(n10054), .A2(n5043), .ZN(n5424) );
  NAND2_X1 U5490 ( .A1(n10548), .A2(n8571), .ZN(n10456) );
  OR2_X1 U5491 ( .A1(n10456), .A2(n10457), .ZN(n5425) );
  AND2_X1 U5492 ( .A1(n9976), .A2(n9975), .ZN(n10457) );
  INV_X1 U5493 ( .A(n5406), .ZN(n5404) );
  INV_X1 U5494 ( .A(n5407), .ZN(n5402) );
  INV_X1 U5495 ( .A(n5393), .ZN(n5392) );
  OAI21_X1 U5496 ( .B1(n8431), .B2(n5394), .A(n8493), .ZN(n5393) );
  AND2_X1 U5497 ( .A1(n9969), .A2(n9970), .ZN(n10052) );
  NAND2_X1 U5498 ( .A1(n6682), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6701) );
  OR2_X1 U5499 ( .A1(n6701), .A2(n6700), .ZN(n6719) );
  AOI21_X1 U5500 ( .B1(n8427), .B2(n8426), .A(n8425), .ZN(n10914) );
  NAND2_X1 U5501 ( .A1(n10914), .A2(n10913), .ZN(n10916) );
  AND2_X1 U5502 ( .A1(n8044), .A2(n5184), .ZN(n5421) );
  NAND2_X1 U5503 ( .A1(n6570), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6596) );
  AND4_X1 U5504 ( .A1(n6630), .A2(n6629), .A3(n6628), .A4(n6627), .ZN(n8160)
         );
  OAI21_X1 U5505 ( .B1(n10040), .B2(n7901), .A(n5124), .ZN(n7903) );
  OR2_X1 U5506 ( .A1(n10765), .A2(n7902), .ZN(n7905) );
  NAND2_X1 U5507 ( .A1(n9928), .A2(n9933), .ZN(n10042) );
  NAND2_X1 U5508 ( .A1(n7836), .A2(n9922), .ZN(n9925) );
  NOR2_X1 U5509 ( .A1(n10760), .A2(n10781), .ZN(n10762) );
  NAND2_X1 U5510 ( .A1(n7985), .A2(n9839), .ZN(n9886) );
  NAND2_X1 U5511 ( .A1(n7847), .A2(n9836), .ZN(n7848) );
  XNOR2_X1 U5512 ( .A(n10107), .B(n7980), .ZN(n10039) );
  AND2_X1 U5513 ( .A1(n6952), .A2(n10033), .ZN(n10769) );
  AND2_X1 U5514 ( .A1(n10291), .A2(n10290), .ZN(n10482) );
  NAND2_X1 U5515 ( .A1(n6755), .A2(n6754), .ZN(n10543) );
  INV_X1 U5516 ( .A(n10827), .ZN(n11029) );
  AND2_X1 U5517 ( .A1(n6927), .A2(n6928), .ZN(n10587) );
  XNOR2_X1 U5518 ( .A(n6160), .B(n6159), .ZN(n9808) );
  AND2_X1 U5519 ( .A1(n6120), .A2(n6132), .ZN(n6121) );
  OR2_X1 U5520 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  NAND2_X1 U5521 ( .A1(n6121), .A2(SI_29_), .ZN(n6133) );
  NAND2_X1 U5522 ( .A1(n6119), .A2(n6118), .ZN(n6132) );
  AOI21_X1 U5523 ( .B1(n6132), .B2(n9471), .A(n6135), .ZN(n5448) );
  INV_X1 U5524 ( .A(n6132), .ZN(n5449) );
  INV_X1 U5525 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9668) );
  INV_X1 U5526 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9669) );
  XNOR2_X1 U5527 ( .A(n6114), .B(n6113), .ZN(n8545) );
  NAND2_X1 U5528 ( .A1(n5467), .A2(n6099), .ZN(n6114) );
  NAND2_X1 U5529 ( .A1(n6084), .A2(n5472), .ZN(n5467) );
  NAND3_X1 U5530 ( .A1(n5544), .A2(n6380), .A3(n6576), .ZN(n6381) );
  XNOR2_X1 U5531 ( .A(n6082), .B(n6081), .ZN(n8445) );
  AND2_X1 U5532 ( .A1(n6377), .A2(n5547), .ZN(n5546) );
  AND2_X1 U5533 ( .A1(n5544), .A2(n6576), .ZN(n6388) );
  OAI21_X1 U5534 ( .B1(n6050), .B2(n6049), .A(n6048), .ZN(n6065) );
  OAI211_X1 U5535 ( .C1(n5855), .C2(n5289), .A(n5286), .B(n5284), .ZN(n7236)
         );
  INV_X1 U5536 ( .A(n5287), .ZN(n5286) );
  OAI21_X1 U5537 ( .B1(n5557), .B2(n5289), .A(n5288), .ZN(n5287) );
  XNOR2_X1 U5538 ( .A(n5793), .B(n5792), .ZN(n7229) );
  AND2_X1 U5539 ( .A1(n5791), .A2(n5805), .ZN(n5793) );
  XNOR2_X1 U5540 ( .A(n5235), .B(n5807), .ZN(n7223) );
  NAND2_X1 U5541 ( .A1(n5831), .A2(n5804), .ZN(n5235) );
  NAND2_X1 U5542 ( .A1(n5751), .A2(n5749), .ZN(n5730) );
  XNOR2_X1 U5543 ( .A(n5719), .B(n9499), .ZN(n5717) );
  XNOR2_X1 U5544 ( .A(n5693), .B(n9503), .ZN(n5691) );
  NAND2_X1 U5545 ( .A1(n5675), .A2(n5674), .ZN(n5676) );
  NAND2_X1 U5546 ( .A1(n5234), .A2(n5619), .ZN(n5630) );
  NAND2_X1 U5547 ( .A1(n8685), .A2(n7004), .ZN(n7962) );
  NAND2_X1 U5548 ( .A1(n6086), .A2(n6085), .ZN(n9167) );
  NAND2_X1 U5549 ( .A1(n5308), .A2(n8648), .ZN(n10728) );
  AND2_X1 U5550 ( .A1(n10729), .A2(n6986), .ZN(n5308) );
  OAI21_X1 U5551 ( .B1(n8528), .B2(n8526), .A(n8525), .ZN(n8561) );
  NAND2_X1 U5552 ( .A1(n5342), .A2(n10727), .ZN(n5439) );
  NAND2_X1 U5553 ( .A1(n6979), .A2(n6978), .ZN(n8639) );
  NAND2_X1 U5554 ( .A1(n7049), .A2(n8693), .ZN(n8698) );
  NAND2_X1 U5555 ( .A1(n5273), .A2(n5270), .ZN(n8858) );
  INV_X1 U5556 ( .A(n5271), .ZN(n5270) );
  OAI21_X1 U5557 ( .B1(n5272), .B2(n5276), .A(n8559), .ZN(n5271) );
  INV_X1 U5558 ( .A(n9075), .ZN(n9034) );
  NAND2_X1 U5559 ( .A1(n6096), .A2(n6095), .ZN(n9000) );
  OR2_X1 U5560 ( .A1(n6090), .A2(n7756), .ZN(n5612) );
  OR2_X1 U5561 ( .A1(n5819), .A2(n7306), .ZN(n5611) );
  OR2_X1 U5562 ( .A1(n6090), .A2(n7704), .ZN(n5599) );
  NAND2_X1 U5563 ( .A1(n5637), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5598) );
  OR2_X1 U5564 ( .A1(n5819), .A2(n5595), .ZN(n5600) );
  NAND2_X1 U5565 ( .A1(n7417), .A2(n7418), .ZN(n7447) );
  NOR2_X1 U5566 ( .A1(n7490), .A2(n7489), .ZN(n7488) );
  NOR2_X1 U5567 ( .A1(n7666), .A2(n7667), .ZN(n7767) );
  INV_X1 U5568 ( .A(n8076), .ZN(n10846) );
  NAND2_X1 U5569 ( .A1(n6433), .A2(n6432), .ZN(n10508) );
  AOI21_X1 U5570 ( .B1(n10275), .B2(n10274), .A(n10273), .ZN(n11034) );
  XNOR2_X1 U5571 ( .A(n5120), .B(n5119), .ZN(n10480) );
  INV_X1 U5572 ( .A(n10062), .ZN(n5119) );
  INV_X1 U5573 ( .A(n8795), .ZN(n5120) );
  NAND2_X1 U5574 ( .A1(n6859), .A2(n6858), .ZN(n10348) );
  AOI21_X1 U5575 ( .B1(n5157), .B2(n10024), .A(n9926), .ZN(n5156) );
  NAND2_X1 U5576 ( .A1(n9925), .A2(n10020), .ZN(n5155) );
  OAI21_X1 U5577 ( .B1(n10766), .B2(n9924), .A(n9923), .ZN(n5157) );
  NAND2_X1 U5578 ( .A1(n9939), .A2(n9940), .ZN(n5149) );
  AOI21_X1 U5579 ( .B1(n9936), .B2(n10020), .A(n10044), .ZN(n5150) );
  NAND2_X1 U5580 ( .A1(n9935), .A2(n10024), .ZN(n5151) );
  NAND2_X1 U5581 ( .A1(n10047), .A2(n9943), .ZN(n5147) );
  AND2_X1 U5582 ( .A1(n9968), .A2(n10052), .ZN(n5141) );
  AND2_X1 U5583 ( .A1(n5132), .A2(n5069), .ZN(n5131) );
  NAND2_X1 U5584 ( .A1(n5136), .A2(n5133), .ZN(n5132) );
  AOI21_X1 U5585 ( .B1(n10003), .B2(n10002), .A(n5154), .ZN(n5153) );
  NAND2_X1 U5586 ( .A1(n10006), .A2(n10341), .ZN(n5154) );
  NAND2_X1 U5587 ( .A1(n5294), .A2(n5297), .ZN(n5292) );
  OR2_X1 U5588 ( .A1(n8594), .A2(n8885), .ZN(n6301) );
  AOI21_X1 U5589 ( .B1(n5250), .B2(n5251), .A(n5064), .ZN(n5248) );
  NOR2_X1 U5590 ( .A1(n8099), .A2(n5241), .ZN(n5240) );
  INV_X1 U5591 ( .A(n5812), .ZN(n5241) );
  NOR2_X1 U5592 ( .A1(n8257), .A2(n10905), .ZN(n5335) );
  INV_X1 U5593 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5400) );
  NAND2_X1 U5594 ( .A1(n5471), .A2(n6099), .ZN(n5470) );
  INV_X1 U5595 ( .A(n6113), .ZN(n5471) );
  NAND2_X1 U5596 ( .A1(n6049), .A2(n6048), .ZN(n5462) );
  NOR2_X1 U5597 ( .A1(n6066), .A2(n5465), .ZN(n5464) );
  INV_X1 U5598 ( .A(n6048), .ZN(n5465) );
  INV_X1 U5599 ( .A(n5557), .ZN(n5456) );
  AND3_X1 U5600 ( .A1(n5306), .A2(n5829), .A3(n5830), .ZN(n5305) );
  INV_X1 U5601 ( .A(n5767), .ZN(n5475) );
  AND2_X1 U5602 ( .A1(n5832), .A2(n5828), .ZN(n5835) );
  OAI21_X1 U5603 ( .B1(n5034), .B2(n5300), .A(n5299), .ZN(n5774) );
  NAND2_X1 U5604 ( .A1(n5034), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n5299) );
  AND2_X1 U5605 ( .A1(n5804), .A2(n5806), .ZN(n5830) );
  NOR2_X1 U5606 ( .A1(n5552), .A2(n5551), .ZN(n5758) );
  AND2_X1 U5607 ( .A1(n8740), .A2(n5071), .ZN(n5321) );
  NOR2_X1 U5608 ( .A1(n8594), .A2(n5341), .ZN(n5340) );
  AOI21_X1 U5609 ( .B1(n5363), .B2(n5361), .A(n5360), .ZN(n5359) );
  INV_X1 U5610 ( .A(n6313), .ZN(n5360) );
  NOR2_X1 U5611 ( .A1(n5365), .A2(n5366), .ZN(n5361) );
  INV_X1 U5612 ( .A(n8991), .ZN(n8658) );
  NOR2_X1 U5613 ( .A1(n5333), .A2(n9194), .ZN(n5331) );
  INV_X1 U5614 ( .A(n8536), .ZN(n5255) );
  OR2_X1 U5615 ( .A1(n9216), .A2(n8651), .ZN(n6254) );
  INV_X1 U5616 ( .A(n5871), .ZN(n5261) );
  INV_X1 U5617 ( .A(n8509), .ZN(n5263) );
  NAND2_X1 U5618 ( .A1(n10949), .A2(n8703), .ZN(n5482) );
  AND2_X1 U5619 ( .A1(n8269), .A2(n5482), .ZN(n5479) );
  NAND2_X1 U5620 ( .A1(n6219), .A2(n5242), .ZN(n8274) );
  NAND2_X1 U5621 ( .A1(n6216), .A2(n6219), .ZN(n5242) );
  OR2_X1 U5622 ( .A1(n5766), .A2(n10879), .ZN(n8242) );
  NAND2_X1 U5623 ( .A1(n8250), .A2(n5335), .ZN(n8604) );
  NAND2_X1 U5624 ( .A1(n8250), .A2(n10896), .ZN(n8280) );
  NOR2_X1 U5625 ( .A1(n8198), .A2(n10879), .ZN(n8250) );
  NOR2_X1 U5626 ( .A1(n10802), .A2(n10806), .ZN(n7792) );
  NAND2_X1 U5627 ( .A1(n5569), .A2(n5510), .ZN(n5509) );
  INV_X1 U5628 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5510) );
  INV_X1 U5629 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5566) );
  OR3_X1 U5630 ( .A1(n5781), .A2(P2_IR_REG_9__SCAN_IN), .A3(
        P2_IR_REG_10__SCAN_IN), .ZN(n5794) );
  OR2_X1 U5631 ( .A1(n5763), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5781) );
  INV_X1 U5632 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5709) );
  INV_X1 U5633 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5232) );
  INV_X1 U5634 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5230) );
  INV_X1 U5635 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5231) );
  OAI21_X1 U5636 ( .B1(n5526), .B2(n5213), .A(n5080), .ZN(n5212) );
  INV_X1 U5637 ( .A(n9776), .ZN(n5213) );
  NOR2_X1 U5638 ( .A1(n9765), .A2(n5535), .ZN(n5534) );
  INV_X1 U5639 ( .A(n6807), .ZN(n5535) );
  OAI21_X1 U5640 ( .B1(n5540), .B2(n5542), .A(n6751), .ZN(n5539) );
  AND2_X1 U5641 ( .A1(n5536), .A2(n5228), .ZN(n5227) );
  INV_X1 U5642 ( .A(n5540), .ZN(n5536) );
  NAND2_X1 U5643 ( .A1(n5227), .A2(n5229), .ZN(n5224) );
  NOR2_X1 U5644 ( .A1(n8448), .A2(n8449), .ZN(n5229) );
  AND2_X1 U5645 ( .A1(n6810), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6825) );
  AND2_X1 U5646 ( .A1(n10271), .A2(n10090), .ZN(n10031) );
  INV_X1 U5647 ( .A(n8804), .ZN(n5389) );
  INV_X1 U5648 ( .A(n8787), .ZN(n5415) );
  NOR2_X1 U5649 ( .A1(n5415), .A2(n5411), .ZN(n5410) );
  INV_X1 U5650 ( .A(n5419), .ZN(n5411) );
  NOR2_X1 U5651 ( .A1(n10368), .A2(n10348), .ZN(n5344) );
  NOR2_X1 U5652 ( .A1(n6796), .A2(n9713), .ZN(n6810) );
  NAND2_X1 U5653 ( .A1(n5355), .A2(n10442), .ZN(n5354) );
  OR2_X1 U5654 ( .A1(n6778), .A2(n6777), .ZN(n6796) );
  NOR2_X1 U5655 ( .A1(n10538), .A2(n10543), .ZN(n5355) );
  INV_X1 U5656 ( .A(n5395), .ZN(n5394) );
  AND2_X1 U5657 ( .A1(n8430), .A2(n9952), .ZN(n5395) );
  NAND2_X1 U5658 ( .A1(n10049), .A2(n8429), .ZN(n5408) );
  NAND2_X1 U5659 ( .A1(n8047), .A2(n9942), .ZN(n8048) );
  NAND2_X1 U5660 ( .A1(n10102), .A2(n10861), .ZN(n9938) );
  INV_X1 U5661 ( .A(n10760), .ZN(n5347) );
  AND2_X1 U5662 ( .A1(n5345), .A2(n10846), .ZN(n5346) );
  INV_X1 U5663 ( .A(n5348), .ZN(n5345) );
  INV_X1 U5664 ( .A(n7902), .ZN(n5124) );
  NAND2_X1 U5665 ( .A1(n7899), .A2(n10764), .ZN(n5348) );
  NAND2_X1 U5666 ( .A1(n8053), .A2(n5039), .ZN(n8473) );
  NOR2_X1 U5667 ( .A1(n6100), .A2(n5473), .ZN(n5472) );
  INV_X1 U5668 ( .A(n6083), .ZN(n5473) );
  INV_X1 U5669 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9657) );
  AOI21_X1 U5670 ( .B1(n5912), .B2(n5453), .A(n5088), .ZN(n5452) );
  NAND2_X1 U5671 ( .A1(n5872), .A2(n5459), .ZN(n5288) );
  AND2_X1 U5672 ( .A1(n5557), .A2(n5872), .ZN(n5285) );
  AND2_X1 U5673 ( .A1(n5805), .A2(n5775), .ZN(n5833) );
  AND2_X1 U5674 ( .A1(n5775), .A2(n5298), .ZN(n5828) );
  INV_X1 U5675 ( .A(n5792), .ZN(n5298) );
  NAND2_X1 U5676 ( .A1(n5836), .A2(n5779), .ZN(n5827) );
  OR2_X1 U5677 ( .A1(n5768), .A2(n5767), .ZN(n5831) );
  NAND2_X1 U5678 ( .A1(n5760), .A2(n9490), .ZN(n5804) );
  OAI211_X1 U5679 ( .C1(n5677), .C2(n5239), .A(n5717), .B(n5238), .ZN(n5751)
         );
  INV_X1 U5680 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9404) );
  OAI21_X1 U5681 ( .B1(n5034), .B2(n5652), .A(n5651), .ZN(n5669) );
  NAND2_X1 U5682 ( .A1(n5034), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5651) );
  INV_X1 U5683 ( .A(SI_1_), .ZN(n9510) );
  NAND2_X1 U5684 ( .A1(n5682), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5703) );
  NOR2_X1 U5685 ( .A1(n5436), .A2(n5435), .ZN(n5434) );
  INV_X1 U5686 ( .A(n8846), .ZN(n5435) );
  INV_X1 U5687 ( .A(n7098), .ZN(n5438) );
  NAND2_X1 U5688 ( .A1(n5701), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5724) );
  INV_X1 U5689 ( .A(n5703), .ZN(n5701) );
  NAND2_X1 U5690 ( .A1(n6034), .A2(n6033), .ZN(n6057) );
  INV_X1 U5691 ( .A(n6036), .ZN(n6034) );
  INV_X1 U5692 ( .A(n5041), .ZN(n5276) );
  NAND2_X1 U5693 ( .A1(n8526), .A2(n8525), .ZN(n5272) );
  NOR2_X1 U5694 ( .A1(n5276), .A2(n5275), .ZN(n5274) );
  AND2_X1 U5695 ( .A1(n5441), .A2(n5281), .ZN(n5280) );
  NAND2_X1 U5696 ( .A1(n8822), .A2(n5282), .ZN(n5281) );
  AND2_X1 U5697 ( .A1(n7082), .A2(n7076), .ZN(n5441) );
  INV_X1 U5698 ( .A(n7071), .ZN(n5282) );
  INV_X1 U5699 ( .A(n8822), .ZN(n5283) );
  NAND2_X1 U5700 ( .A1(n5065), .A2(n8832), .ZN(n8833) );
  AND2_X1 U5701 ( .A1(n7654), .A2(n7653), .ZN(n7656) );
  AND2_X1 U5702 ( .A1(n7656), .A2(n7655), .ZN(n7763) );
  NOR2_X1 U5703 ( .A1(n7767), .A2(n5101), .ZN(n7771) );
  AND2_X1 U5704 ( .A1(n7768), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U5705 ( .A1(n7771), .A2(n7770), .ZN(n7929) );
  NAND2_X1 U5706 ( .A1(n8403), .A2(n8402), .ZN(n8406) );
  OR2_X1 U5707 ( .A1(n8917), .A2(n8916), .ZN(n5105) );
  AND2_X1 U5708 ( .A1(n9002), .A2(n5337), .ZN(n8963) );
  AND2_X1 U5709 ( .A1(n5340), .A2(n5338), .ZN(n5337) );
  INV_X1 U5710 ( .A(n5341), .ZN(n5339) );
  NAND2_X1 U5711 ( .A1(n9002), .A2(n8987), .ZN(n8981) );
  AND2_X1 U5712 ( .A1(n6088), .A2(n6074), .ZN(n9003) );
  NAND2_X1 U5713 ( .A1(n9010), .A2(n9017), .ZN(n9011) );
  NAND2_X1 U5714 ( .A1(n6020), .A2(n6019), .ZN(n9054) );
  OR2_X1 U5715 ( .A1(n9117), .A2(n5330), .ZN(n9051) );
  NAND2_X1 U5716 ( .A1(n9057), .A2(n5331), .ZN(n5330) );
  NOR2_X1 U5717 ( .A1(n9117), .A2(n5329), .ZN(n9063) );
  INV_X1 U5718 ( .A(n5331), .ZN(n5329) );
  INV_X1 U5719 ( .A(n5960), .ZN(n5958) );
  OR2_X1 U5720 ( .A1(n5933), .A2(n5932), .ZN(n5960) );
  AOI21_X1 U5721 ( .B1(n9126), .B2(n9135), .A(n5107), .ZN(n9113) );
  NOR2_X1 U5722 ( .A1(n9216), .A2(n9109), .ZN(n5107) );
  NAND2_X1 U5723 ( .A1(n6254), .A2(n6253), .ZN(n9135) );
  NAND2_X1 U5724 ( .A1(n8650), .A2(n8649), .ZN(n9126) );
  NAND2_X1 U5725 ( .A1(n5919), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5933) );
  INV_X1 U5726 ( .A(n5920), .ZN(n5919) );
  NAND2_X1 U5727 ( .A1(n8537), .A2(n8536), .ZN(n8650) );
  NAND2_X1 U5728 ( .A1(n8417), .A2(n10999), .ZN(n8518) );
  AND2_X1 U5729 ( .A1(n5264), .A2(n6237), .ZN(n8511) );
  NAND2_X1 U5730 ( .A1(n8387), .A2(n5871), .ZN(n5264) );
  OR2_X1 U5731 ( .A1(n5862), .A2(n9520), .ZN(n5881) );
  INV_X1 U5732 ( .A(n8888), .ZN(n8687) );
  NAND2_X1 U5733 ( .A1(n5111), .A2(n5477), .ZN(n8322) );
  NAND2_X1 U5734 ( .A1(n5478), .A2(n5482), .ZN(n5477) );
  NAND2_X1 U5735 ( .A1(n8270), .A2(n5479), .ZN(n5111) );
  INV_X1 U5736 ( .A(n5480), .ZN(n5478) );
  AND2_X1 U5737 ( .A1(n5376), .A2(n5825), .ZN(n8315) );
  NAND2_X1 U5738 ( .A1(n5784), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5847) );
  OR2_X1 U5739 ( .A1(n5818), .A2(n7172), .ZN(n5799) );
  OR2_X1 U5740 ( .A1(n5816), .A2(n5815), .ZN(n5818) );
  INV_X1 U5741 ( .A(n5242), .ZN(n8264) );
  NAND2_X1 U5742 ( .A1(n5723), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5741) );
  INV_X1 U5743 ( .A(n5724), .ZN(n5723) );
  NAND2_X1 U5744 ( .A1(n5740), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5816) );
  INV_X1 U5745 ( .A(n5741), .ZN(n5740) );
  OR2_X1 U5746 ( .A1(n8191), .A2(n8190), .ZN(n8273) );
  NAND2_X1 U5747 ( .A1(n7942), .A2(n5738), .ZN(n7940) );
  NAND2_X1 U5748 ( .A1(n5369), .A2(n5700), .ZN(n7880) );
  NAND2_X1 U5749 ( .A1(n5369), .A2(n5367), .ZN(n7942) );
  NOR2_X1 U5750 ( .A1(n7889), .A2(n5368), .ZN(n5367) );
  INV_X1 U5751 ( .A(n5700), .ZN(n5368) );
  NAND2_X1 U5752 ( .A1(n10795), .A2(n5681), .ZN(n7787) );
  NAND2_X1 U5753 ( .A1(n6320), .A2(n7884), .ZN(n7804) );
  NAND2_X1 U5754 ( .A1(n5325), .A2(n10752), .ZN(n10802) );
  NAND2_X1 U5755 ( .A1(n7716), .A2(n6190), .ZN(n7613) );
  NOR2_X1 U5756 ( .A1(n7752), .A2(n8641), .ZN(n7753) );
  INV_X1 U5757 ( .A(n7745), .ZN(n5356) );
  NAND2_X1 U5758 ( .A1(n5356), .A2(n7748), .ZN(n7747) );
  AND2_X1 U5759 ( .A1(n8903), .A2(n7783), .ZN(n7607) );
  NAND2_X1 U5760 ( .A1(n6032), .A2(n6031), .ZN(n9182) );
  AND2_X1 U5761 ( .A1(n7428), .A2(n7427), .ZN(n10904) );
  OAI21_X1 U5762 ( .B1(n5899), .B2(n5509), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5950) );
  INV_X1 U5763 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5357) );
  OAI22_X1 U5764 ( .A1(n5210), .A2(n5208), .B1(n5212), .B2(n5214), .ZN(n6857)
         );
  AND2_X1 U5765 ( .A1(n5527), .A2(n9776), .ZN(n5214) );
  NAND2_X1 U5766 ( .A1(n9788), .A2(n5209), .ZN(n5208) );
  INV_X1 U5767 ( .A(n5212), .ZN(n5209) );
  INV_X1 U5768 ( .A(n5534), .ZN(n5533) );
  AOI21_X1 U5769 ( .B1(n5534), .B2(n5532), .A(n5531), .ZN(n5530) );
  INV_X1 U5770 ( .A(n9766), .ZN(n5531) );
  INV_X1 U5771 ( .A(n9711), .ZN(n5532) );
  NAND2_X1 U5772 ( .A1(n9737), .A2(n5541), .ZN(n5540) );
  NAND2_X1 U5773 ( .A1(n8547), .A2(n8551), .ZN(n5541) );
  OR2_X1 U5774 ( .A1(n8547), .A2(n8551), .ZN(n5542) );
  NAND2_X1 U5775 ( .A1(n6544), .A2(n6548), .ZN(n7633) );
  NAND2_X1 U5776 ( .A1(n6856), .A2(n5521), .ZN(n5519) );
  INV_X1 U5777 ( .A(n6857), .ZN(n5520) );
  NAND2_X1 U5778 ( .A1(n5207), .A2(n6470), .ZN(n5206) );
  OR2_X1 U5779 ( .A1(n6806), .A2(n6805), .ZN(n6807) );
  NAND2_X1 U5780 ( .A1(n9710), .A2(n9711), .ZN(n9709) );
  AOI21_X1 U5781 ( .B1(n5527), .B2(n5533), .A(n5097), .ZN(n5526) );
  AND2_X1 U5782 ( .A1(n5530), .A2(n5528), .ZN(n5527) );
  INV_X1 U5783 ( .A(n9718), .ZN(n5528) );
  NAND2_X1 U5784 ( .A1(n9784), .A2(n9788), .ZN(n9710) );
  AND2_X1 U5785 ( .A1(n5513), .A2(n5073), .ZN(n5512) );
  NAND2_X1 U5786 ( .A1(n6713), .A2(n6712), .ZN(n8548) );
  NAND2_X1 U5787 ( .A1(n5225), .A2(n8449), .ZN(n6713) );
  NAND2_X1 U5788 ( .A1(n8548), .A2(n8547), .ZN(n9738) );
  NAND2_X1 U5789 ( .A1(n5144), .A2(n10022), .ZN(n5143) );
  AND4_X1 U5790 ( .A1(n6602), .A2(n6601), .A3(n6600), .A4(n6599), .ZN(n7909)
         );
  NAND2_X1 U5791 ( .A1(n6645), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6446) );
  INV_X1 U5792 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6371) );
  OR2_X1 U5793 ( .A1(n10645), .A2(n5081), .ZN(n7362) );
  OAI22_X1 U5794 ( .A1(n7362), .A2(n7363), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n7361), .ZN(n7364) );
  OR2_X1 U5795 ( .A1(n10660), .A2(n10659), .ZN(n5160) );
  OR3_X1 U5796 ( .A1(n6631), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n6640) );
  AND2_X1 U5797 ( .A1(n5176), .A2(n5175), .ZN(n8182) );
  NAND2_X1 U5798 ( .A1(n8179), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5175) );
  AND2_X1 U5799 ( .A1(n5067), .A2(n5173), .ZN(n10199) );
  AND2_X1 U5800 ( .A1(n9825), .A2(n10015), .ZN(n10282) );
  NAND2_X1 U5801 ( .A1(n10325), .A2(n10306), .ZN(n10303) );
  NAND2_X1 U5802 ( .A1(n10319), .A2(n10296), .ZN(n5196) );
  NAND2_X1 U5803 ( .A1(n10315), .A2(n8804), .ZN(n10319) );
  AND4_X1 U5804 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n10322)
         );
  AND2_X1 U5805 ( .A1(n6860), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6862) );
  AND2_X1 U5806 ( .A1(n6862), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U5807 ( .A1(n5344), .A2(n5343), .ZN(n10334) );
  INV_X1 U5808 ( .A(n5344), .ZN(n10349) );
  AND2_X1 U5809 ( .A1(n10409), .A2(n10394), .ZN(n10388) );
  NAND2_X1 U5810 ( .A1(n10388), .A2(n10374), .ZN(n10368) );
  INV_X1 U5811 ( .A(n5186), .ZN(n5185) );
  OAI21_X1 U5812 ( .B1(n5191), .B2(n5187), .A(n9988), .ZN(n5186) );
  INV_X1 U5813 ( .A(n5188), .ZN(n5187) );
  INV_X1 U5814 ( .A(n10034), .ZN(n10383) );
  NAND2_X1 U5815 ( .A1(n5190), .A2(n9862), .ZN(n10400) );
  NAND2_X1 U5816 ( .A1(n5190), .A2(n5188), .ZN(n10402) );
  NAND2_X1 U5817 ( .A1(n10443), .A2(n9984), .ZN(n10420) );
  AND2_X1 U5818 ( .A1(n9983), .A2(n9984), .ZN(n10445) );
  INV_X1 U5819 ( .A(n5114), .ZN(n5113) );
  OAI21_X1 U5820 ( .B1(n5115), .B2(n8571), .A(n5423), .ZN(n5114) );
  INV_X1 U5821 ( .A(n5424), .ZN(n5115) );
  NOR2_X1 U5822 ( .A1(n10559), .A2(n5353), .ZN(n10437) );
  INV_X1 U5823 ( .A(n5355), .ZN(n5353) );
  NOR2_X1 U5824 ( .A1(n10559), .A2(n10543), .ZN(n10461) );
  NAND2_X1 U5825 ( .A1(n8575), .A2(n9972), .ZN(n10452) );
  AND4_X1 U5826 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n10555)
         );
  OR2_X1 U5827 ( .A1(n6719), .A2(n10184), .ZN(n6736) );
  AND4_X1 U5828 ( .A1(n6741), .A2(n6740), .A3(n6739), .A4(n6738), .ZN(n10453)
         );
  NAND2_X1 U5829 ( .A1(n5396), .A2(n5395), .ZN(n8494) );
  NAND2_X1 U5830 ( .A1(n10916), .A2(n5405), .ZN(n8488) );
  INV_X1 U5831 ( .A(n5408), .ZN(n5405) );
  NAND2_X1 U5832 ( .A1(n5396), .A2(n9952), .ZN(n8433) );
  NAND2_X1 U5833 ( .A1(n8053), .A2(n5038), .ZN(n10919) );
  AND4_X1 U5834 ( .A1(n6687), .A2(n6686), .A3(n6685), .A4(n6684), .ZN(n10926)
         );
  NAND2_X1 U5835 ( .A1(n8053), .A2(n5037), .ZN(n10918) );
  AND4_X1 U5836 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(n8428)
         );
  NAND2_X1 U5837 ( .A1(n8048), .A2(n10047), .ZN(n8158) );
  NAND2_X1 U5838 ( .A1(n5180), .A2(n5178), .ZN(n10922) );
  AOI21_X1 U5839 ( .B1(n5181), .B2(n5184), .A(n5179), .ZN(n5178) );
  AOI21_X1 U5840 ( .B1(n10047), .B2(n5183), .A(n5182), .ZN(n5181) );
  AND2_X1 U5841 ( .A1(n8053), .A2(n10888), .ZN(n8163) );
  NAND2_X1 U5842 ( .A1(n8042), .A2(n10101), .ZN(n5422) );
  NAND2_X1 U5843 ( .A1(n8000), .A2(n7908), .ZN(n8043) );
  OR2_X1 U5844 ( .A1(n6596), .A2(n6407), .ZN(n6625) );
  NAND2_X1 U5845 ( .A1(n7914), .A2(n9938), .ZN(n5384) );
  NAND2_X1 U5846 ( .A1(n7914), .A2(n5383), .ZN(n8047) );
  AND2_X1 U5847 ( .A1(n9940), .A2(n9938), .ZN(n5383) );
  NAND2_X1 U5848 ( .A1(n7998), .A2(n10044), .ZN(n8000) );
  NAND2_X1 U5849 ( .A1(n9937), .A2(n9938), .ZN(n10044) );
  NAND2_X1 U5850 ( .A1(n5347), .A2(n5346), .ZN(n8071) );
  NAND2_X1 U5851 ( .A1(n7912), .A2(n8062), .ZN(n8064) );
  NOR2_X1 U5852 ( .A1(n10760), .A2(n5348), .ZN(n8072) );
  AND2_X1 U5853 ( .A1(n9894), .A2(n9930), .ZN(n10040) );
  AND2_X1 U5854 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6531) );
  NAND3_X1 U5855 ( .A1(n6505), .A2(n5556), .A3(n6504), .ZN(n8118) );
  OR2_X1 U5856 ( .A1(n9819), .A2(n7186), .ZN(n6504) );
  AOI21_X1 U5857 ( .B1(n7858), .B2(n8124), .A(n10785), .ZN(n6428) );
  NAND2_X1 U5858 ( .A1(n9811), .A2(n9810), .ZN(n10473) );
  NAND2_X1 U5859 ( .A1(n6890), .A2(n6889), .ZN(n10488) );
  NAND2_X1 U5860 ( .A1(n6794), .A2(n6793), .ZN(n10532) );
  NAND2_X1 U5861 ( .A1(n6607), .A2(n6606), .ZN(n8125) );
  AND2_X1 U5862 ( .A1(n7381), .A2(n10081), .ZN(n10827) );
  AND2_X1 U5863 ( .A1(n9669), .A2(n9673), .ZN(n5386) );
  AND2_X1 U5864 ( .A1(n6133), .A2(n6123), .ZN(n8791) );
  XNOR2_X1 U5865 ( .A(n6101), .B(n6097), .ZN(n8506) );
  NAND2_X1 U5866 ( .A1(n6084), .A2(n6083), .ZN(n6101) );
  NAND2_X1 U5867 ( .A1(n6944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6387) );
  OAI21_X1 U5868 ( .B1(n6014), .B2(n6013), .A(n6015), .ZN(n6028) );
  AND2_X1 U5869 ( .A1(n6029), .A2(n6018), .ZN(n6027) );
  INV_X1 U5870 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6424) );
  INV_X1 U5871 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U5872 ( .A1(n5451), .A2(n5913), .ZN(n5929) );
  OR2_X1 U5873 ( .A1(n5911), .A2(n5912), .ZN(n5451) );
  XNOR2_X1 U5874 ( .A(n5669), .B(n9504), .ZN(n5673) );
  NAND2_X1 U5875 ( .A1(n5233), .A2(n5633), .ZN(n5648) );
  OAI21_X1 U5876 ( .B1(n5034), .B2(n7195), .A(n5607), .ZN(n5616) );
  INV_X1 U5877 ( .A(n7894), .ZN(n10853) );
  XNOR2_X1 U5878 ( .A(n8754), .B(n7037), .ZN(n8740) );
  NAND2_X1 U5879 ( .A1(n8719), .A2(n7084), .ZN(n8725) );
  NAND2_X1 U5880 ( .A1(n8096), .A2(n7020), .ZN(n7160) );
  OAI211_X1 U5881 ( .C1(n5311), .C2(n5313), .A(n6977), .B(n5309), .ZN(n7545)
         );
  NAND2_X1 U5882 ( .A1(n5310), .A2(n5312), .ZN(n5309) );
  INV_X1 U5883 ( .A(n5312), .ZN(n5311) );
  XNOR2_X1 U5884 ( .A(n6980), .B(n8636), .ZN(n7546) );
  NAND2_X1 U5885 ( .A1(n7072), .A2(n7071), .ZN(n8823) );
  NAND2_X1 U5886 ( .A1(n6055), .A2(n6054), .ZN(n9178) );
  NAND2_X1 U5887 ( .A1(n5902), .A2(n5901), .ZN(n9229) );
  NAND2_X1 U5888 ( .A1(n8698), .A2(n7053), .ZN(n8461) );
  XNOR2_X1 U5889 ( .A(n7091), .B(n7089), .ZN(n8847) );
  NAND2_X1 U5890 ( .A1(n7961), .A2(n7010), .ZN(n5293) );
  NAND2_X1 U5891 ( .A1(n5972), .A2(n5971), .ZN(n9204) );
  NAND2_X1 U5892 ( .A1(n5442), .A2(n7076), .ZN(n8868) );
  NAND2_X1 U5893 ( .A1(n8823), .A2(n8822), .ZN(n5442) );
  INV_X1 U5894 ( .A(n8891), .ZN(n8703) );
  NAND2_X1 U5895 ( .A1(n6982), .A2(n8637), .ZN(n8648) );
  NOR2_X1 U5896 ( .A1(n8458), .A2(n5302), .ZN(n5301) );
  INV_X1 U5897 ( .A(n7053), .ZN(n5302) );
  NAND2_X1 U5898 ( .A1(n7000), .A2(n8678), .ZN(n8685) );
  NAND2_X1 U5899 ( .A1(n5307), .A2(n5057), .ZN(n7000) );
  AND2_X1 U5900 ( .A1(n5307), .A2(n5042), .ZN(n8775) );
  NAND2_X1 U5901 ( .A1(n8833), .A2(n7098), .ZN(n8875) );
  NAND2_X1 U5902 ( .A1(n6072), .A2(n6071), .ZN(n9173) );
  AOI21_X1 U5903 ( .B1(n8729), .B2(n7045), .A(n5553), .ZN(n8762) );
  NOR2_X1 U5904 ( .A1(n7044), .A2(n7043), .ZN(n5553) );
  NOR2_X1 U5905 ( .A1(n6342), .A2(n5555), .ZN(n6346) );
  NAND4_X1 U5906 ( .A1(n5626), .A2(n5625), .A3(n5624), .A4(n5623), .ZN(n8900)
         );
  NAND2_X1 U5907 ( .A1(n7299), .A2(n7298), .ZN(n7313) );
  NAND2_X1 U5908 ( .A1(n7313), .A2(n5106), .ZN(n7315) );
  NAND2_X1 U5909 ( .A1(n7302), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5106) );
  AND2_X1 U5910 ( .A1(n7447), .A2(n5103), .ZN(n7490) );
  NAND2_X1 U5911 ( .A1(n7448), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5103) );
  NOR2_X1 U5912 ( .A1(n7475), .A2(n5079), .ZN(n7479) );
  NOR2_X1 U5913 ( .A1(n7479), .A2(n7478), .ZN(n7536) );
  NOR2_X1 U5914 ( .A1(n7536), .A2(n5100), .ZN(n7540) );
  AND2_X1 U5915 ( .A1(n7537), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U5916 ( .A1(n7663), .A2(n7662), .ZN(n7667) );
  INV_X1 U5917 ( .A(n5899), .ZN(n5508) );
  INV_X1 U5918 ( .A(n5105), .ZN(n8923) );
  NAND2_X1 U5919 ( .A1(n5105), .A2(n5104), .ZN(n8925) );
  NAND2_X1 U5920 ( .A1(n8924), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5104) );
  NOR2_X1 U5921 ( .A1(n8925), .A2(n8926), .ZN(n8942) );
  NAND2_X1 U5922 ( .A1(n6163), .A2(n6162), .ZN(n9148) );
  AOI21_X1 U5923 ( .B1(n5487), .B2(n5491), .A(n5090), .ZN(n5485) );
  AOI21_X1 U5924 ( .B1(n5382), .B2(n10798), .A(n5379), .ZN(n9165) );
  NAND2_X1 U5925 ( .A1(n5381), .A2(n5380), .ZN(n5379) );
  NAND2_X1 U5926 ( .A1(n8976), .A2(n9139), .ZN(n5381) );
  NAND2_X1 U5927 ( .A1(n5486), .A2(n5490), .ZN(n8970) );
  AND2_X1 U5928 ( .A1(n8994), .A2(n8993), .ZN(n9170) );
  NAND2_X1 U5929 ( .A1(n9035), .A2(n5365), .ZN(n5358) );
  NOR2_X1 U5930 ( .A1(n9020), .A2(n9019), .ZN(n9018) );
  NOR2_X1 U5931 ( .A1(n9035), .A2(n6045), .ZN(n9020) );
  NAND2_X1 U5932 ( .A1(n9187), .A2(n5549), .ZN(n9029) );
  INV_X1 U5933 ( .A(n9054), .ZN(n9057) );
  NAND2_X1 U5934 ( .A1(n5373), .A2(n5035), .ZN(n9044) );
  INV_X1 U5935 ( .A(n5246), .ZN(n9088) );
  AOI21_X1 U5936 ( .B1(n9108), .B2(n5247), .A(n5249), .ZN(n5246) );
  NAND2_X1 U5937 ( .A1(n9094), .A2(n5554), .ZN(n9081) );
  OAI21_X1 U5938 ( .B1(n9108), .B2(n9112), .A(n6258), .ZN(n9101) );
  NAND2_X1 U5939 ( .A1(n8417), .A2(n5326), .ZN(n9128) );
  NAND2_X1 U5940 ( .A1(n5256), .A2(n5257), .ZN(n8534) );
  NAND2_X1 U5941 ( .A1(n5501), .A2(n5503), .ZN(n8516) );
  NAND2_X1 U5942 ( .A1(n5502), .A2(n8510), .ZN(n5501) );
  AND2_X1 U5943 ( .A1(n8412), .A2(n8411), .ZN(n8515) );
  NAND2_X1 U5944 ( .A1(n5861), .A2(n5860), .ZN(n8744) );
  NAND2_X1 U5945 ( .A1(n7236), .A2(n6161), .ZN(n5861) );
  NAND2_X1 U5946 ( .A1(n8319), .A2(n5483), .ZN(n8601) );
  NAND2_X1 U5947 ( .A1(n5737), .A2(n5736), .ZN(n10868) );
  CLKBUF_X1 U5948 ( .A(n8422), .Z(n10815) );
  INV_X1 U5949 ( .A(n5578), .ZN(n9698) );
  XNOR2_X1 U5950 ( .A(n5577), .B(n5576), .ZN(n8592) );
  OR2_X1 U5951 ( .A1(n5592), .A2(n5645), .ZN(n5594) );
  NAND2_X1 U5952 ( .A1(n6357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5591) );
  INV_X1 U5953 ( .A(n7588), .ZN(n7811) );
  INV_X1 U5954 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5652) );
  AND4_X1 U5955 ( .A1(n6558), .A2(n6557), .A3(n6556), .A4(n6555), .ZN(n8067)
         );
  NAND2_X1 U5956 ( .A1(n5205), .A2(n6638), .ZN(n8229) );
  NAND2_X1 U5957 ( .A1(n5203), .A2(n6639), .ZN(n8230) );
  OR2_X1 U5958 ( .A1(n6497), .A2(n7989), .ZN(n6482) );
  INV_X1 U5959 ( .A(n8118), .ZN(n10719) );
  NOR2_X1 U5960 ( .A1(n5217), .A2(n7146), .ZN(n5216) );
  INV_X1 U5961 ( .A(n5218), .ZN(n5217) );
  NAND2_X1 U5962 ( .A1(n5529), .A2(n5530), .ZN(n9720) );
  OR2_X1 U5963 ( .A1(n9710), .A2(n5533), .ZN(n5529) );
  NAND2_X1 U5964 ( .A1(n5516), .A2(n5513), .ZN(n9731) );
  AND4_X1 U5965 ( .A1(n6783), .A2(n6782), .A3(n6781), .A4(n6780), .ZN(n10454)
         );
  AND4_X1 U5966 ( .A1(n6442), .A2(n6441), .A3(n6440), .A4(n6439), .ZN(n10387)
         );
  AND4_X1 U5967 ( .A1(n6590), .A2(n6589), .A3(n6588), .A4(n6587), .ZN(n8066)
         );
  NAND2_X1 U5968 ( .A1(n9709), .A2(n6807), .ZN(n9769) );
  NAND2_X1 U5969 ( .A1(n5211), .A2(n5526), .ZN(n9778) );
  NAND2_X1 U5970 ( .A1(n9710), .A2(n5527), .ZN(n5211) );
  NAND2_X1 U5971 ( .A1(n6843), .A2(n6842), .ZN(n10515) );
  NAND2_X1 U5972 ( .A1(n6639), .A2(n8231), .ZN(n5201) );
  NAND2_X1 U5973 ( .A1(n6643), .A2(n6642), .ZN(n10564) );
  AND4_X1 U5974 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n10556)
         );
  AND4_X1 U5975 ( .A1(n6575), .A2(n6574), .A3(n6573), .A4(n6572), .ZN(n8022)
         );
  NOR2_X2 U5976 ( .A1(n6951), .A2(n6961), .ZN(n9756) );
  AND4_X1 U5977 ( .A1(n6417), .A2(n6416), .A3(n6415), .A4(n6414), .ZN(n10321)
         );
  AOI21_X1 U5978 ( .B1(n5516), .B2(n5512), .A(n5036), .ZN(n9796) );
  NAND2_X1 U5979 ( .A1(n6876), .A2(n6875), .ZN(n10493) );
  NAND2_X1 U5980 ( .A1(n8445), .A2(n9807), .ZN(n6876) );
  AND4_X1 U5981 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(n9830)
         );
  INV_X1 U5982 ( .A(n9753), .ZN(n9803) );
  OAI21_X1 U5983 ( .B1(n8548), .B2(n8547), .A(n8551), .ZN(n9739) );
  INV_X1 U5984 ( .A(n8066), .ZN(n10102) );
  OR2_X1 U5985 ( .A1(n7251), .A2(P1_U3084), .ZN(n10106) );
  NAND2_X1 U5986 ( .A1(n6795), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U5987 ( .A1(n6644), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6466) );
  NOR2_X1 U5988 ( .A1(n10173), .A2(n5161), .ZN(n10660) );
  NOR2_X1 U5989 ( .A1(n5162), .A2(n7918), .ZN(n5161) );
  INV_X1 U5990 ( .A(n10177), .ZN(n5162) );
  INV_X1 U5991 ( .A(n5160), .ZN(n10658) );
  INV_X1 U5992 ( .A(n5176), .ZN(n8178) );
  XNOR2_X1 U5993 ( .A(n10195), .B(n10194), .ZN(n10190) );
  INV_X1 U5994 ( .A(n5173), .ZN(n10196) );
  OAI21_X1 U5995 ( .B1(n10263), .B2(n10264), .A(n5165), .ZN(n5164) );
  INV_X1 U5996 ( .A(n10262), .ZN(n5165) );
  NOR2_X1 U5997 ( .A1(n10254), .A2(n5169), .ZN(n5168) );
  AND2_X1 U5998 ( .A1(n10255), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5169) );
  AND2_X1 U5999 ( .A1(n5399), .A2(n5398), .ZN(n10479) );
  AOI22_X1 U6000 ( .A1(n10297), .A2(n10768), .B1(n10265), .B2(n10091), .ZN(
        n5398) );
  NAND2_X1 U6001 ( .A1(n8811), .A2(n10930), .ZN(n5399) );
  NAND2_X1 U6002 ( .A1(n6906), .A2(n6905), .ZN(n10481) );
  AOI21_X1 U6003 ( .B1(n5195), .B2(n10930), .A(n5193), .ZN(n10490) );
  INV_X1 U6004 ( .A(n5194), .ZN(n5193) );
  XNOR2_X1 U6005 ( .A(n5196), .B(n10012), .ZN(n5195) );
  AOI22_X1 U6006 ( .A1(n10297), .A2(n10769), .B1(n10768), .B2(n10298), .ZN(
        n5194) );
  NAND2_X1 U6007 ( .A1(n5412), .A2(n8787), .ZN(n10314) );
  NAND2_X1 U6008 ( .A1(n5418), .A2(n5416), .ZN(n5412) );
  NAND2_X1 U6009 ( .A1(n8803), .A2(n10005), .ZN(n10340) );
  NAND2_X1 U6010 ( .A1(n5418), .A2(n8785), .ZN(n10333) );
  NAND2_X1 U6011 ( .A1(n8784), .A2(n8783), .ZN(n10347) );
  INV_X1 U6012 ( .A(n10515), .ZN(n10394) );
  NAND2_X1 U6013 ( .A1(n6824), .A2(n6823), .ZN(n10518) );
  AND2_X1 U6014 ( .A1(n5429), .A2(n5074), .ZN(n10398) );
  NAND2_X1 U6015 ( .A1(n5429), .A2(n5428), .ZN(n10397) );
  NAND2_X1 U6016 ( .A1(n6809), .A2(n6808), .ZN(n10526) );
  NAND2_X1 U6017 ( .A1(n5425), .A2(n5424), .ZN(n8778) );
  INV_X1 U6018 ( .A(n5401), .ZN(n8570) );
  AOI21_X1 U6019 ( .B1(n10916), .B2(n5402), .A(n5404), .ZN(n5401) );
  NAND2_X1 U6020 ( .A1(n6718), .A2(n6717), .ZN(n8569) );
  NAND2_X1 U6021 ( .A1(n6699), .A2(n6698), .ZN(n9831) );
  NAND2_X1 U6022 ( .A1(n6634), .A2(n6633), .ZN(n8155) );
  OAI211_X1 U6023 ( .C1(n6503), .C2(n7276), .A(n6580), .B(n6579), .ZN(n8076)
         );
  OR2_X1 U6024 ( .A1(n7192), .A2(n9819), .ZN(n5431) );
  AND2_X1 U6025 ( .A1(n6540), .A2(n5070), .ZN(n5430) );
  AND2_X1 U6026 ( .A1(n11019), .A2(n7921), .ZN(n10433) );
  NAND2_X1 U6027 ( .A1(n10588), .A2(n7829), .ZN(n11014) );
  OAI21_X1 U6028 ( .B1(n6503), .B2(n6461), .A(n6460), .ZN(n8014) );
  INV_X1 U6029 ( .A(n11012), .ZN(n10413) );
  AND2_X1 U6030 ( .A1(n11023), .A2(n11033), .ZN(n10470) );
  AOI211_X1 U6031 ( .C1(n11034), .C2(n11033), .A(n11032), .B(n11031), .ZN(
        n11039) );
  NAND2_X1 U6032 ( .A1(n6136), .A2(n6157), .ZN(n9820) );
  OR2_X1 U6033 ( .A1(n10591), .A2(n6577), .ZN(n6401) );
  OAI21_X1 U6034 ( .B1(n6381), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5158) );
  XNOR2_X1 U6035 ( .A(n6382), .B(n9673), .ZN(n8508) );
  NAND2_X1 U6036 ( .A1(n6381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U6037 ( .A1(n6395), .A2(n6394), .ZN(n8312) );
  XNOR2_X1 U6038 ( .A(n6028), .B(n6027), .ZN(n8138) );
  NAND2_X1 U6039 ( .A1(n5123), .A2(n5671), .ZN(n5122) );
  XNOR2_X1 U6040 ( .A(n5692), .B(n5691), .ZN(n7192) );
  AND2_X1 U6041 ( .A1(n5677), .A2(n5676), .ZN(n5692) );
  NAND2_X1 U6042 ( .A1(n6450), .A2(n5170), .ZN(n7259) );
  INV_X1 U6043 ( .A(n5171), .ZN(n5170) );
  OAI21_X1 U6044 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_1__SCAN_IN), .A(
        n5172), .ZN(n5171) );
  OR2_X1 U6045 ( .A1(n7130), .A2(n5439), .ZN(n7144) );
  NAND2_X1 U6046 ( .A1(n8903), .A2(n5312), .ZN(n7514) );
  OAI21_X1 U6047 ( .B1(n5166), .B2(n10657), .A(n5163), .ZN(P1_U3260) );
  XNOR2_X1 U6048 ( .A(n5168), .B(n5167), .ZN(n5166) );
  INV_X1 U6049 ( .A(n5164), .ZN(n5163) );
  INV_X1 U6050 ( .A(n10257), .ZN(n5167) );
  OAI21_X1 U6051 ( .B1(n10480), .B2(n11021), .A(n5116), .ZN(P1_U3355) );
  INV_X1 U6052 ( .A(n5117), .ZN(n5116) );
  OAI21_X1 U6053 ( .B1(n10479), .B2(n10465), .A(n5118), .ZN(n5117) );
  AOI21_X1 U6054 ( .B1(n10477), .B2(n10470), .A(n8812), .ZN(n5118) );
  OR2_X1 U6055 ( .A1(n8744), .A2(n8747), .ZN(n6237) );
  AND2_X1 U6056 ( .A1(n9046), .A2(n6272), .ZN(n5035) );
  AND2_X1 U6057 ( .A1(n6874), .A2(n6873), .ZN(n5036) );
  AND2_X1 U6058 ( .A1(n8509), .A2(n6240), .ZN(n8514) );
  AND2_X1 U6059 ( .A1(n8168), .A2(n10888), .ZN(n5037) );
  AND2_X1 U6060 ( .A1(n5037), .A2(n5350), .ZN(n5038) );
  AND2_X1 U6061 ( .A1(n9945), .A2(n9944), .ZN(n10047) );
  INV_X1 U6062 ( .A(n10047), .ZN(n5184) );
  INV_X1 U6063 ( .A(n5491), .ZN(n5490) );
  OAI22_X1 U6064 ( .A1(n8989), .A2(n5494), .B1(n9000), .B2(n9167), .ZN(n5491)
         );
  AND2_X1 U6065 ( .A1(n5038), .A2(n5349), .ZN(n5039) );
  OR2_X1 U6066 ( .A1(n9182), .A2(n6044), .ZN(n6288) );
  NAND2_X1 U6067 ( .A1(n10032), .A2(n10033), .ZN(n5145) );
  NAND2_X1 U6068 ( .A1(n5783), .A2(n5782), .ZN(n8609) );
  AND2_X1 U6069 ( .A1(n5335), .A2(n10949), .ZN(n5040) );
  NAND2_X1 U6070 ( .A1(n5508), .A2(n5569), .ZN(n5915) );
  NAND2_X1 U6071 ( .A1(n5955), .A2(n5954), .ZN(n9211) );
  NAND2_X1 U6072 ( .A1(n5604), .A2(n5603), .ZN(n7314) );
  NAND2_X2 U6073 ( .A1(n7701), .A2(n8039), .ZN(n6308) );
  NAND2_X1 U6074 ( .A1(n8784), .A2(n5419), .ZN(n5418) );
  NAND3_X1 U6075 ( .A1(n6514), .A2(n6513), .A3(n6512), .ZN(n7834) );
  NAND2_X1 U6076 ( .A1(n7064), .A2(n7065), .ZN(n5041) );
  OR2_X1 U6077 ( .A1(n8771), .A2(n6995), .ZN(n5042) );
  NAND3_X1 U6078 ( .A1(n6925), .A2(n6928), .A3(n6396), .ZN(n6418) );
  NOR2_X1 U6079 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6449) );
  NAND4_X1 U6080 ( .A1(n6467), .A2(n6466), .A3(n6465), .A4(n6464), .ZN(n6469)
         );
  OR2_X1 U6081 ( .A1(n10543), .A2(n10093), .ZN(n5043) );
  OAI211_X1 U6082 ( .C1(n6503), .C2(n7207), .A(n6592), .B(n6591), .ZN(n8009)
         );
  OR2_X1 U6083 ( .A1(n9204), .A2(n8653), .ZN(n6263) );
  NOR2_X1 U6084 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5602) );
  INV_X1 U6085 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5593) );
  NOR2_X1 U6086 ( .A1(n6856), .A2(n5521), .ZN(n5044) );
  AND2_X1 U6087 ( .A1(n6559), .A2(n9404), .ZN(n6576) );
  AND2_X1 U6088 ( .A1(n5627), .A2(n5628), .ZN(n5644) );
  NAND2_X1 U6089 ( .A1(n6449), .A2(n9620), .ZN(n6487) );
  AOI21_X1 U6090 ( .B1(n9108), .B2(n5248), .A(n5244), .ZN(n5243) );
  XNOR2_X1 U6091 ( .A(n6401), .B(n9668), .ZN(n6405) );
  OR2_X1 U6092 ( .A1(n9086), .A2(n9102), .ZN(n5045) );
  NAND4_X1 U6093 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n10730)
         );
  INV_X1 U6094 ( .A(n10730), .ZN(n5112) );
  AND2_X1 U6095 ( .A1(n5358), .A2(n5363), .ZN(n5046) );
  OR2_X1 U6096 ( .A1(n6857), .A2(n6856), .ZN(n5047) );
  AND4_X1 U6097 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n5048) );
  INV_X1 U6098 ( .A(n6470), .ZN(n6854) );
  NOR2_X1 U6099 ( .A1(n7154), .A2(n6419), .ZN(n6470) );
  NAND2_X1 U6100 ( .A1(n5986), .A2(n5985), .ZN(n9199) );
  OR3_X1 U6101 ( .A1(n6339), .A2(n7588), .A3(n7428), .ZN(n5049) );
  AND2_X1 U6102 ( .A1(n9946), .A2(n10046), .ZN(n5050) );
  AND2_X1 U6103 ( .A1(n10019), .A2(n10018), .ZN(n5051) );
  INV_X1 U6104 ( .A(n8892), .ZN(n8320) );
  NOR2_X1 U6105 ( .A1(n7540), .A2(n7539), .ZN(n5052) );
  NOR2_X1 U6106 ( .A1(n7496), .A2(n6918), .ZN(n5053) );
  NAND2_X1 U6107 ( .A1(n6775), .A2(n6774), .ZN(n10538) );
  AND2_X1 U6108 ( .A1(n9037), .A2(n5549), .ZN(n5054) );
  NAND2_X1 U6109 ( .A1(n6314), .A2(n6313), .ZN(n8659) );
  INV_X1 U6110 ( .A(n8659), .ZN(n5493) );
  NOR2_X1 U6111 ( .A1(n5870), .A2(n5263), .ZN(n5262) );
  AND2_X1 U6112 ( .A1(n5589), .A2(n5590), .ZN(n5055) );
  AND2_X1 U6113 ( .A1(n10518), .A2(n10422), .ZN(n5056) );
  AND2_X1 U6114 ( .A1(n5042), .A2(n6999), .ZN(n5057) );
  OR2_X1 U6115 ( .A1(n10488), .A2(n10322), .ZN(n9919) );
  INV_X1 U6116 ( .A(n6314), .ZN(n5366) );
  OR2_X1 U6117 ( .A1(n9173), .A2(n8658), .ZN(n6314) );
  AND2_X1 U6118 ( .A1(n8654), .A2(n5554), .ZN(n5058) );
  AND2_X1 U6119 ( .A1(n10538), .A2(n10446), .ZN(n5059) );
  INV_X1 U6120 ( .A(n8594), .ZN(n9156) );
  NAND2_X1 U6121 ( .A1(n6125), .A2(n6124), .ZN(n8594) );
  OR2_X1 U6122 ( .A1(n9194), .A2(n8827), .ZN(n6272) );
  NAND2_X1 U6123 ( .A1(n6176), .A2(n6175), .ZN(n8974) );
  INV_X1 U6124 ( .A(n8974), .ZN(n8969) );
  NOR2_X1 U6125 ( .A1(n8874), .A2(n5438), .ZN(n5437) );
  INV_X1 U6126 ( .A(n5437), .ZN(n5436) );
  AND2_X1 U6127 ( .A1(n5873), .A2(SI_14_), .ZN(n5060) );
  NAND2_X1 U6128 ( .A1(n5386), .A2(n9666), .ZN(n5061) );
  NOR2_X1 U6129 ( .A1(n5899), .A2(n5506), .ZN(n6145) );
  NAND2_X1 U6130 ( .A1(n8313), .A2(n8314), .ZN(n5062) );
  AND2_X1 U6131 ( .A1(n10012), .A2(n10011), .ZN(n5063) );
  OR2_X1 U6132 ( .A1(n9178), .A2(n8851), .ZN(n6178) );
  NOR2_X1 U6133 ( .A1(n9199), .A2(n9068), .ZN(n5064) );
  NAND2_X1 U6134 ( .A1(n5240), .A2(n5813), .ZN(n6219) );
  INV_X1 U6135 ( .A(n10826), .ZN(n7899) );
  AND2_X1 U6136 ( .A1(n8831), .A2(n7097), .ZN(n5065) );
  OR2_X1 U6137 ( .A1(n5910), .A2(n5909), .ZN(n5066) );
  AND2_X1 U6138 ( .A1(n6576), .A2(n5546), .ZN(n6397) );
  NAND2_X1 U6139 ( .A1(n9173), .A2(n8658), .ZN(n6313) );
  AND2_X1 U6140 ( .A1(n9942), .A2(n9941), .ZN(n9940) );
  INV_X1 U6141 ( .A(n5499), .ZN(n5498) );
  NAND2_X1 U6142 ( .A1(n5503), .A2(n5500), .ZN(n5499) );
  INV_X1 U6143 ( .A(n5145), .ZN(n5144) );
  OR2_X1 U6144 ( .A1(n10195), .A2(n10194), .ZN(n5067) );
  AND2_X1 U6145 ( .A1(n10043), .A2(n7908), .ZN(n5068) );
  AND2_X1 U6146 ( .A1(n10457), .A2(n9974), .ZN(n5069) );
  NAND2_X1 U6147 ( .A1(n6139), .A2(n6138), .ZN(n8965) );
  INV_X1 U6148 ( .A(n8965), .ZN(n5338) );
  OR2_X1 U6149 ( .A1(n6503), .A2(n7257), .ZN(n5070) );
  AND2_X1 U6150 ( .A1(n7033), .A2(n7034), .ZN(n5071) );
  AND2_X1 U6151 ( .A1(n6133), .A2(n6132), .ZN(n5072) );
  INV_X1 U6152 ( .A(n5694), .ZN(n5239) );
  NAND2_X1 U6153 ( .A1(n9729), .A2(n9728), .ZN(n5073) );
  INV_X1 U6154 ( .A(n8430), .ZN(n10049) );
  AND2_X1 U6155 ( .A1(n9953), .A2(n9832), .ZN(n8430) );
  OR2_X1 U6156 ( .A1(n10526), .A2(n10447), .ZN(n5074) );
  OR2_X1 U6157 ( .A1(n5835), .A2(n5834), .ZN(n5075) );
  NAND2_X1 U6158 ( .A1(n8027), .A2(n6623), .ZN(n5205) );
  XOR2_X1 U6159 ( .A(n6924), .B(n6923), .Z(n5076) );
  INV_X1 U6160 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5547) );
  AND2_X1 U6161 ( .A1(n8417), .A2(n5328), .ZN(n5077) );
  NAND2_X1 U6162 ( .A1(n10007), .A2(n10005), .ZN(n5391) );
  NAND2_X1 U6163 ( .A1(n6003), .A2(n6002), .ZN(n9194) );
  XOR2_X1 U6164 ( .A(n9831), .B(n10096), .Z(n5078) );
  AND2_X1 U6165 ( .A1(n7476), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5079) );
  OAI21_X1 U6166 ( .B1(n10548), .B2(n5115), .A(n5113), .ZN(n10435) );
  XNOR2_X1 U6167 ( .A(n5873), .B(n9484), .ZN(n5872) );
  NAND2_X1 U6168 ( .A1(n9919), .A2(n9920), .ZN(n10300) );
  OR2_X1 U6169 ( .A1(n6853), .A2(n6852), .ZN(n5080) );
  XNOR2_X1 U6170 ( .A(n6387), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6925) );
  AND2_X1 U6171 ( .A1(n10650), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5081) );
  INV_X1 U6172 ( .A(n5856), .ZN(n5459) );
  NAND2_X1 U6173 ( .A1(n5931), .A2(n5930), .ZN(n9216) );
  INV_X1 U6174 ( .A(n9784), .ZN(n5210) );
  NAND2_X1 U6175 ( .A1(n6384), .A2(n6383), .ZN(n10500) );
  INV_X1 U6176 ( .A(n10500), .ZN(n5343) );
  NAND2_X1 U6177 ( .A1(n6288), .A2(n6282), .ZN(n9037) );
  INV_X1 U6178 ( .A(n9037), .ZN(n5269) );
  AND2_X1 U6179 ( .A1(n8319), .A2(n5480), .ZN(n5082) );
  NAND2_X1 U6180 ( .A1(n5918), .A2(n5917), .ZN(n9223) );
  OR2_X1 U6181 ( .A1(n8381), .A2(n8382), .ZN(n8412) );
  NAND2_X1 U6182 ( .A1(n5316), .A2(n5571), .ZN(n6353) );
  AND2_X1 U6183 ( .A1(n10916), .A2(n8429), .ZN(n5083) );
  NAND2_X1 U6184 ( .A1(n6103), .A2(n6102), .ZN(n9162) );
  INV_X1 U6185 ( .A(n9162), .ZN(n5342) );
  NAND2_X1 U6186 ( .A1(n5878), .A2(n5877), .ZN(n8760) );
  NOR3_X1 U6187 ( .A1(n10559), .A2(n10526), .A3(n5354), .ZN(n5351) );
  INV_X1 U6188 ( .A(n8713), .ZN(n10964) );
  OR2_X1 U6189 ( .A1(n10964), .A2(n8733), .ZN(n5084) );
  AOI21_X1 U6190 ( .B1(n8548), .B2(n5542), .A(n5540), .ZN(n5537) );
  INV_X1 U6191 ( .A(n5352), .ZN(n10438) );
  NOR2_X1 U6192 ( .A1(n10559), .A2(n5354), .ZN(n5352) );
  OR2_X1 U6193 ( .A1(n10417), .A2(n9986), .ZN(n5429) );
  NAND2_X1 U6194 ( .A1(n8250), .A2(n5040), .ZN(n5336) );
  AND2_X1 U6195 ( .A1(n8569), .A2(n10095), .ZN(n5085) );
  AND2_X1 U6196 ( .A1(n5501), .A2(n5498), .ZN(n5086) );
  INV_X1 U6197 ( .A(n5332), .ZN(n9082) );
  NOR2_X1 U6198 ( .A1(n9117), .A2(n5333), .ZN(n5332) );
  INV_X1 U6199 ( .A(n9140), .ZN(n8652) );
  NAND2_X1 U6200 ( .A1(n5425), .A2(n5043), .ZN(n5087) );
  AND2_X1 U6201 ( .A1(n5927), .A2(SI_17_), .ZN(n5088) );
  NOR2_X1 U6202 ( .A1(n6887), .A2(n6888), .ZN(n5089) );
  AND2_X1 U6203 ( .A1(n5342), .A2(n8817), .ZN(n5090) );
  AND2_X1 U6204 ( .A1(n5326), .A2(n9134), .ZN(n5091) );
  AND2_X1 U6205 ( .A1(n6693), .A2(n5226), .ZN(n5092) );
  NOR2_X1 U6206 ( .A1(n5204), .A2(n5202), .ZN(n5093) );
  INV_X1 U6207 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5645) );
  AND2_X1 U6208 ( .A1(n9977), .A2(n9978), .ZN(n5094) );
  AND2_X1 U6209 ( .A1(n7102), .A2(n7101), .ZN(n5095) );
  XNOR2_X1 U6210 ( .A(n5594), .B(n5593), .ZN(n6364) );
  INV_X1 U6211 ( .A(n10046), .ZN(n5179) );
  AND2_X1 U6212 ( .A1(n5293), .A2(n8148), .ZN(n5096) );
  INV_X1 U6213 ( .A(n8525), .ZN(n5275) );
  AND2_X1 U6214 ( .A1(n6841), .A2(n6840), .ZN(n5097) );
  NAND2_X1 U6215 ( .A1(n5422), .A2(n8044), .ZN(n8045) );
  NAND2_X1 U6216 ( .A1(n7753), .A2(n7739), .ZN(n7728) );
  INV_X1 U6217 ( .A(n7728), .ZN(n5325) );
  NAND2_X1 U6218 ( .A1(n5422), .A2(n5421), .ZN(n8157) );
  INV_X1 U6219 ( .A(n5159), .ZN(n10684) );
  NAND2_X1 U6220 ( .A1(n5160), .A2(n7682), .ZN(n5159) );
  NAND2_X1 U6221 ( .A1(n5644), .A2(n5324), .ZN(n5899) );
  AND2_X1 U6222 ( .A1(n6621), .A2(n6620), .ZN(n5098) );
  INV_X1 U6223 ( .A(n5825), .ZN(n5377) );
  AND2_X1 U6224 ( .A1(n8648), .A2(n6986), .ZN(n5099) );
  NAND2_X1 U6225 ( .A1(n6428), .A2(n7155), .ZN(n7857) );
  NAND2_X1 U6226 ( .A1(n6661), .A2(n6660), .ZN(n10917) );
  INV_X1 U6227 ( .A(n10917), .ZN(n5350) );
  NAND4_X1 U6228 ( .A1(n6448), .A2(n6447), .A3(n6446), .A4(n6445), .ZN(n10107)
         );
  NAND2_X1 U6229 ( .A1(n6681), .A2(n6680), .ZN(n8478) );
  INV_X1 U6230 ( .A(n8478), .ZN(n5349) );
  AND2_X1 U6231 ( .A1(n6495), .A2(n7567), .ZN(n7521) );
  AND2_X1 U6232 ( .A1(n7036), .A2(n7783), .ZN(n5312) );
  NOR2_X1 U6233 ( .A1(n6381), .A2(n5061), .ZN(n10591) );
  INV_X1 U6234 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5300) );
  INV_X1 U6235 ( .A(n10812), .ZN(n9004) );
  INV_X1 U6236 ( .A(n10260), .ZN(n10785) );
  XNOR2_X1 U6237 ( .A(n6425), .B(n6424), .ZN(n8124) );
  MUX2_X1 U6238 ( .A(n7707), .B(P2_REG2_REG_1__SCAN_IN), .S(n7314), .Z(n7299)
         );
  AOI21_X2 U6239 ( .B1(n8998), .B2(n8659), .A(n5489), .ZN(n8980) );
  NAND2_X2 U6240 ( .A1(n5110), .A2(n5109), .ZN(n8998) );
  NAND2_X1 U6241 ( .A1(n6187), .A2(n7614), .ZN(n7745) );
  NAND2_X1 U6242 ( .A1(n8641), .A2(n5112), .ZN(n7614) );
  OAI211_X1 U6243 ( .C1(n7286), .C2(n7332), .A(n5621), .B(n5620), .ZN(n8641)
         );
  NAND2_X1 U6244 ( .A1(n10435), .A2(n8779), .ZN(n8781) );
  NAND3_X1 U6245 ( .A1(n5466), .A2(n5122), .A3(n5121), .ZN(n5237) );
  NAND3_X1 U6246 ( .A1(n5233), .A2(n5671), .A3(n5633), .ZN(n5121) );
  INV_X1 U6247 ( .A(n5647), .ZN(n5123) );
  NAND2_X1 U6248 ( .A1(n5648), .A2(n5647), .ZN(n5672) );
  NAND2_X1 U6249 ( .A1(n5672), .A2(n5671), .ZN(n5677) );
  NAND2_X1 U6250 ( .A1(n8000), .A2(n5068), .ZN(n8042) );
  INV_X1 U6251 ( .A(n8043), .ZN(n7910) );
  NAND2_X2 U6252 ( .A1(n5126), .A2(n5125), .ZN(n5650) );
  NAND3_X1 U6253 ( .A1(n5126), .A2(n5125), .A3(n5587), .ZN(n5606) );
  NAND3_X1 U6254 ( .A1(n5400), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5125) );
  NAND3_X1 U6255 ( .A1(n5232), .A2(n5231), .A3(n5230), .ZN(n5126) );
  NAND4_X1 U6256 ( .A1(n5130), .A2(n5129), .A3(n5128), .A4(n5127), .ZN(n6376)
         );
  OR2_X1 U6257 ( .A1(n9958), .A2(n5135), .ZN(n5134) );
  NAND2_X1 U6258 ( .A1(n5140), .A2(n5094), .ZN(n9982) );
  OAI21_X1 U6259 ( .B1(n5051), .B2(n5146), .A(n10028), .ZN(n10072) );
  OR2_X1 U6260 ( .A1(n10028), .A2(n5145), .ZN(n5142) );
  OAI211_X1 U6261 ( .C1(n5051), .C2(n5143), .A(n10068), .B(n5142), .ZN(n10066)
         );
  INV_X1 U6262 ( .A(n10022), .ZN(n5146) );
  AOI21_X1 U6263 ( .B1(n5151), .B2(n5150), .A(n5149), .ZN(n5148) );
  NAND2_X1 U6264 ( .A1(n5156), .A2(n5155), .ZN(n9931) );
  NAND2_X4 U6265 ( .A1(n8508), .A2(n6952), .ZN(n6503) );
  MUX2_X1 U6266 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7979), .S(n7259), .Z(n10109)
         );
  NAND3_X1 U6267 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6268 ( .A1(n8047), .A2(n5181), .ZN(n5180) );
  OAI21_X1 U6269 ( .B1(n10443), .B2(n5187), .A(n5185), .ZN(n10384) );
  NAND2_X1 U6270 ( .A1(n5199), .A2(n9845), .ZN(n10766) );
  INV_X1 U6271 ( .A(n9845), .ZN(n5198) );
  NAND2_X1 U6272 ( .A1(n8027), .A2(n5093), .ZN(n5200) );
  NAND2_X1 U6273 ( .A1(n5200), .A2(n5201), .ZN(n8207) );
  NAND2_X1 U6274 ( .A1(n6518), .A2(n5206), .ZN(n6519) );
  NAND2_X1 U6275 ( .A1(n5516), .A2(n5219), .ZN(n5215) );
  NAND2_X1 U6276 ( .A1(n5215), .A2(n5218), .ZN(n7147) );
  NAND2_X1 U6277 ( .A1(n5222), .A2(n5223), .ZN(n9745) );
  NAND3_X1 U6278 ( .A1(n6694), .A2(n6693), .A3(n5227), .ZN(n5222) );
  NAND2_X1 U6279 ( .A1(n6694), .A2(n5092), .ZN(n5225) );
  INV_X1 U6280 ( .A(n8448), .ZN(n5226) );
  NAND2_X1 U6281 ( .A1(n8448), .A2(n8449), .ZN(n5228) );
  NAND2_X1 U6282 ( .A1(n8451), .A2(n8448), .ZN(n6712) );
  NAND2_X1 U6283 ( .A1(n6694), .A2(n6693), .ZN(n8451) );
  NAND2_X1 U6284 ( .A1(n5630), .A2(n5631), .ZN(n5233) );
  NAND2_X1 U6285 ( .A1(n5616), .A2(n5617), .ZN(n5234) );
  NAND2_X1 U6286 ( .A1(n5236), .A2(n5694), .ZN(n5238) );
  INV_X1 U6287 ( .A(n5466), .ZN(n5236) );
  NAND2_X1 U6288 ( .A1(n5237), .A2(n5694), .ZN(n5718) );
  INV_X1 U6289 ( .A(n5243), .ZN(n9071) );
  NOR2_X1 U6290 ( .A1(n9036), .A2(n9037), .ZN(n9035) );
  OAI21_X1 U6291 ( .B1(n9036), .B2(n5268), .A(n5267), .ZN(n8990) );
  NAND2_X1 U6292 ( .A1(n8528), .A2(n5274), .ZN(n5273) );
  OAI21_X1 U6293 ( .B1(n7072), .B2(n5283), .A(n5280), .ZN(n8865) );
  NAND2_X1 U6294 ( .A1(n7072), .A2(n5280), .ZN(n5279) );
  NAND2_X1 U6295 ( .A1(n5855), .A2(n5285), .ZN(n5284) );
  NAND2_X1 U6296 ( .A1(n7961), .A2(n5294), .ZN(n5291) );
  NAND2_X1 U6297 ( .A1(n5291), .A2(n5290), .ZN(n7159) );
  NAND2_X1 U6298 ( .A1(n8698), .A2(n5301), .ZN(n7059) );
  NAND3_X1 U6299 ( .A1(n5304), .A2(n5075), .A3(n5303), .ZN(n5837) );
  NAND2_X1 U6300 ( .A1(n5305), .A2(n5767), .ZN(n5303) );
  NAND2_X1 U6301 ( .A1(n5759), .A2(n5305), .ZN(n5304) );
  NAND2_X1 U6302 ( .A1(n5476), .A2(n5475), .ZN(n5306) );
  NOR2_X1 U6303 ( .A1(n6167), .A2(n5318), .ZN(n5592) );
  NAND2_X1 U6304 ( .A1(n5316), .A2(n5315), .ZN(n5575) );
  INV_X1 U6305 ( .A(n6167), .ZN(n5316) );
  INV_X1 U6306 ( .A(n5495), .ZN(n5317) );
  NAND2_X2 U6307 ( .A1(n6677), .A2(n8289), .ZN(n8333) );
  NAND2_X1 U6308 ( .A1(n7059), .A2(n8459), .ZN(n8528) );
  NAND2_X1 U6309 ( .A1(n9843), .A2(n7833), .ZN(n7985) );
  NAND2_X2 U6310 ( .A1(n7286), .A2(n7182), .ZN(n6137) );
  OR3_X2 U6311 ( .A1(n7149), .A2(n5076), .A3(n6948), .ZN(n6974) );
  XNOR2_X1 U6312 ( .A(n7112), .B(n7111), .ZN(n7130) );
  OAI211_X2 U6313 ( .C1(n6137), .C2(n7194), .A(n5323), .B(n5322), .ZN(n7606)
         );
  OR2_X1 U6314 ( .A1(n7286), .A2(n7314), .ZN(n5322) );
  NAND2_X4 U6315 ( .A1(n7286), .A2(n5034), .ZN(n5695) );
  NAND2_X4 U6316 ( .A1(n6363), .A2(n6364), .ZN(n7286) );
  NAND2_X1 U6317 ( .A1(n6145), .A2(n6147), .ZN(n6167) );
  NOR2_X1 U6318 ( .A1(n9117), .A2(n9204), .ZN(n9096) );
  INV_X1 U6319 ( .A(n5336), .ZN(n8605) );
  AND2_X1 U6320 ( .A1(n9002), .A2(n5339), .ZN(n8971) );
  NAND2_X1 U6321 ( .A1(n9002), .A2(n5340), .ZN(n8964) );
  NOR2_X2 U6322 ( .A1(n10334), .A2(n10493), .ZN(n10325) );
  INV_X1 U6323 ( .A(n5351), .ZN(n10427) );
  AND2_X1 U6324 ( .A1(n6390), .A2(n6381), .ZN(n6928) );
  OAI21_X1 U6325 ( .B1(n7748), .B2(n5356), .A(n7747), .ZN(n7749) );
  NAND4_X1 U6326 ( .A1(n6319), .A2(n6318), .A3(n10797), .A4(n5356), .ZN(n6321)
         );
  NAND2_X1 U6327 ( .A1(n6186), .A2(n5356), .ZN(n6189) );
  NAND2_X1 U6328 ( .A1(n5370), .A2(n5371), .ZN(n9036) );
  NAND2_X1 U6329 ( .A1(n9071), .A2(n5035), .ZN(n5370) );
  NOR2_X1 U6330 ( .A1(n9069), .A2(n6012), .ZN(n9045) );
  NAND2_X1 U6331 ( .A1(n7940), .A2(n5374), .ZN(n5376) );
  NOR2_X1 U6332 ( .A1(n9165), .A2(n10817), .ZN(n8977) );
  XNOR2_X1 U6333 ( .A(n8975), .B(n8974), .ZN(n5382) );
  NAND2_X1 U6334 ( .A1(n5384), .A2(n10043), .ZN(n7915) );
  NAND2_X1 U6335 ( .A1(n8803), .A2(n9872), .ZN(n10315) );
  OAI21_X1 U6336 ( .B1(n10922), .B2(n5394), .A(n5392), .ZN(n8495) );
  NAND2_X1 U6337 ( .A1(n8784), .A2(n5410), .ZN(n5409) );
  INV_X1 U6338 ( .A(n5425), .ZN(n10455) );
  NAND2_X1 U6339 ( .A1(n10417), .A2(n5428), .ZN(n5427) );
  NAND2_X1 U6340 ( .A1(n8847), .A2(n8846), .ZN(n8832) );
  OAI211_X1 U6341 ( .C1(n8831), .C2(n5436), .A(n5433), .B(n5432), .ZN(n8815)
         );
  AOI21_X1 U6342 ( .B1(n8835), .B2(n5437), .A(n5095), .ZN(n5432) );
  NAND2_X1 U6343 ( .A1(n8847), .A2(n5434), .ZN(n5433) );
  INV_X1 U6344 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5614) );
  OAI21_X1 U6345 ( .B1(n6121), .B2(n5449), .A(n5448), .ZN(n6157) );
  NAND3_X1 U6346 ( .A1(n5447), .A2(n5446), .A3(n6156), .ZN(n6160) );
  NAND2_X1 U6347 ( .A1(n5448), .A2(n5449), .ZN(n5446) );
  NAND2_X1 U6348 ( .A1(n6121), .A2(n5448), .ZN(n5447) );
  NAND2_X1 U6349 ( .A1(n5911), .A2(n5453), .ZN(n5450) );
  NAND2_X1 U6350 ( .A1(n5450), .A2(n5452), .ZN(n5942) );
  NAND2_X1 U6351 ( .A1(n6050), .A2(n5464), .ZN(n5463) );
  NAND2_X1 U6352 ( .A1(n8998), .A2(n5487), .ZN(n5484) );
  NAND2_X1 U6353 ( .A1(n5484), .A2(n5485), .ZN(n8662) );
  NAND2_X1 U6354 ( .A1(n8998), .A2(n5492), .ZN(n5486) );
  NAND2_X2 U6355 ( .A1(n9050), .A2(n9049), .ZN(n9187) );
  INV_X1 U6356 ( .A(n8412), .ZN(n5502) );
  NAND2_X1 U6357 ( .A1(n6857), .A2(n6856), .ZN(n9701) );
  INV_X1 U6358 ( .A(n9702), .ZN(n5521) );
  OR2_X1 U6359 ( .A1(n6872), .A2(n6871), .ZN(n5522) );
  NAND2_X1 U6360 ( .A1(n6621), .A2(n5523), .ZN(n8030) );
  NAND3_X1 U6361 ( .A1(n8030), .A2(n8029), .A3(n8028), .ZN(n8027) );
  NAND2_X1 U6362 ( .A1(n6576), .A2(n6377), .ZN(n6426) );
  NAND2_X1 U6363 ( .A1(n5751), .A2(n5750), .ZN(n5759) );
  NAND2_X1 U6364 ( .A1(n6342), .A2(n6168), .ZN(n6341) );
  INV_X1 U6365 ( .A(n7545), .ZN(n6978) );
  NAND2_X1 U6366 ( .A1(n6082), .A2(n6081), .ZN(n6084) );
  NAND2_X1 U6367 ( .A1(n5034), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5607) );
  XNOR2_X1 U6368 ( .A(n6065), .B(n6066), .ZN(n8308) );
  INV_X1 U6369 ( .A(n6355), .ZN(n6356) );
  INV_X1 U6370 ( .A(n8901), .ZN(n7605) );
  INV_X1 U6371 ( .A(n6497), .ZN(n6644) );
  OR2_X1 U6372 ( .A1(n7804), .A2(n7802), .ZN(n7886) );
  OR2_X1 U6373 ( .A1(n7800), .A2(n10793), .ZN(n7802) );
  NAND2_X1 U6374 ( .A1(n10107), .A2(n6434), .ZN(n6454) );
  OR2_X1 U6375 ( .A1(n10281), .A2(n10280), .ZN(n10485) );
  AOI21_X1 U6376 ( .B1(n10297), .B2(n10481), .A(n10281), .ZN(n8795) );
  OR2_X1 U6377 ( .A1(n5638), .A2(n5596), .ZN(n5597) );
  NAND2_X1 U6378 ( .A1(n7723), .A2(n7722), .ZN(n7725) );
  NAND2_X1 U6379 ( .A1(n6494), .A2(n6492), .ZN(n7567) );
  NAND2_X4 U6380 ( .A1(n9698), .A2(n5579), .ZN(n5819) );
  XNOR2_X1 U6381 ( .A(n6522), .B(n6520), .ZN(n6524) );
  INV_X1 U6382 ( .A(n7567), .ZN(n6523) );
  NOR2_X1 U6383 ( .A1(n6473), .A2(n5053), .ZN(n6475) );
  NAND2_X1 U6384 ( .A1(n6524), .A2(n6523), .ZN(n7569) );
  INV_X1 U6385 ( .A(n9822), .ZN(n6792) );
  OR2_X1 U6386 ( .A1(n9822), .A2(n7181), .ZN(n6490) );
  OR2_X1 U6387 ( .A1(n6910), .A2(n10134), .ZN(n6483) );
  INV_X1 U6388 ( .A(n6910), .ZN(n6795) );
  OR2_X1 U6389 ( .A1(n6910), .A2(n6444), .ZN(n6445) );
  OAI211_X1 U6390 ( .C1(n6503), .C2(n7200), .A(n6562), .B(n6561), .ZN(n10826)
         );
  NAND2_X1 U6391 ( .A1(n6503), .A2(n10598), .ZN(n6460) );
  INV_X2 U6392 ( .A(n6484), .ZN(n6434) );
  OAI21_X1 U6393 ( .B1(n7149), .B2(n7148), .A(n9756), .ZN(n7153) );
  AND2_X1 U6394 ( .A1(n8723), .A2(n10904), .ZN(n10733) );
  AND2_X1 U6395 ( .A1(n6469), .A2(n6915), .ZN(n5548) );
  OR2_X1 U6396 ( .A1(n9057), .A2(n9034), .ZN(n5549) );
  OR2_X1 U6397 ( .A1(n10306), .A2(n9753), .ZN(n5550) );
  NOR2_X1 U6398 ( .A1(n5757), .A2(n5756), .ZN(n5551) );
  NOR2_X1 U6399 ( .A1(n5754), .A2(n5753), .ZN(n5552) );
  OR2_X1 U6400 ( .A1(n7433), .A2(n9004), .ZN(n5555) );
  OR2_X1 U6401 ( .A1(n6503), .A2(n7258), .ZN(n5556) );
  AND2_X1 U6402 ( .A1(n5856), .A2(n5840), .ZN(n5557) );
  INV_X1 U6403 ( .A(n7889), .ZN(n5722) );
  NOR2_X1 U6404 ( .A1(n10052), .A2(n8489), .ZN(n5559) );
  AND2_X1 U6405 ( .A1(n8901), .A2(n7606), .ZN(n5560) );
  INV_X1 U6406 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6461) );
  INV_X1 U6407 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5565) );
  INV_X1 U6408 ( .A(n5827), .ZN(n5832) );
  AND2_X1 U6409 ( .A1(n10004), .A2(n10351), .ZN(n10001) );
  AND2_X1 U6410 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  NAND2_X1 U6411 ( .A1(n6153), .A2(n5338), .ZN(n6154) );
  INV_X1 U6412 ( .A(n6057), .ZN(n6056) );
  INV_X1 U6413 ( .A(n7613), .ZN(n6318) );
  INV_X2 U6414 ( .A(n6854), .ZN(n6922) );
  OR2_X1 U6415 ( .A1(n6494), .A2(n6492), .ZN(n6495) );
  INV_X1 U6416 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6551) );
  AND2_X1 U6417 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n6409), .ZN(n6860) );
  NAND2_X1 U6418 ( .A1(n10764), .A2(n10104), .ZN(n9923) );
  INV_X1 U6419 ( .A(n5993), .ZN(n5995) );
  INV_X1 U6420 ( .A(n5888), .ZN(n5889) );
  INV_X1 U6421 ( .A(n7161), .ZN(n7025) );
  INV_X1 U6422 ( .A(n8867), .ZN(n7082) );
  OR2_X1 U6423 ( .A1(n5695), .A2(n7184), .ZN(n5621) );
  OR2_X1 U6424 ( .A1(n6104), .A2(n7133), .ZN(n6126) );
  OR2_X1 U6425 ( .A1(n6073), .A2(n9565), .ZN(n6088) );
  OR2_X1 U6426 ( .A1(n6004), .A2(n9557), .ZN(n6036) );
  NAND2_X1 U6427 ( .A1(n5879), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5903) );
  OAI21_X1 U6428 ( .B1(n8975), .B2(n6112), .A(n6175), .ZN(n8663) );
  NAND2_X1 U6429 ( .A1(n5958), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5974) );
  OR2_X1 U6430 ( .A1(n5903), .A2(n9323), .ZN(n5920) );
  INV_X1 U6431 ( .A(n6137), .ZN(n6161) );
  INV_X1 U6432 ( .A(n8660), .ZN(n8661) );
  INV_X1 U6433 ( .A(n6826), .ZN(n6845) );
  NOR2_X1 U6434 ( .A1(n6625), .A2(n8234), .ZN(n6663) );
  OR2_X1 U6435 ( .A1(n6831), .A2(n7246), .ZN(n6500) );
  NOR2_X1 U6436 ( .A1(n6736), .A2(n6735), .ZN(n6757) );
  NAND2_X1 U6437 ( .A1(n10086), .A2(n9916), .ZN(n7155) );
  AND2_X1 U6438 ( .A1(n9922), .A2(n9923), .ZN(n10765) );
  NAND2_X1 U6439 ( .A1(n6469), .A2(n8014), .ZN(n7970) );
  INV_X1 U6440 ( .A(n5872), .ZN(n5874) );
  INV_X1 U6441 ( .A(n9000), .ZN(n8879) );
  AND2_X1 U6442 ( .A1(n6126), .A2(n6105), .ZN(n8972) );
  OR2_X1 U6443 ( .A1(n9182), .A2(n8886), .ZN(n8657) );
  AND2_X1 U6444 ( .A1(n8649), .A2(n6248), .ZN(n8536) );
  INV_X1 U6445 ( .A(n10732), .ZN(n7739) );
  NAND2_X1 U6446 ( .A1(n7725), .A2(n7724), .ZN(n10791) );
  OR2_X1 U6447 ( .A1(n7423), .A2(n7422), .ZN(n7695) );
  INV_X1 U6448 ( .A(n10404), .ZN(n9722) );
  AOI21_X1 U6449 ( .B1(n10500), .B2(n6434), .A(n6431), .ZN(n9728) );
  XNOR2_X1 U6450 ( .A(n6519), .B(n6850), .ZN(n6527) );
  NAND2_X1 U6451 ( .A1(n9786), .A2(n9785), .ZN(n9784) );
  NOR2_X1 U6452 ( .A1(n10683), .A2(n10684), .ZN(n10681) );
  INV_X1 U6453 ( .A(n10508), .ZN(n10374) );
  OR2_X1 U6454 ( .A1(n7383), .A2(n10076), .ZN(n10990) );
  NAND2_X1 U6455 ( .A1(n5804), .A2(n5762), .ZN(n5767) );
  NOR2_X1 U6456 ( .A1(n7140), .A2(n10742), .ZN(n7141) );
  AND2_X1 U6457 ( .A1(n8840), .A2(n9137), .ZN(n10731) );
  NAND2_X1 U6458 ( .A1(n7031), .A2(n7168), .ZN(n8729) );
  OR2_X1 U6459 ( .A1(n8984), .A2(n6090), .ZN(n6096) );
  NAND2_X1 U6460 ( .A1(n6178), .A2(n6177), .ZN(n9019) );
  INV_X1 U6461 ( .A(n9133), .ZN(n9122) );
  INV_X1 U6462 ( .A(n10904), .ZN(n10998) );
  AND2_X1 U6463 ( .A1(n6361), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7700) );
  INV_X1 U6464 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5628) );
  AND4_X1 U6465 ( .A1(n6914), .A2(n6913), .A3(n6912), .A4(n6911), .ZN(n8790)
         );
  AND4_X1 U6466 ( .A1(n6835), .A2(n6834), .A3(n6833), .A4(n6832), .ZN(n10385)
         );
  NOR2_X1 U6467 ( .A1(n9918), .A2(n9910), .ZN(n10062) );
  OAI21_X1 U6468 ( .B1(n10314), .B2(n10316), .A(n10313), .ZN(n10492) );
  OAI22_X1 U6469 ( .A1(n10382), .A2(n8782), .B1(n10404), .B2(n10515), .ZN(
        n10367) );
  AND2_X1 U6470 ( .A1(n7264), .A2(n10033), .ZN(n10768) );
  INV_X1 U6471 ( .A(n10990), .ZN(n11033) );
  AOI21_X1 U6472 ( .B1(n10286), .B2(n10930), .A(n10285), .ZN(n10484) );
  AND2_X1 U6473 ( .A1(n6418), .A2(n6946), .ZN(n10588) );
  INV_X1 U6474 ( .A(n9916), .ZN(n6947) );
  XNOR2_X1 U6475 ( .A(n5731), .B(n9498), .ZN(n5753) );
  XNOR2_X1 U6476 ( .A(n5649), .B(n9509), .ZN(n5647) );
  NOR2_X1 U6477 ( .A1(n7142), .A2(n7141), .ZN(n7143) );
  OR2_X1 U6478 ( .A1(n6367), .A2(n6366), .ZN(n6368) );
  OR3_X1 U6479 ( .A1(n5964), .A2(n5963), .A3(n5962), .ZN(n9140) );
  INV_X1 U6480 ( .A(n11007), .ZN(n11006) );
  INV_X1 U6481 ( .A(n11011), .ZN(n11008) );
  INV_X1 U6482 ( .A(n10532), .ZN(n10442) );
  OR2_X1 U6483 ( .A1(n9764), .A2(n11029), .ZN(n9753) );
  AND4_X1 U6484 ( .A1(n6960), .A2(n6959), .A3(n6958), .A4(n6957), .ZN(n10284)
         );
  INV_X1 U6485 ( .A(n9830), .ZN(n10096) );
  INV_X1 U6486 ( .A(n7909), .ZN(n10101) );
  INV_X1 U6487 ( .A(n11036), .ZN(n11035) );
  INV_X1 U6488 ( .A(n11040), .ZN(n11037) );
  INV_X1 U6489 ( .A(n10600), .ZN(n10601) );
  INV_X1 U6490 ( .A(n10106), .ZN(P1_U4006) );
  NOR2_X1 U6491 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5564) );
  NAND4_X1 U6492 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .ZN(n5568)
         );
  NAND4_X1 U6493 ( .A1(n5709), .A2(n5841), .A3(n5566), .A4(n5565), .ZN(n5567)
         );
  NOR3_X1 U6494 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n5570) );
  NOR3_X1 U6495 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n5571) );
  INV_X1 U6496 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5572) );
  INV_X1 U6497 ( .A(n5575), .ZN(n5573) );
  INV_X1 U6498 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U6499 ( .A1(n5573), .A2(n5576), .ZN(n9690) );
  XNOR2_X2 U6500 ( .A(n5574), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U6501 ( .A1(n5575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5577) );
  INV_X1 U6502 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7289) );
  OR2_X1 U6503 ( .A1(n5819), .A2(n7289), .ZN(n5584) );
  NAND2_X2 U6504 ( .A1(n5578), .A2(n5031), .ZN(n5957) );
  NAND2_X1 U6505 ( .A1(n5637), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5583) );
  INV_X1 U6506 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7779) );
  INV_X1 U6507 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5580) );
  OR2_X1 U6508 ( .A1(n5638), .A2(n5580), .ZN(n5581) );
  NAND2_X1 U6509 ( .A1(n7182), .A2(SI_0_), .ZN(n5586) );
  INV_X1 U6510 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U6511 ( .A1(n5586), .A2(n5585), .ZN(n5588) );
  AND2_X1 U6512 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5587) );
  AND2_X1 U6513 ( .A1(n5588), .A2(n5606), .ZN(n9700) );
  MUX2_X1 U6514 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9700), .S(n7286), .Z(n7783) );
  INV_X1 U6515 ( .A(n7783), .ZN(n7513) );
  INV_X1 U6516 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5595) );
  INV_X1 U6517 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7704) );
  INV_X1 U6518 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U6519 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5601) );
  MUX2_X1 U6520 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5601), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5604) );
  INV_X1 U6521 ( .A(n5602), .ZN(n5603) );
  INV_X1 U6522 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7195) );
  AND2_X1 U6523 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U6524 ( .A1(n5650), .A2(n5605), .ZN(n6458) );
  NAND2_X1 U6525 ( .A1(n6458), .A2(n5606), .ZN(n5618) );
  XNOR2_X1 U6526 ( .A(n5618), .B(n9510), .ZN(n5617) );
  XNOR2_X1 U6527 ( .A(n5617), .B(n5616), .ZN(n7194) );
  INV_X1 U6528 ( .A(n7606), .ZN(n7710) );
  NAND2_X1 U6529 ( .A1(n8901), .A2(n7710), .ZN(n6316) );
  NAND2_X1 U6530 ( .A1(n7584), .A2(n6316), .ZN(n5608) );
  OR2_X1 U6531 ( .A1(n8901), .A2(n7710), .ZN(n6317) );
  NAND2_X1 U6532 ( .A1(n5608), .A2(n6317), .ZN(n7748) );
  NAND2_X1 U6533 ( .A1(n5637), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5613) );
  INV_X1 U6534 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7756) );
  INV_X1 U6535 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7306) );
  INV_X1 U6536 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5609) );
  OR2_X1 U6537 ( .A1(n5638), .A2(n5609), .ZN(n5610) );
  OR2_X1 U6538 ( .A1(n5602), .A2(n5645), .ZN(n5615) );
  XNOR2_X1 U6539 ( .A(n5615), .B(n5614), .ZN(n7332) );
  INV_X1 U6540 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7184) );
  NAND2_X1 U6541 ( .A1(n5618), .A2(SI_1_), .ZN(n5619) );
  MUX2_X1 U6542 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5650), .Z(n5632) );
  INV_X1 U6543 ( .A(SI_2_), .ZN(n9508) );
  XNOR2_X1 U6544 ( .A(n5632), .B(n9508), .ZN(n5631) );
  XNOR2_X1 U6545 ( .A(n5630), .B(n5631), .ZN(n7183) );
  OR2_X1 U6546 ( .A1(n6137), .A2(n7183), .ZN(n5620) );
  NAND2_X1 U6547 ( .A1(n10730), .A2(n7609), .ZN(n6187) );
  NAND2_X1 U6548 ( .A1(n7747), .A2(n7614), .ZN(n5636) );
  NAND2_X1 U6549 ( .A1(n5637), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5626) );
  OR2_X1 U6550 ( .A1(n6090), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5625) );
  INV_X1 U6551 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7323) );
  OR2_X1 U6552 ( .A1(n5819), .A2(n7323), .ZN(n5624) );
  INV_X1 U6553 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5622) );
  OR2_X1 U6554 ( .A1(n5638), .A2(n5622), .ZN(n5623) );
  OR2_X1 U6555 ( .A1(n5627), .A2(n5645), .ZN(n5629) );
  XNOR2_X1 U6556 ( .A(n5629), .B(n5628), .ZN(n7348) );
  INV_X1 U6557 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7187) );
  OR2_X1 U6558 ( .A1(n5695), .A2(n7187), .ZN(n5635) );
  NAND2_X1 U6559 ( .A1(n5632), .A2(SI_2_), .ZN(n5633) );
  MUX2_X1 U6560 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5034), .Z(n5649) );
  INV_X1 U6561 ( .A(SI_3_), .ZN(n9509) );
  XNOR2_X1 U6562 ( .A(n5648), .B(n5647), .ZN(n7186) );
  OR2_X1 U6563 ( .A1(n6137), .A2(n7186), .ZN(n5634) );
  OAI211_X1 U6564 ( .C1(n7286), .C2(n7348), .A(n5635), .B(n5634), .ZN(n10732)
         );
  NAND2_X1 U6565 ( .A1(n8900), .A2(n7739), .ZN(n6190) );
  NAND2_X1 U6566 ( .A1(n5636), .A2(n6318), .ZN(n7612) );
  NAND2_X1 U6567 ( .A1(n7612), .A2(n7716), .ZN(n5657) );
  NAND2_X1 U6568 ( .A1(n5637), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5643) );
  XNOR2_X1 U6569 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7726) );
  OR2_X1 U6570 ( .A1(n6090), .A2(n7726), .ZN(n5642) );
  INV_X1 U6571 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7407) );
  OR2_X1 U6572 ( .A1(n5819), .A2(n7407), .ZN(n5641) );
  INV_X1 U6573 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5639) );
  OR2_X1 U6574 ( .A1(n5638), .A2(n5639), .ZN(n5640) );
  NAND4_X1 U6575 ( .A1(n5643), .A2(n5642), .A3(n5641), .A4(n5640), .ZN(n8899)
         );
  OR2_X1 U6576 ( .A1(n5644), .A2(n5645), .ZN(n5646) );
  INV_X1 U6577 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5666) );
  XNOR2_X1 U6578 ( .A(n5646), .B(n5666), .ZN(n7416) );
  NAND2_X1 U6579 ( .A1(n5649), .A2(SI_3_), .ZN(n5670) );
  NAND2_X1 U6580 ( .A1(n5672), .A2(n5670), .ZN(n5653) );
  INV_X1 U6581 ( .A(SI_4_), .ZN(n9504) );
  XNOR2_X1 U6582 ( .A(n5653), .B(n5673), .ZN(n7189) );
  OR2_X1 U6583 ( .A1(n6137), .A2(n7189), .ZN(n5655) );
  OR2_X1 U6584 ( .A1(n5695), .A2(n5652), .ZN(n5654) );
  OAI211_X1 U6585 ( .C1(n7286), .C2(n7416), .A(n5655), .B(n5654), .ZN(n7727)
         );
  INV_X1 U6586 ( .A(n7727), .ZN(n10752) );
  XNOR2_X1 U6587 ( .A(n8899), .B(n10752), .ZN(n7724) );
  INV_X1 U6588 ( .A(n7724), .ZN(n5656) );
  NAND2_X1 U6589 ( .A1(n5657), .A2(n5656), .ZN(n7715) );
  INV_X1 U6590 ( .A(n8899), .ZN(n10737) );
  NAND2_X1 U6591 ( .A1(n10737), .A2(n7727), .ZN(n5658) );
  NAND2_X1 U6592 ( .A1(n7715), .A2(n5658), .ZN(n10796) );
  INV_X2 U6593 ( .A(n5638), .ZN(n5814) );
  NAND2_X1 U6594 ( .A1(n5814), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5665) );
  INV_X1 U6595 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5659) );
  OR2_X1 U6596 ( .A1(n5957), .A2(n5659), .ZN(n5664) );
  NAND3_X1 U6597 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5683) );
  INV_X1 U6598 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U6599 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5660) );
  NAND2_X1 U6600 ( .A1(n9543), .A2(n5660), .ZN(n5661) );
  NAND2_X1 U6601 ( .A1(n5683), .A2(n5661), .ZN(n10808) );
  OR2_X1 U6602 ( .A1(n6090), .A2(n10808), .ZN(n5663) );
  INV_X1 U6603 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7408) );
  OR2_X1 U6604 ( .A1(n5819), .A2(n7408), .ZN(n5662) );
  NAND2_X1 U6605 ( .A1(n5644), .A2(n5666), .ZN(n5712) );
  NAND2_X1 U6606 ( .A1(n5712), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5667) );
  INV_X1 U6607 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U6608 ( .A1(n5667), .A2(n5710), .ZN(n5689) );
  OR2_X1 U6609 ( .A1(n5667), .A2(n5710), .ZN(n5668) );
  NAND2_X1 U6610 ( .A1(n5689), .A2(n5668), .ZN(n7446) );
  NAND2_X1 U6611 ( .A1(n5669), .A2(SI_4_), .ZN(n5675) );
  AND2_X1 U6612 ( .A1(n5670), .A2(n5675), .ZN(n5671) );
  INV_X1 U6613 ( .A(n5673), .ZN(n5674) );
  MUX2_X1 U6614 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5034), .Z(n5693) );
  INV_X1 U6615 ( .A(SI_5_), .ZN(n9503) );
  OR2_X1 U6616 ( .A1(n6137), .A2(n7192), .ZN(n5679) );
  INV_X1 U6617 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7193) );
  OR2_X1 U6618 ( .A1(n5695), .A2(n7193), .ZN(n5678) );
  INV_X1 U6619 ( .A(n10806), .ZN(n10820) );
  NAND2_X1 U6620 ( .A1(n8898), .A2(n10820), .ZN(n5680) );
  NAND2_X1 U6621 ( .A1(n5681), .A2(n5680), .ZN(n10793) );
  INV_X1 U6622 ( .A(n10793), .ZN(n10797) );
  NAND2_X1 U6623 ( .A1(n10796), .A2(n10797), .ZN(n10795) );
  NAND2_X1 U6624 ( .A1(n5814), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5688) );
  INV_X1 U6625 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7791) );
  OR2_X1 U6626 ( .A1(n5957), .A2(n7791), .ZN(n5687) );
  INV_X1 U6627 ( .A(n5683), .ZN(n5682) );
  INV_X1 U6628 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U6629 ( .A1(n5683), .A2(n9564), .ZN(n5684) );
  NAND2_X1 U6630 ( .A1(n5703), .A2(n5684), .ZN(n8675) );
  OR2_X1 U6631 ( .A1(n6090), .A2(n8675), .ZN(n5686) );
  INV_X1 U6632 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7436) );
  OR2_X1 U6633 ( .A1(n5819), .A2(n7436), .ZN(n5685) );
  NAND4_X1 U6634 ( .A1(n5688), .A2(n5687), .A3(n5686), .A4(n5685), .ZN(n8897)
         );
  NAND2_X1 U6635 ( .A1(n5689), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5690) );
  XNOR2_X1 U6636 ( .A(n5690), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7493) );
  INV_X1 U6637 ( .A(n7493), .ZN(n7196) );
  NAND2_X1 U6638 ( .A1(n5693), .A2(SI_5_), .ZN(n5694) );
  MUX2_X1 U6639 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5034), .Z(n5719) );
  INV_X1 U6640 ( .A(SI_6_), .ZN(n9499) );
  XNOR2_X1 U6641 ( .A(n5718), .B(n5717), .ZN(n7199) );
  OR2_X1 U6642 ( .A1(n6137), .A2(n7199), .ZN(n5697) );
  INV_X1 U6643 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7197) );
  OR2_X1 U6644 ( .A1(n5695), .A2(n7197), .ZN(n5696) );
  OAI211_X1 U6645 ( .C1(n7286), .C2(n7196), .A(n5697), .B(n5696), .ZN(n7796)
         );
  INV_X1 U6646 ( .A(n7796), .ZN(n10838) );
  NAND2_X1 U6647 ( .A1(n8897), .A2(n10838), .ZN(n5698) );
  INV_X1 U6648 ( .A(n8897), .ZN(n5699) );
  NAND2_X1 U6649 ( .A1(n5699), .A2(n7796), .ZN(n5700) );
  NAND2_X1 U6650 ( .A1(n5814), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5708) );
  INV_X1 U6651 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7892) );
  OR2_X1 U6652 ( .A1(n5957), .A2(n7892), .ZN(n5707) );
  INV_X1 U6653 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6654 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NAND2_X1 U6655 ( .A1(n5724), .A2(n5704), .ZN(n7966) );
  OR2_X1 U6656 ( .A1(n6090), .A2(n7966), .ZN(n5706) );
  INV_X1 U6657 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7439) );
  OR2_X1 U6658 ( .A1(n5819), .A2(n7439), .ZN(n5705) );
  NAND4_X1 U6659 ( .A1(n5708), .A2(n5707), .A3(n5706), .A4(n5705), .ZN(n8896)
         );
  NAND2_X1 U6660 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  NOR2_X1 U6661 ( .A1(n5712), .A2(n5711), .ZN(n5715) );
  OR2_X1 U6662 ( .A1(n5715), .A2(n5645), .ZN(n5713) );
  MUX2_X1 U6663 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5713), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5716) );
  INV_X1 U6664 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U6665 ( .A1(n5715), .A2(n5714), .ZN(n5763) );
  NAND2_X1 U6666 ( .A1(n5716), .A2(n5763), .ZN(n7445) );
  NAND2_X1 U6667 ( .A1(n5719), .A2(SI_6_), .ZN(n5749) );
  MUX2_X1 U6668 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5034), .Z(n5731) );
  INV_X1 U6669 ( .A(SI_7_), .ZN(n9498) );
  XNOR2_X1 U6670 ( .A(n5730), .B(n5753), .ZN(n7202) );
  OR2_X1 U6671 ( .A1(n7202), .A2(n6137), .ZN(n5721) );
  INV_X1 U6672 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7203) );
  OR2_X1 U6673 ( .A1(n5695), .A2(n7203), .ZN(n5720) );
  OAI211_X1 U6674 ( .C1(n7286), .C2(n7445), .A(n5721), .B(n5720), .ZN(n7894)
         );
  OR2_X1 U6675 ( .A1(n8896), .A2(n10853), .ZN(n6204) );
  NAND2_X1 U6676 ( .A1(n8896), .A2(n10853), .ZN(n7941) );
  NAND2_X1 U6677 ( .A1(n6204), .A2(n7941), .ZN(n7889) );
  NAND2_X1 U6678 ( .A1(n5814), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5729) );
  INV_X1 U6679 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7948) );
  OR2_X1 U6680 ( .A1(n5957), .A2(n7948), .ZN(n5728) );
  INV_X1 U6681 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U6682 ( .A1(n5724), .A2(n9528), .ZN(n5725) );
  NAND2_X1 U6683 ( .A1(n5741), .A2(n5725), .ZN(n8146) );
  OR2_X1 U6684 ( .A1(n6090), .A2(n8146), .ZN(n5727) );
  INV_X1 U6685 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7440) );
  OR2_X1 U6686 ( .A1(n5819), .A2(n7440), .ZN(n5726) );
  NAND4_X1 U6687 ( .A1(n5729), .A2(n5728), .A3(n5727), .A4(n5726), .ZN(n8895)
         );
  NAND2_X1 U6688 ( .A1(n5730), .A2(n5753), .ZN(n5732) );
  NAND2_X1 U6689 ( .A1(n5731), .A2(SI_7_), .ZN(n5748) );
  NAND2_X1 U6690 ( .A1(n5732), .A2(n5748), .ZN(n5734) );
  MUX2_X1 U6691 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5034), .Z(n5747) );
  INV_X1 U6692 ( .A(SI_8_), .ZN(n5733) );
  XNOR2_X1 U6693 ( .A(n5747), .B(n5733), .ZN(n5756) );
  XNOR2_X1 U6694 ( .A(n5734), .B(n5756), .ZN(n7206) );
  OR2_X1 U6695 ( .A1(n7206), .A2(n6137), .ZN(n5737) );
  NAND2_X1 U6696 ( .A1(n5763), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5735) );
  XNOR2_X1 U6697 ( .A(n5735), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7476) );
  AOI22_X1 U6698 ( .A1(n5953), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5952), .B2(
        n7476), .ZN(n5736) );
  OR2_X1 U6699 ( .A1(n8895), .A2(n10868), .ZN(n6206) );
  NAND2_X1 U6700 ( .A1(n8895), .A2(n10868), .ZN(n8187) );
  NAND2_X1 U6701 ( .A1(n6206), .A2(n8187), .ZN(n7956) );
  AND2_X1 U6702 ( .A1(n7956), .A2(n7941), .ZN(n5738) );
  INV_X1 U6703 ( .A(n8895), .ZN(n8094) );
  NAND2_X1 U6704 ( .A1(n8094), .A2(n10868), .ZN(n5739) );
  NAND2_X1 U6705 ( .A1(n5814), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5746) );
  INV_X1 U6706 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8197) );
  OR2_X1 U6707 ( .A1(n5957), .A2(n8197), .ZN(n5745) );
  INV_X1 U6708 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U6709 ( .A1(n5741), .A2(n9552), .ZN(n5742) );
  NAND2_X1 U6710 ( .A1(n5816), .A2(n5742), .ZN(n8196) );
  OR2_X1 U6711 ( .A1(n6090), .A2(n8196), .ZN(n5744) );
  INV_X1 U6712 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7470) );
  OR2_X1 U6713 ( .A1(n5819), .A2(n7470), .ZN(n5743) );
  NAND4_X1 U6714 ( .A1(n5746), .A2(n5745), .A3(n5744), .A4(n5743), .ZN(n8894)
         );
  INV_X1 U6715 ( .A(n8894), .ZN(n5766) );
  NAND2_X1 U6716 ( .A1(n5747), .A2(SI_8_), .ZN(n5755) );
  AND2_X1 U6717 ( .A1(n5749), .A2(n5752), .ZN(n5750) );
  INV_X1 U6718 ( .A(n5752), .ZN(n5754) );
  INV_X1 U6719 ( .A(n5755), .ZN(n5757) );
  INV_X1 U6720 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7211) );
  INV_X1 U6721 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9383) );
  MUX2_X1 U6722 ( .A(n7211), .B(n9383), .S(n5034), .Z(n5760) );
  INV_X1 U6723 ( .A(SI_9_), .ZN(n9490) );
  INV_X1 U6724 ( .A(n5760), .ZN(n5761) );
  NAND2_X1 U6725 ( .A1(n5761), .A2(SI_9_), .ZN(n5762) );
  XNOR2_X1 U6726 ( .A(n5768), .B(n5767), .ZN(n7208) );
  NAND2_X1 U6727 ( .A1(n7208), .A2(n6161), .ZN(n5765) );
  NAND2_X1 U6728 ( .A1(n5781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U6729 ( .A(n5809), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7537) );
  AOI22_X1 U6730 ( .A1(n5953), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5952), .B2(
        n7537), .ZN(n5764) );
  NAND2_X1 U6731 ( .A1(n5766), .A2(n10879), .ZN(n6217) );
  NAND2_X1 U6732 ( .A1(n8242), .A2(n6217), .ZN(n8190) );
  INV_X1 U6733 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5769) );
  INV_X1 U6734 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9384) );
  MUX2_X1 U6735 ( .A(n5769), .B(n9384), .S(n5034), .Z(n5771) );
  INV_X1 U6736 ( .A(SI_10_), .ZN(n5770) );
  NAND2_X1 U6737 ( .A1(n5771), .A2(n5770), .ZN(n5806) );
  NAND2_X1 U6738 ( .A1(n5831), .A2(n5830), .ZN(n5791) );
  INV_X1 U6739 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U6740 ( .A1(n5772), .A2(SI_10_), .ZN(n5805) );
  NAND2_X1 U6741 ( .A1(n5774), .A2(SI_11_), .ZN(n5775) );
  AND2_X1 U6742 ( .A1(n5791), .A2(n5833), .ZN(n5776) );
  INV_X1 U6743 ( .A(SI_11_), .ZN(n5773) );
  NOR2_X1 U6744 ( .A1(n5776), .A2(n5828), .ZN(n5780) );
  INV_X1 U6745 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7239) );
  INV_X1 U6746 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9382) );
  MUX2_X1 U6747 ( .A(n7239), .B(n9382), .S(n5034), .Z(n5777) );
  INV_X1 U6748 ( .A(SI_12_), .ZN(n9489) );
  INV_X1 U6749 ( .A(n5777), .ZN(n5778) );
  NAND2_X1 U6750 ( .A1(n5778), .A2(SI_12_), .ZN(n5779) );
  XNOR2_X1 U6751 ( .A(n5780), .B(n5827), .ZN(n7234) );
  NAND2_X1 U6752 ( .A1(n7234), .A2(n6161), .ZN(n5783) );
  OAI21_X1 U6753 ( .B1(n5794), .B2(P2_IR_REG_11__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5858) );
  XNOR2_X1 U6754 ( .A(n5858), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7768) );
  AOI22_X1 U6755 ( .A1(n5953), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5952), .B2(
        n7768), .ZN(n5782) );
  NAND2_X1 U6756 ( .A1(n5814), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5790) );
  INV_X1 U6757 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8603) );
  OR2_X1 U6758 ( .A1(n5957), .A2(n8603), .ZN(n5789) );
  INV_X1 U6759 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5815) );
  INV_X1 U6760 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7172) );
  INV_X1 U6761 ( .A(n5799), .ZN(n5784) );
  INV_X1 U6762 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U6763 ( .A1(n5799), .A2(n9536), .ZN(n5785) );
  NAND2_X1 U6764 ( .A1(n5847), .A2(n5785), .ZN(n8602) );
  OR2_X1 U6765 ( .A1(n6090), .A2(n8602), .ZN(n5788) );
  INV_X1 U6766 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5786) );
  OR2_X1 U6767 ( .A1(n5819), .A2(n5786), .ZN(n5787) );
  NAND4_X1 U6768 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n8891)
         );
  NAND2_X1 U6769 ( .A1(n8609), .A2(n8703), .ZN(n6222) );
  NAND2_X1 U6770 ( .A1(n7229), .A2(n6161), .ZN(n5797) );
  NAND2_X1 U6771 ( .A1(n5794), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  XNOR2_X1 U6772 ( .A(n5795), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7652) );
  AOI22_X1 U6773 ( .A1(n5953), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5952), .B2(
        n7652), .ZN(n5796) );
  NAND2_X1 U6774 ( .A1(n5814), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5803) );
  INV_X1 U6775 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7660) );
  OR2_X1 U6776 ( .A1(n5957), .A2(n7660), .ZN(n5802) );
  NAND2_X1 U6777 ( .A1(n5818), .A2(n7172), .ZN(n5798) );
  NAND2_X1 U6778 ( .A1(n5799), .A2(n5798), .ZN(n8283) );
  OR2_X1 U6779 ( .A1(n6090), .A2(n8283), .ZN(n5801) );
  INV_X1 U6780 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7555) );
  OR2_X1 U6781 ( .A1(n5819), .A2(n7555), .ZN(n5800) );
  NAND4_X1 U6782 ( .A1(n5803), .A2(n5802), .A3(n5801), .A4(n5800), .ZN(n8892)
         );
  NAND2_X1 U6783 ( .A1(n10905), .A2(n8320), .ZN(n8611) );
  AND2_X1 U6784 ( .A1(n6222), .A2(n8611), .ZN(n6227) );
  AND2_X1 U6785 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  NAND2_X1 U6786 ( .A1(n7223), .A2(n6161), .ZN(n5813) );
  INV_X1 U6787 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U6788 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  NAND2_X1 U6789 ( .A1(n5810), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5811) );
  XNOR2_X1 U6790 ( .A(n5811), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7556) );
  AOI22_X1 U6791 ( .A1(n5953), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5952), .B2(
        n7556), .ZN(n5812) );
  NAND2_X1 U6792 ( .A1(n5814), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5823) );
  INV_X1 U6793 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8249) );
  OR2_X1 U6794 ( .A1(n5957), .A2(n8249), .ZN(n5822) );
  NAND2_X1 U6795 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  NAND2_X1 U6796 ( .A1(n5818), .A2(n5817), .ZN(n8248) );
  OR2_X1 U6797 ( .A1(n6090), .A2(n8248), .ZN(n5821) );
  INV_X1 U6798 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7530) );
  OR2_X1 U6799 ( .A1(n5819), .A2(n7530), .ZN(n5820) );
  NAND4_X1 U6800 ( .A1(n5823), .A2(n5822), .A3(n5821), .A4(n5820), .ZN(n8893)
         );
  INV_X1 U6801 ( .A(n8893), .ZN(n8099) );
  NAND2_X1 U6802 ( .A1(n8257), .A2(n8099), .ZN(n6216) );
  NAND2_X1 U6803 ( .A1(n6227), .A2(n8274), .ZN(n5824) );
  OR2_X1 U6804 ( .A1(n8190), .A2(n5824), .ZN(n5826) );
  AND2_X1 U6805 ( .A1(n8242), .A2(n6219), .ZN(n8272) );
  OR2_X1 U6806 ( .A1(n5824), .A2(n8272), .ZN(n5825) );
  INV_X1 U6807 ( .A(n5835), .ZN(n5829) );
  INV_X1 U6808 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7232) );
  INV_X1 U6809 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9603) );
  MUX2_X1 U6810 ( .A(n7232), .B(n9603), .S(n5034), .Z(n5838) );
  INV_X1 U6811 ( .A(SI_13_), .ZN(n9485) );
  NAND2_X1 U6812 ( .A1(n5838), .A2(n9485), .ZN(n5856) );
  INV_X1 U6813 ( .A(n5838), .ZN(n5839) );
  NAND2_X1 U6814 ( .A1(n5839), .A2(SI_13_), .ZN(n5840) );
  XNOR2_X1 U6815 ( .A(n5855), .B(n5557), .ZN(n7227) );
  NAND2_X1 U6816 ( .A1(n7227), .A2(n6161), .ZN(n5845) );
  NAND2_X1 U6817 ( .A1(n5858), .A2(n5841), .ZN(n5842) );
  NAND2_X1 U6818 ( .A1(n5842), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5843) );
  XNOR2_X1 U6819 ( .A(n5843), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7930) );
  AOI22_X1 U6820 ( .A1(n5953), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5952), .B2(
        n7930), .ZN(n5844) );
  NAND2_X1 U6821 ( .A1(n5845), .A2(n5844), .ZN(n8713) );
  NAND2_X1 U6822 ( .A1(n5814), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5853) );
  INV_X1 U6823 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8324) );
  OR2_X1 U6824 ( .A1(n5957), .A2(n8324), .ZN(n5852) );
  INV_X1 U6825 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U6826 ( .A1(n5847), .A2(n9337), .ZN(n5848) );
  NAND2_X1 U6827 ( .A1(n5862), .A2(n5848), .ZN(n8706) );
  OR2_X1 U6828 ( .A1(n6090), .A2(n8706), .ZN(n5851) );
  INV_X1 U6829 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5849) );
  OR2_X1 U6830 ( .A1(n5819), .A2(n5849), .ZN(n5850) );
  NAND4_X1 U6831 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n8890)
         );
  INV_X1 U6832 ( .A(n8890), .ZN(n8733) );
  OR2_X1 U6833 ( .A1(n8713), .A2(n8733), .ZN(n6233) );
  NAND2_X1 U6834 ( .A1(n8713), .A2(n8733), .ZN(n8386) );
  NAND2_X1 U6835 ( .A1(n6233), .A2(n8386), .ZN(n8321) );
  INV_X1 U6836 ( .A(n8321), .ZN(n8313) );
  OR2_X1 U6837 ( .A1(n8609), .A2(n8703), .ZN(n6225) );
  OR2_X1 U6838 ( .A1(n10905), .A2(n8320), .ZN(n8610) );
  NAND2_X1 U6839 ( .A1(n6225), .A2(n8610), .ZN(n5854) );
  NAND2_X1 U6840 ( .A1(n5854), .A2(n6222), .ZN(n8314) );
  MUX2_X1 U6841 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5034), .Z(n5873) );
  INV_X1 U6842 ( .A(SI_14_), .ZN(n9484) );
  OAI21_X1 U6843 ( .B1(P2_IR_REG_12__SCAN_IN), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U6844 ( .A1(n5858), .A2(n5857), .ZN(n5875) );
  INV_X1 U6845 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5859) );
  XNOR2_X1 U6846 ( .A(n5875), .B(n5859), .ZN(n8215) );
  AOI22_X1 U6847 ( .A1(n5953), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5952), .B2(
        n8215), .ZN(n5860) );
  NAND2_X1 U6848 ( .A1(n5814), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5868) );
  INV_X1 U6849 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8383) );
  OR2_X1 U6850 ( .A1(n5957), .A2(n8383), .ZN(n5867) );
  INV_X1 U6851 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U6852 ( .A1(n5862), .A2(n9520), .ZN(n5863) );
  NAND2_X1 U6853 ( .A1(n5881), .A2(n5863), .ZN(n8736) );
  OR2_X1 U6854 ( .A1(n6090), .A2(n8736), .ZN(n5866) );
  INV_X1 U6855 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5864) );
  OR2_X1 U6856 ( .A1(n5819), .A2(n5864), .ZN(n5865) );
  NAND4_X1 U6857 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(n8889)
         );
  NAND2_X1 U6858 ( .A1(n8744), .A2(n8747), .ZN(n6236) );
  INV_X1 U6859 ( .A(n8382), .ZN(n8388) );
  INV_X1 U6860 ( .A(n8386), .ZN(n5869) );
  NOR2_X1 U6861 ( .A1(n8388), .A2(n5869), .ZN(n5871) );
  INV_X1 U6862 ( .A(n6237), .ZN(n5870) );
  MUX2_X1 U6863 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5034), .Z(n5891) );
  XNOR2_X1 U6864 ( .A(n5890), .B(n5888), .ZN(n7373) );
  NAND2_X1 U6865 ( .A1(n7373), .A2(n6161), .ZN(n5878) );
  OAI21_X1 U6866 ( .B1(n5875), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5876) );
  XNOR2_X1 U6867 ( .A(n5876), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8394) );
  AOI22_X1 U6868 ( .A1(n5953), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5952), .B2(
        n8394), .ZN(n5877) );
  NAND2_X1 U6869 ( .A1(n5814), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5887) );
  INV_X1 U6870 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8418) );
  OR2_X1 U6871 ( .A1(n5957), .A2(n8418), .ZN(n5886) );
  INV_X1 U6872 ( .A(n5881), .ZN(n5879) );
  INV_X1 U6873 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U6874 ( .A1(n5881), .A2(n5880), .ZN(n5882) );
  NAND2_X1 U6875 ( .A1(n5903), .A2(n5882), .ZN(n8752) );
  OR2_X1 U6876 ( .A1(n6090), .A2(n8752), .ZN(n5885) );
  INV_X1 U6877 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5883) );
  OR2_X1 U6878 ( .A1(n5819), .A2(n5883), .ZN(n5884) );
  NAND4_X1 U6879 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n8888)
         );
  NAND2_X1 U6880 ( .A1(n5891), .A2(SI_15_), .ZN(n5892) );
  INV_X1 U6881 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5894) );
  INV_X1 U6882 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9600) );
  MUX2_X1 U6883 ( .A(n5894), .B(n9600), .S(n5034), .Z(n5896) );
  INV_X1 U6884 ( .A(SI_16_), .ZN(n5895) );
  NAND2_X1 U6885 ( .A1(n5896), .A2(n5895), .ZN(n5913) );
  INV_X1 U6886 ( .A(n5896), .ZN(n5897) );
  NAND2_X1 U6887 ( .A1(n5897), .A2(SI_16_), .ZN(n5898) );
  NAND2_X1 U6888 ( .A1(n5913), .A2(n5898), .ZN(n5912) );
  XNOR2_X1 U6889 ( .A(n5911), .B(n5912), .ZN(n7401) );
  NAND2_X1 U6890 ( .A1(n7401), .A2(n6161), .ZN(n5902) );
  NAND2_X1 U6891 ( .A1(n5899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U6892 ( .A(n5900), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8914) );
  AOI22_X1 U6893 ( .A1(n5953), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5952), .B2(
        n8914), .ZN(n5901) );
  NAND2_X1 U6894 ( .A1(n5814), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5908) );
  INV_X1 U6895 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8520) );
  OR2_X1 U6896 ( .A1(n5957), .A2(n8520), .ZN(n5907) );
  INV_X1 U6897 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U6898 ( .A1(n5903), .A2(n9323), .ZN(n5904) );
  NAND2_X1 U6899 ( .A1(n5920), .A2(n5904), .ZN(n8690) );
  OR2_X1 U6900 ( .A1(n6090), .A2(n8690), .ZN(n5906) );
  INV_X1 U6901 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8905) );
  OR2_X1 U6902 ( .A1(n5819), .A2(n8905), .ZN(n5905) );
  NAND4_X1 U6903 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(n8887)
         );
  INV_X1 U6904 ( .A(n8887), .ZN(n8414) );
  NAND2_X1 U6905 ( .A1(n9229), .A2(n8414), .ZN(n6242) );
  INV_X1 U6906 ( .A(n6242), .ZN(n5910) );
  NAND2_X1 U6907 ( .A1(n8760), .A2(n8687), .ZN(n6240) );
  INV_X1 U6908 ( .A(n6240), .ZN(n5909) );
  OR2_X1 U6909 ( .A1(n9229), .A2(n8414), .ZN(n6243) );
  MUX2_X1 U6910 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5034), .Z(n5927) );
  INV_X1 U6911 ( .A(SI_17_), .ZN(n5914) );
  XNOR2_X1 U6912 ( .A(n5927), .B(n5914), .ZN(n5926) );
  XNOR2_X1 U6913 ( .A(n5929), .B(n5926), .ZN(n7502) );
  NAND2_X1 U6914 ( .A1(n7502), .A2(n6161), .ZN(n5918) );
  NAND2_X1 U6915 ( .A1(n5915), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5916) );
  XNOR2_X1 U6916 ( .A(n5916), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8924) );
  AOI22_X1 U6917 ( .A1(n5953), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5952), .B2(
        n8924), .ZN(n5917) );
  NAND2_X1 U6918 ( .A1(n5814), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5925) );
  INV_X1 U6919 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8540) );
  OR2_X1 U6920 ( .A1(n5957), .A2(n8540), .ZN(n5924) );
  INV_X1 U6921 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U6922 ( .A1(n5920), .A2(n9327), .ZN(n5921) );
  NAND2_X1 U6923 ( .A1(n5933), .A2(n5921), .ZN(n8539) );
  OR2_X1 U6924 ( .A1(n6090), .A2(n8539), .ZN(n5923) );
  INV_X1 U6925 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8931) );
  OR2_X1 U6926 ( .A1(n5819), .A2(n8931), .ZN(n5922) );
  NAND4_X1 U6927 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n9138)
         );
  NAND2_X1 U6928 ( .A1(n9223), .A2(n9138), .ZN(n6248) );
  INV_X1 U6929 ( .A(n9138), .ZN(n6247) );
  INV_X1 U6930 ( .A(n5926), .ZN(n5928) );
  MUX2_X1 U6931 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5034), .Z(n5943) );
  XNOR2_X1 U6932 ( .A(n5943), .B(SI_18_), .ZN(n5940) );
  XNOR2_X1 U6933 ( .A(n5942), .B(n5940), .ZN(n7579) );
  NAND2_X1 U6934 ( .A1(n7579), .A2(n6161), .ZN(n5931) );
  XNOR2_X1 U6935 ( .A(n5950), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8939) );
  AOI22_X1 U6936 ( .A1(n5953), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5952), .B2(
        n8939), .ZN(n5930) );
  NAND2_X1 U6937 ( .A1(n5814), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5938) );
  INV_X1 U6938 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8944) );
  OR2_X1 U6939 ( .A1(n5957), .A2(n8944), .ZN(n5937) );
  INV_X1 U6940 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U6941 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  NAND2_X1 U6942 ( .A1(n5960), .A2(n5934), .ZN(n9129) );
  OR2_X1 U6943 ( .A1(n6090), .A2(n9129), .ZN(n5936) );
  INV_X1 U6944 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8933) );
  OR2_X1 U6945 ( .A1(n5819), .A2(n8933), .ZN(n5935) );
  NAND4_X1 U6946 ( .A1(n5938), .A2(n5937), .A3(n5936), .A4(n5935), .ZN(n9109)
         );
  INV_X1 U6947 ( .A(n9109), .ZN(n8651) );
  NAND2_X1 U6948 ( .A1(n9216), .A2(n8651), .ZN(n6253) );
  INV_X1 U6949 ( .A(n9135), .ZN(n9125) );
  INV_X1 U6950 ( .A(n6254), .ZN(n5939) );
  INV_X1 U6951 ( .A(n5940), .ZN(n5941) );
  NAND2_X1 U6952 ( .A1(n5943), .A2(SI_18_), .ZN(n5944) );
  INV_X1 U6953 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7627) );
  INV_X1 U6954 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7625) );
  MUX2_X1 U6955 ( .A(n7627), .B(n7625), .S(n5034), .Z(n5946) );
  INV_X1 U6956 ( .A(SI_19_), .ZN(n9268) );
  NAND2_X1 U6957 ( .A1(n5946), .A2(n9268), .ZN(n5967) );
  INV_X1 U6958 ( .A(n5946), .ZN(n5947) );
  NAND2_X1 U6959 ( .A1(n5947), .A2(SI_19_), .ZN(n5948) );
  NAND2_X1 U6960 ( .A1(n5967), .A2(n5948), .ZN(n5965) );
  XNOR2_X1 U6961 ( .A(n5966), .B(n5965), .ZN(n7624) );
  NAND2_X1 U6962 ( .A1(n7624), .A2(n6161), .ZN(n5955) );
  INV_X1 U6963 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U6964 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  NAND2_X1 U6965 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6166) );
  XNOR2_X1 U6966 ( .A(n6166), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U6967 ( .A1(n5953), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10812), 
        .B2(n5952), .ZN(n5954) );
  INV_X1 U6968 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U6969 ( .A1(n5814), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5956) );
  OAI21_X1 U6970 ( .B1(n5957), .B2(n9116), .A(n5956), .ZN(n5964) );
  INV_X1 U6971 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U6972 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  NAND2_X1 U6973 ( .A1(n5974), .A2(n5961), .ZN(n9115) );
  NOR2_X1 U6974 ( .A1(n9115), .A2(n6090), .ZN(n5963) );
  INV_X1 U6975 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8950) );
  NOR2_X1 U6976 ( .A1(n5819), .A2(n8950), .ZN(n5962) );
  NAND2_X1 U6977 ( .A1(n9211), .A2(n8652), .ZN(n6259) );
  NAND2_X1 U6978 ( .A1(n6258), .A2(n6259), .ZN(n9112) );
  INV_X1 U6979 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7810) );
  INV_X1 U6980 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9592) );
  MUX2_X1 U6981 ( .A(n7810), .B(n9592), .S(n5034), .Z(n5968) );
  INV_X1 U6982 ( .A(SI_20_), .ZN(n9453) );
  NAND2_X1 U6983 ( .A1(n5968), .A2(n9453), .ZN(n5983) );
  INV_X1 U6984 ( .A(n5968), .ZN(n5969) );
  NAND2_X1 U6985 ( .A1(n5969), .A2(SI_20_), .ZN(n5970) );
  XNOR2_X1 U6986 ( .A(n5982), .B(n5981), .ZN(n7809) );
  NAND2_X1 U6987 ( .A1(n7809), .A2(n6161), .ZN(n5972) );
  OR2_X1 U6988 ( .A1(n5695), .A2(n7810), .ZN(n5971) );
  INV_X1 U6989 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5980) );
  INV_X1 U6990 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U6991 ( .A1(n5974), .A2(n9556), .ZN(n5975) );
  NAND2_X1 U6992 ( .A1(n5987), .A2(n5975), .ZN(n8859) );
  OR2_X1 U6993 ( .A1(n8859), .A2(n6090), .ZN(n5979) );
  NAND2_X1 U6994 ( .A1(n5637), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U6995 ( .A1(n5814), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5976) );
  AND2_X1 U6996 ( .A1(n5977), .A2(n5976), .ZN(n5978) );
  OAI211_X1 U6997 ( .C1(n5819), .C2(n5980), .A(n5979), .B(n5978), .ZN(n9110)
         );
  INV_X1 U6998 ( .A(n9110), .ZN(n8653) );
  NAND2_X1 U6999 ( .A1(n9204), .A2(n8653), .ZN(n6262) );
  NAND2_X1 U7000 ( .A1(n6263), .A2(n6262), .ZN(n9100) );
  INV_X1 U7001 ( .A(n9100), .ZN(n6329) );
  MUX2_X1 U7002 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5034), .Z(n5996) );
  INV_X1 U7003 ( .A(SI_21_), .ZN(n9267) );
  XNOR2_X1 U7004 ( .A(n5996), .B(n9267), .ZN(n5994) );
  XNOR2_X1 U7005 ( .A(n5993), .B(n5994), .ZN(n7823) );
  NAND2_X1 U7006 ( .A1(n7823), .A2(n6161), .ZN(n5986) );
  INV_X1 U7007 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7824) );
  OR2_X1 U7008 ( .A1(n5695), .A2(n7824), .ZN(n5985) );
  INV_X1 U7009 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5992) );
  INV_X1 U7010 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U7011 ( .A1(n5987), .A2(n9318), .ZN(n5988) );
  NAND2_X1 U7012 ( .A1(n6004), .A2(n5988), .ZN(n8824) );
  OR2_X1 U7013 ( .A1(n8824), .A2(n6090), .ZN(n5991) );
  INV_X1 U7014 ( .A(n5819), .ZN(n5989) );
  AOI22_X1 U7015 ( .A1(n5989), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5637), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5990) );
  OAI211_X1 U7016 ( .C1(n5638), .C2(n5992), .A(n5991), .B(n5990), .ZN(n9102)
         );
  INV_X1 U7017 ( .A(n9102), .ZN(n9068) );
  INV_X1 U7018 ( .A(n9199), .ZN(n9086) );
  NAND2_X1 U7019 ( .A1(n5995), .A2(n5994), .ZN(n5998) );
  NAND2_X1 U7020 ( .A1(n5996), .A2(SI_21_), .ZN(n5997) );
  INV_X1 U7021 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8041) );
  INV_X1 U7022 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9588) );
  MUX2_X1 U7023 ( .A(n8041), .B(n9588), .S(n5034), .Z(n5999) );
  INV_X1 U7024 ( .A(SI_22_), .ZN(n9476) );
  NAND2_X1 U7025 ( .A1(n5999), .A2(n9476), .ZN(n6015) );
  INV_X1 U7026 ( .A(n5999), .ZN(n6000) );
  NAND2_X1 U7027 ( .A1(n6000), .A2(SI_22_), .ZN(n6001) );
  NAND2_X1 U7028 ( .A1(n6015), .A2(n6001), .ZN(n6013) );
  XNOR2_X1 U7029 ( .A(n6014), .B(n6013), .ZN(n8038) );
  NAND2_X1 U7030 ( .A1(n8038), .A2(n6161), .ZN(n6003) );
  OR2_X1 U7031 ( .A1(n5695), .A2(n8041), .ZN(n6002) );
  INV_X1 U7032 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U7033 ( .A1(n6004), .A2(n9557), .ZN(n6005) );
  AND2_X1 U7034 ( .A1(n6036), .A2(n6005), .ZN(n9064) );
  INV_X1 U7035 ( .A(n6090), .ZN(n6131) );
  NAND2_X1 U7036 ( .A1(n9064), .A2(n6131), .ZN(n6011) );
  INV_X1 U7037 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7038 ( .A1(n5637), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7039 ( .A1(n5814), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6006) );
  OAI211_X1 U7040 ( .C1(n5819), .C2(n6008), .A(n6007), .B(n6006), .ZN(n6009)
         );
  INV_X1 U7041 ( .A(n6009), .ZN(n6010) );
  NAND2_X1 U7042 ( .A1(n6011), .A2(n6010), .ZN(n9089) );
  INV_X1 U7043 ( .A(n9089), .ZN(n8827) );
  NAND2_X1 U7044 ( .A1(n9194), .A2(n8827), .ZN(n6273) );
  NAND2_X1 U7045 ( .A1(n6272), .A2(n6273), .ZN(n9072) );
  INV_X1 U7046 ( .A(n6272), .ZN(n6012) );
  INV_X1 U7047 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8141) );
  INV_X1 U7048 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9367) );
  MUX2_X1 U7049 ( .A(n8141), .B(n9367), .S(n5034), .Z(n6016) );
  INV_X1 U7050 ( .A(SI_23_), .ZN(n9468) );
  NAND2_X1 U7051 ( .A1(n6016), .A2(n9468), .ZN(n6029) );
  INV_X1 U7052 ( .A(n6016), .ZN(n6017) );
  NAND2_X1 U7053 ( .A1(n6017), .A2(SI_23_), .ZN(n6018) );
  NAND2_X1 U7054 ( .A1(n8138), .A2(n6161), .ZN(n6020) );
  OR2_X1 U7055 ( .A1(n5695), .A2(n8141), .ZN(n6019) );
  XNOR2_X1 U7056 ( .A(n6036), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U7057 ( .A1(n9055), .A2(n6131), .ZN(n6026) );
  INV_X1 U7058 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7059 ( .A1(n5637), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7060 ( .A1(n5814), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6021) );
  OAI211_X1 U7061 ( .C1(n6023), .C2(n5819), .A(n6022), .B(n6021), .ZN(n6024)
         );
  INV_X1 U7062 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U7063 ( .A1(n6026), .A2(n6025), .ZN(n9075) );
  NAND2_X1 U7064 ( .A1(n9054), .A2(n9034), .ZN(n6281) );
  NAND2_X1 U7065 ( .A1(n6280), .A2(n6281), .ZN(n9049) );
  INV_X1 U7066 ( .A(n9049), .ZN(n9046) );
  MUX2_X1 U7067 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n5034), .Z(n6047) );
  INV_X1 U7068 ( .A(SI_24_), .ZN(n9470) );
  XNOR2_X1 U7069 ( .A(n6047), .B(n9470), .ZN(n6046) );
  XNOR2_X1 U7070 ( .A(n6050), .B(n6046), .ZN(n8204) );
  NAND2_X1 U7071 ( .A1(n8204), .A2(n6161), .ZN(n6032) );
  INV_X1 U7072 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8205) );
  OR2_X1 U7073 ( .A1(n5695), .A2(n8205), .ZN(n6031) );
  AND2_X1 U7074 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n6033) );
  INV_X1 U7075 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6035) );
  INV_X1 U7076 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8850) );
  OAI21_X1 U7077 ( .B1(n6036), .B2(n6035), .A(n8850), .ZN(n6037) );
  NAND2_X1 U7078 ( .A1(n6057), .A2(n6037), .ZN(n9030) );
  OR2_X1 U7079 ( .A1(n9030), .A2(n6090), .ZN(n6043) );
  INV_X1 U7080 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7081 ( .A1(n5637), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7082 ( .A1(n5814), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6038) );
  OAI211_X1 U7083 ( .C1(n5819), .C2(n6040), .A(n6039), .B(n6038), .ZN(n6041)
         );
  INV_X1 U7084 ( .A(n6041), .ZN(n6042) );
  NAND2_X1 U7085 ( .A1(n6043), .A2(n6042), .ZN(n8886) );
  INV_X1 U7086 ( .A(n8886), .ZN(n6044) );
  NAND2_X1 U7087 ( .A1(n9182), .A2(n6044), .ZN(n6282) );
  INV_X1 U7088 ( .A(n6288), .ZN(n6045) );
  INV_X1 U7089 ( .A(n6046), .ZN(n6049) );
  NAND2_X1 U7090 ( .A1(n6047), .A2(SI_24_), .ZN(n6048) );
  INV_X1 U7091 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8310) );
  INV_X1 U7092 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9361) );
  MUX2_X1 U7093 ( .A(n8310), .B(n9361), .S(n5034), .Z(n6051) );
  INV_X1 U7094 ( .A(SI_25_), .ZN(n9469) );
  NAND2_X1 U7095 ( .A1(n6051), .A2(n9469), .ZN(n6067) );
  INV_X1 U7096 ( .A(n6051), .ZN(n6052) );
  NAND2_X1 U7097 ( .A1(n6052), .A2(SI_25_), .ZN(n6053) );
  NAND2_X1 U7098 ( .A1(n6067), .A2(n6053), .ZN(n6066) );
  NAND2_X1 U7099 ( .A1(n8308), .A2(n6161), .ZN(n6055) );
  OR2_X1 U7100 ( .A1(n5695), .A2(n8310), .ZN(n6054) );
  INV_X1 U7101 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U7102 ( .A1(n6057), .A2(n9322), .ZN(n6058) );
  NAND2_X1 U7103 ( .A1(n6073), .A2(n6058), .ZN(n9014) );
  OR2_X1 U7104 ( .A1(n9014), .A2(n6090), .ZN(n6064) );
  INV_X1 U7105 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7106 ( .A1(n5637), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7107 ( .A1(n5814), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6059) );
  OAI211_X1 U7108 ( .C1(n6061), .C2(n5819), .A(n6060), .B(n6059), .ZN(n6062)
         );
  INV_X1 U7109 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7110 ( .A1(n6064), .A2(n6063), .ZN(n9040) );
  INV_X1 U7111 ( .A(n9040), .ZN(n8851) );
  NAND2_X1 U7112 ( .A1(n9178), .A2(n8851), .ZN(n6177) );
  INV_X1 U7113 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8446) );
  INV_X1 U7114 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9580) );
  MUX2_X1 U7115 ( .A(n8446), .B(n9580), .S(n5034), .Z(n6068) );
  INV_X1 U7116 ( .A(SI_26_), .ZN(n9259) );
  NAND2_X1 U7117 ( .A1(n6068), .A2(n9259), .ZN(n6083) );
  INV_X1 U7118 ( .A(n6068), .ZN(n6069) );
  NAND2_X1 U7119 ( .A1(n6069), .A2(SI_26_), .ZN(n6070) );
  AND2_X1 U7120 ( .A1(n6083), .A2(n6070), .ZN(n6081) );
  NAND2_X1 U7121 ( .A1(n8445), .A2(n6161), .ZN(n6072) );
  OR2_X1 U7122 ( .A1(n5695), .A2(n8446), .ZN(n6071) );
  INV_X1 U7123 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U7124 ( .A1(n6073), .A2(n9565), .ZN(n6074) );
  NAND2_X1 U7125 ( .A1(n9003), .A2(n6131), .ZN(n6080) );
  INV_X1 U7126 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7127 ( .A1(n5637), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7128 ( .A1(n5814), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6075) );
  OAI211_X1 U7129 ( .C1(n5819), .C2(n6077), .A(n6076), .B(n6075), .ZN(n6078)
         );
  INV_X1 U7130 ( .A(n6078), .ZN(n6079) );
  NAND2_X1 U7131 ( .A1(n6080), .A2(n6079), .ZN(n8991) );
  MUX2_X1 U7132 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n5034), .Z(n6098) );
  INV_X1 U7133 ( .A(SI_27_), .ZN(n9463) );
  XNOR2_X1 U7134 ( .A(n6098), .B(n9463), .ZN(n6097) );
  NAND2_X1 U7135 ( .A1(n8506), .A2(n6161), .ZN(n6086) );
  INV_X1 U7136 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8776) );
  OR2_X1 U7137 ( .A1(n5695), .A2(n8776), .ZN(n6085) );
  INV_X1 U7138 ( .A(n6088), .ZN(n6087) );
  NAND2_X1 U7139 ( .A1(n6087), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6104) );
  INV_X1 U7140 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U7141 ( .A1(n6088), .A2(n9303), .ZN(n6089) );
  NAND2_X1 U7142 ( .A1(n6104), .A2(n6089), .ZN(n8984) );
  INV_X1 U7143 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7144 ( .A1(n5637), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7145 ( .A1(n5814), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6091) );
  OAI211_X1 U7146 ( .C1(n6093), .C2(n5819), .A(n6092), .B(n6091), .ZN(n6094)
         );
  INV_X1 U7147 ( .A(n6094), .ZN(n6095) );
  NAND2_X1 U7148 ( .A1(n9167), .A2(n8879), .ZN(n6296) );
  INV_X1 U7149 ( .A(n6097), .ZN(n6100) );
  NAND2_X1 U7150 ( .A1(n6098), .A2(SI_27_), .ZN(n6099) );
  MUX2_X1 U7151 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5034), .Z(n6115) );
  XNOR2_X1 U7152 ( .A(n6115), .B(SI_28_), .ZN(n6113) );
  NAND2_X1 U7153 ( .A1(n8545), .A2(n6161), .ZN(n6103) );
  INV_X1 U7154 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8546) );
  OR2_X1 U7155 ( .A1(n5695), .A2(n8546), .ZN(n6102) );
  INV_X1 U7156 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U7157 ( .A1(n6104), .A2(n7133), .ZN(n6105) );
  NAND2_X1 U7158 ( .A1(n8972), .A2(n6131), .ZN(n6111) );
  INV_X1 U7159 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7160 ( .A1(n5637), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7161 ( .A1(n5814), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6106) );
  OAI211_X1 U7162 ( .C1(n6108), .C2(n5819), .A(n6107), .B(n6106), .ZN(n6109)
         );
  INV_X1 U7163 ( .A(n6109), .ZN(n6110) );
  NAND2_X1 U7164 ( .A1(n6111), .A2(n6110), .ZN(n8992) );
  INV_X1 U7165 ( .A(n6176), .ZN(n6112) );
  NAND2_X1 U7166 ( .A1(n9162), .A2(n8817), .ZN(n6175) );
  INV_X1 U7167 ( .A(n6115), .ZN(n6116) );
  INV_X1 U7168 ( .A(SI_28_), .ZN(n9258) );
  NAND2_X1 U7169 ( .A1(n6116), .A2(n9258), .ZN(n6117) );
  MUX2_X1 U7170 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5034), .Z(n6118) );
  INV_X1 U7171 ( .A(n6121), .ZN(n6122) );
  INV_X1 U7172 ( .A(SI_29_), .ZN(n9471) );
  NAND2_X1 U7173 ( .A1(n6122), .A2(n9471), .ZN(n6123) );
  NAND2_X1 U7174 ( .A1(n8791), .A2(n6161), .ZN(n6125) );
  INV_X1 U7175 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8591) );
  OR2_X1 U7176 ( .A1(n5695), .A2(n8591), .ZN(n6124) );
  INV_X1 U7177 ( .A(n6126), .ZN(n8668) );
  INV_X1 U7178 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7179 ( .A1(n5637), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7180 ( .A1(n5814), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6127) );
  OAI211_X1 U7181 ( .C1(n6129), .C2(n5819), .A(n6128), .B(n6127), .ZN(n6130)
         );
  AOI21_X1 U7182 ( .B1(n8668), .B2(n6131), .A(n6130), .ZN(n8885) );
  NAND2_X1 U7183 ( .A1(n8594), .A2(n8885), .ZN(n6302) );
  OAI21_X1 U7184 ( .B1(n8663), .B2(n8661), .A(n6301), .ZN(n6153) );
  MUX2_X1 U7185 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7182), .Z(n6134) );
  NAND2_X1 U7186 ( .A1(n6134), .A2(SI_30_), .ZN(n6156) );
  OAI21_X1 U7187 ( .B1(SI_30_), .B2(n6134), .A(n6156), .ZN(n6135) );
  NAND2_X1 U7188 ( .A1(n5072), .A2(n6135), .ZN(n6136) );
  INV_X1 U7189 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9697) );
  OR2_X1 U7190 ( .A1(n5695), .A2(n9697), .ZN(n6138) );
  NAND2_X1 U7191 ( .A1(n5637), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6144) );
  INV_X1 U7192 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7193 ( .A1(n5819), .A2(n6140), .ZN(n6143) );
  INV_X1 U7194 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6141) );
  OR2_X1 U7195 ( .A1(n5638), .A2(n6141), .ZN(n6142) );
  AND3_X1 U7196 ( .A1(n6144), .A2(n6143), .A3(n6142), .ZN(n8665) );
  NOR2_X1 U7197 ( .A1(n8965), .A2(n8665), .ZN(n6171) );
  INV_X1 U7198 ( .A(n6145), .ZN(n6146) );
  NAND2_X1 U7199 ( .A1(n6146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6148) );
  XNOR2_X1 U7200 ( .A(n6148), .B(n6147), .ZN(n7825) );
  INV_X1 U7201 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7202 ( .A1(n5637), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6151) );
  INV_X1 U7203 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6149) );
  OR2_X1 U7204 ( .A1(n5638), .A2(n6149), .ZN(n6150) );
  OAI211_X1 U7205 ( .C1(n5819), .C2(n6152), .A(n6151), .B(n6150), .ZN(n8884)
         );
  OAI22_X1 U7206 ( .A1(n6153), .A2(n6171), .B1(n7825), .B2(n8884), .ZN(n6155)
         );
  NAND2_X1 U7207 ( .A1(n6155), .A2(n6154), .ZN(n6164) );
  MUX2_X1 U7208 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7182), .Z(n6158) );
  XNOR2_X1 U7209 ( .A(n6158), .B(SI_31_), .ZN(n6159) );
  NAND2_X1 U7210 ( .A1(n9808), .A2(n6161), .ZN(n6163) );
  INV_X1 U7211 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9692) );
  OR2_X1 U7212 ( .A1(n5695), .A2(n9692), .ZN(n6162) );
  INV_X1 U7213 ( .A(n8884), .ZN(n8598) );
  NAND2_X1 U7214 ( .A1(n8965), .A2(n8665), .ZN(n6303) );
  AND2_X1 U7215 ( .A1(n9148), .A2(n8598), .ZN(n6170) );
  INV_X1 U7216 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6165) );
  INV_X1 U7217 ( .A(n7825), .ZN(n6365) );
  NAND2_X1 U7218 ( .A1(n7588), .A2(n6365), .ZN(n7433) );
  NAND2_X1 U7219 ( .A1(n7811), .A2(n9004), .ZN(n7427) );
  NAND2_X1 U7220 ( .A1(n6167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6344) );
  INV_X1 U7221 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6343) );
  XNOR2_X1 U7222 ( .A(n6344), .B(n6343), .ZN(n8039) );
  NAND2_X1 U7223 ( .A1(n8039), .A2(n7825), .ZN(n7702) );
  OR2_X2 U7224 ( .A1(n7427), .A2(n7702), .ZN(n7036) );
  OAI21_X1 U7225 ( .B1(n10812), .B2(n7433), .A(n7036), .ZN(n6168) );
  AND2_X1 U7226 ( .A1(n6365), .A2(n10812), .ZN(n7701) );
  NAND2_X1 U7227 ( .A1(n6333), .A2(n6274), .ZN(n6174) );
  INV_X1 U7228 ( .A(n6170), .ZN(n6172) );
  INV_X1 U7229 ( .A(n6171), .ZN(n6304) );
  NAND2_X1 U7230 ( .A1(n6172), .A2(n6304), .ZN(n6334) );
  NAND2_X1 U7231 ( .A1(n6334), .A2(n6308), .ZN(n6173) );
  NAND2_X1 U7232 ( .A1(n6174), .A2(n6173), .ZN(n6312) );
  MUX2_X1 U7233 ( .A(n6176), .B(n6175), .S(n6308), .Z(n6300) );
  NAND2_X1 U7234 ( .A1(n6313), .A2(n6177), .ZN(n6180) );
  NAND2_X1 U7235 ( .A1(n6314), .A2(n6178), .ZN(n6179) );
  MUX2_X1 U7236 ( .A(n6180), .B(n6179), .S(n6308), .Z(n6294) );
  AND2_X1 U7237 ( .A1(n8903), .A2(n7513), .ZN(n6315) );
  INV_X1 U7238 ( .A(n6315), .ZN(n6182) );
  NAND2_X1 U7239 ( .A1(n6316), .A2(n6182), .ZN(n6181) );
  NAND2_X1 U7240 ( .A1(n6181), .A2(n6317), .ZN(n6185) );
  AND3_X1 U7241 ( .A1(n6316), .A2(n6182), .A3(n6365), .ZN(n6183) );
  NOR2_X1 U7242 ( .A1(n7748), .A2(n6183), .ZN(n6184) );
  MUX2_X1 U7243 ( .A(n6185), .B(n6184), .S(n6308), .Z(n6186) );
  MUX2_X1 U7244 ( .A(n7614), .B(n6187), .S(n6308), .Z(n6188) );
  NAND3_X1 U7245 ( .A1(n6189), .A2(n6318), .A3(n6188), .ZN(n6192) );
  MUX2_X1 U7246 ( .A(n7716), .B(n6190), .S(n6274), .Z(n6191) );
  AOI21_X1 U7247 ( .B1(n6192), .B2(n6191), .A(n7724), .ZN(n6196) );
  NOR2_X1 U7248 ( .A1(n8899), .A2(n6274), .ZN(n6194) );
  AND2_X1 U7249 ( .A1(n8899), .A2(n6274), .ZN(n6193) );
  MUX2_X1 U7250 ( .A(n6194), .B(n6193), .S(n10752), .Z(n6195) );
  OAI21_X1 U7251 ( .B1(n6196), .B2(n6195), .A(n10797), .ZN(n6203) );
  OR2_X1 U7252 ( .A1(n8898), .A2(n10806), .ZN(n7799) );
  MUX2_X1 U7253 ( .A(n10806), .B(n8898), .S(n6308), .Z(n6197) );
  INV_X1 U7254 ( .A(n6197), .ZN(n6198) );
  MUX2_X1 U7255 ( .A(n8897), .B(n7796), .S(n6308), .Z(n6199) );
  NAND2_X1 U7256 ( .A1(n8897), .A2(n7796), .ZN(n7884) );
  AOI22_X1 U7257 ( .A1(n7799), .A2(n6198), .B1(n6199), .B2(n7884), .ZN(n6202)
         );
  OR2_X1 U7258 ( .A1(n8897), .A2(n7796), .ZN(n6320) );
  INV_X1 U7259 ( .A(n6320), .ZN(n6200) );
  OAI21_X1 U7260 ( .B1(n6200), .B2(n6199), .A(n5722), .ZN(n6201) );
  AOI21_X1 U7261 ( .B1(n6203), .B2(n6202), .A(n6201), .ZN(n6209) );
  MUX2_X1 U7262 ( .A(n6204), .B(n7941), .S(n6274), .Z(n6205) );
  INV_X1 U7263 ( .A(n6205), .ZN(n6208) );
  INV_X1 U7264 ( .A(n6206), .ZN(n6207) );
  MUX2_X1 U7265 ( .A(n8895), .B(n10868), .S(n6308), .Z(n6210) );
  OAI22_X1 U7266 ( .A1(n6209), .A2(n6208), .B1(n6207), .B2(n6210), .ZN(n6212)
         );
  NAND2_X1 U7267 ( .A1(n6210), .A2(n8187), .ZN(n6211) );
  NAND2_X1 U7268 ( .A1(n6212), .A2(n6211), .ZN(n6215) );
  AND2_X1 U7269 ( .A1(n6216), .A2(n6217), .ZN(n6213) );
  MUX2_X1 U7270 ( .A(n8242), .B(n6213), .S(n6308), .Z(n6214) );
  NAND2_X1 U7271 ( .A1(n6214), .A2(n6219), .ZN(n6218) );
  AOI21_X1 U7272 ( .B1(n6215), .B2(n8242), .A(n6218), .ZN(n6224) );
  OAI211_X1 U7273 ( .C1(n6218), .C2(n6217), .A(n6216), .B(n8611), .ZN(n6221)
         );
  NAND2_X1 U7274 ( .A1(n8610), .A2(n6219), .ZN(n6220) );
  MUX2_X1 U7275 ( .A(n6221), .B(n6220), .S(n6308), .Z(n6223) );
  INV_X1 U7276 ( .A(n8614), .ZN(n6323) );
  OR3_X1 U7277 ( .A1(n6224), .A2(n6223), .A3(n6323), .ZN(n6232) );
  INV_X1 U7278 ( .A(n6225), .ZN(n6226) );
  NOR2_X1 U7279 ( .A1(n6227), .A2(n6226), .ZN(n6229) );
  INV_X1 U7280 ( .A(n8314), .ZN(n6228) );
  MUX2_X1 U7281 ( .A(n6229), .B(n6228), .S(n6274), .Z(n6230) );
  NOR2_X1 U7282 ( .A1(n6230), .A2(n8321), .ZN(n6231) );
  NAND2_X1 U7283 ( .A1(n6232), .A2(n6231), .ZN(n6235) );
  MUX2_X1 U7284 ( .A(n6233), .B(n8386), .S(n6274), .Z(n6234) );
  NAND3_X1 U7285 ( .A1(n6235), .A2(n8382), .A3(n6234), .ZN(n6239) );
  MUX2_X1 U7286 ( .A(n6237), .B(n6236), .S(n6308), .Z(n6238) );
  INV_X1 U7287 ( .A(n8514), .ZN(n8510) );
  AOI21_X1 U7288 ( .B1(n6239), .B2(n6238), .A(n8510), .ZN(n6246) );
  MUX2_X1 U7289 ( .A(n8509), .B(n6240), .S(n6308), .Z(n6241) );
  NAND2_X1 U7290 ( .A1(n6241), .A2(n8517), .ZN(n6245) );
  MUX2_X1 U7291 ( .A(n6243), .B(n6242), .S(n6274), .Z(n6244) );
  OAI21_X1 U7292 ( .B1(n6246), .B2(n6245), .A(n6244), .ZN(n6252) );
  INV_X1 U7293 ( .A(n9223), .ZN(n8595) );
  MUX2_X1 U7294 ( .A(n6247), .B(n8595), .S(n6308), .Z(n6250) );
  INV_X1 U7295 ( .A(n6250), .ZN(n6249) );
  NAND2_X1 U7296 ( .A1(n6249), .A2(n6248), .ZN(n6251) );
  AOI22_X1 U7297 ( .A1(n6252), .A2(n6251), .B1(n6250), .B2(n8649), .ZN(n6256)
         );
  MUX2_X1 U7298 ( .A(n6254), .B(n6253), .S(n6274), .Z(n6255) );
  OAI21_X1 U7299 ( .B1(n6256), .B2(n9135), .A(n6255), .ZN(n6257) );
  INV_X1 U7300 ( .A(n9112), .ZN(n9107) );
  NAND2_X1 U7301 ( .A1(n6257), .A2(n9107), .ZN(n6261) );
  MUX2_X1 U7302 ( .A(n6259), .B(n6258), .S(n6308), .Z(n6260) );
  NAND3_X1 U7303 ( .A1(n6261), .A2(n6329), .A3(n6260), .ZN(n6265) );
  MUX2_X1 U7304 ( .A(n6263), .B(n6262), .S(n6308), .Z(n6264) );
  NAND2_X1 U7305 ( .A1(n6265), .A2(n6264), .ZN(n6270) );
  NAND2_X1 U7306 ( .A1(n9199), .A2(n9102), .ZN(n6327) );
  INV_X1 U7307 ( .A(n6327), .ZN(n6266) );
  NAND2_X1 U7308 ( .A1(n6270), .A2(n6266), .ZN(n6268) );
  MUX2_X1 U7309 ( .A(n9102), .B(n9199), .S(n6274), .Z(n6267) );
  NAND2_X1 U7310 ( .A1(n6268), .A2(n6267), .ZN(n6269) );
  OAI21_X1 U7311 ( .B1(n6270), .B2(n8655), .A(n6269), .ZN(n6271) );
  INV_X1 U7312 ( .A(n9072), .ZN(n9061) );
  NAND2_X1 U7313 ( .A1(n6271), .A2(n9061), .ZN(n6279) );
  NAND2_X1 U7314 ( .A1(n6280), .A2(n6272), .ZN(n6276) );
  INV_X1 U7315 ( .A(n6273), .ZN(n6275) );
  MUX2_X1 U7316 ( .A(n6276), .B(n6275), .S(n6274), .Z(n6277) );
  INV_X1 U7317 ( .A(n6277), .ZN(n6278) );
  NAND3_X1 U7318 ( .A1(n6279), .A2(n6281), .A3(n6278), .ZN(n6287) );
  NAND2_X1 U7319 ( .A1(n6288), .A2(n6280), .ZN(n6284) );
  NAND2_X1 U7320 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  MUX2_X1 U7321 ( .A(n6284), .B(n6283), .S(n6308), .Z(n6285) );
  INV_X1 U7322 ( .A(n6285), .ZN(n6286) );
  NAND2_X1 U7323 ( .A1(n6287), .A2(n6286), .ZN(n6291) );
  OAI21_X1 U7324 ( .B1(n6308), .B2(n8886), .A(n6288), .ZN(n6289) );
  OAI21_X1 U7325 ( .B1(n6308), .B2(n9182), .A(n6289), .ZN(n6290) );
  AOI21_X1 U7326 ( .B1(n6291), .B2(n6290), .A(n9019), .ZN(n6293) );
  MUX2_X1 U7327 ( .A(n6314), .B(n6313), .S(n6308), .Z(n6292) );
  OAI211_X1 U7328 ( .C1(n6294), .C2(n6293), .A(n8989), .B(n6292), .ZN(n6298)
         );
  MUX2_X1 U7329 ( .A(n6296), .B(n6295), .S(n6308), .Z(n6297) );
  NAND3_X1 U7330 ( .A1(n8969), .A2(n6298), .A3(n6297), .ZN(n6299) );
  NAND3_X1 U7331 ( .A1(n8660), .A2(n6300), .A3(n6299), .ZN(n6307) );
  MUX2_X1 U7332 ( .A(n6302), .B(n6301), .S(n6308), .Z(n6306) );
  NAND2_X1 U7333 ( .A1(n6304), .A2(n6303), .ZN(n6305) );
  AOI21_X1 U7334 ( .B1(n6307), .B2(n6306), .A(n6305), .ZN(n6311) );
  MUX2_X1 U7335 ( .A(n8884), .B(n9148), .S(n6308), .Z(n6310) );
  NOR2_X1 U7336 ( .A1(n9148), .A2(n8884), .ZN(n6309) );
  OR2_X1 U7337 ( .A1(n6315), .A2(n7584), .ZN(n7781) );
  NAND2_X1 U7338 ( .A1(n6317), .A2(n6316), .ZN(n7586) );
  NOR3_X1 U7339 ( .A1(n7781), .A2(n7811), .A3(n7586), .ZN(n6319) );
  INV_X1 U7340 ( .A(n7804), .ZN(n7797) );
  NOR4_X1 U7341 ( .A1(n6321), .A2(n7724), .A3(n7797), .A4(n7889), .ZN(n6322)
         );
  INV_X1 U7342 ( .A(n8190), .ZN(n8192) );
  NAND4_X1 U7343 ( .A1(n6322), .A2(n8192), .A3(n8264), .A4(n7956), .ZN(n6324)
         );
  NAND2_X1 U7344 ( .A1(n8610), .A2(n8611), .ZN(n8276) );
  NOR4_X1 U7345 ( .A1(n8321), .A2(n6324), .A3(n6323), .A4(n8276), .ZN(n6325)
         );
  NAND4_X1 U7346 ( .A1(n8517), .A2(n8514), .A3(n8382), .A4(n6325), .ZN(n6326)
         );
  NOR4_X1 U7347 ( .A1(n9112), .A2(n9135), .A3(n8536), .A4(n6326), .ZN(n6328)
         );
  NAND2_X1 U7348 ( .A1(n8655), .A2(n6327), .ZN(n9087) );
  NAND4_X1 U7349 ( .A1(n9061), .A2(n6329), .A3(n6328), .A4(n9087), .ZN(n6330)
         );
  NOR4_X1 U7350 ( .A1(n9019), .A2(n9037), .A3(n9049), .A4(n6330), .ZN(n6331)
         );
  NAND4_X1 U7351 ( .A1(n8969), .A2(n8989), .A3(n5493), .A4(n6331), .ZN(n6332)
         );
  NOR4_X1 U7352 ( .A1(n6334), .A2(n6333), .A3(n8661), .A4(n6332), .ZN(n6335)
         );
  XNOR2_X1 U7353 ( .A(n6335), .B(n10812), .ZN(n6336) );
  AOI211_X1 U7354 ( .C1(n7811), .C2(n6338), .A(n6365), .B(n6336), .ZN(n6337)
         );
  INV_X1 U7355 ( .A(n6337), .ZN(n6340) );
  OR2_X1 U7356 ( .A1(n8039), .A2(n9004), .ZN(n7432) );
  XOR2_X1 U7357 ( .A(n7432), .B(n6338), .Z(n6339) );
  INV_X1 U7358 ( .A(n7702), .ZN(n7428) );
  NAND3_X1 U7359 ( .A1(n6341), .A2(n6340), .A3(n5049), .ZN(n6347) );
  NAND2_X1 U7360 ( .A1(n6344), .A2(n6343), .ZN(n6345) );
  NAND2_X1 U7361 ( .A1(n6345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6349) );
  INV_X1 U7362 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6348) );
  XNOR2_X1 U7363 ( .A(n6349), .B(n6348), .ZN(n7179) );
  OR2_X1 U7364 ( .A1(n7179), .A2(P2_U3152), .ZN(n8139) );
  INV_X1 U7365 ( .A(n8139), .ZN(n7220) );
  OAI21_X1 U7366 ( .B1(n6347), .B2(n6346), .A(n7220), .ZN(n6369) );
  NAND2_X1 U7367 ( .A1(n6349), .A2(n6348), .ZN(n6350) );
  NAND2_X1 U7368 ( .A1(n6350), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6352) );
  INV_X1 U7369 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6351) );
  XNOR2_X1 U7370 ( .A(n6352), .B(n6351), .ZN(n8206) );
  INV_X1 U7371 ( .A(n8206), .ZN(n6360) );
  NAND2_X1 U7372 ( .A1(n6353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6354) );
  XNOR2_X1 U7373 ( .A(n6354), .B(n5572), .ZN(n8309) );
  INV_X1 U7374 ( .A(n8309), .ZN(n6359) );
  NAND2_X1 U7375 ( .A1(n6356), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6358) );
  AND2_X1 U7376 ( .A1(n6358), .A2(n6357), .ZN(n7115) );
  NAND3_X1 U7377 ( .A1(n6360), .A2(n6359), .A3(n7115), .ZN(n7282) );
  NAND2_X1 U7378 ( .A1(n7282), .A2(n7179), .ZN(n7136) );
  INV_X1 U7379 ( .A(n7136), .ZN(n6361) );
  INV_X1 U7380 ( .A(n7427), .ZN(n6362) );
  NAND2_X1 U7381 ( .A1(n7700), .A2(n6362), .ZN(n7131) );
  INV_X1 U7382 ( .A(n6364), .ZN(n7297) );
  INV_X1 U7383 ( .A(n8039), .ZN(n6975) );
  AND2_X1 U7384 ( .A1(n6975), .A2(n6365), .ZN(n7429) );
  AND2_X2 U7385 ( .A1(n7297), .A2(n7429), .ZN(n9137) );
  INV_X1 U7386 ( .A(n9137), .ZN(n9067) );
  NOR3_X1 U7387 ( .A1(n7131), .A2(n6363), .A3(n9067), .ZN(n6367) );
  OAI21_X1 U7388 ( .B1(n8139), .B2(n6975), .A(P2_B_REG_SCAN_IN), .ZN(n6366) );
  NAND2_X1 U7389 ( .A1(n6369), .A2(n6368), .ZN(P2_U3244) );
  NAND2_X1 U7390 ( .A1(n6371), .A2(n9625), .ZN(n6372) );
  INV_X1 U7391 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6374) );
  INV_X1 U7392 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6373) );
  NAND4_X1 U7393 ( .A1(n6374), .A2(n6373), .A3(n9640), .A4(n9653), .ZN(n6375)
         );
  INV_X1 U7394 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6379) );
  NOR2_X1 U7395 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6378) );
  AND2_X1 U7396 ( .A1(n6379), .A2(n6391), .ZN(n6380) );
  INV_X1 U7397 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6577) );
  INV_X1 U7398 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U7399 ( .A1(n8308), .A2(n9807), .ZN(n6384) );
  NAND2_X4 U7400 ( .A1(n6503), .A2(n7182), .ZN(n9822) );
  OR2_X1 U7401 ( .A1(n9822), .A2(n9361), .ZN(n6383) );
  NAND2_X1 U7402 ( .A1(n6397), .A2(n6385), .ZN(n6386) );
  NAND2_X1 U7403 ( .A1(n6386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6945) );
  INV_X1 U7404 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U7405 ( .A1(n6945), .A2(n9431), .ZN(n6944) );
  NAND2_X1 U7406 ( .A1(n6391), .A2(n6388), .ZN(n6394) );
  NAND2_X1 U7407 ( .A1(n6394), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6389) );
  MUX2_X1 U7408 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6389), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6390) );
  NAND2_X1 U7409 ( .A1(n6391), .A2(n6397), .ZN(n6392) );
  NAND2_X1 U7410 ( .A1(n6392), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6393) );
  MUX2_X1 U7411 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6393), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6395) );
  INV_X1 U7412 ( .A(n8312), .ZN(n6396) );
  INV_X1 U7413 ( .A(n6418), .ZN(n7154) );
  INV_X1 U7414 ( .A(n6397), .ZN(n6398) );
  NAND2_X1 U7415 ( .A1(n6400), .A2(n9657), .ZN(n6399) );
  XNOR2_X1 U7416 ( .A(n6400), .B(P1_IR_REG_20__SCAN_IN), .ZN(n10076) );
  INV_X1 U7417 ( .A(n10076), .ZN(n7822) );
  INV_X1 U7418 ( .A(n7858), .ZN(n6419) );
  NAND2_X1 U7419 ( .A1(n10500), .A2(n6922), .ZN(n6421) );
  NAND2_X1 U7420 ( .A1(n6402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6403) );
  INV_X1 U7421 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U7422 ( .A1(n5033), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6417) );
  INV_X1 U7423 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6404) );
  OR2_X1 U7424 ( .A1(n6831), .A2(n6404), .ZN(n6416) );
  NAND2_X4 U7425 ( .A1(n6413), .A2(n6406), .ZN(n6910) );
  NAND2_X1 U7426 ( .A1(n6531), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U7427 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n6407) );
  INV_X1 U7428 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8234) );
  AND2_X1 U7429 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n6408) );
  INV_X1 U7430 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6700) );
  INV_X1 U7431 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10184) );
  INV_X1 U7432 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U7433 ( .A1(n6757), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6778) );
  INV_X1 U7434 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6777) );
  INV_X1 U7435 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U7436 ( .A1(n6825), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U7437 ( .A1(n6845), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6844) );
  INV_X1 U7438 ( .A(n6844), .ZN(n6409) );
  INV_X1 U7439 ( .A(n6878), .ZN(n6412) );
  INV_X1 U7440 ( .A(n6862), .ZN(n6410) );
  INV_X1 U7441 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U7442 ( .A1(n6410), .A2(n9732), .ZN(n6411) );
  NAND2_X1 U7443 ( .A1(n6412), .A2(n6411), .ZN(n10336) );
  OR2_X1 U7444 ( .A1(n6910), .A2(n10336), .ZN(n6415) );
  INV_X1 U7445 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10337) );
  OR2_X1 U7446 ( .A1(n9815), .A2(n10337), .ZN(n6414) );
  INV_X1 U7447 ( .A(n10321), .ZN(n10358) );
  NAND2_X1 U7448 ( .A1(n6418), .A2(n6419), .ZN(n6484) );
  NAND2_X1 U7449 ( .A1(n10358), .A2(n6434), .ZN(n6420) );
  NAND2_X1 U7450 ( .A1(n6421), .A2(n6420), .ZN(n6429) );
  NAND2_X1 U7451 ( .A1(n6422), .A2(n9426), .ZN(n6423) );
  NAND2_X1 U7452 ( .A1(n6423), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U7453 ( .A1(n6426), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6427) );
  XNOR2_X1 U7454 ( .A(n6427), .B(n5547), .ZN(n10260) );
  XNOR2_X1 U7455 ( .A(n6429), .B(n6918), .ZN(n9729) );
  INV_X1 U7456 ( .A(n9729), .ZN(n6874) );
  AND2_X1 U7457 ( .A1(n7822), .A2(n10260), .ZN(n10083) );
  NAND2_X1 U7458 ( .A1(n8124), .A2(n10083), .ZN(n6430) );
  NOR2_X1 U7459 ( .A1(n10321), .A2(n6901), .ZN(n6431) );
  INV_X1 U7460 ( .A(n9728), .ZN(n6873) );
  NAND2_X1 U7461 ( .A1(n8138), .A2(n9807), .ZN(n6433) );
  OR2_X1 U7462 ( .A1(n9822), .A2(n9367), .ZN(n6432) );
  NAND2_X1 U7463 ( .A1(n5033), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6442) );
  INV_X1 U7464 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6435) );
  OR2_X1 U7465 ( .A1(n6831), .A2(n6435), .ZN(n6441) );
  INV_X1 U7466 ( .A(n6860), .ZN(n6437) );
  INV_X1 U7467 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U7468 ( .A1(n9704), .A2(n6844), .ZN(n6436) );
  NAND2_X1 U7469 ( .A1(n6437), .A2(n6436), .ZN(n10371) );
  OR2_X1 U7470 ( .A1(n6910), .A2(n10371), .ZN(n6440) );
  INV_X1 U7471 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6438) );
  OR2_X1 U7472 ( .A1(n9815), .A2(n6438), .ZN(n6439) );
  NOR2_X1 U7473 ( .A1(n10387), .A2(n6901), .ZN(n6443) );
  AOI21_X1 U7474 ( .B1(n10508), .B2(n6434), .A(n6443), .ZN(n9702) );
  NAND2_X1 U7475 ( .A1(n6644), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U7476 ( .A1(n5032), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6447) );
  INV_X1 U7477 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6444) );
  INV_X1 U7478 ( .A(n6449), .ZN(n6450) );
  OR2_X1 U7479 ( .A1(n9819), .A2(n7194), .ZN(n6452) );
  INV_X1 U7480 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7180) );
  OR2_X1 U7481 ( .A1(n9822), .A2(n7180), .ZN(n6451) );
  NAND2_X1 U7482 ( .A1(n7980), .A2(n6922), .ZN(n6453) );
  NAND2_X1 U7483 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  XNOR2_X1 U7484 ( .A(n6455), .B(n6850), .ZN(n6476) );
  INV_X1 U7485 ( .A(SI_0_), .ZN(n6457) );
  INV_X1 U7486 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6456) );
  OAI21_X1 U7487 ( .B1(n7182), .B2(n6457), .A(n6456), .ZN(n6459) );
  AND2_X1 U7488 ( .A1(n6459), .A2(n6458), .ZN(n10598) );
  NOR2_X1 U7489 ( .A1(n6418), .A2(n6461), .ZN(n6462) );
  INV_X1 U7490 ( .A(n6463), .ZN(n6468) );
  NAND2_X1 U7491 ( .A1(n5032), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U7492 ( .A1(n6645), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U7493 ( .A1(n6469), .A2(n6434), .ZN(n6472) );
  AOI22_X1 U7494 ( .A1(n8014), .A2(n6470), .B1(n7154), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U7495 ( .A1(n6472), .A2(n6471), .ZN(n7496) );
  NAND2_X1 U7496 ( .A1(n7497), .A2(n7496), .ZN(n7499) );
  INV_X1 U7497 ( .A(n7499), .ZN(n6473) );
  NAND2_X1 U7498 ( .A1(n6476), .A2(n6475), .ZN(n7505) );
  AND2_X1 U7499 ( .A1(n7980), .A2(n6434), .ZN(n6474) );
  AOI21_X1 U7500 ( .B1(n10107), .B2(n6915), .A(n6474), .ZN(n7506) );
  NAND2_X1 U7501 ( .A1(n7505), .A2(n7506), .ZN(n6479) );
  INV_X1 U7502 ( .A(n6475), .ZN(n6478) );
  INV_X1 U7503 ( .A(n6476), .ZN(n6477) );
  NAND2_X1 U7504 ( .A1(n6478), .A2(n6477), .ZN(n7504) );
  NAND2_X1 U7505 ( .A1(n6479), .A2(n7504), .ZN(n7522) );
  INV_X1 U7506 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10134) );
  INV_X1 U7507 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U7508 ( .A1(n5033), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6481) );
  INV_X1 U7509 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10710) );
  OR2_X1 U7510 ( .A1(n6831), .A2(n10710), .ZN(n6480) );
  AND4_X2 U7511 ( .A1(n6483), .A2(n6482), .A3(n6481), .A4(n6480), .ZN(n7831)
         );
  NOR2_X1 U7512 ( .A1(n6449), .A2(n6577), .ZN(n6485) );
  MUX2_X1 U7513 ( .A(n6577), .B(n6485), .S(P1_IR_REG_2__SCAN_IN), .Z(n6486) );
  INV_X1 U7514 ( .A(n6486), .ZN(n6488) );
  AND2_X1 U7515 ( .A1(n6488), .A2(n6487), .ZN(n10130) );
  INV_X1 U7516 ( .A(n10130), .ZN(n7244) );
  INV_X1 U7517 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7181) );
  OR2_X1 U7518 ( .A1(n9819), .A2(n7183), .ZN(n6489) );
  INV_X1 U7519 ( .A(n7994), .ZN(n7850) );
  XNOR2_X1 U7520 ( .A(n6491), .B(n6918), .ZN(n6494) );
  OAI22_X1 U7521 ( .A1(n7831), .A2(n6901), .B1(n7850), .B2(n6920), .ZN(n6493)
         );
  INV_X1 U7522 ( .A(n6493), .ZN(n6492) );
  INV_X1 U7523 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6496) );
  OR2_X1 U7524 ( .A1(n6497), .A2(n6496), .ZN(n6501) );
  INV_X1 U7525 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7246) );
  OR2_X1 U7526 ( .A1(n6910), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U7527 ( .A1(n5033), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6498) );
  INV_X1 U7528 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7185) );
  OR2_X1 U7529 ( .A1(n9822), .A2(n7185), .ZN(n6505) );
  NAND2_X1 U7530 ( .A1(n6487), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6502) );
  XNOR2_X1 U7531 ( .A(n6502), .B(n6370), .ZN(n7258) );
  NAND3_X1 U7532 ( .A1(n7522), .A2(n7521), .A3(n6524), .ZN(n7570) );
  NAND2_X1 U7533 ( .A1(n5033), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U7534 ( .A1(n6645), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6509) );
  AND2_X1 U7535 ( .A1(n6510), .A2(n6509), .ZN(n6514) );
  NAND2_X1 U7536 ( .A1(n6644), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6513) );
  NOR2_X1 U7537 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6511) );
  NOR2_X1 U7538 ( .A1(n6531), .A2(n6511), .ZN(n8628) );
  NAND2_X1 U7539 ( .A1(n6795), .A2(n8628), .ZN(n6512) );
  NAND2_X1 U7540 ( .A1(n7834), .A2(n6434), .ZN(n6518) );
  INV_X1 U7541 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7188) );
  OR2_X1 U7542 ( .A1(n9822), .A2(n7188), .ZN(n6517) );
  NAND2_X1 U7543 ( .A1(n6515), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6537) );
  XNOR2_X1 U7544 ( .A(n6537), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10155) );
  INV_X1 U7545 ( .A(n10155), .ZN(n7190) );
  OR2_X1 U7546 ( .A1(n6503), .A2(n7190), .ZN(n6516) );
  XNOR2_X1 U7547 ( .A(n6527), .B(n6528), .ZN(n8621) );
  INV_X1 U7548 ( .A(n6520), .ZN(n6521) );
  NAND2_X1 U7549 ( .A1(n6522), .A2(n6521), .ZN(n8622) );
  AND2_X1 U7550 ( .A1(n8621), .A2(n8622), .ZN(n6525) );
  NAND2_X1 U7551 ( .A1(n7570), .A2(n6526), .ZN(n6544) );
  INV_X1 U7552 ( .A(n6527), .ZN(n6529) );
  OR2_X1 U7553 ( .A1(n6529), .A2(n6528), .ZN(n6547) );
  NAND2_X1 U7554 ( .A1(n6544), .A2(n6547), .ZN(n6542) );
  INV_X1 U7555 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6530) );
  OR2_X1 U7556 ( .A1(n9815), .A2(n6530), .ZN(n6536) );
  OAI21_X1 U7557 ( .B1(n6531), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6552), .ZN(
        n10778) );
  OR2_X1 U7558 ( .A1(n6910), .A2(n10778), .ZN(n6535) );
  NAND2_X1 U7559 ( .A1(n5033), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6534) );
  INV_X1 U7560 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6532) );
  OR2_X1 U7561 ( .A1(n9813), .A2(n6532), .ZN(n6533) );
  NAND4_X1 U7562 ( .A1(n6536), .A2(n6535), .A3(n6534), .A4(n6533), .ZN(n10104)
         );
  NAND2_X1 U7563 ( .A1(n6537), .A2(n9625), .ZN(n6538) );
  NAND2_X1 U7564 ( .A1(n6538), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6539) );
  XNOR2_X1 U7565 ( .A(n6539), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7275) );
  INV_X1 U7566 ( .A(n7275), .ZN(n7257) );
  INV_X1 U7567 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7191) );
  OR2_X1 U7568 ( .A1(n9822), .A2(n7191), .ZN(n6540) );
  OAI22_X1 U7569 ( .A1(n8625), .A2(n6920), .B1(n10764), .B2(n6854), .ZN(n6541)
         );
  XNOR2_X1 U7570 ( .A(n6541), .B(n6850), .ZN(n6545) );
  NAND2_X1 U7571 ( .A1(n6542), .A2(n6545), .ZN(n7632) );
  OAI22_X1 U7572 ( .A1(n8625), .A2(n6901), .B1(n10764), .B2(n6920), .ZN(n7634)
         );
  INV_X1 U7573 ( .A(n7634), .ZN(n6543) );
  NAND2_X1 U7574 ( .A1(n7632), .A2(n6543), .ZN(n6549) );
  INV_X1 U7575 ( .A(n6545), .ZN(n6546) );
  AND2_X1 U7576 ( .A1(n6547), .A2(n6546), .ZN(n6548) );
  NAND2_X1 U7577 ( .A1(n6549), .A2(n7633), .ZN(n7644) );
  NAND2_X1 U7578 ( .A1(n5033), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6558) );
  INV_X1 U7579 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6550) );
  OR2_X1 U7580 ( .A1(n9813), .A2(n6550), .ZN(n6557) );
  AND2_X1 U7581 ( .A1(n6552), .A2(n6551), .ZN(n6553) );
  OR2_X1 U7582 ( .A1(n6553), .A2(n6570), .ZN(n7843) );
  OR2_X1 U7583 ( .A1(n6910), .A2(n7843), .ZN(n6556) );
  INV_X1 U7584 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6554) );
  OR2_X1 U7585 ( .A1(n9815), .A2(n6554), .ZN(n6555) );
  OR2_X1 U7586 ( .A1(n6559), .A2(n6577), .ZN(n6560) );
  XNOR2_X1 U7587 ( .A(n6560), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10650) );
  INV_X1 U7588 ( .A(n10650), .ZN(n7200) );
  OR2_X1 U7589 ( .A1(n9819), .A2(n7199), .ZN(n6562) );
  INV_X1 U7590 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7198) );
  OR2_X1 U7591 ( .A1(n9822), .A2(n7198), .ZN(n6561) );
  OAI22_X1 U7592 ( .A1(n8067), .A2(n6920), .B1(n7899), .B2(n6854), .ZN(n6563)
         );
  XNOR2_X1 U7593 ( .A(n6563), .B(n6918), .ZN(n6565) );
  OAI22_X1 U7594 ( .A1(n8067), .A2(n6901), .B1(n7899), .B2(n6920), .ZN(n6566)
         );
  INV_X1 U7595 ( .A(n6566), .ZN(n6564) );
  NAND2_X1 U7596 ( .A1(n6565), .A2(n6564), .ZN(n6569) );
  INV_X1 U7597 ( .A(n6565), .ZN(n6567) );
  NAND2_X1 U7598 ( .A1(n6567), .A2(n6566), .ZN(n6568) );
  AND2_X1 U7599 ( .A1(n6569), .A2(n6568), .ZN(n7645) );
  NAND2_X1 U7600 ( .A1(n5033), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6575) );
  INV_X1 U7601 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7271) );
  OR2_X1 U7602 ( .A1(n9813), .A2(n7271), .ZN(n6574) );
  OR2_X1 U7603 ( .A1(n6570), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U7604 ( .A1(n6596), .A2(n6571), .ZN(n8073) );
  OR2_X1 U7605 ( .A1(n6910), .A2(n8073), .ZN(n6573) );
  INV_X1 U7606 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8074) );
  OR2_X1 U7607 ( .A1(n9815), .A2(n8074), .ZN(n6572) );
  OR2_X1 U7608 ( .A1(n6576), .A2(n6577), .ZN(n6578) );
  INV_X1 U7609 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9629) );
  XNOR2_X1 U7610 ( .A(n6578), .B(n9629), .ZN(n7276) );
  OR2_X1 U7611 ( .A1(n9819), .A2(n7202), .ZN(n6580) );
  INV_X1 U7612 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7201) );
  OR2_X1 U7613 ( .A1(n9822), .A2(n7201), .ZN(n6579) );
  OAI22_X1 U7614 ( .A1(n8022), .A2(n6920), .B1(n10846), .B2(n6854), .ZN(n6581)
         );
  XNOR2_X1 U7615 ( .A(n6581), .B(n6918), .ZN(n6584) );
  OAI22_X1 U7616 ( .A1(n8022), .A2(n6901), .B1(n10846), .B2(n6920), .ZN(n6582)
         );
  XNOR2_X1 U7617 ( .A(n6584), .B(n6582), .ZN(n7814) );
  INV_X1 U7618 ( .A(n6582), .ZN(n6583) );
  NAND2_X1 U7619 ( .A1(n6584), .A2(n6583), .ZN(n6619) );
  NAND2_X1 U7620 ( .A1(n5033), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6590) );
  INV_X1 U7621 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6585) );
  OR2_X1 U7622 ( .A1(n6831), .A2(n6585), .ZN(n6589) );
  INV_X1 U7623 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6595) );
  XNOR2_X1 U7624 ( .A(n6596), .B(n6595), .ZN(n8021) );
  OR2_X1 U7625 ( .A1(n6910), .A2(n8021), .ZN(n6588) );
  INV_X1 U7626 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6586) );
  OR2_X1 U7627 ( .A1(n9815), .A2(n6586), .ZN(n6587) );
  NAND2_X1 U7628 ( .A1(n6576), .A2(n9629), .ZN(n6631) );
  NAND2_X1 U7629 ( .A1(n6631), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6603) );
  XNOR2_X1 U7630 ( .A(n6603), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7681) );
  INV_X1 U7631 ( .A(n7681), .ZN(n7207) );
  OR2_X1 U7632 ( .A1(n7206), .A2(n9819), .ZN(n6592) );
  INV_X1 U7633 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7205) );
  OR2_X1 U7634 ( .A1(n9822), .A2(n7205), .ZN(n6591) );
  INV_X1 U7635 ( .A(n8009), .ZN(n10861) );
  OAI22_X1 U7636 ( .A1(n8066), .A2(n6901), .B1(n10861), .B2(n6920), .ZN(n6616)
         );
  AND2_X1 U7637 ( .A1(n6619), .A2(n6616), .ZN(n6593) );
  NAND2_X1 U7638 ( .A1(n5033), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6602) );
  INV_X1 U7639 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7918) );
  OR2_X1 U7640 ( .A1(n9815), .A2(n7918), .ZN(n6601) );
  INV_X1 U7641 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6594) );
  OAI21_X1 U7642 ( .B1(n6596), .B2(n6595), .A(n6594), .ZN(n6597) );
  NAND2_X1 U7643 ( .A1(n6597), .A2(n6625), .ZN(n8033) );
  OR2_X1 U7644 ( .A1(n6910), .A2(n8033), .ZN(n6600) );
  INV_X1 U7645 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6598) );
  OR2_X1 U7646 ( .A1(n9813), .A2(n6598), .ZN(n6599) );
  NAND2_X1 U7647 ( .A1(n7208), .A2(n9807), .ZN(n6607) );
  INV_X1 U7648 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U7649 ( .A1(n6603), .A2(n9630), .ZN(n6604) );
  NAND2_X1 U7650 ( .A1(n6604), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6605) );
  XNOR2_X1 U7651 ( .A(n6605), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U7652 ( .A1(n6792), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7243), .B2(
        n10177), .ZN(n6606) );
  NAND2_X1 U7653 ( .A1(n8125), .A2(n6922), .ZN(n6608) );
  OAI21_X1 U7654 ( .B1(n7909), .B2(n6920), .A(n6608), .ZN(n6609) );
  XNOR2_X1 U7655 ( .A(n6609), .B(n6918), .ZN(n6611) );
  AND2_X1 U7656 ( .A1(n8125), .A2(n6434), .ZN(n6610) );
  AOI21_X1 U7657 ( .B1(n10101), .B2(n6915), .A(n6610), .ZN(n6612) );
  NAND2_X1 U7658 ( .A1(n6611), .A2(n6612), .ZN(n6623) );
  INV_X1 U7659 ( .A(n6611), .ZN(n6614) );
  INV_X1 U7660 ( .A(n6612), .ZN(n6613) );
  NAND2_X1 U7661 ( .A1(n6614), .A2(n6613), .ZN(n6615) );
  AND2_X1 U7662 ( .A1(n6623), .A2(n6615), .ZN(n8028) );
  INV_X1 U7663 ( .A(n6616), .ZN(n6618) );
  AND2_X1 U7664 ( .A1(n7814), .A2(n6618), .ZN(n6617) );
  NAND2_X1 U7665 ( .A1(n7813), .A2(n6617), .ZN(n6621) );
  OR2_X1 U7666 ( .A1(n6616), .A2(n6619), .ZN(n6620) );
  OAI22_X1 U7667 ( .A1(n8066), .A2(n6920), .B1(n10861), .B2(n6854), .ZN(n6622)
         );
  XNOR2_X1 U7668 ( .A(n6622), .B(n6850), .ZN(n8018) );
  NAND2_X1 U7669 ( .A1(n5033), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6630) );
  INV_X1 U7670 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6624) );
  OR2_X1 U7671 ( .A1(n9813), .A2(n6624), .ZN(n6629) );
  AND2_X1 U7672 ( .A1(n6625), .A2(n8234), .ZN(n6626) );
  OR2_X1 U7673 ( .A1(n6626), .A2(n6663), .ZN(n8235) );
  OR2_X1 U7674 ( .A1(n6910), .A2(n8235), .ZN(n6628) );
  INV_X1 U7675 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8055) );
  OR2_X1 U7676 ( .A1(n9815), .A2(n8055), .ZN(n6627) );
  NAND2_X1 U7677 ( .A1(n7223), .A2(n9807), .ZN(n6634) );
  NAND2_X1 U7678 ( .A1(n6640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6632) );
  XNOR2_X1 U7679 ( .A(n6632), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U7680 ( .A1(n6792), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7243), .B2(
        n10663), .ZN(n6633) );
  NAND2_X1 U7681 ( .A1(n8155), .A2(n6922), .ZN(n6635) );
  OAI21_X1 U7682 ( .B1(n8160), .B2(n6920), .A(n6635), .ZN(n6636) );
  XNOR2_X1 U7683 ( .A(n6636), .B(n6918), .ZN(n6638) );
  NAND2_X1 U7684 ( .A1(n8155), .A2(n6434), .ZN(n6637) );
  OAI21_X1 U7685 ( .B1(n8160), .B2(n6901), .A(n6637), .ZN(n8231) );
  INV_X1 U7686 ( .A(n6638), .ZN(n6639) );
  NAND2_X1 U7687 ( .A1(n7229), .A2(n9807), .ZN(n6643) );
  NOR2_X1 U7688 ( .A1(n6640), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6659) );
  OR2_X1 U7689 ( .A1(n6659), .A2(n6577), .ZN(n6641) );
  XNOR2_X1 U7690 ( .A(n6641), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7683) );
  AOI22_X1 U7691 ( .A1(n6792), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7243), .B2(
        n7683), .ZN(n6642) );
  NAND2_X1 U7692 ( .A1(n10564), .A2(n6922), .ZN(n6651) );
  NAND2_X1 U7693 ( .A1(n6644), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6649) );
  XNOR2_X1 U7694 ( .A(n6663), .B(P1_REG3_REG_11__SCAN_IN), .ZN(n8209) );
  OR2_X1 U7695 ( .A1(n6910), .A2(n8209), .ZN(n6648) );
  NAND2_X1 U7696 ( .A1(n5033), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U7697 ( .A1(n6645), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6646) );
  NAND4_X1 U7698 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n10099)
         );
  NAND2_X1 U7699 ( .A1(n10099), .A2(n6434), .ZN(n6650) );
  NAND2_X1 U7700 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  XNOR2_X1 U7701 ( .A(n6652), .B(n6850), .ZN(n6656) );
  AND2_X1 U7702 ( .A1(n10099), .A2(n6915), .ZN(n6653) );
  AOI21_X1 U7703 ( .B1(n10564), .B2(n6434), .A(n6653), .ZN(n6654) );
  XNOR2_X1 U7704 ( .A(n6656), .B(n6654), .ZN(n8208) );
  NAND2_X1 U7705 ( .A1(n8207), .A2(n8208), .ZN(n6658) );
  INV_X1 U7706 ( .A(n6654), .ZN(n6655) );
  NAND2_X1 U7707 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  NAND2_X1 U7708 ( .A1(n6658), .A2(n6657), .ZN(n8287) );
  NAND2_X1 U7709 ( .A1(n7234), .A2(n9807), .ZN(n6661) );
  INV_X1 U7710 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U7711 ( .A1(n6659), .A2(n9638), .ZN(n6715) );
  NAND2_X1 U7712 ( .A1(n6715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6678) );
  XNOR2_X1 U7713 ( .A(n6678), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7869) );
  AOI22_X1 U7714 ( .A1(n6792), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7243), .B2(
        n7869), .ZN(n6660) );
  NAND2_X1 U7715 ( .A1(n10917), .A2(n6922), .ZN(n6670) );
  NAND2_X1 U7716 ( .A1(n6644), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6668) );
  INV_X1 U7717 ( .A(n5033), .ZN(n6829) );
  INV_X1 U7718 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6662) );
  OR2_X1 U7719 ( .A1(n6829), .A2(n6662), .ZN(n6667) );
  AOI21_X1 U7720 ( .B1(n6663), .B2(P1_REG3_REG_11__SCAN_IN), .A(
        P1_REG3_REG_12__SCAN_IN), .ZN(n6664) );
  OR2_X1 U7721 ( .A1(n6682), .A2(n6664), .ZN(n10941) );
  OR2_X1 U7722 ( .A1(n6910), .A2(n10941), .ZN(n6666) );
  INV_X1 U7723 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7675) );
  OR2_X1 U7724 ( .A1(n9813), .A2(n7675), .ZN(n6665) );
  INV_X1 U7725 ( .A(n8428), .ZN(n10098) );
  NAND2_X1 U7726 ( .A1(n10098), .A2(n6434), .ZN(n6669) );
  NAND2_X1 U7727 ( .A1(n6670), .A2(n6669), .ZN(n6671) );
  XNOR2_X1 U7728 ( .A(n6671), .B(n6918), .ZN(n6673) );
  NOR2_X1 U7729 ( .A1(n8428), .A2(n6901), .ZN(n6672) );
  AOI21_X1 U7730 ( .B1(n10917), .B2(n6434), .A(n6672), .ZN(n6674) );
  NAND2_X1 U7731 ( .A1(n6673), .A2(n6674), .ZN(n8288) );
  NAND2_X1 U7732 ( .A1(n8287), .A2(n8288), .ZN(n6677) );
  INV_X1 U7733 ( .A(n6673), .ZN(n6676) );
  INV_X1 U7734 ( .A(n6674), .ZN(n6675) );
  NAND2_X1 U7735 ( .A1(n6676), .A2(n6675), .ZN(n8289) );
  NAND2_X1 U7736 ( .A1(n7227), .A2(n9807), .ZN(n6681) );
  INV_X1 U7737 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U7738 ( .A1(n6678), .A2(n9639), .ZN(n6679) );
  NAND2_X1 U7739 ( .A1(n6679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6695) );
  XNOR2_X1 U7740 ( .A(n6695), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8179) );
  AOI22_X1 U7741 ( .A1(n6792), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7243), .B2(
        n8179), .ZN(n6680) );
  NAND2_X1 U7742 ( .A1(n8478), .A2(n6922), .ZN(n6689) );
  NAND2_X1 U7743 ( .A1(n5033), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6687) );
  INV_X1 U7744 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7863) );
  OR2_X1 U7745 ( .A1(n9813), .A2(n7863), .ZN(n6686) );
  OR2_X1 U7746 ( .A1(n6682), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6683) );
  NAND2_X1 U7747 ( .A1(n6701), .A2(n6683), .ZN(n8437) );
  OR2_X1 U7748 ( .A1(n6910), .A2(n8437), .ZN(n6685) );
  INV_X1 U7749 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8438) );
  OR2_X1 U7750 ( .A1(n9815), .A2(n8438), .ZN(n6684) );
  INV_X1 U7751 ( .A(n10926), .ZN(n10097) );
  NAND2_X1 U7752 ( .A1(n10097), .A2(n6434), .ZN(n6688) );
  NAND2_X1 U7753 ( .A1(n6689), .A2(n6688), .ZN(n6690) );
  XNOR2_X1 U7754 ( .A(n6690), .B(n6850), .ZN(n8331) );
  NAND2_X1 U7755 ( .A1(n8478), .A2(n6434), .ZN(n6692) );
  NAND2_X1 U7756 ( .A1(n10097), .A2(n6915), .ZN(n6691) );
  NAND2_X1 U7757 ( .A1(n6692), .A2(n6691), .ZN(n8330) );
  OAI21_X1 U7758 ( .B1(n8333), .B2(n8331), .A(n8330), .ZN(n6694) );
  NAND2_X1 U7759 ( .A1(n8333), .A2(n8331), .ZN(n6693) );
  NAND2_X1 U7760 ( .A1(n7236), .A2(n9807), .ZN(n6699) );
  INV_X1 U7761 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U7762 ( .A1(n6695), .A2(n9412), .ZN(n6696) );
  NAND2_X1 U7763 ( .A1(n6696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6697) );
  XNOR2_X1 U7764 ( .A(n6697), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U7765 ( .A1(n6792), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7243), .B2(
        n10189), .ZN(n6698) );
  NAND2_X1 U7766 ( .A1(n9831), .A2(n6922), .ZN(n6708) );
  NAND2_X1 U7767 ( .A1(n5033), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6706) );
  INV_X1 U7768 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8472) );
  OR2_X1 U7769 ( .A1(n9815), .A2(n8472), .ZN(n6705) );
  NAND2_X1 U7770 ( .A1(n6701), .A2(n6700), .ZN(n6702) );
  NAND2_X1 U7771 ( .A1(n6719), .A2(n6702), .ZN(n8471) );
  OR2_X1 U7772 ( .A1(n6910), .A2(n8471), .ZN(n6704) );
  INV_X1 U7773 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8171) );
  OR2_X1 U7774 ( .A1(n9813), .A2(n8171), .ZN(n6703) );
  NAND2_X1 U7775 ( .A1(n10096), .A2(n6434), .ZN(n6707) );
  NAND2_X1 U7776 ( .A1(n6708), .A2(n6707), .ZN(n6709) );
  XNOR2_X1 U7777 ( .A(n6709), .B(n6850), .ZN(n8448) );
  NAND2_X1 U7778 ( .A1(n9831), .A2(n6434), .ZN(n6711) );
  NAND2_X1 U7779 ( .A1(n10096), .A2(n6915), .ZN(n6710) );
  NAND2_X1 U7780 ( .A1(n6711), .A2(n6710), .ZN(n8449) );
  NAND2_X1 U7781 ( .A1(n7373), .A2(n9807), .ZN(n6718) );
  NAND3_X1 U7782 ( .A1(n9640), .A2(n9412), .A3(n9639), .ZN(n6714) );
  OR2_X1 U7783 ( .A1(n6715), .A2(n6714), .ZN(n6731) );
  NAND2_X1 U7784 ( .A1(n6731), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6716) );
  XNOR2_X1 U7785 ( .A(n6716), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U7786 ( .A1(n6792), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7243), .B2(
        n10205), .ZN(n6717) );
  NAND2_X1 U7787 ( .A1(n8569), .A2(n6922), .ZN(n6727) );
  NAND2_X1 U7788 ( .A1(n5033), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6725) );
  INV_X1 U7789 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8499) );
  OR2_X1 U7790 ( .A1(n9815), .A2(n8499), .ZN(n6724) );
  NAND2_X1 U7791 ( .A1(n6719), .A2(n10184), .ZN(n6720) );
  NAND2_X1 U7792 ( .A1(n6736), .A2(n6720), .ZN(n8554) );
  OR2_X1 U7793 ( .A1(n6910), .A2(n8554), .ZN(n6723) );
  INV_X1 U7794 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6721) );
  OR2_X1 U7795 ( .A1(n9813), .A2(n6721), .ZN(n6722) );
  INV_X1 U7796 ( .A(n10555), .ZN(n10095) );
  NAND2_X1 U7797 ( .A1(n10095), .A2(n6434), .ZN(n6726) );
  NAND2_X1 U7798 ( .A1(n6727), .A2(n6726), .ZN(n6728) );
  XNOR2_X1 U7799 ( .A(n6728), .B(n6850), .ZN(n8547) );
  NAND2_X1 U7800 ( .A1(n8569), .A2(n6434), .ZN(n6730) );
  NAND2_X1 U7801 ( .A1(n10095), .A2(n6915), .ZN(n6729) );
  NAND2_X1 U7802 ( .A1(n6730), .A2(n6729), .ZN(n8551) );
  NAND2_X1 U7803 ( .A1(n7401), .A2(n9807), .ZN(n6733) );
  OAI21_X1 U7804 ( .B1(n6731), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6752) );
  XNOR2_X1 U7805 ( .A(n6752), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U7806 ( .A1(n6792), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7243), .B2(
        n10222), .ZN(n6732) );
  NAND2_X1 U7807 ( .A1(n10557), .A2(n6922), .ZN(n6743) );
  NAND2_X1 U7808 ( .A1(n6644), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6741) );
  INV_X1 U7809 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6734) );
  OR2_X1 U7810 ( .A1(n6829), .A2(n6734), .ZN(n6740) );
  AND2_X1 U7811 ( .A1(n6736), .A2(n6735), .ZN(n6737) );
  OR2_X1 U7812 ( .A1(n6737), .A2(n6757), .ZN(n11015) );
  OR2_X1 U7813 ( .A1(n6910), .A2(n11015), .ZN(n6739) );
  INV_X1 U7814 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10224) );
  OR2_X1 U7815 ( .A1(n9813), .A2(n10224), .ZN(n6738) );
  INV_X1 U7816 ( .A(n10453), .ZN(n10094) );
  NAND2_X1 U7817 ( .A1(n10094), .A2(n6434), .ZN(n6742) );
  NAND2_X1 U7818 ( .A1(n6743), .A2(n6742), .ZN(n6744) );
  XNOR2_X1 U7819 ( .A(n6744), .B(n6918), .ZN(n6746) );
  NOR2_X1 U7820 ( .A1(n10453), .A2(n6901), .ZN(n6745) );
  AOI21_X1 U7821 ( .B1(n10557), .B2(n6434), .A(n6745), .ZN(n6747) );
  NAND2_X1 U7822 ( .A1(n6746), .A2(n6747), .ZN(n6751) );
  INV_X1 U7823 ( .A(n6746), .ZN(n6749) );
  INV_X1 U7824 ( .A(n6747), .ZN(n6748) );
  NAND2_X1 U7825 ( .A1(n6749), .A2(n6748), .ZN(n6750) );
  AND2_X1 U7826 ( .A1(n6751), .A2(n6750), .ZN(n9737) );
  NAND2_X1 U7827 ( .A1(n7502), .A2(n9807), .ZN(n6755) );
  INV_X1 U7828 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U7829 ( .A1(n6752), .A2(n9648), .ZN(n6753) );
  NAND2_X1 U7830 ( .A1(n6753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6771) );
  XNOR2_X1 U7831 ( .A(n6771), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U7832 ( .A1(n6792), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7243), .B2(
        n10238), .ZN(n6754) );
  NAND2_X1 U7833 ( .A1(n10543), .A2(n6922), .ZN(n6764) );
  NAND2_X1 U7834 ( .A1(n6644), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6762) );
  INV_X1 U7835 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n6756) );
  OR2_X1 U7836 ( .A1(n6829), .A2(n6756), .ZN(n6761) );
  OR2_X1 U7837 ( .A1(n6757), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U7838 ( .A1(n6778), .A2(n6758), .ZN(n10462) );
  OR2_X1 U7839 ( .A1(n6910), .A2(n10462), .ZN(n6760) );
  INV_X1 U7840 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10233) );
  OR2_X1 U7841 ( .A1(n9813), .A2(n10233), .ZN(n6759) );
  INV_X1 U7842 ( .A(n10556), .ZN(n10093) );
  NAND2_X1 U7843 ( .A1(n10093), .A2(n6434), .ZN(n6763) );
  NAND2_X1 U7844 ( .A1(n6764), .A2(n6763), .ZN(n6765) );
  XNOR2_X1 U7845 ( .A(n6765), .B(n6850), .ZN(n6767) );
  NOR2_X1 U7846 ( .A1(n10556), .A2(n6901), .ZN(n6766) );
  AOI21_X1 U7847 ( .B1(n10543), .B2(n6434), .A(n6766), .ZN(n6768) );
  XNOR2_X1 U7848 ( .A(n6767), .B(n6768), .ZN(n9747) );
  NAND2_X1 U7849 ( .A1(n9745), .A2(n9747), .ZN(n9746) );
  INV_X1 U7850 ( .A(n6767), .ZN(n6769) );
  NAND2_X1 U7851 ( .A1(n6769), .A2(n6768), .ZN(n6770) );
  NAND2_X1 U7852 ( .A1(n7579), .A2(n9807), .ZN(n6775) );
  INV_X1 U7853 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U7854 ( .A1(n6771), .A2(n9649), .ZN(n6772) );
  NAND2_X1 U7855 ( .A1(n6772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6773) );
  XNOR2_X1 U7856 ( .A(n6773), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U7857 ( .A1(n6792), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7243), .B2(
        n10255), .ZN(n6774) );
  NAND2_X1 U7858 ( .A1(n10538), .A2(n6922), .ZN(n6785) );
  NAND2_X1 U7859 ( .A1(n6644), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6783) );
  INV_X1 U7860 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n6776) );
  OR2_X1 U7861 ( .A1(n6829), .A2(n6776), .ZN(n6782) );
  NAND2_X1 U7862 ( .A1(n6778), .A2(n6777), .ZN(n6779) );
  NAND2_X1 U7863 ( .A1(n6796), .A2(n6779), .ZN(n9789) );
  OR2_X1 U7864 ( .A1(n6910), .A2(n9789), .ZN(n6781) );
  INV_X1 U7865 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10230) );
  OR2_X1 U7866 ( .A1(n9813), .A2(n10230), .ZN(n6780) );
  INV_X1 U7867 ( .A(n10454), .ZN(n10446) );
  NAND2_X1 U7868 ( .A1(n10446), .A2(n6434), .ZN(n6784) );
  NAND2_X1 U7869 ( .A1(n6785), .A2(n6784), .ZN(n6786) );
  XNOR2_X1 U7870 ( .A(n6786), .B(n6850), .ZN(n6789) );
  NOR2_X1 U7871 ( .A1(n10454), .A2(n6901), .ZN(n6787) );
  AOI21_X1 U7872 ( .B1(n10538), .B2(n6434), .A(n6787), .ZN(n9785) );
  INV_X1 U7873 ( .A(n6788), .ZN(n6791) );
  INV_X1 U7874 ( .A(n6789), .ZN(n6790) );
  NAND2_X1 U7875 ( .A1(n6791), .A2(n6790), .ZN(n9788) );
  NAND2_X1 U7876 ( .A1(n7624), .A2(n9807), .ZN(n6794) );
  AOI22_X1 U7877 ( .A1(n6792), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10785), 
        .B2(n7243), .ZN(n6793) );
  NAND2_X1 U7878 ( .A1(n10532), .A2(n6922), .ZN(n6803) );
  NAND2_X1 U7879 ( .A1(n5033), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U7880 ( .A1(n6645), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6800) );
  AND2_X1 U7881 ( .A1(n6796), .A2(n9713), .ZN(n6797) );
  NOR2_X1 U7882 ( .A1(n6810), .A2(n6797), .ZN(n10440) );
  NAND2_X1 U7883 ( .A1(n6795), .A2(n10440), .ZN(n6799) );
  NAND2_X1 U7884 ( .A1(n6644), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6798) );
  NAND4_X1 U7885 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n10421)
         );
  NAND2_X1 U7886 ( .A1(n10421), .A2(n6434), .ZN(n6802) );
  NAND2_X1 U7887 ( .A1(n6803), .A2(n6802), .ZN(n6804) );
  XNOR2_X1 U7888 ( .A(n6804), .B(n6850), .ZN(n6806) );
  INV_X1 U7889 ( .A(n10421), .ZN(n9790) );
  OAI22_X1 U7890 ( .A1(n10442), .A2(n6920), .B1(n9790), .B2(n6901), .ZN(n6805)
         );
  XOR2_X1 U7891 ( .A(n6806), .B(n6805), .Z(n9711) );
  NAND2_X1 U7892 ( .A1(n7809), .A2(n9807), .ZN(n6809) );
  OR2_X1 U7893 ( .A1(n9822), .A2(n9592), .ZN(n6808) );
  NAND2_X1 U7894 ( .A1(n10526), .A2(n6922), .ZN(n6817) );
  NAND2_X1 U7895 ( .A1(n5033), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U7896 ( .A1(n6644), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6814) );
  NOR2_X1 U7897 ( .A1(n6810), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6811) );
  OR2_X1 U7898 ( .A1(n6825), .A2(n6811), .ZN(n9771) );
  INV_X1 U7899 ( .A(n9771), .ZN(n10428) );
  NAND2_X1 U7900 ( .A1(n6795), .A2(n10428), .ZN(n6813) );
  NAND2_X1 U7901 ( .A1(n6645), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6812) );
  NAND4_X1 U7902 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n10447)
         );
  NAND2_X1 U7903 ( .A1(n10447), .A2(n6434), .ZN(n6816) );
  NAND2_X1 U7904 ( .A1(n6817), .A2(n6816), .ZN(n6818) );
  XNOR2_X1 U7905 ( .A(n6818), .B(n6850), .ZN(n6822) );
  NAND2_X1 U7906 ( .A1(n10526), .A2(n6434), .ZN(n6820) );
  NAND2_X1 U7907 ( .A1(n10447), .A2(n6915), .ZN(n6819) );
  NAND2_X1 U7908 ( .A1(n6820), .A2(n6819), .ZN(n6821) );
  NOR2_X1 U7909 ( .A1(n6822), .A2(n6821), .ZN(n9765) );
  NAND2_X1 U7910 ( .A1(n6822), .A2(n6821), .ZN(n9766) );
  NAND2_X1 U7911 ( .A1(n7823), .A2(n9807), .ZN(n6824) );
  INV_X1 U7912 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8633) );
  OR2_X1 U7913 ( .A1(n9822), .A2(n8633), .ZN(n6823) );
  NAND2_X1 U7914 ( .A1(n10518), .A2(n6922), .ZN(n6837) );
  OR2_X1 U7915 ( .A1(n6825), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6827) );
  AND2_X1 U7916 ( .A1(n6827), .A2(n6826), .ZN(n9723) );
  NAND2_X1 U7917 ( .A1(n9723), .A2(n6795), .ZN(n6835) );
  INV_X1 U7918 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n10411) );
  OR2_X1 U7919 ( .A1(n9815), .A2(n10411), .ZN(n6834) );
  INV_X1 U7920 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n6828) );
  OR2_X1 U7921 ( .A1(n6829), .A2(n6828), .ZN(n6833) );
  INV_X1 U7922 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6830) );
  OR2_X1 U7923 ( .A1(n6831), .A2(n6830), .ZN(n6832) );
  INV_X1 U7924 ( .A(n10385), .ZN(n10422) );
  NAND2_X1 U7925 ( .A1(n10422), .A2(n6434), .ZN(n6836) );
  NAND2_X1 U7926 ( .A1(n6837), .A2(n6836), .ZN(n6838) );
  XNOR2_X1 U7927 ( .A(n6838), .B(n6918), .ZN(n6841) );
  NOR2_X1 U7928 ( .A1(n10385), .A2(n6901), .ZN(n6839) );
  AOI21_X1 U7929 ( .B1(n10518), .B2(n6434), .A(n6839), .ZN(n6840) );
  NOR2_X1 U7930 ( .A1(n6841), .A2(n6840), .ZN(n9718) );
  NAND2_X1 U7931 ( .A1(n8038), .A2(n9807), .ZN(n6843) );
  OR2_X1 U7932 ( .A1(n9822), .A2(n9588), .ZN(n6842) );
  NAND2_X1 U7933 ( .A1(n6644), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6849) );
  OAI21_X1 U7934 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n6845), .A(n6844), .ZN(
        n10390) );
  OR2_X1 U7935 ( .A1(n6910), .A2(n10390), .ZN(n6848) );
  NAND2_X1 U7936 ( .A1(n5033), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6847) );
  NAND2_X1 U7937 ( .A1(n6645), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6846) );
  NAND4_X1 U7938 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n10404)
         );
  OAI22_X1 U7939 ( .A1(n10394), .A2(n6854), .B1(n9722), .B2(n6920), .ZN(n6851)
         );
  XNOR2_X1 U7940 ( .A(n6851), .B(n6850), .ZN(n6853) );
  OAI22_X1 U7941 ( .A1(n10394), .A2(n6920), .B1(n9722), .B2(n6901), .ZN(n6852)
         );
  NAND2_X1 U7942 ( .A1(n6853), .A2(n6852), .ZN(n9776) );
  OAI22_X1 U7943 ( .A1(n10374), .A2(n6854), .B1(n10387), .B2(n6920), .ZN(n6855) );
  XNOR2_X1 U7944 ( .A(n6855), .B(n6850), .ZN(n6856) );
  NAND2_X1 U7945 ( .A1(n8204), .A2(n9807), .ZN(n6859) );
  INV_X1 U7946 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8226) );
  OR2_X1 U7947 ( .A1(n9822), .A2(n8226), .ZN(n6858) );
  NAND2_X1 U7948 ( .A1(n6644), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U7949 ( .A1(n5033), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6865) );
  NOR2_X1 U7950 ( .A1(n6860), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6861) );
  NOR2_X1 U7951 ( .A1(n6862), .A2(n6861), .ZN(n10362) );
  NAND2_X1 U7952 ( .A1(n6795), .A2(n10362), .ZN(n6864) );
  NAND2_X1 U7953 ( .A1(n6645), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6863) );
  NAND4_X1 U7954 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n10378)
         );
  AOI22_X1 U7955 ( .A1(n10348), .A2(n6434), .B1(n6915), .B2(n10378), .ZN(n6870) );
  NAND2_X1 U7956 ( .A1(n10348), .A2(n6922), .ZN(n6868) );
  NAND2_X1 U7957 ( .A1(n10378), .A2(n6434), .ZN(n6867) );
  NAND2_X1 U7958 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  XNOR2_X1 U7959 ( .A(n6869), .B(n6850), .ZN(n6872) );
  XOR2_X1 U7960 ( .A(n6870), .B(n6872), .Z(n9754) );
  INV_X1 U7961 ( .A(n6870), .ZN(n6871) );
  OR2_X1 U7962 ( .A1(n9822), .A2(n9580), .ZN(n6875) );
  NAND2_X1 U7963 ( .A1(n10493), .A2(n6922), .ZN(n6884) );
  NAND2_X1 U7964 ( .A1(n5033), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6882) );
  INV_X1 U7965 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6877) );
  OR2_X1 U7966 ( .A1(n9813), .A2(n6877), .ZN(n6881) );
  NAND2_X1 U7967 ( .A1(n6878), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6892) );
  OAI21_X1 U7968 ( .B1(n6878), .B2(P1_REG3_REG_26__SCAN_IN), .A(n6892), .ZN(
        n10327) );
  OR2_X1 U7969 ( .A1(n6910), .A2(n10327), .ZN(n6880) );
  INV_X1 U7970 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10328) );
  OR2_X1 U7971 ( .A1(n9815), .A2(n10328), .ZN(n6879) );
  INV_X1 U7972 ( .A(n10344), .ZN(n10298) );
  NAND2_X1 U7973 ( .A1(n10298), .A2(n6434), .ZN(n6883) );
  NAND2_X1 U7974 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  XNOR2_X1 U7975 ( .A(n6885), .B(n6918), .ZN(n6887) );
  NOR2_X1 U7976 ( .A1(n10344), .A2(n6901), .ZN(n6886) );
  AOI21_X1 U7977 ( .B1(n10493), .B2(n6434), .A(n6886), .ZN(n6888) );
  XNOR2_X1 U7978 ( .A(n6887), .B(n6888), .ZN(n9795) );
  NAND2_X1 U7979 ( .A1(n8506), .A2(n9807), .ZN(n6890) );
  INV_X1 U7980 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8507) );
  OR2_X1 U7981 ( .A1(n9822), .A2(n8507), .ZN(n6889) );
  NAND2_X1 U7982 ( .A1(n10488), .A2(n6922), .ZN(n6899) );
  NAND2_X1 U7983 ( .A1(n5033), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6897) );
  INV_X1 U7984 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6891) );
  OR2_X1 U7985 ( .A1(n9813), .A2(n6891), .ZN(n6896) );
  INV_X1 U7986 ( .A(n6892), .ZN(n6893) );
  NAND2_X1 U7987 ( .A1(n6893), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6908) );
  OAI21_X1 U7988 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n6893), .A(n6908), .ZN(
        n10307) );
  OR2_X1 U7989 ( .A1(n6910), .A2(n10307), .ZN(n6895) );
  INV_X1 U7990 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10308) );
  OR2_X1 U7991 ( .A1(n9815), .A2(n10308), .ZN(n6894) );
  INV_X1 U7992 ( .A(n10322), .ZN(n10092) );
  NAND2_X1 U7993 ( .A1(n10092), .A2(n6434), .ZN(n6898) );
  NAND2_X1 U7994 ( .A1(n6899), .A2(n6898), .ZN(n6900) );
  XNOR2_X1 U7995 ( .A(n6900), .B(n6918), .ZN(n6904) );
  NOR2_X1 U7996 ( .A1(n10322), .A2(n6901), .ZN(n6902) );
  AOI21_X1 U7997 ( .B1(n10488), .B2(n6434), .A(n6902), .ZN(n6903) );
  NAND2_X1 U7998 ( .A1(n6904), .A2(n6903), .ZN(n6949) );
  OAI21_X1 U7999 ( .B1(n6904), .B2(n6903), .A(n6949), .ZN(n7146) );
  NAND2_X1 U8000 ( .A1(n8545), .A2(n9807), .ZN(n6906) );
  INV_X1 U8001 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8567) );
  OR2_X1 U8002 ( .A1(n9822), .A2(n8567), .ZN(n6905) );
  NAND2_X1 U8003 ( .A1(n10481), .A2(n6434), .ZN(n6917) );
  NAND2_X1 U8004 ( .A1(n5033), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6914) );
  INV_X1 U8005 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6907) );
  OR2_X1 U8006 ( .A1(n9813), .A2(n6907), .ZN(n6913) );
  INV_X1 U8007 ( .A(n6908), .ZN(n6909) );
  NAND2_X1 U8008 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n6909), .ZN(n8796) );
  OAI21_X1 U8009 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n6909), .A(n8796), .ZN(
        n10287) );
  OR2_X1 U8010 ( .A1(n6910), .A2(n10287), .ZN(n6912) );
  INV_X1 U8011 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10288) );
  OR2_X1 U8012 ( .A1(n9815), .A2(n10288), .ZN(n6911) );
  NAND2_X1 U8013 ( .A1(n10297), .A2(n6915), .ZN(n6916) );
  NAND2_X1 U8014 ( .A1(n6917), .A2(n6916), .ZN(n6919) );
  XNOR2_X1 U8015 ( .A(n6919), .B(n6918), .ZN(n6924) );
  NOR2_X1 U8016 ( .A1(n8790), .A2(n6920), .ZN(n6921) );
  AOI21_X1 U8017 ( .B1(n10481), .B2(n6922), .A(n6921), .ZN(n6923) );
  NAND2_X1 U8018 ( .A1(n8312), .A2(P1_B_REG_SCAN_IN), .ZN(n6926) );
  MUX2_X1 U8019 ( .A(n6926), .B(P1_B_REG_SCAN_IN), .S(n6925), .Z(n6927) );
  INV_X1 U8020 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U8021 ( .A1(n10587), .A2(n9446), .ZN(n6930) );
  INV_X1 U8022 ( .A(n6928), .ZN(n8468) );
  NAND2_X1 U8023 ( .A1(n8468), .A2(n8312), .ZN(n6929) );
  NAND2_X1 U8024 ( .A1(n6930), .A2(n6929), .ZN(n7379) );
  INV_X1 U8025 ( .A(n7379), .ZN(n10586) );
  NOR4_X1 U8026 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6934) );
  NOR4_X1 U8027 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6933) );
  NOR4_X1 U8028 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6932) );
  NOR4_X1 U8029 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6931) );
  NAND4_X1 U8030 ( .A1(n6934), .A2(n6933), .A3(n6932), .A4(n6931), .ZN(n6940)
         );
  NOR2_X1 U8031 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n6938) );
  NOR4_X1 U8032 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6937) );
  NOR4_X1 U8033 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6936) );
  NOR4_X1 U8034 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6935) );
  NAND4_X1 U8035 ( .A1(n6938), .A2(n6937), .A3(n6936), .A4(n6935), .ZN(n6939)
         );
  OAI21_X1 U8036 ( .B1(n6940), .B2(n6939), .A(n10587), .ZN(n7378) );
  AND2_X1 U8037 ( .A1(n10586), .A2(n7378), .ZN(n7827) );
  INV_X1 U8038 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U8039 ( .A1(n10587), .A2(n6941), .ZN(n6942) );
  INV_X1 U8040 ( .A(n6925), .ZN(n8228) );
  NAND2_X1 U8041 ( .A1(n8468), .A2(n8228), .ZN(n10590) );
  NAND2_X1 U8042 ( .A1(n6942), .A2(n10590), .ZN(n7387) );
  INV_X1 U8043 ( .A(n7387), .ZN(n6943) );
  NAND2_X1 U8044 ( .A1(n7827), .A2(n6943), .ZN(n7495) );
  OAI21_X1 U8045 ( .B1(n6945), .B2(n9431), .A(n6944), .ZN(n8135) );
  AND2_X1 U8046 ( .A1(n8135), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6946) );
  INV_X1 U8047 ( .A(n10588), .ZN(n10585) );
  OR2_X1 U8048 ( .A1(n7495), .A2(n10585), .ZN(n6951) );
  NAND2_X1 U8049 ( .A1(n8124), .A2(n6947), .ZN(n7383) );
  INV_X1 U8050 ( .A(n7383), .ZN(n7381) );
  INV_X1 U8051 ( .A(n10083), .ZN(n10081) );
  INV_X1 U8052 ( .A(n7155), .ZN(n10033) );
  OR2_X1 U8053 ( .A1(n10827), .A2(n10033), .ZN(n6961) );
  NAND2_X1 U8054 ( .A1(n6949), .A2(n9756), .ZN(n6948) );
  NAND3_X1 U8055 ( .A1(n7149), .A2(n5076), .A3(n9756), .ZN(n6973) );
  INV_X1 U8056 ( .A(n6949), .ZN(n6950) );
  NAND3_X1 U8057 ( .A1(n5076), .A2(n6950), .A3(n9756), .ZN(n6971) );
  NOR2_X1 U8058 ( .A1(n7383), .A2(n7822), .ZN(n10780) );
  OAI211_X1 U8059 ( .C1(n10033), .C2(n10780), .A(n7495), .B(n10588), .ZN(n6966) );
  OR2_X1 U8060 ( .A1(n7155), .A2(n10083), .ZN(n6962) );
  NAND2_X1 U8061 ( .A1(n10588), .A2(n6962), .ZN(n7386) );
  INV_X1 U8062 ( .A(n7386), .ZN(n7377) );
  NAND2_X1 U8063 ( .A1(n6966), .A2(n7377), .ZN(n9764) );
  NOR2_X1 U8064 ( .A1(n6951), .A2(n10081), .ZN(n6954) );
  INV_X1 U8065 ( .A(n6952), .ZN(n7264) );
  NAND2_X1 U8066 ( .A1(n6954), .A2(n10768), .ZN(n9800) );
  INV_X1 U8067 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6953) );
  OAI22_X1 U8068 ( .A1(n9800), .A2(n10322), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6953), .ZN(n6969) );
  NAND2_X1 U8069 ( .A1(n6954), .A2(n10769), .ZN(n9798) );
  NAND2_X1 U8070 ( .A1(n5033), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6960) );
  INV_X1 U8071 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6955) );
  OR2_X1 U8072 ( .A1(n9813), .A2(n6955), .ZN(n6959) );
  OR2_X1 U8073 ( .A1(n6910), .A2(n8796), .ZN(n6958) );
  INV_X1 U8074 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6956) );
  OR2_X1 U8075 ( .A1(n9815), .A2(n6956), .ZN(n6957) );
  INV_X1 U8076 ( .A(n6961), .ZN(n6964) );
  NAND3_X1 U8077 ( .A1(n6418), .A2(n8135), .A3(n6962), .ZN(n6963) );
  AOI21_X1 U8078 ( .B1(n7495), .B2(n6964), .A(n6963), .ZN(n6965) );
  OR2_X1 U8079 ( .A1(n6965), .A2(P1_U3084), .ZN(n6967) );
  AND2_X2 U8080 ( .A1(n6967), .A2(n6966), .ZN(n9799) );
  OAI22_X1 U8081 ( .A1(n9798), .A2(n10284), .B1(n9799), .B2(n10287), .ZN(n6968) );
  AOI211_X1 U8082 ( .C1(n10481), .C2(n9803), .A(n6969), .B(n6968), .ZN(n6970)
         );
  AND2_X1 U8083 ( .A1(n6971), .A2(n6970), .ZN(n6972) );
  NAND3_X1 U8084 ( .A1(n6974), .A2(n6973), .A3(n6972), .ZN(P1_U3218) );
  NAND2_X1 U8085 ( .A1(n8901), .A2(n7036), .ZN(n6980) );
  NAND2_X1 U8086 ( .A1(n6975), .A2(n9004), .ZN(n7426) );
  NAND2_X1 U8087 ( .A1(n7426), .A2(n7825), .ZN(n6976) );
  INV_X1 U8088 ( .A(n7546), .ZN(n6979) );
  NAND2_X1 U8089 ( .A1(n7513), .A2(n7109), .ZN(n6977) );
  NAND2_X1 U8090 ( .A1(n6980), .A2(n8636), .ZN(n6981) );
  NAND2_X1 U8091 ( .A1(n8639), .A2(n6981), .ZN(n6982) );
  NAND2_X1 U8092 ( .A1(n10730), .A2(n7036), .ZN(n6985) );
  INV_X2 U8093 ( .A(n7109), .ZN(n7103) );
  XNOR2_X1 U8094 ( .A(n8641), .B(n7103), .ZN(n6983) );
  XNOR2_X1 U8095 ( .A(n6985), .B(n6983), .ZN(n8637) );
  INV_X1 U8096 ( .A(n6983), .ZN(n6984) );
  NAND2_X1 U8097 ( .A1(n6985), .A2(n6984), .ZN(n6986) );
  AND2_X1 U8098 ( .A1(n8900), .A2(n7036), .ZN(n6987) );
  XNOR2_X1 U8099 ( .A(n10732), .B(n7103), .ZN(n6988) );
  NAND2_X1 U8100 ( .A1(n6987), .A2(n6988), .ZN(n6991) );
  INV_X1 U8101 ( .A(n6987), .ZN(n6989) );
  INV_X1 U8102 ( .A(n6988), .ZN(n7592) );
  NAND2_X1 U8103 ( .A1(n6989), .A2(n7592), .ZN(n6990) );
  AND2_X1 U8104 ( .A1(n6991), .A2(n6990), .ZN(n10729) );
  NAND2_X1 U8105 ( .A1(n8899), .A2(n7036), .ZN(n6994) );
  XNOR2_X1 U8106 ( .A(n7727), .B(n7103), .ZN(n6993) );
  XNOR2_X1 U8107 ( .A(n6994), .B(n6993), .ZN(n7604) );
  AND2_X1 U8108 ( .A1(n7604), .A2(n6991), .ZN(n7595) );
  NAND2_X1 U8109 ( .A1(n8898), .A2(n7036), .ZN(n6998) );
  XNOR2_X1 U8110 ( .A(n10806), .B(n7103), .ZN(n6997) );
  XNOR2_X1 U8111 ( .A(n6998), .B(n6997), .ZN(n6992) );
  AND2_X1 U8112 ( .A1(n7595), .A2(n6992), .ZN(n6996) );
  INV_X1 U8113 ( .A(n6992), .ZN(n8771) );
  INV_X1 U8114 ( .A(n6993), .ZN(n8768) );
  NAND2_X1 U8115 ( .A1(n6994), .A2(n8768), .ZN(n6995) );
  INV_X1 U8116 ( .A(n6997), .ZN(n8679) );
  NAND2_X1 U8117 ( .A1(n6998), .A2(n8679), .ZN(n6999) );
  NAND2_X1 U8118 ( .A1(n8897), .A2(n7036), .ZN(n7003) );
  XNOR2_X1 U8119 ( .A(n7796), .B(n7103), .ZN(n7001) );
  XNOR2_X1 U8120 ( .A(n7003), .B(n7001), .ZN(n8678) );
  INV_X1 U8121 ( .A(n7001), .ZN(n7002) );
  NAND2_X1 U8122 ( .A1(n7003), .A2(n7002), .ZN(n7004) );
  AND2_X1 U8123 ( .A1(n8896), .A2(n7036), .ZN(n7005) );
  XNOR2_X1 U8124 ( .A(n7894), .B(n7103), .ZN(n8147) );
  NAND2_X1 U8125 ( .A1(n7005), .A2(n8147), .ZN(n7010) );
  INV_X1 U8126 ( .A(n7005), .ZN(n7007) );
  INV_X1 U8127 ( .A(n8147), .ZN(n7006) );
  NAND2_X1 U8128 ( .A1(n7007), .A2(n7006), .ZN(n7008) );
  NAND2_X1 U8129 ( .A1(n7010), .A2(n7008), .ZN(n7963) );
  INV_X1 U8130 ( .A(n7963), .ZN(n7009) );
  XNOR2_X1 U8131 ( .A(n10868), .B(n7103), .ZN(n7011) );
  AND2_X1 U8132 ( .A1(n8895), .A2(n7036), .ZN(n7012) );
  NAND2_X1 U8133 ( .A1(n7011), .A2(n7012), .ZN(n7015) );
  INV_X1 U8134 ( .A(n7011), .ZN(n8093) );
  INV_X1 U8135 ( .A(n7012), .ZN(n7013) );
  NAND2_X1 U8136 ( .A1(n8093), .A2(n7013), .ZN(n7014) );
  AND2_X1 U8137 ( .A1(n7015), .A2(n7014), .ZN(n8148) );
  XNOR2_X1 U8138 ( .A(n10879), .B(n7103), .ZN(n7017) );
  NAND2_X1 U8139 ( .A1(n8894), .A2(n7036), .ZN(n7018) );
  XNOR2_X1 U8140 ( .A(n7017), .B(n7018), .ZN(n8106) );
  AND2_X1 U8141 ( .A1(n8106), .A2(n7015), .ZN(n7016) );
  INV_X1 U8142 ( .A(n7017), .ZN(n7019) );
  NAND2_X1 U8143 ( .A1(n7019), .A2(n7018), .ZN(n7020) );
  XNOR2_X1 U8144 ( .A(n8257), .B(n7103), .ZN(n7167) );
  AND2_X1 U8145 ( .A1(n8893), .A2(n7036), .ZN(n7021) );
  NAND2_X1 U8146 ( .A1(n7167), .A2(n7021), .ZN(n7026) );
  INV_X1 U8147 ( .A(n7167), .ZN(n7023) );
  INV_X1 U8148 ( .A(n7021), .ZN(n7022) );
  NAND2_X1 U8149 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  NAND2_X1 U8150 ( .A1(n7026), .A2(n7024), .ZN(n7161) );
  NAND2_X1 U8151 ( .A1(n7159), .A2(n7026), .ZN(n7031) );
  XNOR2_X1 U8152 ( .A(n10905), .B(n7103), .ZN(n7027) );
  AND2_X1 U8153 ( .A1(n8892), .A2(n7036), .ZN(n7028) );
  NAND2_X1 U8154 ( .A1(n7027), .A2(n7028), .ZN(n7032) );
  INV_X1 U8155 ( .A(n7027), .ZN(n8296) );
  INV_X1 U8156 ( .A(n7028), .ZN(n7029) );
  NAND2_X1 U8157 ( .A1(n8296), .A2(n7029), .ZN(n7030) );
  AND2_X1 U8158 ( .A1(n7032), .A2(n7030), .ZN(n7168) );
  XNOR2_X1 U8159 ( .A(n8609), .B(n7103), .ZN(n8707) );
  NAND2_X1 U8160 ( .A1(n8891), .A2(n7036), .ZN(n7040) );
  XNOR2_X1 U8161 ( .A(n8707), .B(n7040), .ZN(n8307) );
  AND2_X1 U8162 ( .A1(n8307), .A2(n7032), .ZN(n8299) );
  NAND2_X1 U8163 ( .A1(n8889), .A2(n7036), .ZN(n7037) );
  XNOR2_X1 U8164 ( .A(n8713), .B(n7103), .ZN(n8738) );
  INV_X1 U8165 ( .A(n8738), .ZN(n7033) );
  NAND2_X1 U8166 ( .A1(n8890), .A2(n7036), .ZN(n7034) );
  XNOR2_X1 U8167 ( .A(n8738), .B(n7034), .ZN(n8709) );
  AND2_X1 U8168 ( .A1(n8709), .A2(n8740), .ZN(n7035) );
  AND2_X1 U8169 ( .A1(n8299), .A2(n7039), .ZN(n8728) );
  XNOR2_X1 U8170 ( .A(n8760), .B(n7103), .ZN(n8691) );
  NAND2_X1 U8171 ( .A1(n8888), .A2(n7036), .ZN(n7046) );
  XNOR2_X1 U8172 ( .A(n8691), .B(n7046), .ZN(n8756) );
  AND2_X1 U8173 ( .A1(n8728), .A2(n8756), .ZN(n7045) );
  INV_X1 U8174 ( .A(n8756), .ZN(n7044) );
  INV_X1 U8175 ( .A(n8754), .ZN(n7038) );
  NAND2_X1 U8176 ( .A1(n7038), .A2(n7037), .ZN(n7042) );
  INV_X1 U8177 ( .A(n8707), .ZN(n7041) );
  NAND2_X1 U8178 ( .A1(n7041), .A2(n7040), .ZN(n8699) );
  INV_X1 U8179 ( .A(n8691), .ZN(n7047) );
  NAND2_X1 U8180 ( .A1(n7047), .A2(n7046), .ZN(n7048) );
  NAND2_X1 U8181 ( .A1(n8762), .A2(n7048), .ZN(n7049) );
  XNOR2_X1 U8182 ( .A(n9229), .B(n7103), .ZN(n7050) );
  NAND2_X1 U8183 ( .A1(n8887), .A2(n7036), .ZN(n7051) );
  XNOR2_X1 U8184 ( .A(n7050), .B(n7051), .ZN(n8693) );
  INV_X1 U8185 ( .A(n7050), .ZN(n7052) );
  NAND2_X1 U8186 ( .A1(n7052), .A2(n7051), .ZN(n7053) );
  XNOR2_X1 U8187 ( .A(n9223), .B(n7109), .ZN(n7055) );
  NAND2_X1 U8188 ( .A1(n9138), .A2(n7036), .ZN(n7056) );
  AND2_X1 U8189 ( .A1(n7055), .A2(n7056), .ZN(n8458) );
  INV_X1 U8190 ( .A(n8458), .ZN(n7054) );
  INV_X1 U8191 ( .A(n7055), .ZN(n7058) );
  INV_X1 U8192 ( .A(n7056), .ZN(n7057) );
  NAND2_X1 U8193 ( .A1(n7058), .A2(n7057), .ZN(n8459) );
  XNOR2_X1 U8194 ( .A(n9216), .B(n7103), .ZN(n7060) );
  AND2_X1 U8195 ( .A1(n9109), .A2(n7036), .ZN(n7061) );
  AND2_X1 U8196 ( .A1(n7060), .A2(n7061), .ZN(n8526) );
  INV_X1 U8197 ( .A(n7060), .ZN(n7063) );
  INV_X1 U8198 ( .A(n7061), .ZN(n7062) );
  NAND2_X1 U8199 ( .A1(n7063), .A2(n7062), .ZN(n8525) );
  XNOR2_X1 U8200 ( .A(n9211), .B(n7109), .ZN(n7064) );
  NAND2_X1 U8201 ( .A1(n9140), .A2(n7036), .ZN(n7065) );
  INV_X1 U8202 ( .A(n7064), .ZN(n7067) );
  INV_X1 U8203 ( .A(n7065), .ZN(n7066) );
  NAND2_X1 U8204 ( .A1(n7067), .A2(n7066), .ZN(n8559) );
  XNOR2_X1 U8205 ( .A(n9204), .B(n7103), .ZN(n7070) );
  NAND2_X1 U8206 ( .A1(n9110), .A2(n7036), .ZN(n7068) );
  XNOR2_X1 U8207 ( .A(n7070), .B(n7068), .ZN(n8857) );
  NAND2_X1 U8208 ( .A1(n8858), .A2(n8857), .ZN(n7072) );
  INV_X1 U8209 ( .A(n7068), .ZN(n7069) );
  NAND2_X1 U8210 ( .A1(n7070), .A2(n7069), .ZN(n7071) );
  XNOR2_X1 U8211 ( .A(n9199), .B(n7103), .ZN(n7075) );
  NAND2_X1 U8212 ( .A1(n9102), .A2(n7036), .ZN(n7073) );
  XNOR2_X1 U8213 ( .A(n7075), .B(n7073), .ZN(n8822) );
  INV_X1 U8214 ( .A(n7073), .ZN(n7074) );
  NAND2_X1 U8215 ( .A1(n7075), .A2(n7074), .ZN(n7076) );
  XNOR2_X1 U8216 ( .A(n9194), .B(n7109), .ZN(n7077) );
  NAND2_X1 U8217 ( .A1(n9089), .A2(n7036), .ZN(n7078) );
  NAND2_X1 U8218 ( .A1(n7077), .A2(n7078), .ZN(n7083) );
  INV_X1 U8219 ( .A(n7077), .ZN(n7080) );
  INV_X1 U8220 ( .A(n7078), .ZN(n7079) );
  NAND2_X1 U8221 ( .A1(n7080), .A2(n7079), .ZN(n7081) );
  NAND2_X1 U8222 ( .A1(n7083), .A2(n7081), .ZN(n8867) );
  XNOR2_X1 U8223 ( .A(n9054), .B(n7103), .ZN(n7085) );
  NAND2_X1 U8224 ( .A1(n9075), .A2(n7036), .ZN(n7084) );
  INV_X1 U8225 ( .A(n7085), .ZN(n7086) );
  NAND2_X1 U8226 ( .A1(n7087), .A2(n7086), .ZN(n7088) );
  XNOR2_X1 U8227 ( .A(n9182), .B(n7103), .ZN(n7089) );
  AND2_X1 U8228 ( .A1(n8886), .A2(n7036), .ZN(n8846) );
  INV_X1 U8229 ( .A(n7089), .ZN(n7090) );
  XNOR2_X1 U8230 ( .A(n9178), .B(n7109), .ZN(n7092) );
  NAND2_X1 U8231 ( .A1(n9040), .A2(n7036), .ZN(n7093) );
  NAND2_X1 U8232 ( .A1(n7092), .A2(n7093), .ZN(n7098) );
  INV_X1 U8233 ( .A(n7092), .ZN(n7095) );
  INV_X1 U8234 ( .A(n7093), .ZN(n7094) );
  NAND2_X1 U8235 ( .A1(n7095), .A2(n7094), .ZN(n7096) );
  NAND2_X1 U8236 ( .A1(n7098), .A2(n7096), .ZN(n8835) );
  INV_X1 U8237 ( .A(n8835), .ZN(n7097) );
  XNOR2_X1 U8238 ( .A(n9173), .B(n7109), .ZN(n7099) );
  NAND2_X1 U8239 ( .A1(n8991), .A2(n7036), .ZN(n7100) );
  XNOR2_X1 U8240 ( .A(n7099), .B(n7100), .ZN(n8874) );
  INV_X1 U8241 ( .A(n7099), .ZN(n7102) );
  INV_X1 U8242 ( .A(n7100), .ZN(n7101) );
  XNOR2_X1 U8243 ( .A(n9167), .B(n7103), .ZN(n7106) );
  NAND2_X1 U8244 ( .A1(n9000), .A2(n7036), .ZN(n7104) );
  XNOR2_X1 U8245 ( .A(n7106), .B(n7104), .ZN(n8814) );
  NAND2_X1 U8246 ( .A1(n8815), .A2(n8814), .ZN(n7108) );
  INV_X1 U8247 ( .A(n7104), .ZN(n7105) );
  NAND2_X1 U8248 ( .A1(n7106), .A2(n7105), .ZN(n7107) );
  NAND2_X1 U8249 ( .A1(n7108), .A2(n7107), .ZN(n7112) );
  NAND2_X1 U8250 ( .A1(n8992), .A2(n7036), .ZN(n7110) );
  MUX2_X1 U8251 ( .A(n8992), .B(n7110), .S(n7109), .Z(n7111) );
  XNOR2_X1 U8252 ( .A(n8206), .B(P2_B_REG_SCAN_IN), .ZN(n7113) );
  NAND2_X1 U8253 ( .A1(n7113), .A2(n8309), .ZN(n7114) );
  NAND2_X1 U8254 ( .A1(n7114), .A2(n7115), .ZN(n7212) );
  OR2_X1 U8255 ( .A1(n7212), .A2(P2_D_REG_0__SCAN_IN), .ZN(n7116) );
  INV_X1 U8256 ( .A(n7115), .ZN(n8447) );
  NAND2_X1 U8257 ( .A1(n8206), .A2(n8447), .ZN(n7216) );
  NAND2_X1 U8258 ( .A1(n7116), .A2(n7216), .ZN(n7693) );
  OR2_X1 U8259 ( .A1(n7212), .A2(P2_D_REG_1__SCAN_IN), .ZN(n7117) );
  NAND2_X1 U8260 ( .A1(n8447), .A2(n8309), .ZN(n7213) );
  NAND2_X1 U8261 ( .A1(n7117), .A2(n7213), .ZN(n7692) );
  NOR2_X1 U8262 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n7121) );
  NOR4_X1 U8263 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n7120) );
  NOR4_X1 U8264 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n7119) );
  NOR4_X1 U8265 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n7118) );
  NAND4_X1 U8266 ( .A1(n7121), .A2(n7120), .A3(n7119), .A4(n7118), .ZN(n7127)
         );
  NOR4_X1 U8267 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n7125) );
  NOR4_X1 U8268 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n7124) );
  NOR4_X1 U8269 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n7123) );
  NOR4_X1 U8270 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n7122) );
  NAND4_X1 U8271 ( .A1(n7125), .A2(n7124), .A3(n7123), .A4(n7122), .ZN(n7126)
         );
  NOR2_X1 U8272 ( .A1(n7127), .A2(n7126), .ZN(n7128) );
  NOR2_X1 U8273 ( .A1(n7212), .A2(n7128), .ZN(n7423) );
  OR3_X1 U8274 ( .A1(n7693), .A2(n7692), .A3(n7423), .ZN(n7132) );
  INV_X1 U8275 ( .A(n7429), .ZN(n7281) );
  NAND3_X1 U8276 ( .A1(n7700), .A2(n10998), .A3(n7281), .ZN(n7129) );
  NOR2_X2 U8277 ( .A1(n7132), .A2(n7129), .ZN(n10727) );
  AND3_X1 U8278 ( .A1(n7811), .A2(n10812), .A3(n8039), .ZN(n10901) );
  NAND2_X1 U8279 ( .A1(n10901), .A2(n7825), .ZN(n7698) );
  NAND2_X1 U8280 ( .A1(n7132), .A2(n7698), .ZN(n7138) );
  AND2_X1 U8281 ( .A1(n7138), .A2(n7700), .ZN(n8723) );
  AOI21_X1 U8282 ( .B1(n7130), .B2(n10727), .A(n10733), .ZN(n7145) );
  NOR2_X1 U8283 ( .A1(n7132), .A2(n7131), .ZN(n8840) );
  AND2_X1 U8284 ( .A1(n6364), .A2(n7429), .ZN(n9139) );
  INV_X1 U8285 ( .A(n9139), .ZN(n8415) );
  INV_X1 U8286 ( .A(n8415), .ZN(n8837) );
  NAND2_X1 U8287 ( .A1(n8840), .A2(n8837), .ZN(n10736) );
  OAI22_X1 U8288 ( .A1(n8885), .A2(n10736), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7133), .ZN(n7134) );
  AOI21_X1 U8289 ( .B1(n10731), .B2(n9000), .A(n7134), .ZN(n7135) );
  INV_X1 U8290 ( .A(n7135), .ZN(n7142) );
  INV_X1 U8291 ( .A(n8972), .ZN(n7140) );
  AND2_X1 U8292 ( .A1(n7429), .A2(n7427), .ZN(n7421) );
  NOR2_X1 U8293 ( .A1(n7136), .A2(n7421), .ZN(n7137) );
  NAND2_X1 U8294 ( .A1(n7138), .A2(n7137), .ZN(n7139) );
  NAND2_X1 U8295 ( .A1(n7139), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10742) );
  OAI211_X1 U8296 ( .C1(n7145), .C2(n5342), .A(n7144), .B(n7143), .ZN(P2_U3222) );
  AND2_X1 U8297 ( .A1(n7147), .A2(n7146), .ZN(n7148) );
  NOR2_X1 U8298 ( .A1(n9800), .A2(n10344), .ZN(n7151) );
  OAI22_X1 U8299 ( .A1(n9798), .A2(n8790), .B1(n9799), .B2(n10307), .ZN(n7150)
         );
  AOI211_X1 U8300 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3084), .A(n7151), 
        .B(n7150), .ZN(n7152) );
  INV_X1 U8301 ( .A(n10488), .ZN(n10306) );
  NAND3_X1 U8302 ( .A1(n7153), .A2(n7152), .A3(n5550), .ZN(P1_U3212) );
  NAND2_X1 U8303 ( .A1(n7154), .A2(n8135), .ZN(n7251) );
  NAND2_X1 U8304 ( .A1(n6418), .A2(n7155), .ZN(n7156) );
  NAND2_X1 U8305 ( .A1(n7156), .A2(n8135), .ZN(n7157) );
  NAND2_X1 U8306 ( .A1(n6503), .A2(n7157), .ZN(n7158) );
  NAND2_X1 U8307 ( .A1(n7158), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U8308 ( .A(n10727), .ZN(n8882) );
  INV_X1 U8309 ( .A(n7159), .ZN(n7169) );
  AOI211_X1 U8310 ( .C1(n7161), .C2(n7160), .A(n8882), .B(n7169), .ZN(n7166)
         );
  AND2_X1 U8311 ( .A1(n10733), .A2(n8257), .ZN(n7165) );
  NOR2_X1 U8312 ( .A1(n10742), .A2(n8248), .ZN(n7164) );
  NAND2_X1 U8313 ( .A1(n10731), .A2(n8894), .ZN(n7162) );
  NAND2_X1 U8314 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7533) );
  OAI211_X1 U8315 ( .C1(n8320), .C2(n10736), .A(n7162), .B(n7533), .ZN(n7163)
         );
  OR4_X1 U8316 ( .A1(n7166), .A2(n7165), .A3(n7164), .A4(n7163), .ZN(P2_U3219)
         );
  AND2_X1 U8317 ( .A1(n10727), .A2(n7036), .ZN(n8845) );
  NAND3_X1 U8318 ( .A1(n7167), .A2(n8845), .A3(n8893), .ZN(n7171) );
  OAI21_X1 U8319 ( .B1(n7169), .B2(n7168), .A(n10727), .ZN(n7170) );
  INV_X1 U8320 ( .A(n8729), .ZN(n8298) );
  AOI21_X1 U8321 ( .B1(n7171), .B2(n7170), .A(n8298), .ZN(n7178) );
  AND2_X1 U8322 ( .A1(n10905), .A2(n10733), .ZN(n7177) );
  NOR2_X1 U8323 ( .A1(n10742), .A2(n8283), .ZN(n7176) );
  NAND2_X1 U8324 ( .A1(n10731), .A2(n8893), .ZN(n7174) );
  NOR2_X1 U8325 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7172), .ZN(n7554) );
  INV_X1 U8326 ( .A(n7554), .ZN(n7173) );
  OAI211_X1 U8327 ( .C1(n8703), .C2(n10736), .A(n7174), .B(n7173), .ZN(n7175)
         );
  OR4_X1 U8328 ( .A1(n7178), .A2(n7177), .A3(n7176), .A4(n7175), .ZN(P2_U3238)
         );
  NAND2_X1 U8329 ( .A1(n7179), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7215) );
  OR2_X2 U8330 ( .A1(n7282), .A2(n7215), .ZN(n8902) );
  INV_X1 U8331 ( .A(n8902), .ZN(P2_U3966) );
  AND2_X1 U8332 ( .A1(n5034), .A2(P1_U3084), .ZN(n8134) );
  INV_X2 U8333 ( .A(n8134), .ZN(n10596) );
  OAI222_X1 U8334 ( .A1(n7259), .A2(P1_U3084), .B1(n10596), .B2(n7194), .C1(
        n7180), .C2(n8813), .ZN(P1_U3352) );
  OAI222_X1 U8335 ( .A1(n8813), .A2(n7181), .B1(n10596), .B2(n7183), .C1(n7244), .C2(P1_U3084), .ZN(P1_U3351) );
  AND2_X1 U8336 ( .A1(n5034), .A2(P2_U3152), .ZN(n7581) );
  INV_X2 U8337 ( .A(n7581), .ZN(n9696) );
  NAND2_X1 U8338 ( .A1(n7182), .A2(P2_U3152), .ZN(n9699) );
  OAI222_X1 U8339 ( .A1(n9696), .A2(n7184), .B1(n9699), .B2(n7183), .C1(
        P2_U3152), .C2(n7332), .ZN(P2_U3356) );
  OAI222_X1 U8340 ( .A1(n8813), .A2(n7185), .B1(n10596), .B2(n7186), .C1(n7258), .C2(P1_U3084), .ZN(P1_U3350) );
  OAI222_X1 U8341 ( .A1(n9696), .A2(n7187), .B1(n9699), .B2(n7186), .C1(
        P2_U3152), .C2(n7348), .ZN(P2_U3355) );
  OAI222_X1 U8342 ( .A1(n9696), .A2(n5652), .B1(n9699), .B2(n7189), .C1(
        P2_U3152), .C2(n7416), .ZN(P2_U3354) );
  OAI222_X1 U8343 ( .A1(n7190), .A2(P1_U3084), .B1(n10596), .B2(n7189), .C1(
        n7188), .C2(n8813), .ZN(P1_U3349) );
  OAI222_X1 U8344 ( .A1(n7257), .A2(P1_U3084), .B1(n10596), .B2(n7192), .C1(
        n7191), .C2(n8813), .ZN(P1_U3348) );
  OAI222_X1 U8345 ( .A1(n9696), .A2(n7193), .B1(n9699), .B2(n7192), .C1(
        P2_U3152), .C2(n7446), .ZN(P2_U3353) );
  INV_X1 U8346 ( .A(n9699), .ZN(n8137) );
  INV_X1 U8347 ( .A(n8137), .ZN(n8593) );
  OAI222_X1 U8348 ( .A1(n9696), .A2(n7195), .B1(n8593), .B2(n7194), .C1(
        P2_U3152), .C2(n7314), .ZN(P2_U3357) );
  OAI222_X1 U8349 ( .A1(n9696), .A2(n7197), .B1(n9699), .B2(n7199), .C1(
        P2_U3152), .C2(n7196), .ZN(P2_U3352) );
  OAI222_X1 U8350 ( .A1(n7200), .A2(P1_U3084), .B1(n10596), .B2(n7199), .C1(
        n7198), .C2(n8813), .ZN(P1_U3347) );
  OAI222_X1 U8351 ( .A1(n7276), .A2(P1_U3084), .B1(n10596), .B2(n7202), .C1(
        n7201), .C2(n8813), .ZN(P1_U3346) );
  OAI222_X1 U8352 ( .A1(n9696), .A2(n7203), .B1(n9699), .B2(n7202), .C1(
        P2_U3152), .C2(n7445), .ZN(P2_U3351) );
  INV_X1 U8353 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7204) );
  INV_X1 U8354 ( .A(n7476), .ZN(n7469) );
  OAI222_X1 U8355 ( .A1(n9696), .A2(n7204), .B1(n9699), .B2(n7206), .C1(
        P2_U3152), .C2(n7469), .ZN(P2_U3350) );
  OAI222_X1 U8356 ( .A1(n7207), .A2(P1_U3084), .B1(n10596), .B2(n7206), .C1(
        n7205), .C2(n8813), .ZN(P1_U3345) );
  INV_X1 U8357 ( .A(n7208), .ZN(n7210) );
  INV_X1 U8358 ( .A(n8813), .ZN(n10594) );
  AOI22_X1 U8359 ( .A1(n10177), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10594), .ZN(n7209) );
  OAI21_X1 U8360 ( .B1(n7210), .B2(n10596), .A(n7209), .ZN(P1_U3344) );
  INV_X1 U8361 ( .A(n7537), .ZN(n7529) );
  OAI222_X1 U8362 ( .A1(n9696), .A2(n7211), .B1(n8593), .B2(n7210), .C1(
        P2_U3152), .C2(n7529), .ZN(P2_U3349) );
  NAND2_X1 U8363 ( .A1(n7700), .A2(n7212), .ZN(n10602) );
  INV_X1 U8364 ( .A(n10602), .ZN(n7217) );
  OAI22_X1 U8365 ( .A1(n7217), .A2(P2_D_REG_1__SCAN_IN), .B1(n7213), .B2(n7215), .ZN(n7214) );
  INV_X1 U8366 ( .A(n7214), .ZN(P2_U3438) );
  OAI22_X1 U8367 ( .A1(n7217), .A2(P2_D_REG_0__SCAN_IN), .B1(n7216), .B2(n7215), .ZN(n7218) );
  INV_X1 U8368 ( .A(n7218), .ZN(P2_U3437) );
  NAND2_X1 U8369 ( .A1(n7700), .A2(n7429), .ZN(n7219) );
  NAND2_X1 U8370 ( .A1(n7219), .A2(n7286), .ZN(n7222) );
  OR2_X1 U8371 ( .A1(n7700), .A2(n7220), .ZN(n7221) );
  NAND2_X1 U8372 ( .A1(n7222), .A2(n7221), .ZN(n8929) );
  INV_X1 U8373 ( .A(n8929), .ZN(n8953) );
  NOR2_X1 U8374 ( .A1(n8953), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8375 ( .A(n7223), .ZN(n7226) );
  AOI22_X1 U8376 ( .A1(n7556), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n7581), .ZN(n7224) );
  OAI21_X1 U8377 ( .B1(n7226), .B2(n9699), .A(n7224), .ZN(P2_U3348) );
  NAND2_X1 U8378 ( .A1(n8902), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7225) );
  OAI21_X1 U8379 ( .B1(n8665), .B2(n8902), .A(n7225), .ZN(P2_U3582) );
  INV_X1 U8380 ( .A(n10663), .ZN(n7671) );
  OAI222_X1 U8381 ( .A1(P1_U3084), .A2(n7671), .B1(n10596), .B2(n7226), .C1(
        n9384), .C2(n8813), .ZN(P1_U3343) );
  INV_X1 U8382 ( .A(n7227), .ZN(n7233) );
  AOI22_X1 U8383 ( .A1(n8179), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10594), .ZN(n7228) );
  OAI21_X1 U8384 ( .B1(n7233), .B2(n10596), .A(n7228), .ZN(P1_U3340) );
  INV_X1 U8385 ( .A(n7229), .ZN(n7231) );
  INV_X1 U8386 ( .A(n7652), .ZN(n7661) );
  OAI222_X1 U8387 ( .A1(n8593), .A2(n7231), .B1(n7661), .B2(P2_U3152), .C1(
        n5300), .C2(n9696), .ZN(P2_U3347) );
  INV_X1 U8388 ( .A(n7683), .ZN(n10694) );
  INV_X1 U8389 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7230) );
  OAI222_X1 U8390 ( .A1(P1_U3084), .A2(n10694), .B1(n10596), .B2(n7231), .C1(
        n7230), .C2(n8813), .ZN(P1_U3342) );
  INV_X1 U8391 ( .A(n7930), .ZN(n7925) );
  OAI222_X1 U8392 ( .A1(n8593), .A2(n7233), .B1(n7925), .B2(P2_U3152), .C1(
        n7232), .C2(n9696), .ZN(P2_U3345) );
  INV_X1 U8393 ( .A(n7234), .ZN(n7238) );
  AOI22_X1 U8394 ( .A1(n7869), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10594), .ZN(n7235) );
  OAI21_X1 U8395 ( .B1(n7238), .B2(n10596), .A(n7235), .ZN(P1_U3341) );
  INV_X1 U8396 ( .A(n10189), .ZN(n10182) );
  INV_X1 U8397 ( .A(n7236), .ZN(n7240) );
  INV_X1 U8398 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7237) );
  OAI222_X1 U8399 ( .A1(P1_U3084), .A2(n10182), .B1(n10596), .B2(n7240), .C1(
        n7237), .C2(n8813), .ZN(P1_U3339) );
  INV_X1 U8400 ( .A(n7768), .ZN(n7764) );
  OAI222_X1 U8401 ( .A1(n9696), .A2(n7239), .B1(n9699), .B2(n7238), .C1(
        P2_U3152), .C2(n7764), .ZN(P2_U3346) );
  INV_X1 U8402 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7241) );
  INV_X1 U8403 ( .A(n8215), .ZN(n8221) );
  OAI222_X1 U8404 ( .A1(n9696), .A2(n7241), .B1(P2_U3152), .B2(n8221), .C1(
        n7240), .C2(n9699), .ZN(P2_U3344) );
  AOI21_X1 U8405 ( .B1(n10033), .B2(n8135), .A(P1_U3084), .ZN(n7242) );
  NAND2_X1 U8406 ( .A1(n7251), .A2(n7242), .ZN(n7256) );
  OR2_X1 U8407 ( .A1(n7243), .A2(n7256), .ZN(n10643) );
  INV_X1 U8408 ( .A(n8508), .ZN(n10640) );
  NOR2_X2 U8409 ( .A1(n10643), .A2(n10640), .ZN(n10689) );
  AOI22_X1 U8410 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n7257), .B1(n7275), .B2(
        n6532), .ZN(n7250) );
  INV_X1 U8411 ( .A(n7259), .ZN(n10111) );
  INV_X1 U8412 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7392) );
  INV_X1 U8413 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U8414 ( .A1(P1_REG1_REG_1__SCAN_IN), .A2(n7259), .B1(n10111), .B2(
        n10702), .ZN(n10113) );
  NOR3_X1 U8415 ( .A1(n6461), .A2(n7392), .A3(n10113), .ZN(n10112) );
  AOI21_X1 U8416 ( .B1(n10111), .B2(P1_REG1_REG_1__SCAN_IN), .A(n10112), .ZN(
        n10133) );
  AOI22_X1 U8417 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(n7244), .B1(n10130), .B2(
        n10710), .ZN(n10132) );
  NOR2_X1 U8418 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  AND2_X1 U8419 ( .A1(n10130), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7245) );
  OR2_X1 U8420 ( .A1(n10131), .A2(n7245), .ZN(n10147) );
  XNOR2_X1 U8421 ( .A(n7258), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n10148) );
  NAND2_X1 U8422 ( .A1(n10147), .A2(n10148), .ZN(n10146) );
  OAI21_X1 U8423 ( .B1(n7258), .B2(n7246), .A(n10146), .ZN(n10157) );
  NOR2_X1 U8424 ( .A1(n10155), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7247) );
  AOI21_X1 U8425 ( .B1(n10155), .B2(P1_REG1_REG_4__SCAN_IN), .A(n7247), .ZN(
        n10159) );
  INV_X1 U8426 ( .A(n10159), .ZN(n7248) );
  OR2_X1 U8427 ( .A1(n10157), .A2(n7248), .ZN(n10158) );
  OAI21_X1 U8428 ( .B1(n10155), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10158), .ZN(
        n7249) );
  NOR2_X1 U8429 ( .A1(n7250), .A2(n7249), .ZN(n7269) );
  AOI21_X1 U8430 ( .B1(n7250), .B2(n7249), .A(n7269), .ZN(n7255) );
  INV_X1 U8431 ( .A(n7251), .ZN(n7252) );
  OR2_X1 U8432 ( .A1(P1_U3083), .A2(n7252), .ZN(n10679) );
  INV_X1 U8433 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7253) );
  NAND2_X1 U8434 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7637) );
  OAI21_X1 U8435 ( .B1(n10679), .B2(n7253), .A(n7637), .ZN(n7254) );
  AOI21_X1 U8436 ( .B1(n10689), .B2(n7255), .A(n7254), .ZN(n7268) );
  NOR2_X1 U8437 ( .A1(n7256), .A2(n8508), .ZN(n10675) );
  NAND2_X1 U8438 ( .A1(n10675), .A2(n7264), .ZN(n10657) );
  INV_X1 U8439 ( .A(n10657), .ZN(n10690) );
  AOI22_X1 U8440 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n7275), .B1(n7257), .B2(
        n6530), .ZN(n7263) );
  INV_X1 U8441 ( .A(n7258), .ZN(n10144) );
  XOR2_X1 U8442 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7258), .Z(n10141) );
  NAND2_X1 U8443 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10121) );
  INV_X1 U8444 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7979) );
  NOR2_X1 U8445 ( .A1(n10121), .A2(n10109), .ZN(n10108) );
  AOI21_X1 U8446 ( .B1(n10111), .B2(P1_REG2_REG_1__SCAN_IN), .A(n10108), .ZN(
        n10128) );
  NAND2_X1 U8447 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n10130), .ZN(n7260) );
  OAI21_X1 U8448 ( .B1(n10130), .B2(P1_REG2_REG_2__SCAN_IN), .A(n7260), .ZN(
        n10127) );
  NOR2_X1 U8449 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  AOI21_X1 U8450 ( .B1(n10130), .B2(P1_REG2_REG_2__SCAN_IN), .A(n10126), .ZN(
        n10142) );
  NOR2_X1 U8451 ( .A1(n10141), .A2(n10142), .ZN(n10140) );
  AOI21_X1 U8452 ( .B1(n10144), .B2(P1_REG2_REG_3__SCAN_IN), .A(n10140), .ZN(
        n10154) );
  NOR2_X1 U8453 ( .A1(n10155), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7261) );
  AOI21_X1 U8454 ( .B1(n10155), .B2(P1_REG2_REG_4__SCAN_IN), .A(n7261), .ZN(
        n10153) );
  NAND2_X1 U8455 ( .A1(n10154), .A2(n10153), .ZN(n10152) );
  OAI21_X1 U8456 ( .B1(n10155), .B2(P1_REG2_REG_4__SCAN_IN), .A(n10152), .ZN(
        n7262) );
  NAND2_X1 U8457 ( .A1(n7263), .A2(n7262), .ZN(n7274) );
  OAI21_X1 U8458 ( .B1(n7263), .B2(n7262), .A(n7274), .ZN(n7266) );
  INV_X1 U8459 ( .A(n10675), .ZN(n7265) );
  NOR2_X2 U8460 ( .A1(n7265), .A2(n7264), .ZN(n10672) );
  AOI22_X1 U8461 ( .A1(n10690), .A2(n7266), .B1(n10672), .B2(n7275), .ZN(n7267) );
  NAND2_X1 U8462 ( .A1(n7268), .A2(n7267), .ZN(P1_U3246) );
  AOI21_X1 U8463 ( .B1(n7275), .B2(P1_REG1_REG_5__SCAN_IN), .A(n7269), .ZN(
        n10653) );
  NAND2_X1 U8464 ( .A1(n10650), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7270) );
  OAI21_X1 U8465 ( .B1(n10650), .B2(P1_REG1_REG_6__SCAN_IN), .A(n7270), .ZN(
        n10652) );
  NOR2_X1 U8466 ( .A1(n10653), .A2(n10652), .ZN(n10651) );
  AOI21_X1 U8467 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10650), .A(n10651), .ZN(
        n7354) );
  XNOR2_X1 U8468 ( .A(n7276), .B(n7271), .ZN(n7355) );
  XNOR2_X1 U8469 ( .A(n7354), .B(n7355), .ZN(n7280) );
  INV_X1 U8470 ( .A(n10689), .ZN(n10264) );
  INV_X1 U8471 ( .A(n10679), .ZN(n10667) );
  INV_X1 U8472 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7272) );
  NOR2_X1 U8473 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7272), .ZN(n7815) );
  AOI21_X1 U8474 ( .B1(n10667), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7815), .ZN(
        n7279) );
  XNOR2_X1 U8475 ( .A(n7276), .B(n8074), .ZN(n7363) );
  NAND2_X1 U8476 ( .A1(n10650), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7273) );
  OAI21_X1 U8477 ( .B1(n10650), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7273), .ZN(
        n10646) );
  OAI21_X1 U8478 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7275), .A(n7274), .ZN(
        n10647) );
  XNOR2_X1 U8479 ( .A(n7363), .B(n7362), .ZN(n7277) );
  INV_X1 U8480 ( .A(n7276), .ZN(n7361) );
  AOI22_X1 U8481 ( .A1(n10690), .A2(n7277), .B1(n10672), .B2(n7361), .ZN(n7278) );
  OAI211_X1 U8482 ( .C1(n7280), .C2(n10264), .A(n7279), .B(n7278), .ZN(
        P1_U3248) );
  NAND2_X1 U8483 ( .A1(n7700), .A2(n7281), .ZN(n7285) );
  OAI21_X1 U8484 ( .B1(n7282), .B2(P2_U3152), .A(n8139), .ZN(n7283) );
  INV_X1 U8485 ( .A(n7283), .ZN(n7284) );
  NAND2_X1 U8486 ( .A1(n7285), .A2(n7284), .ZN(n7287) );
  NAND2_X1 U8487 ( .A1(n7287), .A2(n7286), .ZN(n7290) );
  NAND2_X1 U8488 ( .A1(n7290), .A2(n8902), .ZN(n7296) );
  AND2_X1 U8489 ( .A1(n6364), .A2(n7296), .ZN(n8959) );
  INV_X1 U8490 ( .A(n8959), .ZN(n7563) );
  NAND2_X1 U8491 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n7292) );
  MUX2_X1 U8492 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n5595), .S(n7314), .Z(n7291)
         );
  INV_X1 U8493 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7288) );
  NOR3_X1 U8494 ( .A1(n7291), .A2(n7289), .A3(n7288), .ZN(n7309) );
  INV_X1 U8495 ( .A(n6363), .ZN(n7295) );
  OR2_X1 U8496 ( .A1(n7290), .A2(n7295), .ZN(n8957) );
  AOI211_X1 U8497 ( .C1(n7292), .C2(n7291), .A(n7309), .B(n8957), .ZN(n7294)
         );
  INV_X1 U8498 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8340) );
  OAI22_X1 U8499 ( .A1(n8929), .A2(n8340), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7704), .ZN(n7293) );
  NOR2_X1 U8500 ( .A1(n7294), .A2(n7293), .ZN(n7301) );
  INV_X1 U8501 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7707) );
  AND2_X1 U8502 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7298) );
  AND2_X1 U8503 ( .A1(n7296), .A2(n7295), .ZN(n7394) );
  NAND2_X1 U8504 ( .A1(n7394), .A2(n7297), .ZN(n8961) );
  INV_X1 U8505 ( .A(n8961), .ZN(n7936) );
  OAI211_X1 U8506 ( .C1(n7299), .C2(n7298), .A(n7936), .B(n7313), .ZN(n7300)
         );
  OAI211_X1 U8507 ( .C1(n7563), .C2(n7314), .A(n7301), .B(n7300), .ZN(P2_U3246) );
  NOR2_X1 U8508 ( .A1(n7756), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7312) );
  INV_X1 U8509 ( .A(n7309), .ZN(n7304) );
  INV_X1 U8510 ( .A(n7314), .ZN(n7302) );
  NAND2_X1 U8511 ( .A1(n7302), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7305) );
  MUX2_X1 U8512 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7306), .S(n7332), .Z(n7303)
         );
  AOI21_X1 U8513 ( .B1(n7304), .B2(n7305), .A(n7303), .ZN(n7326) );
  INV_X1 U8514 ( .A(n7305), .ZN(n7308) );
  MUX2_X1 U8515 ( .A(n7306), .B(P2_REG1_REG_2__SCAN_IN), .S(n7332), .Z(n7307)
         );
  NOR3_X1 U8516 ( .A1(n7309), .A2(n7308), .A3(n7307), .ZN(n7310) );
  NOR3_X1 U8517 ( .A1(n8957), .A2(n7326), .A3(n7310), .ZN(n7311) );
  AOI211_X1 U8518 ( .C1(n8953), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n7312), .B(
        n7311), .ZN(n7318) );
  XNOR2_X1 U8519 ( .A(n7332), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7316) );
  NAND2_X1 U8520 ( .A1(n7315), .A2(n7316), .ZN(n7330) );
  OAI211_X1 U8521 ( .C1(n7316), .C2(n7315), .A(n7936), .B(n7330), .ZN(n7317)
         );
  OAI211_X1 U8522 ( .C1(n7563), .C2(n7332), .A(n7318), .B(n7317), .ZN(P2_U3247) );
  INV_X1 U8523 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7735) );
  NOR2_X1 U8524 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7735), .ZN(n7329) );
  INV_X1 U8525 ( .A(n7326), .ZN(n7321) );
  INV_X1 U8526 ( .A(n7332), .ZN(n7319) );
  NAND2_X1 U8527 ( .A1(n7319), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7322) );
  MUX2_X1 U8528 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7323), .S(n7348), .Z(n7320)
         );
  AOI21_X1 U8529 ( .B1(n7321), .B2(n7322), .A(n7320), .ZN(n7343) );
  INV_X1 U8530 ( .A(n7322), .ZN(n7325) );
  MUX2_X1 U8531 ( .A(n7323), .B(P2_REG1_REG_3__SCAN_IN), .S(n7348), .Z(n7324)
         );
  NOR3_X1 U8532 ( .A1(n7326), .A2(n7325), .A3(n7324), .ZN(n7327) );
  NOR3_X1 U8533 ( .A1(n8957), .A2(n7343), .A3(n7327), .ZN(n7328) );
  AOI211_X1 U8534 ( .C1(n8953), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n7329), .B(
        n7328), .ZN(n7336) );
  XNOR2_X1 U8535 ( .A(n7348), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n7334) );
  INV_X1 U8536 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7331) );
  OAI21_X1 U8537 ( .B1(n7332), .B2(n7331), .A(n7330), .ZN(n7333) );
  NAND2_X1 U8538 ( .A1(n7333), .A2(n7334), .ZN(n7347) );
  OAI211_X1 U8539 ( .C1(n7334), .C2(n7333), .A(n7936), .B(n7347), .ZN(n7335)
         );
  OAI211_X1 U8540 ( .C1(n7563), .C2(n7348), .A(n7336), .B(n7335), .ZN(P2_U3248) );
  NAND2_X1 U8541 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7596) );
  INV_X1 U8542 ( .A(n7596), .ZN(n7346) );
  INV_X1 U8543 ( .A(n7343), .ZN(n7339) );
  INV_X1 U8544 ( .A(n7348), .ZN(n7337) );
  NAND2_X1 U8545 ( .A1(n7337), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7340) );
  MUX2_X1 U8546 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7407), .S(n7416), .Z(n7338)
         );
  AOI21_X1 U8547 ( .B1(n7339), .B2(n7340), .A(n7338), .ZN(n7405) );
  INV_X1 U8548 ( .A(n7340), .ZN(n7342) );
  MUX2_X1 U8549 ( .A(n7407), .B(P2_REG1_REG_4__SCAN_IN), .S(n7416), .Z(n7341)
         );
  NOR3_X1 U8550 ( .A1(n7343), .A2(n7342), .A3(n7341), .ZN(n7344) );
  NOR3_X1 U8551 ( .A1(n8957), .A2(n7405), .A3(n7344), .ZN(n7345) );
  AOI211_X1 U8552 ( .C1(n8953), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7346), .B(
        n7345), .ZN(n7353) );
  XNOR2_X1 U8553 ( .A(n7416), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7351) );
  INV_X1 U8554 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7349) );
  OAI21_X1 U8555 ( .B1(n7349), .B2(n7348), .A(n7347), .ZN(n7350) );
  NAND2_X1 U8556 ( .A1(n7350), .A2(n7351), .ZN(n7414) );
  OAI211_X1 U8557 ( .C1(n7351), .C2(n7350), .A(n7936), .B(n7414), .ZN(n7352)
         );
  OAI211_X1 U8558 ( .C1(n7563), .C2(n7416), .A(n7353), .B(n7352), .ZN(P2_U3249) );
  INV_X1 U8559 ( .A(n7354), .ZN(n7356) );
  OAI22_X1 U8560 ( .A1(n7356), .A2(n7355), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n7361), .ZN(n7359) );
  NOR2_X1 U8561 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7681), .ZN(n7357) );
  AOI21_X1 U8562 ( .B1(n7681), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7357), .ZN(
        n7358) );
  NAND2_X1 U8563 ( .A1(n7358), .A2(n7359), .ZN(n7673) );
  OAI21_X1 U8564 ( .B1(n7359), .B2(n7358), .A(n7673), .ZN(n7371) );
  INV_X1 U8565 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7369) );
  NOR2_X1 U8566 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7681), .ZN(n7360) );
  AOI21_X1 U8567 ( .B1(n7681), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7360), .ZN(
        n7365) );
  NAND2_X1 U8568 ( .A1(n7365), .A2(n7364), .ZN(n7680) );
  OAI21_X1 U8569 ( .B1(n7365), .B2(n7364), .A(n7680), .ZN(n7366) );
  AOI22_X1 U8570 ( .A1(n10690), .A2(n7366), .B1(n10672), .B2(n7681), .ZN(n7368) );
  AND2_X1 U8571 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8024) );
  INV_X1 U8572 ( .A(n8024), .ZN(n7367) );
  OAI211_X1 U8573 ( .C1(n7369), .C2(n10679), .A(n7368), .B(n7367), .ZN(n7370)
         );
  AOI21_X1 U8574 ( .B1(n7371), .B2(n10689), .A(n7370), .ZN(n7372) );
  INV_X1 U8575 ( .A(n7372), .ZN(P1_U3249) );
  INV_X1 U8576 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7374) );
  INV_X1 U8577 ( .A(n7373), .ZN(n7376) );
  INV_X1 U8578 ( .A(n8394), .ZN(n8401) );
  OAI222_X1 U8579 ( .A1(n9696), .A2(n7374), .B1(n8593), .B2(n7376), .C1(
        P2_U3152), .C2(n8401), .ZN(P2_U3343) );
  INV_X1 U8580 ( .A(n10205), .ZN(n10194) );
  INV_X1 U8581 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7375) );
  OAI222_X1 U8582 ( .A1(n10194), .A2(P1_U3084), .B1(n10596), .B2(n7376), .C1(
        n7375), .C2(n8813), .ZN(P1_U3338) );
  AND2_X1 U8583 ( .A1(n7377), .A2(n7387), .ZN(n7826) );
  OR2_X1 U8584 ( .A1(n10990), .A2(n10260), .ZN(n7828) );
  AND3_X1 U8585 ( .A1(n7379), .A2(n7378), .A3(n7828), .ZN(n7389) );
  AND2_X2 U8586 ( .A1(n7826), .A2(n7389), .ZN(n11040) );
  INV_X1 U8587 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7385) );
  INV_X1 U8588 ( .A(n8014), .ZN(n9835) );
  INV_X1 U8589 ( .A(n6469), .ZN(n7973) );
  INV_X1 U8590 ( .A(n7970), .ZN(n7380) );
  AOI21_X1 U8591 ( .B1(n7973), .B2(n9835), .A(n7380), .ZN(n10038) );
  NOR2_X1 U8592 ( .A1(n10033), .A2(n7381), .ZN(n7382) );
  AOI22_X1 U8593 ( .A1(n10038), .A2(n7382), .B1(n10769), .B2(n10107), .ZN(
        n8017) );
  OAI21_X1 U8594 ( .B1(n9835), .B2(n7383), .A(n8017), .ZN(n7390) );
  NAND2_X1 U8595 ( .A1(n7390), .A2(n11040), .ZN(n7384) );
  OAI21_X1 U8596 ( .B1(n11040), .B2(n7385), .A(n7384), .ZN(P1_U3454) );
  NOR2_X1 U8597 ( .A1(n7387), .A2(n7386), .ZN(n7388) );
  AND2_X2 U8598 ( .A1(n7389), .A2(n7388), .ZN(n11036) );
  NAND2_X1 U8599 ( .A1(n7390), .A2(n11036), .ZN(n7391) );
  OAI21_X1 U8600 ( .B1(n11036), .B2(n7392), .A(n7391), .ZN(P1_U3523) );
  INV_X1 U8601 ( .A(n8957), .ZN(n8907) );
  AOI22_X1 U8602 ( .A1(n7936), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n8907), .ZN(n7398) );
  INV_X1 U8603 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U8604 ( .A1(n7394), .A2(n7393), .ZN(n7395) );
  OAI211_X1 U8605 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n8957), .A(n7563), .B(
        n7395), .ZN(n7396) );
  INV_X1 U8606 ( .A(n7396), .ZN(n7397) );
  MUX2_X1 U8607 ( .A(n7398), .B(n7397), .S(P2_IR_REG_0__SCAN_IN), .Z(n7400) );
  NAND2_X1 U8608 ( .A1(n8953), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n7399) );
  OAI211_X1 U8609 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7779), .A(n7400), .B(n7399), .ZN(P2_U3245) );
  INV_X1 U8610 ( .A(n7401), .ZN(n7404) );
  AOI22_X1 U8611 ( .A1(n8914), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n7581), .ZN(n7402) );
  OAI21_X1 U8612 ( .B1(n7404), .B2(n9699), .A(n7402), .ZN(P2_U3342) );
  AOI22_X1 U8613 ( .A1(n10222), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10594), .ZN(n7403) );
  OAI21_X1 U8614 ( .B1(n7404), .B2(n10596), .A(n7403), .ZN(P1_U3337) );
  NOR2_X1 U8615 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9543), .ZN(n7413) );
  INV_X1 U8616 ( .A(n7405), .ZN(n7406) );
  OAI21_X1 U8617 ( .B1(n7416), .B2(n7407), .A(n7406), .ZN(n7410) );
  MUX2_X1 U8618 ( .A(n7408), .B(P2_REG1_REG_5__SCAN_IN), .S(n7446), .Z(n7409)
         );
  NAND2_X1 U8619 ( .A1(n7409), .A2(n7410), .ZN(n7437) );
  OAI211_X1 U8620 ( .C1(n7410), .C2(n7409), .A(n8907), .B(n7437), .ZN(n7411)
         );
  INV_X1 U8621 ( .A(n7411), .ZN(n7412) );
  AOI211_X1 U8622 ( .C1(n8953), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7413), .B(
        n7412), .ZN(n7420) );
  MUX2_X1 U8623 ( .A(n5659), .B(P2_REG2_REG_5__SCAN_IN), .S(n7446), .Z(n7418)
         );
  INV_X1 U8624 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7415) );
  OAI21_X1 U8625 ( .B1(n7416), .B2(n7415), .A(n7414), .ZN(n7417) );
  OAI211_X1 U8626 ( .C1(n7418), .C2(n7417), .A(n7936), .B(n7447), .ZN(n7419)
         );
  OAI211_X1 U8627 ( .C1(n7563), .C2(n7446), .A(n7420), .B(n7419), .ZN(P2_U3250) );
  INV_X1 U8628 ( .A(n7421), .ZN(n7516) );
  NAND2_X1 U8629 ( .A1(n7700), .A2(n7516), .ZN(n7422) );
  NAND2_X1 U8630 ( .A1(n7692), .A2(n7698), .ZN(n7424) );
  NOR2_X1 U8631 ( .A1(n7695), .A2(n7424), .ZN(n7621) );
  INV_X1 U8632 ( .A(n7693), .ZN(n7425) );
  AND2_X2 U8633 ( .A1(n7621), .A2(n7425), .ZN(n11007) );
  AND2_X1 U8634 ( .A1(n7427), .A2(n7426), .ZN(n7430) );
  OR3_X1 U8635 ( .A1(n7430), .A2(n7429), .A3(n7428), .ZN(n8247) );
  INV_X1 U8636 ( .A(n10901), .ZN(n7431) );
  NAND2_X1 U8637 ( .A1(n8247), .A2(n7431), .ZN(n11004) );
  AND2_X1 U8638 ( .A1(n7433), .A2(n7432), .ZN(n9070) );
  OAI21_X1 U8639 ( .B1(n11004), .B2(n10798), .A(n7781), .ZN(n7434) );
  NAND2_X1 U8640 ( .A1(n8901), .A2(n8837), .ZN(n7778) );
  OAI211_X1 U8641 ( .C1(n7513), .C2(n7702), .A(n7434), .B(n7778), .ZN(n7630)
         );
  NAND2_X1 U8642 ( .A1(n7630), .A2(n11007), .ZN(n7435) );
  OAI21_X1 U8643 ( .B1(n11007), .B2(n7289), .A(n7435), .ZN(P2_U3520) );
  INV_X1 U8644 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7444) );
  NAND2_X1 U8645 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n7493), .ZN(n7438) );
  MUX2_X1 U8646 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7436), .S(n7493), .Z(n7485)
         );
  OAI21_X1 U8647 ( .B1(n7446), .B2(n7408), .A(n7437), .ZN(n7484) );
  NAND2_X1 U8648 ( .A1(n7485), .A2(n7484), .ZN(n7483) );
  NAND2_X1 U8649 ( .A1(n7438), .A2(n7483), .ZN(n7458) );
  MUX2_X1 U8650 ( .A(n7439), .B(P2_REG1_REG_7__SCAN_IN), .S(n7445), .Z(n7457)
         );
  NAND2_X1 U8651 ( .A1(n7458), .A2(n7457), .ZN(n7456) );
  OAI21_X1 U8652 ( .B1(n7439), .B2(n7445), .A(n7456), .ZN(n7442) );
  MUX2_X1 U8653 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7440), .S(n7476), .Z(n7441)
         );
  NAND2_X1 U8654 ( .A1(n7441), .A2(n7442), .ZN(n7468) );
  OAI211_X1 U8655 ( .C1(n7442), .C2(n7441), .A(n8907), .B(n7468), .ZN(n7443)
         );
  NAND2_X1 U8656 ( .A1(P2_U3152), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8144) );
  OAI211_X1 U8657 ( .C1(n8929), .C2(n7444), .A(n7443), .B(n8144), .ZN(n7454)
         );
  INV_X1 U8658 ( .A(n7445), .ZN(n7466) );
  XNOR2_X1 U8659 ( .A(n7445), .B(n7892), .ZN(n7462) );
  INV_X1 U8660 ( .A(n7446), .ZN(n7448) );
  NAND2_X1 U8661 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n7493), .ZN(n7449) );
  OAI21_X1 U8662 ( .B1(n7493), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7449), .ZN(
        n7489) );
  AOI21_X1 U8663 ( .B1(n7493), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7488), .ZN(
        n7463) );
  NOR2_X1 U8664 ( .A1(n7462), .A2(n7463), .ZN(n7461) );
  AOI21_X1 U8665 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7466), .A(n7461), .ZN(
        n7452) );
  NAND2_X1 U8666 ( .A1(n7476), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7450) );
  OAI21_X1 U8667 ( .B1(n7476), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7450), .ZN(
        n7451) );
  NOR2_X1 U8668 ( .A1(n7452), .A2(n7451), .ZN(n7475) );
  AOI211_X1 U8669 ( .C1(n7452), .C2(n7451), .A(n7475), .B(n8961), .ZN(n7453)
         );
  AOI211_X1 U8670 ( .C1(n8959), .C2(n7476), .A(n7454), .B(n7453), .ZN(n7455)
         );
  INV_X1 U8671 ( .A(n7455), .ZN(P2_U3253) );
  INV_X1 U8672 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7460) );
  OAI211_X1 U8673 ( .C1(n7458), .C2(n7457), .A(n8907), .B(n7456), .ZN(n7459)
         );
  NAND2_X1 U8674 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7964) );
  OAI211_X1 U8675 ( .C1(n8929), .C2(n7460), .A(n7459), .B(n7964), .ZN(n7465)
         );
  AOI211_X1 U8676 ( .C1(n7463), .C2(n7462), .A(n7461), .B(n8961), .ZN(n7464)
         );
  AOI211_X1 U8677 ( .C1(n8959), .C2(n7466), .A(n7465), .B(n7464), .ZN(n7467)
         );
  INV_X1 U8678 ( .A(n7467), .ZN(P2_U3252) );
  INV_X1 U8679 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7474) );
  OAI21_X1 U8680 ( .B1(n7469), .B2(n7440), .A(n7468), .ZN(n7472) );
  MUX2_X1 U8681 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7470), .S(n7537), .Z(n7471)
         );
  NAND2_X1 U8682 ( .A1(n7471), .A2(n7472), .ZN(n7528) );
  OAI211_X1 U8683 ( .C1(n7472), .C2(n7471), .A(n8907), .B(n7528), .ZN(n7473)
         );
  NAND2_X1 U8684 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8097) );
  OAI211_X1 U8685 ( .C1(n8929), .C2(n7474), .A(n7473), .B(n8097), .ZN(n7481)
         );
  NAND2_X1 U8686 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n7537), .ZN(n7477) );
  OAI21_X1 U8687 ( .B1(n7537), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7477), .ZN(
        n7478) );
  AOI211_X1 U8688 ( .C1(n7479), .C2(n7478), .A(n7536), .B(n8961), .ZN(n7480)
         );
  AOI211_X1 U8689 ( .C1(n8959), .C2(n7537), .A(n7481), .B(n7480), .ZN(n7482)
         );
  INV_X1 U8690 ( .A(n7482), .ZN(P2_U3254) );
  INV_X1 U8691 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7487) );
  OAI211_X1 U8692 ( .C1(n7485), .C2(n7484), .A(n8907), .B(n7483), .ZN(n7486)
         );
  NAND2_X1 U8693 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8674) );
  OAI211_X1 U8694 ( .C1(n8929), .C2(n7487), .A(n7486), .B(n8674), .ZN(n7492)
         );
  AOI211_X1 U8695 ( .C1(n7490), .C2(n7489), .A(n7488), .B(n8961), .ZN(n7491)
         );
  AOI211_X1 U8696 ( .C1(n8959), .C2(n7493), .A(n7492), .B(n7491), .ZN(n7494)
         );
  INV_X1 U8697 ( .A(n7494), .ZN(P2_U3251) );
  AOI21_X1 U8698 ( .B1(n11029), .B2(n7495), .A(n9764), .ZN(n7523) );
  INV_X1 U8699 ( .A(n7523), .ZN(n7509) );
  INV_X1 U8700 ( .A(n9798), .ZN(n8454) );
  AOI22_X1 U8701 ( .A1(n7509), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n8454), .B2(
        n10107), .ZN(n7501) );
  OR2_X1 U8702 ( .A1(n7497), .A2(n7496), .ZN(n7498) );
  NAND2_X1 U8703 ( .A1(n7499), .A2(n7498), .ZN(n10120) );
  AOI22_X1 U8704 ( .A1(n10120), .A2(n9756), .B1(n8014), .B2(n9803), .ZN(n7500)
         );
  NAND2_X1 U8705 ( .A1(n7501), .A2(n7500), .ZN(P1_U3230) );
  INV_X1 U8706 ( .A(n7502), .ZN(n7520) );
  AOI22_X1 U8707 ( .A1(n10238), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10594), .ZN(n7503) );
  OAI21_X1 U8708 ( .B1(n7520), .B2(n10596), .A(n7503), .ZN(P1_U3336) );
  NAND2_X1 U8709 ( .A1(n7505), .A2(n7504), .ZN(n7507) );
  XNOR2_X1 U8710 ( .A(n7507), .B(n7506), .ZN(n7512) );
  INV_X1 U8711 ( .A(n9756), .ZN(n9805) );
  AND2_X1 U8712 ( .A1(n7980), .A2(n10827), .ZN(n10696) );
  INV_X1 U8713 ( .A(n9764), .ZN(n7508) );
  AOI22_X1 U8714 ( .A1(n8454), .A2(n7832), .B1(n10696), .B2(n7508), .ZN(n7511)
         );
  INV_X1 U8715 ( .A(n9800), .ZN(n9750) );
  AOI22_X1 U8716 ( .A1(n7509), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9750), .B2(
        n6469), .ZN(n7510) );
  OAI211_X1 U8717 ( .C1(n7512), .C2(n9805), .A(n7511), .B(n7510), .ZN(P1_U3220) );
  INV_X1 U8718 ( .A(n8840), .ZN(n8765) );
  INV_X1 U8719 ( .A(n8845), .ZN(n8769) );
  INV_X1 U8720 ( .A(n8903), .ZN(n7547) );
  OAI22_X1 U8721 ( .A1(n8769), .A2(n7547), .B1(n7513), .B2(n8882), .ZN(n7515)
         );
  AOI22_X1 U8722 ( .A1(n7515), .A2(n7514), .B1(n10733), .B2(n7783), .ZN(n7518)
         );
  NAND2_X1 U8723 ( .A1(n8723), .A2(n7516), .ZN(n8642) );
  NAND2_X1 U8724 ( .A1(n8642), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7517) );
  OAI211_X1 U8725 ( .C1(n8765), .C2(n7778), .A(n7518), .B(n7517), .ZN(P2_U3234) );
  INV_X1 U8726 ( .A(n8924), .ZN(n8932) );
  INV_X1 U8727 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7519) );
  OAI222_X1 U8728 ( .A1(n8593), .A2(n7520), .B1(n8932), .B2(P2_U3152), .C1(
        n7519), .C2(n9696), .ZN(P2_U3341) );
  NAND2_X1 U8729 ( .A1(n7521), .A2(n7522), .ZN(n7568) );
  OAI21_X1 U8730 ( .B1(n7521), .B2(n7522), .A(n7568), .ZN(n7526) );
  NAND2_X1 U8731 ( .A1(n7994), .A2(n10827), .ZN(n10705) );
  OAI22_X1 U8732 ( .A1(n9798), .A2(n6507), .B1(n10705), .B2(n9764), .ZN(n7525)
         );
  OAI22_X1 U8733 ( .A1(n7523), .A2(n10134), .B1(n9800), .B2(n7847), .ZN(n7524)
         );
  AOI211_X1 U8734 ( .C1(n7526), .C2(n9756), .A(n7525), .B(n7524), .ZN(n7527)
         );
  INV_X1 U8735 ( .A(n7527), .ZN(P1_U3235) );
  INV_X1 U8736 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7535) );
  OAI21_X1 U8737 ( .B1(n7529), .B2(n7470), .A(n7528), .ZN(n7532) );
  MUX2_X1 U8738 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7530), .S(n7556), .Z(n7531)
         );
  NAND2_X1 U8739 ( .A1(n7531), .A2(n7532), .ZN(n7557) );
  OAI211_X1 U8740 ( .C1(n7532), .C2(n7531), .A(n8907), .B(n7557), .ZN(n7534)
         );
  OAI211_X1 U8741 ( .C1(n8929), .C2(n7535), .A(n7534), .B(n7533), .ZN(n7542)
         );
  NAND2_X1 U8742 ( .A1(n7556), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7538) );
  OAI21_X1 U8743 ( .B1(n7556), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7538), .ZN(
        n7539) );
  AOI211_X1 U8744 ( .C1(n7540), .C2(n7539), .A(n5052), .B(n8961), .ZN(n7541)
         );
  AOI211_X1 U8745 ( .C1(n8959), .C2(n7556), .A(n7542), .B(n7541), .ZN(n7543)
         );
  INV_X1 U8746 ( .A(n7543), .ZN(P2_U3255) );
  INV_X1 U8747 ( .A(n8639), .ZN(n7544) );
  AOI21_X1 U8748 ( .B1(n7546), .B2(n7545), .A(n7544), .ZN(n7551) );
  INV_X1 U8749 ( .A(n10731), .ZN(n8748) );
  OAI22_X1 U8750 ( .A1(n8748), .A2(n7547), .B1(n5112), .B2(n10736), .ZN(n7549)
         );
  INV_X1 U8751 ( .A(n10733), .ZN(n8856) );
  NOR2_X1 U8752 ( .A1(n8856), .A2(n7710), .ZN(n7548) );
  AOI211_X1 U8753 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(n8642), .A(n7549), .B(
        n7548), .ZN(n7550) );
  OAI21_X1 U8754 ( .B1(n7551), .B2(n8882), .A(n7550), .ZN(P2_U3224) );
  AOI21_X1 U8755 ( .B1(n7556), .B2(P2_REG2_REG_10__SCAN_IN), .A(n5052), .ZN(
        n7553) );
  MUX2_X1 U8756 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7660), .S(n7652), .Z(n7552)
         );
  NAND2_X1 U8757 ( .A1(n7552), .A2(n7553), .ZN(n7663) );
  OAI21_X1 U8758 ( .B1(n7553), .B2(n7552), .A(n7663), .ZN(n7565) );
  AOI21_X1 U8759 ( .B1(n8953), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7554), .ZN(
        n7562) );
  MUX2_X1 U8760 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7555), .S(n7652), .Z(n7560)
         );
  NAND2_X1 U8761 ( .A1(n7556), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U8762 ( .A1(n7558), .A2(n7557), .ZN(n7559) );
  NAND2_X1 U8763 ( .A1(n7560), .A2(n7559), .ZN(n7654) );
  OAI211_X1 U8764 ( .C1(n7560), .C2(n7559), .A(n8907), .B(n7654), .ZN(n7561)
         );
  OAI211_X1 U8765 ( .C1(n7563), .C2(n7661), .A(n7562), .B(n7561), .ZN(n7564)
         );
  AOI21_X1 U8766 ( .B1(n7936), .B2(n7565), .A(n7564), .ZN(n7566) );
  INV_X1 U8767 ( .A(n7566), .ZN(P2_U3256) );
  NAND2_X1 U8768 ( .A1(n7568), .A2(n7567), .ZN(n7571) );
  AND2_X1 U8769 ( .A1(n7570), .A2(n7569), .ZN(n8623) );
  OAI21_X1 U8770 ( .B1(n6524), .B2(n7571), .A(n8623), .ZN(n7576) );
  OAI22_X1 U8771 ( .A1(n9800), .A2(n7831), .B1(n10719), .B2(n9753), .ZN(n7575)
         );
  INV_X1 U8772 ( .A(n7834), .ZN(n7636) );
  OR2_X1 U8773 ( .A1(n9798), .A2(n7636), .ZN(n7573) );
  INV_X1 U8774 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8117) );
  NOR2_X1 U8775 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8117), .ZN(n10145) );
  INV_X1 U8776 ( .A(n10145), .ZN(n7572) );
  OAI211_X1 U8777 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9799), .A(n7573), .B(
        n7572), .ZN(n7574) );
  AOI211_X1 U8778 ( .C1(n7576), .C2(n9756), .A(n7575), .B(n7574), .ZN(n7577)
         );
  INV_X1 U8779 ( .A(n7577), .ZN(P1_U3216) );
  NAND2_X1 U8780 ( .A1(n10106), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7578) );
  OAI21_X1 U8781 ( .B1(n10284), .B2(n10106), .A(n7578), .ZN(P1_U3584) );
  INV_X1 U8782 ( .A(n7579), .ZN(n7583) );
  AOI22_X1 U8783 ( .A1(n10255), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10594), .ZN(n7580) );
  OAI21_X1 U8784 ( .B1(n7583), .B2(n10596), .A(n7580), .ZN(P1_U3335) );
  AOI22_X1 U8785 ( .A1(n8939), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7581), .ZN(n7582) );
  OAI21_X1 U8786 ( .B1(n7583), .B2(n9699), .A(n7582), .ZN(P2_U3340) );
  XOR2_X1 U8787 ( .A(n7586), .B(n7584), .Z(n7585) );
  AOI222_X1 U8788 ( .A1(n10798), .A2(n7585), .B1(n10730), .B2(n9139), .C1(
        n8903), .C2(n9137), .ZN(n7714) );
  XOR2_X1 U8789 ( .A(n7607), .B(n7586), .Z(n7712) );
  OR2_X1 U8790 ( .A1(n7606), .A2(n7783), .ZN(n7752) );
  NAND2_X1 U8791 ( .A1(n7606), .A2(n7783), .ZN(n7587) );
  NAND2_X1 U8792 ( .A1(n7752), .A2(n7587), .ZN(n7705) );
  OR2_X1 U8793 ( .A1(n7588), .A2(n7702), .ZN(n11000) );
  OAI22_X1 U8794 ( .A1(n7705), .A2(n11000), .B1(n7710), .B2(n10998), .ZN(n7589) );
  AOI21_X1 U8795 ( .B1(n7712), .B2(n11004), .A(n7589), .ZN(n7590) );
  NAND2_X1 U8796 ( .A1(n7714), .A2(n7590), .ZN(n7628) );
  NAND2_X1 U8797 ( .A1(n7628), .A2(n11007), .ZN(n7591) );
  OAI21_X1 U8798 ( .B1(n11007), .B2(n5595), .A(n7591), .ZN(P2_U3521) );
  INV_X1 U8799 ( .A(n10728), .ZN(n7594) );
  INV_X1 U8800 ( .A(n8900), .ZN(n7721) );
  NOR3_X1 U8801 ( .A1(n8769), .A2(n7721), .A3(n7592), .ZN(n7593) );
  AOI21_X1 U8802 ( .B1(n7594), .B2(n10727), .A(n7593), .ZN(n7603) );
  NAND2_X1 U8803 ( .A1(n10728), .A2(n7595), .ZN(n8772) );
  INV_X1 U8804 ( .A(n8772), .ZN(n7601) );
  INV_X1 U8805 ( .A(n8898), .ZN(n8680) );
  NAND2_X1 U8806 ( .A1(n10731), .A2(n8900), .ZN(n7597) );
  OAI211_X1 U8807 ( .C1(n8680), .C2(n10736), .A(n7597), .B(n7596), .ZN(n7600)
         );
  NAND2_X1 U8808 ( .A1(n10733), .A2(n7727), .ZN(n7598) );
  OAI21_X1 U8809 ( .B1(n10742), .B2(n7726), .A(n7598), .ZN(n7599) );
  AOI211_X1 U8810 ( .C1(n7601), .C2(n10727), .A(n7600), .B(n7599), .ZN(n7602)
         );
  OAI21_X1 U8811 ( .B1(n7604), .B2(n7603), .A(n7602), .ZN(P2_U3232) );
  INV_X1 U8812 ( .A(n11004), .ZN(n10962) );
  NAND2_X1 U8813 ( .A1(n7605), .A2(n7710), .ZN(n7608) );
  AOI21_X1 U8814 ( .B1(n7608), .B2(n7607), .A(n5560), .ZN(n7746) );
  NAND2_X1 U8815 ( .A1(n7746), .A2(n7745), .ZN(n7744) );
  NAND2_X1 U8816 ( .A1(n5112), .A2(n7609), .ZN(n7610) );
  NAND2_X1 U8817 ( .A1(n7744), .A2(n7610), .ZN(n7611) );
  NAND2_X1 U8818 ( .A1(n7611), .A2(n7613), .ZN(n7723) );
  OAI21_X1 U8819 ( .B1(n7611), .B2(n7613), .A(n7723), .ZN(n7741) );
  INV_X1 U8820 ( .A(n7741), .ZN(n7619) );
  NAND3_X1 U8821 ( .A1(n7747), .A2(n7614), .A3(n7613), .ZN(n7615) );
  NAND2_X1 U8822 ( .A1(n7612), .A2(n7615), .ZN(n7616) );
  AOI222_X1 U8823 ( .A1(n10798), .A2(n7616), .B1(n10730), .B2(n9137), .C1(
        n8899), .C2(n9139), .ZN(n7743) );
  OR2_X1 U8824 ( .A1(n7753), .A2(n7739), .ZN(n7617) );
  AND2_X1 U8825 ( .A1(n7617), .A2(n7728), .ZN(n7736) );
  INV_X1 U8826 ( .A(n11000), .ZN(n10803) );
  AOI22_X1 U8827 ( .A1(n7736), .A2(n10803), .B1(n10904), .B2(n10732), .ZN(
        n7618) );
  OAI211_X1 U8828 ( .C1(n10962), .C2(n7619), .A(n7743), .B(n7618), .ZN(n7622)
         );
  NAND2_X1 U8829 ( .A1(n7622), .A2(n11007), .ZN(n7620) );
  OAI21_X1 U8830 ( .B1(n11007), .B2(n7323), .A(n7620), .ZN(P2_U3523) );
  AND2_X2 U8831 ( .A1(n7621), .A2(n7693), .ZN(n11011) );
  NAND2_X1 U8832 ( .A1(n7622), .A2(n11011), .ZN(n7623) );
  OAI21_X1 U8833 ( .B1(n11011), .B2(n5622), .A(n7623), .ZN(P2_U3460) );
  INV_X1 U8834 ( .A(n7624), .ZN(n7626) );
  OAI222_X1 U8835 ( .A1(n10260), .A2(P1_U3084), .B1(n10596), .B2(n7626), .C1(
        n7625), .C2(n8813), .ZN(P1_U3334) );
  OAI222_X1 U8836 ( .A1(n9696), .A2(n7627), .B1(n8593), .B2(n7626), .C1(n9004), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U8837 ( .A1(n7628), .A2(n11011), .ZN(n7629) );
  OAI21_X1 U8838 ( .B1(n11011), .B2(n5596), .A(n7629), .ZN(P2_U3454) );
  NAND2_X1 U8839 ( .A1(n7630), .A2(n11011), .ZN(n7631) );
  OAI21_X1 U8840 ( .B1(n11011), .B2(n5580), .A(n7631), .ZN(P2_U3451) );
  NAND2_X1 U8841 ( .A1(n7633), .A2(n7632), .ZN(n7635) );
  XNOR2_X1 U8842 ( .A(n7635), .B(n7634), .ZN(n7641) );
  OAI22_X1 U8843 ( .A1(n9800), .A2(n7636), .B1(n10764), .B2(n9753), .ZN(n7640)
         );
  OR2_X1 U8844 ( .A1(n9798), .A2(n8067), .ZN(n7638) );
  OAI211_X1 U8845 ( .C1(n9799), .C2(n10778), .A(n7638), .B(n7637), .ZN(n7639)
         );
  AOI211_X1 U8846 ( .C1(n7641), .C2(n9756), .A(n7640), .B(n7639), .ZN(n7642)
         );
  INV_X1 U8847 ( .A(n7642), .ZN(P1_U3225) );
  OAI21_X1 U8848 ( .B1(n7645), .B2(n7644), .A(n7643), .ZN(n7650) );
  OAI22_X1 U8849 ( .A1(n9798), .A2(n8022), .B1(n7899), .B2(n9753), .ZN(n7649)
         );
  OR2_X1 U8850 ( .A1(n9800), .A2(n8625), .ZN(n7647) );
  AND2_X1 U8851 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10649) );
  INV_X1 U8852 ( .A(n10649), .ZN(n7646) );
  OAI211_X1 U8853 ( .C1(n9799), .C2(n7843), .A(n7647), .B(n7646), .ZN(n7648)
         );
  AOI211_X1 U8854 ( .C1(n7650), .C2(n9756), .A(n7649), .B(n7648), .ZN(n7651)
         );
  INV_X1 U8855 ( .A(n7651), .ZN(P1_U3237) );
  INV_X1 U8856 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U8857 ( .A1(n7652), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7653) );
  MUX2_X1 U8858 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n5786), .S(n7768), .Z(n7655)
         );
  NOR2_X1 U8859 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  OAI21_X1 U8860 ( .B1(n7763), .B2(n7657), .A(n8907), .ZN(n7658) );
  NAND2_X1 U8861 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8300) );
  OAI211_X1 U8862 ( .C1(n8929), .C2(n7659), .A(n7658), .B(n8300), .ZN(n7669)
         );
  NAND2_X1 U8863 ( .A1(n7661), .A2(n7660), .ZN(n7662) );
  OR2_X1 U8864 ( .A1(n7768), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7665) );
  NAND2_X1 U8865 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7768), .ZN(n7664) );
  NAND2_X1 U8866 ( .A1(n7665), .A2(n7664), .ZN(n7666) );
  AOI211_X1 U8867 ( .C1(n7667), .C2(n7666), .A(n7767), .B(n8961), .ZN(n7668)
         );
  AOI211_X1 U8868 ( .C1(n8959), .C2(n7768), .A(n7669), .B(n7668), .ZN(n7670)
         );
  INV_X1 U8869 ( .A(n7670), .ZN(P2_U3257) );
  AOI22_X1 U8870 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n10663), .B1(n7671), .B2(
        n6624), .ZN(n10666) );
  NOR2_X1 U8871 ( .A1(n10177), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7672) );
  AOI21_X1 U8872 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10177), .A(n7672), .ZN(
        n10169) );
  OAI21_X1 U8873 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7681), .A(n7673), .ZN(
        n10170) );
  NAND2_X1 U8874 ( .A1(n10169), .A2(n10170), .ZN(n10168) );
  OAI21_X1 U8875 ( .B1(n10177), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10168), .ZN(
        n10665) );
  NAND2_X1 U8876 ( .A1(n10666), .A2(n10665), .ZN(n10664) );
  OAI21_X1 U8877 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n10663), .A(n10664), .ZN(
        n10686) );
  NAND2_X1 U8878 ( .A1(n7683), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7674) );
  NOR2_X1 U8879 ( .A1(n7683), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10687) );
  AOI21_X1 U8880 ( .B1(n10686), .B2(n7674), .A(n10687), .ZN(n10685) );
  MUX2_X1 U8881 ( .A(n7675), .B(P1_REG1_REG_12__SCAN_IN), .S(n7869), .Z(n7676)
         );
  NOR2_X1 U8882 ( .A1(n10685), .A2(n7676), .ZN(n7864) );
  AOI21_X1 U8883 ( .B1(n10685), .B2(n7676), .A(n7864), .ZN(n7691) );
  INV_X1 U8884 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7678) );
  AND2_X1 U8885 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8293) );
  INV_X1 U8886 ( .A(n8293), .ZN(n7677) );
  OAI21_X1 U8887 ( .B1(n10679), .B2(n7678), .A(n7677), .ZN(n7689) );
  NOR2_X1 U8888 ( .A1(n7683), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10683) );
  NAND2_X1 U8889 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10663), .ZN(n7682) );
  NAND2_X1 U8890 ( .A1(n10177), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7679) );
  OAI21_X1 U8891 ( .B1(n10177), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7679), .ZN(
        n10174) );
  OAI21_X1 U8892 ( .B1(n7681), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7680), .ZN(
        n10175) );
  NOR2_X1 U8893 ( .A1(n10174), .A2(n10175), .ZN(n10173) );
  OAI21_X1 U8894 ( .B1(n10663), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7682), .ZN(
        n10659) );
  AND2_X1 U8895 ( .A1(n7683), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10682) );
  NOR2_X1 U8896 ( .A1(n10681), .A2(n10682), .ZN(n7687) );
  OR2_X1 U8897 ( .A1(n7869), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U8898 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7869), .ZN(n7684) );
  NAND2_X1 U8899 ( .A1(n7685), .A2(n7684), .ZN(n7686) );
  AOI211_X1 U8900 ( .C1(n7687), .C2(n7686), .A(n7868), .B(n10657), .ZN(n7688)
         );
  AOI211_X1 U8901 ( .C1(n10672), .C2(n7869), .A(n7689), .B(n7688), .ZN(n7690)
         );
  OAI21_X1 U8902 ( .B1(n7691), .B2(n10264), .A(n7690), .ZN(P1_U3253) );
  INV_X1 U8903 ( .A(n7692), .ZN(n7694) );
  AND2_X1 U8904 ( .A1(n7694), .A2(n7693), .ZN(n7697) );
  INV_X1 U8905 ( .A(n7695), .ZN(n7696) );
  NAND2_X1 U8906 ( .A1(n7697), .A2(n7696), .ZN(n7703) );
  INV_X1 U8907 ( .A(n7698), .ZN(n7699) );
  NAND2_X1 U8908 ( .A1(n7700), .A2(n7699), .ZN(n10809) );
  NAND2_X1 U8909 ( .A1(n7703), .A2(n10809), .ZN(n8422) );
  INV_X2 U8910 ( .A(n8422), .ZN(n10817) );
  NAND2_X1 U8911 ( .A1(n7701), .A2(n7811), .ZN(n7757) );
  NAND2_X1 U8912 ( .A1(n8247), .A2(n7757), .ZN(n10794) );
  NAND2_X1 U8913 ( .A1(n10815), .A2(n10794), .ZN(n9146) );
  INV_X1 U8914 ( .A(n9146), .ZN(n9114) );
  NOR2_X1 U8915 ( .A1(n7702), .A2(n7811), .ZN(n10805) );
  NAND2_X1 U8916 ( .A1(n10815), .A2(n10805), .ZN(n9133) );
  OR2_X1 U8917 ( .A1(n7703), .A2(n7036), .ZN(n8667) );
  OAI22_X1 U8918 ( .A1(n8667), .A2(n7705), .B1(n7704), .B2(n10809), .ZN(n7706)
         );
  INV_X1 U8919 ( .A(n7706), .ZN(n7709) );
  OR2_X1 U8920 ( .A1(n10815), .A2(n7707), .ZN(n7708) );
  OAI211_X1 U8921 ( .C1(n7710), .C2(n9133), .A(n7709), .B(n7708), .ZN(n7711)
         );
  AOI21_X1 U8922 ( .B1(n9114), .B2(n7712), .A(n7711), .ZN(n7713) );
  OAI21_X1 U8923 ( .B1(n7714), .B2(n10817), .A(n7713), .ZN(P2_U3295) );
  NAND3_X1 U8924 ( .A1(n7612), .A2(n7724), .A3(n7716), .ZN(n7717) );
  NAND2_X1 U8925 ( .A1(n7715), .A2(n7717), .ZN(n7718) );
  NAND2_X1 U8926 ( .A1(n7718), .A2(n10798), .ZN(n7720) );
  AOI22_X1 U8927 ( .A1(n9139), .A2(n8898), .B1(n8900), .B2(n9137), .ZN(n7719)
         );
  NAND2_X1 U8928 ( .A1(n7720), .A2(n7719), .ZN(n10754) );
  INV_X1 U8929 ( .A(n10754), .ZN(n7734) );
  NAND2_X1 U8930 ( .A1(n7721), .A2(n7739), .ZN(n7722) );
  OAI21_X1 U8931 ( .B1(n7725), .B2(n7724), .A(n10791), .ZN(n10756) );
  NOR2_X1 U8932 ( .A1(n7726), .A2(n10809), .ZN(n7730) );
  OAI21_X1 U8933 ( .B1(n5325), .B2(n10752), .A(n10802), .ZN(n10753) );
  NOR2_X1 U8934 ( .A1(n10753), .A2(n8667), .ZN(n7729) );
  AOI211_X1 U8935 ( .C1(n10817), .C2(P2_REG2_REG_4__SCAN_IN), .A(n7730), .B(
        n7729), .ZN(n7731) );
  OAI21_X1 U8936 ( .B1(n10752), .B2(n9133), .A(n7731), .ZN(n7732) );
  AOI21_X1 U8937 ( .B1(n9114), .B2(n10756), .A(n7732), .ZN(n7733) );
  OAI21_X1 U8938 ( .B1(n10817), .B2(n7734), .A(n7733), .ZN(P2_U3292) );
  INV_X1 U8939 ( .A(n8667), .ZN(n9144) );
  INV_X1 U8940 ( .A(n10809), .ZN(n9130) );
  AOI22_X1 U8941 ( .A1(n7736), .A2(n9144), .B1(n9130), .B2(n7735), .ZN(n7738)
         );
  NAND2_X1 U8942 ( .A1(n10817), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7737) );
  OAI211_X1 U8943 ( .C1(n7739), .C2(n9133), .A(n7738), .B(n7737), .ZN(n7740)
         );
  AOI21_X1 U8944 ( .B1(n7741), .B2(n9114), .A(n7740), .ZN(n7742) );
  OAI21_X1 U8945 ( .B1(n7743), .B2(n10817), .A(n7742), .ZN(P2_U3293) );
  OAI21_X1 U8946 ( .B1(n7746), .B2(n7745), .A(n7744), .ZN(n10716) );
  INV_X1 U8947 ( .A(n10716), .ZN(n7758) );
  AOI22_X1 U8948 ( .A1(n9137), .A2(n8901), .B1(n8900), .B2(n8837), .ZN(n7751)
         );
  NAND2_X1 U8949 ( .A1(n7749), .A2(n10798), .ZN(n7750) );
  OAI211_X1 U8950 ( .C1(n7758), .C2(n8247), .A(n7751), .B(n7750), .ZN(n10714)
         );
  INV_X1 U8951 ( .A(n10714), .ZN(n7762) );
  INV_X1 U8952 ( .A(n7752), .ZN(n7755) );
  INV_X1 U8953 ( .A(n7753), .ZN(n7754) );
  OAI21_X1 U8954 ( .B1(n7609), .B2(n7755), .A(n7754), .ZN(n10713) );
  OAI22_X1 U8955 ( .A1(n10713), .A2(n8667), .B1(n7756), .B2(n10809), .ZN(n7760) );
  OR2_X1 U8956 ( .A1(n10817), .A2(n7757), .ZN(n8256) );
  OAI22_X1 U8957 ( .A1(n7758), .A2(n8256), .B1(n7609), .B2(n9133), .ZN(n7759)
         );
  AOI211_X1 U8958 ( .C1(P2_REG2_REG_2__SCAN_IN), .C2(n10817), .A(n7760), .B(
        n7759), .ZN(n7761) );
  OAI21_X1 U8959 ( .B1(n10817), .B2(n7762), .A(n7761), .ZN(P2_U3294) );
  AOI21_X1 U8960 ( .B1(n5786), .B2(n7764), .A(n7763), .ZN(n7766) );
  AOI22_X1 U8961 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7925), .B1(n7930), .B2(
        n5849), .ZN(n7765) );
  NOR2_X1 U8962 ( .A1(n7766), .A2(n7765), .ZN(n7924) );
  AOI21_X1 U8963 ( .B1(n7766), .B2(n7765), .A(n7924), .ZN(n7777) );
  NOR2_X1 U8964 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n7930), .ZN(n7769) );
  AOI21_X1 U8965 ( .B1(n7930), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7769), .ZN(
        n7770) );
  OAI21_X1 U8966 ( .B1(n7771), .B2(n7770), .A(n7929), .ZN(n7772) );
  NAND2_X1 U8967 ( .A1(n7772), .A2(n7936), .ZN(n7776) );
  INV_X1 U8968 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U8969 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8702) );
  OAI21_X1 U8970 ( .B1(n8929), .B2(n7773), .A(n8702), .ZN(n7774) );
  AOI21_X1 U8971 ( .B1(n8959), .B2(n7930), .A(n7774), .ZN(n7775) );
  OAI211_X1 U8972 ( .C1(n7777), .C2(n8957), .A(n7776), .B(n7775), .ZN(P2_U3258) );
  INV_X1 U8973 ( .A(n7781), .ZN(n7786) );
  OAI21_X1 U8974 ( .B1(n10809), .B2(n7779), .A(n7778), .ZN(n7780) );
  AOI21_X1 U8975 ( .B1(n7781), .B2(n10798), .A(n7780), .ZN(n7782) );
  MUX2_X1 U8976 ( .A(n7782), .B(n7393), .S(n10817), .Z(n7785) );
  OAI21_X1 U8977 ( .B1(n9122), .B2(n9144), .A(n7783), .ZN(n7784) );
  OAI211_X1 U8978 ( .C1(n7786), .C2(n9146), .A(n7785), .B(n7784), .ZN(P2_U3296) );
  XNOR2_X1 U8979 ( .A(n7787), .B(n7804), .ZN(n7788) );
  NAND2_X1 U8980 ( .A1(n7788), .A2(n10798), .ZN(n7790) );
  AOI22_X1 U8981 ( .A1(n9137), .A2(n8898), .B1(n8896), .B2(n8837), .ZN(n7789)
         );
  NAND2_X1 U8982 ( .A1(n7790), .A2(n7789), .ZN(n10841) );
  INV_X1 U8983 ( .A(n10841), .ZN(n7808) );
  OAI22_X1 U8984 ( .A1(n10815), .A2(n7791), .B1(n8675), .B2(n10809), .ZN(n7795) );
  AND2_X1 U8985 ( .A1(n7792), .A2(n10838), .ZN(n7891) );
  NOR2_X1 U8986 ( .A1(n7792), .A2(n10838), .ZN(n7793) );
  OR2_X1 U8987 ( .A1(n7891), .A2(n7793), .ZN(n10839) );
  NOR2_X1 U8988 ( .A1(n10839), .A2(n8667), .ZN(n7794) );
  AOI211_X1 U8989 ( .C1(n9122), .C2(n7796), .A(n7795), .B(n7794), .ZN(n7807)
         );
  NAND2_X1 U8990 ( .A1(n10737), .A2(n10752), .ZN(n10790) );
  AND2_X1 U8991 ( .A1(n10790), .A2(n7799), .ZN(n7801) );
  AND2_X1 U8992 ( .A1(n7801), .A2(n7797), .ZN(n7798) );
  NAND2_X1 U8993 ( .A1(n10791), .A2(n7798), .ZN(n7888) );
  INV_X1 U8994 ( .A(n7799), .ZN(n7800) );
  AND2_X1 U8995 ( .A1(n7888), .A2(n7886), .ZN(n10837) );
  NAND2_X1 U8996 ( .A1(n10791), .A2(n7801), .ZN(n7803) );
  AND2_X1 U8997 ( .A1(n7803), .A2(n7802), .ZN(n7805) );
  NAND2_X1 U8998 ( .A1(n7805), .A2(n7804), .ZN(n10836) );
  NAND3_X1 U8999 ( .A1(n10837), .A2(n9114), .A3(n10836), .ZN(n7806) );
  OAI211_X1 U9000 ( .C1(n7808), .C2(n10817), .A(n7807), .B(n7806), .ZN(
        P2_U3290) );
  INV_X1 U9001 ( .A(n7809), .ZN(n7821) );
  OAI222_X1 U9002 ( .A1(n8593), .A2(n7821), .B1(P2_U3152), .B2(n7811), .C1(
        n7810), .C2(n9696), .ZN(P2_U3338) );
  OAI21_X1 U9003 ( .B1(n7814), .B2(n7813), .A(n7812), .ZN(n7819) );
  OAI22_X1 U9004 ( .A1(n9800), .A2(n8067), .B1(n9799), .B2(n8073), .ZN(n7818)
         );
  AOI21_X1 U9005 ( .B1(n8454), .B2(n10102), .A(n7815), .ZN(n7816) );
  OAI21_X1 U9006 ( .B1(n10846), .B2(n9753), .A(n7816), .ZN(n7817) );
  AOI211_X1 U9007 ( .C1(n7819), .C2(n9756), .A(n7818), .B(n7817), .ZN(n7820)
         );
  INV_X1 U9008 ( .A(n7820), .ZN(P1_U3211) );
  OAI222_X1 U9009 ( .A1(P1_U3084), .A2(n7822), .B1(n10596), .B2(n7821), .C1(
        n9592), .C2(n8813), .ZN(P1_U3333) );
  INV_X1 U9010 ( .A(n7823), .ZN(n8634) );
  OAI222_X1 U9011 ( .A1(n8593), .A2(n8634), .B1(P2_U3152), .B2(n7825), .C1(
        n7824), .C2(n9696), .ZN(P2_U3337) );
  NAND2_X1 U9012 ( .A1(n7827), .A2(n7826), .ZN(n7841) );
  INV_X1 U9013 ( .A(n7828), .ZN(n7829) );
  INV_X1 U9014 ( .A(n11019), .ZN(n10789) );
  NAND2_X1 U9015 ( .A1(n8067), .A2(n10826), .ZN(n9930) );
  INV_X1 U9016 ( .A(n8067), .ZN(n10770) );
  NOR2_X1 U9017 ( .A1(n6469), .A2(n9835), .ZN(n7972) );
  NAND2_X1 U9018 ( .A1(n10039), .A2(n7972), .ZN(n7971) );
  INV_X1 U9019 ( .A(n7980), .ZN(n9836) );
  OR2_X1 U9020 ( .A1(n10107), .A2(n9836), .ZN(n7830) );
  NAND2_X1 U9021 ( .A1(n7971), .A2(n7830), .ZN(n9843) );
  NAND2_X1 U9022 ( .A1(n7831), .A2(n7994), .ZN(n9839) );
  INV_X1 U9023 ( .A(n7831), .ZN(n7832) );
  NAND2_X1 U9024 ( .A1(n7832), .A2(n7850), .ZN(n9841) );
  NAND2_X1 U9025 ( .A1(n9839), .A2(n9841), .ZN(n10037) );
  INV_X1 U9026 ( .A(n10037), .ZN(n7833) );
  INV_X1 U9027 ( .A(n6507), .ZN(n10105) );
  NAND2_X1 U9028 ( .A1(n10105), .A2(n10719), .ZN(n8080) );
  NAND2_X1 U9029 ( .A1(n7834), .A2(n10743), .ZN(n9889) );
  AND2_X1 U9030 ( .A1(n8080), .A2(n9889), .ZN(n9885) );
  NAND2_X1 U9031 ( .A1(n6507), .A2(n8118), .ZN(n9888) );
  INV_X1 U9032 ( .A(n9888), .ZN(n8081) );
  OR2_X1 U9033 ( .A1(n7834), .A2(n10743), .ZN(n9887) );
  INV_X1 U9034 ( .A(n9887), .ZN(n7835) );
  AOI21_X1 U9035 ( .B1(n9885), .B2(n8081), .A(n7835), .ZN(n9845) );
  NAND2_X1 U9036 ( .A1(n10766), .A2(n9923), .ZN(n7836) );
  NAND2_X1 U9037 ( .A1(n8625), .A2(n10781), .ZN(n9922) );
  XNOR2_X1 U9038 ( .A(n10040), .B(n9925), .ZN(n7840) );
  NAND2_X1 U9039 ( .A1(n10086), .A2(n10785), .ZN(n7838) );
  NAND2_X1 U9040 ( .A1(n9916), .A2(n10076), .ZN(n7837) );
  NAND2_X1 U9041 ( .A1(n7838), .A2(n7837), .ZN(n10930) );
  INV_X1 U9042 ( .A(n10768), .ZN(n10927) );
  INV_X1 U9043 ( .A(n10769), .ZN(n10925) );
  OAI22_X1 U9044 ( .A1(n8625), .A2(n10927), .B1(n8022), .B2(n10925), .ZN(n7839) );
  AOI21_X1 U9045 ( .B1(n7840), .B2(n10930), .A(n7839), .ZN(n10830) );
  NOR2_X1 U9046 ( .A1(n7841), .A2(n10785), .ZN(n11023) );
  OR2_X1 U9047 ( .A1(n7980), .A2(n8014), .ZN(n7990) );
  NOR2_X1 U9048 ( .A1(n7990), .A2(n7994), .ZN(n8114) );
  NAND2_X1 U9049 ( .A1(n8114), .A2(n10719), .ZN(n8116) );
  OR2_X2 U9050 ( .A1(n8116), .A2(n5207), .ZN(n10760) );
  INV_X1 U9051 ( .A(n10762), .ZN(n7842) );
  AOI21_X1 U9052 ( .B1(n10826), .B2(n7842), .A(n8072), .ZN(n10828) );
  NAND2_X1 U9053 ( .A1(n11019), .A2(n10780), .ZN(n11012) );
  INV_X1 U9054 ( .A(n11019), .ZN(n10465) );
  INV_X1 U9055 ( .A(n7843), .ZN(n7844) );
  INV_X1 U9056 ( .A(n11014), .ZN(n10463) );
  AOI22_X1 U9057 ( .A1(n10465), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7844), .B2(
        n10463), .ZN(n7845) );
  OAI21_X1 U9058 ( .B1(n7899), .B2(n11012), .A(n7845), .ZN(n7861) );
  NAND2_X1 U9059 ( .A1(n10107), .A2(n7980), .ZN(n7846) );
  NAND2_X1 U9060 ( .A1(n7846), .A2(n7970), .ZN(n7849) );
  INV_X1 U9061 ( .A(n10107), .ZN(n7847) );
  NAND2_X1 U9062 ( .A1(n7849), .A2(n7848), .ZN(n7984) );
  NAND2_X1 U9063 ( .A1(n7984), .A2(n10037), .ZN(n7852) );
  NAND2_X1 U9064 ( .A1(n7831), .A2(n7850), .ZN(n7851) );
  NAND2_X1 U9065 ( .A1(n7852), .A2(n7851), .ZN(n8109) );
  NAND2_X1 U9066 ( .A1(n9888), .A2(n8080), .ZN(n10036) );
  NAND2_X1 U9067 ( .A1(n8109), .A2(n10036), .ZN(n8086) );
  NAND2_X1 U9068 ( .A1(n6507), .A2(n10719), .ZN(n8085) );
  OR2_X1 U9069 ( .A1(n7834), .A2(n5207), .ZN(n7853) );
  AND2_X1 U9070 ( .A1(n8085), .A2(n7853), .ZN(n7855) );
  INV_X1 U9071 ( .A(n7853), .ZN(n7854) );
  NAND2_X1 U9072 ( .A1(n9887), .A2(n9889), .ZN(n10035) );
  OR2_X1 U9073 ( .A1(n7904), .A2(n10765), .ZN(n10759) );
  NAND2_X1 U9074 ( .A1(n10104), .A2(n10781), .ZN(n7900) );
  NAND2_X1 U9075 ( .A1(n10759), .A2(n7900), .ZN(n7856) );
  INV_X1 U9076 ( .A(n10040), .ZN(n9926) );
  XNOR2_X1 U9077 ( .A(n7856), .B(n9926), .ZN(n10831) );
  NOR2_X1 U9078 ( .A1(n7858), .A2(n10260), .ZN(n7921) );
  INV_X1 U9079 ( .A(n7921), .ZN(n7859) );
  NAND2_X1 U9080 ( .A1(n7857), .A2(n7859), .ZN(n10776) );
  NAND2_X1 U9081 ( .A1(n11019), .A2(n10776), .ZN(n11021) );
  NOR2_X1 U9082 ( .A1(n10831), .A2(n11021), .ZN(n7860) );
  AOI211_X1 U9083 ( .C1(n10470), .C2(n10828), .A(n7861), .B(n7860), .ZN(n7862)
         );
  OAI21_X1 U9084 ( .B1(n10789), .B2(n10830), .A(n7862), .ZN(P1_U3285) );
  MUX2_X1 U9085 ( .A(n7863), .B(P1_REG1_REG_13__SCAN_IN), .S(n8179), .Z(n7867)
         );
  INV_X1 U9086 ( .A(n7869), .ZN(n7865) );
  AOI21_X1 U9087 ( .B1(n7865), .B2(n7675), .A(n7864), .ZN(n7866) );
  NOR2_X1 U9088 ( .A1(n7866), .A2(n7867), .ZN(n8172) );
  AOI21_X1 U9089 ( .B1(n7867), .B2(n7866), .A(n8172), .ZN(n7879) );
  NAND2_X1 U9090 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n8179), .ZN(n7870) );
  OAI21_X1 U9091 ( .B1(n8179), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7870), .ZN(
        n7871) );
  AOI211_X1 U9092 ( .C1(n7872), .C2(n7871), .A(n8178), .B(n10657), .ZN(n7873)
         );
  AOI21_X1 U9093 ( .B1(n10672), .B2(n8179), .A(n7873), .ZN(n7878) );
  INV_X1 U9094 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7875) );
  INV_X1 U9095 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7874) );
  OR2_X1 U9096 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7874), .ZN(n8335) );
  OAI21_X1 U9097 ( .B1(n10679), .B2(n7875), .A(n8335), .ZN(n7876) );
  INV_X1 U9098 ( .A(n7876), .ZN(n7877) );
  OAI211_X1 U9099 ( .C1(n7879), .C2(n10264), .A(n7878), .B(n7877), .ZN(
        P1_U3254) );
  NAND2_X1 U9100 ( .A1(n7880), .A2(n7889), .ZN(n7881) );
  NAND3_X1 U9101 ( .A1(n7942), .A2(n10798), .A3(n7881), .ZN(n7883) );
  AOI22_X1 U9102 ( .A1(n9139), .A2(n8895), .B1(n8897), .B2(n9137), .ZN(n7882)
         );
  NAND2_X1 U9103 ( .A1(n7883), .A2(n7882), .ZN(n10855) );
  INV_X1 U9104 ( .A(n10855), .ZN(n7898) );
  AND2_X1 U9105 ( .A1(n10837), .A2(n7884), .ZN(n7890) );
  AND2_X1 U9106 ( .A1(n7889), .A2(n7884), .ZN(n7885) );
  AND2_X1 U9107 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  NAND2_X1 U9108 ( .A1(n7888), .A2(n7887), .ZN(n7955) );
  OAI21_X1 U9109 ( .B1(n7890), .B2(n7889), .A(n7955), .ZN(n10857) );
  NAND2_X1 U9110 ( .A1(n7891), .A2(n10853), .ZN(n7949) );
  OAI21_X1 U9111 ( .B1(n7891), .B2(n10853), .A(n7949), .ZN(n10854) );
  OAI22_X1 U9112 ( .A1(n10815), .A2(n7892), .B1(n7966), .B2(n10809), .ZN(n7893) );
  AOI21_X1 U9113 ( .B1(n9122), .B2(n7894), .A(n7893), .ZN(n7895) );
  OAI21_X1 U9114 ( .B1(n10854), .B2(n8667), .A(n7895), .ZN(n7896) );
  AOI21_X1 U9115 ( .B1(n10857), .B2(n9114), .A(n7896), .ZN(n7897) );
  OAI21_X1 U9116 ( .B1(n7898), .B2(n10817), .A(n7897), .ZN(P2_U3289) );
  AND2_X1 U9117 ( .A1(n8067), .A2(n7899), .ZN(n7902) );
  INV_X1 U9118 ( .A(n7900), .ZN(n7901) );
  OAI21_X1 U9119 ( .B1(n7905), .B2(n7904), .A(n7903), .ZN(n7906) );
  INV_X1 U9120 ( .A(n7906), .ZN(n8060) );
  NAND2_X1 U9121 ( .A1(n8022), .A2(n8076), .ZN(n9928) );
  INV_X1 U9122 ( .A(n8022), .ZN(n10103) );
  NAND2_X1 U9123 ( .A1(n10103), .A2(n10846), .ZN(n9933) );
  NOR2_X1 U9124 ( .A1(n10103), .A2(n8076), .ZN(n7907) );
  AOI21_X1 U9125 ( .B1(n8060), .B2(n10042), .A(n7907), .ZN(n7998) );
  NAND2_X1 U9126 ( .A1(n8066), .A2(n8009), .ZN(n9937) );
  NAND2_X1 U9127 ( .A1(n10102), .A2(n8009), .ZN(n7908) );
  NAND2_X1 U9128 ( .A1(n7909), .A2(n8125), .ZN(n9942) );
  INV_X1 U9129 ( .A(n8125), .ZN(n8037) );
  NAND2_X1 U9130 ( .A1(n8037), .A2(n10101), .ZN(n9941) );
  INV_X1 U9131 ( .A(n9940), .ZN(n10043) );
  OAI21_X1 U9132 ( .B1(n7910), .B2(n10043), .A(n8042), .ZN(n8123) );
  INV_X1 U9133 ( .A(n7857), .ZN(n10426) );
  NAND2_X1 U9134 ( .A1(n9930), .A2(n9922), .ZN(n9844) );
  INV_X1 U9135 ( .A(n9923), .ZN(n7911) );
  NAND2_X1 U9136 ( .A1(n9930), .A2(n7911), .ZN(n9884) );
  NAND2_X1 U9137 ( .A1(n9884), .A2(n9894), .ZN(n9848) );
  NOR2_X1 U9138 ( .A1(n9848), .A2(n10042), .ZN(n7912) );
  INV_X1 U9139 ( .A(n9928), .ZN(n9932) );
  NOR2_X1 U9140 ( .A1(n10044), .A2(n9932), .ZN(n7913) );
  NAND2_X1 U9141 ( .A1(n8064), .A2(n7913), .ZN(n7914) );
  INV_X1 U9142 ( .A(n10930), .ZN(n10554) );
  AOI21_X1 U9143 ( .B1(n8047), .B2(n7915), .A(n10554), .ZN(n7917) );
  OAI22_X1 U9144 ( .A1(n8160), .A2(n10925), .B1(n8066), .B2(n10927), .ZN(n7916) );
  AOI211_X1 U9145 ( .C1(n8123), .C2(n10426), .A(n7917), .B(n7916), .ZN(n8128)
         );
  NOR2_X2 U9146 ( .A1(n8006), .A2(n8125), .ZN(n8053) );
  AOI21_X1 U9147 ( .B1(n8125), .B2(n8006), .A(n8053), .ZN(n8126) );
  NOR2_X1 U9148 ( .A1(n11012), .A2(n8037), .ZN(n7920) );
  OAI22_X1 U9149 ( .A1(n11019), .A2(n7918), .B1(n8033), .B2(n11014), .ZN(n7919) );
  AOI211_X1 U9150 ( .C1(n8126), .C2(n10470), .A(n7920), .B(n7919), .ZN(n7923)
         );
  NAND2_X1 U9151 ( .A1(n8123), .A2(n10433), .ZN(n7922) );
  OAI211_X1 U9152 ( .C1(n8128), .C2(n10789), .A(n7923), .B(n7922), .ZN(
        P1_U3282) );
  AOI21_X1 U9153 ( .B1(n5849), .B2(n7925), .A(n7924), .ZN(n7927) );
  AOI22_X1 U9154 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8221), .B1(n8215), .B2(
        n5864), .ZN(n7926) );
  NOR2_X1 U9155 ( .A1(n7927), .A2(n7926), .ZN(n8220) );
  AOI21_X1 U9156 ( .B1(n7927), .B2(n7926), .A(n8220), .ZN(n7939) );
  NOR2_X1 U9157 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8215), .ZN(n7928) );
  AOI21_X1 U9158 ( .B1(n8215), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7928), .ZN(
        n7932) );
  OAI21_X1 U9159 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7930), .A(n7929), .ZN(
        n7931) );
  NAND2_X1 U9160 ( .A1(n7932), .A2(n7931), .ZN(n8214) );
  OAI21_X1 U9161 ( .B1(n7932), .B2(n7931), .A(n8214), .ZN(n7937) );
  INV_X1 U9162 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U9163 ( .A1(n8959), .A2(n8215), .ZN(n7933) );
  NAND2_X1 U9164 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8732) );
  OAI211_X1 U9165 ( .C1(n7934), .C2(n8929), .A(n7933), .B(n8732), .ZN(n7935)
         );
  AOI21_X1 U9166 ( .B1(n7937), .B2(n7936), .A(n7935), .ZN(n7938) );
  OAI21_X1 U9167 ( .B1(n7939), .B2(n8957), .A(n7938), .ZN(P2_U3259) );
  INV_X1 U9168 ( .A(n7940), .ZN(n7944) );
  AOI21_X1 U9169 ( .B1(n7942), .B2(n7941), .A(n7956), .ZN(n7943) );
  OAI21_X1 U9170 ( .B1(n7944), .B2(n7943), .A(n10798), .ZN(n7947) );
  NAND2_X1 U9171 ( .A1(n8894), .A2(n8837), .ZN(n7946) );
  NAND2_X1 U9172 ( .A1(n8896), .A2(n9137), .ZN(n7945) );
  AND2_X1 U9173 ( .A1(n7946), .A2(n7945), .ZN(n8142) );
  NAND2_X1 U9174 ( .A1(n7947), .A2(n8142), .ZN(n10875) );
  INV_X1 U9175 ( .A(n10875), .ZN(n7960) );
  OAI22_X1 U9176 ( .A1(n10815), .A2(n7948), .B1(n8146), .B2(n10809), .ZN(n7952) );
  AOI21_X1 U9177 ( .B1(n7949), .B2(n10868), .A(n11000), .ZN(n7950) );
  AND2_X1 U9178 ( .A1(n10815), .A2(n9004), .ZN(n9025) );
  INV_X1 U9179 ( .A(n9025), .ZN(n9119) );
  NOR2_X1 U9180 ( .A1(n10871), .A2(n9119), .ZN(n7951) );
  AOI211_X1 U9181 ( .C1(n9122), .C2(n10868), .A(n7952), .B(n7951), .ZN(n7959)
         );
  INV_X1 U9182 ( .A(n8896), .ZN(n7953) );
  NAND2_X1 U9183 ( .A1(n7953), .A2(n10853), .ZN(n7954) );
  NAND2_X1 U9184 ( .A1(n7955), .A2(n7954), .ZN(n7957) );
  OR2_X2 U9185 ( .A1(n7957), .A2(n7956), .ZN(n10870) );
  NAND2_X1 U9186 ( .A1(n7957), .A2(n7956), .ZN(n10869) );
  NAND3_X1 U9187 ( .A1(n10870), .A2(n9114), .A3(n10869), .ZN(n7958) );
  OAI211_X1 U9188 ( .C1(n7960), .C2(n10817), .A(n7959), .B(n7958), .ZN(
        P2_U3288) );
  INV_X1 U9189 ( .A(n7961), .ZN(n8149) );
  AOI211_X1 U9190 ( .C1(n7963), .C2(n7962), .A(n8882), .B(n8149), .ZN(n7969)
         );
  NAND2_X1 U9191 ( .A1(n10731), .A2(n8897), .ZN(n7965) );
  OAI211_X1 U9192 ( .C1(n8094), .C2(n10736), .A(n7965), .B(n7964), .ZN(n7968)
         );
  OAI22_X1 U9193 ( .A1(n8856), .A2(n10853), .B1(n7966), .B2(n10742), .ZN(n7967) );
  OR3_X1 U9194 ( .A1(n7969), .A2(n7968), .A3(n7967), .ZN(P2_U3215) );
  XNOR2_X1 U9195 ( .A(n10039), .B(n7970), .ZN(n10699) );
  OAI21_X1 U9196 ( .B1(n7972), .B2(n10039), .A(n7971), .ZN(n7975) );
  OAI22_X1 U9197 ( .A1(n7973), .A2(n10927), .B1(n7831), .B2(n10925), .ZN(n7974) );
  AOI21_X1 U9198 ( .B1(n7975), .B2(n10930), .A(n7974), .ZN(n7976) );
  OAI21_X1 U9199 ( .B1(n10699), .B2(n7857), .A(n7976), .ZN(n10701) );
  OAI211_X1 U9200 ( .C1(n9836), .C2(n9835), .A(n11033), .B(n7990), .ZN(n10698)
         );
  OAI22_X1 U9201 ( .A1(n10698), .A2(n10785), .B1(n6444), .B2(n11014), .ZN(
        n7977) );
  NOR2_X1 U9202 ( .A1(n10701), .A2(n7977), .ZN(n7978) );
  MUX2_X1 U9203 ( .A(n7979), .B(n7978), .S(n11019), .Z(n7983) );
  INV_X1 U9204 ( .A(n10699), .ZN(n7981) );
  AOI22_X1 U9205 ( .A1(n7981), .A2(n10433), .B1(n10413), .B2(n7980), .ZN(n7982) );
  NAND2_X1 U9206 ( .A1(n7983), .A2(n7982), .ZN(P1_U3290) );
  XNOR2_X1 U9207 ( .A(n10037), .B(n7984), .ZN(n10709) );
  INV_X1 U9208 ( .A(n10709), .ZN(n7997) );
  INV_X1 U9209 ( .A(n9843), .ZN(n7987) );
  INV_X1 U9210 ( .A(n7985), .ZN(n7986) );
  AOI21_X1 U9211 ( .B1(n7987), .B2(n10037), .A(n7986), .ZN(n7988) );
  OAI222_X1 U9212 ( .A1(n10925), .A2(n6507), .B1(n10927), .B2(n7847), .C1(
        n10554), .C2(n7988), .ZN(n10707) );
  NAND2_X1 U9213 ( .A1(n10707), .A2(n11019), .ZN(n7996) );
  OAI22_X1 U9214 ( .A1(n11019), .A2(n7989), .B1(n10134), .B2(n11014), .ZN(
        n7993) );
  INV_X1 U9215 ( .A(n10470), .ZN(n8588) );
  AND2_X1 U9216 ( .A1(n7990), .A2(n7994), .ZN(n7991) );
  OR2_X1 U9217 ( .A1(n7991), .A2(n8114), .ZN(n10706) );
  NOR2_X1 U9218 ( .A1(n8588), .A2(n10706), .ZN(n7992) );
  AOI211_X1 U9219 ( .C1(n10413), .C2(n7994), .A(n7993), .B(n7992), .ZN(n7995)
         );
  OAI211_X1 U9220 ( .C1(n11021), .C2(n7997), .A(n7996), .B(n7995), .ZN(
        P1_U3289) );
  OR2_X1 U9221 ( .A1(n7998), .A2(n10044), .ZN(n7999) );
  NAND2_X1 U9222 ( .A1(n8000), .A2(n7999), .ZN(n10860) );
  INV_X1 U9223 ( .A(n10433), .ZN(n10938) );
  AOI22_X1 U9224 ( .A1(n10768), .A2(n10103), .B1(n10101), .B2(n10769), .ZN(
        n8004) );
  NAND2_X1 U9225 ( .A1(n8064), .A2(n9928), .ZN(n8001) );
  XOR2_X1 U9226 ( .A(n10044), .B(n8001), .Z(n8002) );
  NAND2_X1 U9227 ( .A1(n8002), .A2(n10930), .ZN(n8003) );
  OAI211_X1 U9228 ( .C1(n10860), .C2(n7857), .A(n8004), .B(n8003), .ZN(n10863)
         );
  NAND2_X1 U9229 ( .A1(n10863), .A2(n11019), .ZN(n8011) );
  OAI22_X1 U9230 ( .A1(n11019), .A2(n6586), .B1(n8021), .B2(n11014), .ZN(n8008) );
  NAND2_X1 U9231 ( .A1(n8071), .A2(n8009), .ZN(n8005) );
  NAND2_X1 U9232 ( .A1(n8006), .A2(n8005), .ZN(n10862) );
  NOR2_X1 U9233 ( .A1(n10862), .A2(n8588), .ZN(n8007) );
  AOI211_X1 U9234 ( .C1(n10413), .C2(n8009), .A(n8008), .B(n8007), .ZN(n8010)
         );
  OAI211_X1 U9235 ( .C1(n10860), .C2(n10938), .A(n8011), .B(n8010), .ZN(
        P1_U3283) );
  INV_X1 U9236 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10119) );
  INV_X1 U9237 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8012) );
  OAI22_X1 U9238 ( .A1(n11019), .A2(n10119), .B1(n8012), .B2(n11014), .ZN(
        n8013) );
  INV_X1 U9239 ( .A(n8013), .ZN(n8016) );
  OAI21_X1 U9240 ( .B1(n10470), .B2(n10413), .A(n8014), .ZN(n8015) );
  OAI211_X1 U9241 ( .C1(n8017), .C2(n10789), .A(n8016), .B(n8015), .ZN(
        P1_U3291) );
  NAND2_X1 U9242 ( .A1(n5098), .A2(n8029), .ZN(n8019) );
  XNOR2_X1 U9243 ( .A(n8019), .B(n8018), .ZN(n8020) );
  NAND2_X1 U9244 ( .A1(n8020), .A2(n9756), .ZN(n8026) );
  OAI22_X1 U9245 ( .A1(n9800), .A2(n8022), .B1(n9799), .B2(n8021), .ZN(n8023)
         );
  AOI211_X1 U9246 ( .C1(n8454), .C2(n10101), .A(n8024), .B(n8023), .ZN(n8025)
         );
  OAI211_X1 U9247 ( .C1(n10861), .C2(n9753), .A(n8026), .B(n8025), .ZN(
        P1_U3219) );
  INV_X1 U9248 ( .A(n8027), .ZN(n8032) );
  AOI21_X1 U9249 ( .B1(n8030), .B2(n8029), .A(n8028), .ZN(n8031) );
  OAI21_X1 U9250 ( .B1(n8032), .B2(n8031), .A(n9756), .ZN(n8036) );
  INV_X1 U9251 ( .A(n8160), .ZN(n10100) );
  AND2_X1 U9252 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10172) );
  OAI22_X1 U9253 ( .A1(n9800), .A2(n8066), .B1(n9799), .B2(n8033), .ZN(n8034)
         );
  AOI211_X1 U9254 ( .C1(n8454), .C2(n10100), .A(n10172), .B(n8034), .ZN(n8035)
         );
  OAI211_X1 U9255 ( .C1(n8037), .C2(n9753), .A(n8036), .B(n8035), .ZN(P1_U3229) );
  INV_X1 U9256 ( .A(n8038), .ZN(n8040) );
  OAI222_X1 U9257 ( .A1(P1_U3084), .A2(n8124), .B1(n10596), .B2(n8040), .C1(
        n9588), .C2(n8813), .ZN(P1_U3331) );
  OAI222_X1 U9258 ( .A1(n9696), .A2(n8041), .B1(n8593), .B2(n8040), .C1(n8039), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U9259 ( .A1(n8043), .A2(n8125), .ZN(n8044) );
  OR2_X1 U9260 ( .A1(n8160), .A2(n8155), .ZN(n9945) );
  NAND2_X1 U9261 ( .A1(n8155), .A2(n8160), .ZN(n9944) );
  NAND2_X1 U9262 ( .A1(n8045), .A2(n10047), .ZN(n8046) );
  NAND2_X1 U9263 ( .A1(n8157), .A2(n8046), .ZN(n10890) );
  OAI21_X1 U9264 ( .B1(n10047), .B2(n8048), .A(n8158), .ZN(n8049) );
  NAND2_X1 U9265 ( .A1(n8049), .A2(n10930), .ZN(n8051) );
  AOI22_X1 U9266 ( .A1(n10101), .A2(n10768), .B1(n10769), .B2(n10099), .ZN(
        n8050) );
  NAND2_X1 U9267 ( .A1(n8051), .A2(n8050), .ZN(n8052) );
  AOI21_X1 U9268 ( .B1(n10890), .B2(n10426), .A(n8052), .ZN(n10892) );
  INV_X1 U9269 ( .A(n8155), .ZN(n10888) );
  OAI21_X1 U9270 ( .B1(n8053), .B2(n10888), .A(n11033), .ZN(n8054) );
  OR2_X1 U9271 ( .A1(n8054), .A2(n8163), .ZN(n10887) );
  INV_X1 U9272 ( .A(n11023), .ZN(n10937) );
  OAI22_X1 U9273 ( .A1(n11019), .A2(n8055), .B1(n8235), .B2(n11014), .ZN(n8056) );
  AOI21_X1 U9274 ( .B1(n10413), .B2(n8155), .A(n8056), .ZN(n8057) );
  OAI21_X1 U9275 ( .B1(n10887), .B2(n10937), .A(n8057), .ZN(n8058) );
  AOI21_X1 U9276 ( .B1(n10890), .B2(n10433), .A(n8058), .ZN(n8059) );
  OAI21_X1 U9277 ( .B1(n10892), .B2(n10789), .A(n8059), .ZN(P1_U3281) );
  XNOR2_X1 U9278 ( .A(n8060), .B(n10042), .ZN(n10848) );
  INV_X1 U9279 ( .A(n9848), .ZN(n8061) );
  NAND2_X1 U9280 ( .A1(n8062), .A2(n8061), .ZN(n8063) );
  NAND2_X1 U9281 ( .A1(n8063), .A2(n10042), .ZN(n8065) );
  AOI21_X1 U9282 ( .B1(n8065), .B2(n8064), .A(n10554), .ZN(n8069) );
  OAI22_X1 U9283 ( .A1(n8067), .A2(n10927), .B1(n8066), .B2(n10925), .ZN(n8068) );
  OR2_X1 U9284 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  AOI21_X1 U9285 ( .B1(n10848), .B2(n10426), .A(n8070), .ZN(n10850) );
  OAI211_X1 U9286 ( .C1(n8072), .C2(n10846), .A(n11033), .B(n8071), .ZN(n10845) );
  OAI22_X1 U9287 ( .A1(n11019), .A2(n8074), .B1(n8073), .B2(n11014), .ZN(n8075) );
  AOI21_X1 U9288 ( .B1(n10413), .B2(n8076), .A(n8075), .ZN(n8077) );
  OAI21_X1 U9289 ( .B1(n10845), .B2(n10937), .A(n8077), .ZN(n8078) );
  AOI21_X1 U9290 ( .B1(n10848), .B2(n10433), .A(n8078), .ZN(n8079) );
  OAI21_X1 U9291 ( .B1(n10850), .B2(n10465), .A(n8079), .ZN(P1_U3284) );
  OAI21_X1 U9292 ( .B1(n9886), .B2(n8081), .A(n8080), .ZN(n8082) );
  XNOR2_X1 U9293 ( .A(n8082), .B(n10035), .ZN(n8084) );
  OAI22_X1 U9294 ( .A1(n6507), .A2(n10927), .B1(n8625), .B2(n10925), .ZN(n8083) );
  AOI21_X1 U9295 ( .B1(n8084), .B2(n10930), .A(n8083), .ZN(n10748) );
  NAND2_X1 U9296 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  XNOR2_X1 U9297 ( .A(n8087), .B(n10035), .ZN(n10746) );
  INV_X1 U9298 ( .A(n11021), .ZN(n10302) );
  NAND2_X1 U9299 ( .A1(n8116), .A2(n5207), .ZN(n8088) );
  NAND2_X1 U9300 ( .A1(n10760), .A2(n8088), .ZN(n10744) );
  AOI22_X1 U9301 ( .A1(n10465), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n8628), .B2(
        n10463), .ZN(n8090) );
  NAND2_X1 U9302 ( .A1(n10413), .A2(n5207), .ZN(n8089) );
  OAI211_X1 U9303 ( .C1(n10744), .C2(n8588), .A(n8090), .B(n8089), .ZN(n8091)
         );
  AOI21_X1 U9304 ( .B1(n10746), .B2(n10302), .A(n8091), .ZN(n8092) );
  OAI21_X1 U9305 ( .B1(n10748), .B2(n10465), .A(n8092), .ZN(P1_U3287) );
  NOR3_X1 U9306 ( .A1(n8769), .A2(n8094), .A3(n8093), .ZN(n8095) );
  AOI21_X1 U9307 ( .B1(n5096), .B2(n10727), .A(n8095), .ZN(n8105) );
  NOR2_X1 U9308 ( .A1(n8096), .A2(n8882), .ZN(n8103) );
  AND2_X1 U9309 ( .A1(n10733), .A2(n10879), .ZN(n8102) );
  NOR2_X1 U9310 ( .A1(n10742), .A2(n8196), .ZN(n8101) );
  NAND2_X1 U9311 ( .A1(n10731), .A2(n8895), .ZN(n8098) );
  OAI211_X1 U9312 ( .C1(n8099), .C2(n10736), .A(n8098), .B(n8097), .ZN(n8100)
         );
  NOR4_X1 U9313 ( .A1(n8103), .A2(n8102), .A3(n8101), .A4(n8100), .ZN(n8104)
         );
  OAI21_X1 U9314 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(P2_U3233) );
  INV_X1 U9315 ( .A(n10036), .ZN(n8107) );
  XNOR2_X1 U9316 ( .A(n9886), .B(n8107), .ZN(n8108) );
  NAND2_X1 U9317 ( .A1(n8108), .A2(n10930), .ZN(n8113) );
  XNOR2_X1 U9318 ( .A(n8109), .B(n10036), .ZN(n10722) );
  NAND2_X1 U9319 ( .A1(n7834), .A2(n10769), .ZN(n8110) );
  OAI21_X1 U9320 ( .B1(n7831), .B2(n10927), .A(n8110), .ZN(n8111) );
  AOI21_X1 U9321 ( .B1(n10722), .B2(n10426), .A(n8111), .ZN(n8112) );
  AND2_X1 U9322 ( .A1(n8113), .A2(n8112), .ZN(n10724) );
  OR2_X1 U9323 ( .A1(n8114), .A2(n10719), .ZN(n8115) );
  NAND2_X1 U9324 ( .A1(n8116), .A2(n8115), .ZN(n10720) );
  AOI22_X1 U9325 ( .A1(n10465), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10463), .B2(
        n8117), .ZN(n8120) );
  NAND2_X1 U9326 ( .A1(n10413), .A2(n8118), .ZN(n8119) );
  OAI211_X1 U9327 ( .C1(n8588), .C2(n10720), .A(n8120), .B(n8119), .ZN(n8121)
         );
  AOI21_X1 U9328 ( .B1(n10722), .B2(n10433), .A(n8121), .ZN(n8122) );
  OAI21_X1 U9329 ( .B1(n10724), .B2(n10789), .A(n8122), .ZN(P1_U3288) );
  INV_X1 U9330 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8131) );
  INV_X1 U9331 ( .A(n8123), .ZN(n8129) );
  OR2_X1 U9332 ( .A1(n10024), .A2(n10076), .ZN(n10718) );
  AOI22_X1 U9333 ( .A1(n8126), .A2(n11033), .B1(n10827), .B2(n8125), .ZN(n8127) );
  OAI211_X1 U9334 ( .C1(n8129), .C2(n10718), .A(n8128), .B(n8127), .ZN(n8132)
         );
  NAND2_X1 U9335 ( .A1(n8132), .A2(n11040), .ZN(n8130) );
  OAI21_X1 U9336 ( .B1(n11040), .B2(n8131), .A(n8130), .ZN(P1_U3481) );
  NAND2_X1 U9337 ( .A1(n8132), .A2(n11036), .ZN(n8133) );
  OAI21_X1 U9338 ( .B1(n11036), .B2(n6598), .A(n8133), .ZN(P1_U3532) );
  NAND2_X1 U9339 ( .A1(n8138), .A2(n8134), .ZN(n8136) );
  NOR2_X1 U9340 ( .A1(n8135), .A2(P1_U3084), .ZN(n10080) );
  INV_X1 U9341 ( .A(n10080), .ZN(n10085) );
  OAI211_X1 U9342 ( .C1(n9367), .C2(n8813), .A(n8136), .B(n10085), .ZN(
        P1_U3330) );
  NAND2_X1 U9343 ( .A1(n8138), .A2(n8137), .ZN(n8140) );
  OAI211_X1 U9344 ( .C1(n8141), .C2(n9696), .A(n8140), .B(n8139), .ZN(P2_U3335) );
  INV_X1 U9345 ( .A(n8142), .ZN(n8143) );
  NAND2_X1 U9346 ( .A1(n8143), .A2(n8840), .ZN(n8145) );
  OAI211_X1 U9347 ( .C1(n10742), .C2(n8146), .A(n8145), .B(n8144), .ZN(n8153)
         );
  NAND3_X1 U9348 ( .A1(n8845), .A2(n8147), .A3(n8896), .ZN(n8151) );
  OAI21_X1 U9349 ( .B1(n8149), .B2(n8148), .A(n10727), .ZN(n8150) );
  AOI21_X1 U9350 ( .B1(n8151), .B2(n8150), .A(n5096), .ZN(n8152) );
  AOI211_X1 U9351 ( .C1(n10733), .C2(n10868), .A(n8153), .B(n8152), .ZN(n8154)
         );
  INV_X1 U9352 ( .A(n8154), .ZN(P2_U3223) );
  OR2_X1 U9353 ( .A1(n10100), .A2(n8155), .ZN(n8156) );
  XNOR2_X1 U9354 ( .A(n10564), .B(n10099), .ZN(n10046) );
  XNOR2_X1 U9355 ( .A(n8427), .B(n5179), .ZN(n10563) );
  NAND3_X1 U9356 ( .A1(n8158), .A2(n5179), .A3(n9944), .ZN(n8159) );
  AOI21_X1 U9357 ( .B1(n10922), .B2(n8159), .A(n10554), .ZN(n8162) );
  OAI22_X1 U9358 ( .A1(n8428), .A2(n10925), .B1(n8160), .B2(n10927), .ZN(n8161) );
  AOI211_X1 U9359 ( .C1(n10563), .C2(n10426), .A(n8162), .B(n8161), .ZN(n10567) );
  INV_X1 U9360 ( .A(n10564), .ZN(n8168) );
  OR2_X1 U9361 ( .A1(n8163), .A2(n8168), .ZN(n8164) );
  AND2_X1 U9362 ( .A1(n10918), .A2(n8164), .ZN(n10565) );
  NAND2_X1 U9363 ( .A1(n10565), .A2(n10470), .ZN(n8167) );
  INV_X1 U9364 ( .A(n8209), .ZN(n8165) );
  AOI22_X1 U9365 ( .A1(n10465), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8165), .B2(
        n10463), .ZN(n8166) );
  OAI211_X1 U9366 ( .C1(n8168), .C2(n11012), .A(n8167), .B(n8166), .ZN(n8169)
         );
  AOI21_X1 U9367 ( .B1(n10563), .B2(n10433), .A(n8169), .ZN(n8170) );
  OAI21_X1 U9368 ( .B1(n10567), .B2(n10465), .A(n8170), .ZN(P1_U3280) );
  MUX2_X1 U9369 ( .A(n8171), .B(P1_REG1_REG_14__SCAN_IN), .S(n10189), .Z(n8175) );
  INV_X1 U9370 ( .A(n8179), .ZN(n8173) );
  AOI21_X1 U9371 ( .B1(n8173), .B2(n7863), .A(n8172), .ZN(n8174) );
  NOR2_X1 U9372 ( .A1(n8174), .A2(n8175), .ZN(n10181) );
  AOI21_X1 U9373 ( .B1(n8175), .B2(n8174), .A(n10181), .ZN(n8186) );
  INV_X1 U9374 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n8177) );
  AND2_X1 U9375 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8453) );
  INV_X1 U9376 ( .A(n8453), .ZN(n8176) );
  OAI21_X1 U9377 ( .B1(n10679), .B2(n8177), .A(n8176), .ZN(n8184) );
  NAND2_X1 U9378 ( .A1(n10189), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8180) );
  OAI21_X1 U9379 ( .B1(n10189), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8180), .ZN(
        n8181) );
  NOR2_X1 U9380 ( .A1(n8182), .A2(n8181), .ZN(n10188) );
  AOI211_X1 U9381 ( .C1(n8182), .C2(n8181), .A(n10188), .B(n10657), .ZN(n8183)
         );
  AOI211_X1 U9382 ( .C1(n10672), .C2(n10189), .A(n8184), .B(n8183), .ZN(n8185)
         );
  OAI21_X1 U9383 ( .B1(n8186), .B2(n10264), .A(n8185), .ZN(P1_U3255) );
  AND2_X1 U9384 ( .A1(n8190), .A2(n8187), .ZN(n8260) );
  NAND2_X1 U9385 ( .A1(n10870), .A2(n8260), .ZN(n8239) );
  INV_X1 U9386 ( .A(n8239), .ZN(n8189) );
  AOI21_X1 U9387 ( .B1(n10870), .B2(n8187), .A(n8190), .ZN(n8188) );
  NOR2_X1 U9388 ( .A1(n8189), .A2(n8188), .ZN(n10878) );
  AOI22_X1 U9389 ( .A1(n9137), .A2(n8895), .B1(n8893), .B2(n8837), .ZN(n8195)
         );
  INV_X1 U9390 ( .A(n8191), .ZN(n8193) );
  OAI211_X1 U9391 ( .C1(n8193), .C2(n8192), .A(n10798), .B(n8273), .ZN(n8194)
         );
  OAI211_X1 U9392 ( .C1(n10878), .C2(n8247), .A(n8195), .B(n8194), .ZN(n10882)
         );
  NAND2_X1 U9393 ( .A1(n10882), .A2(n10815), .ZN(n8203) );
  OAI22_X1 U9394 ( .A1(n10815), .A2(n8197), .B1(n8196), .B2(n10809), .ZN(n8201) );
  AND2_X1 U9395 ( .A1(n8198), .A2(n10879), .ZN(n8199) );
  OR2_X1 U9396 ( .A1(n8199), .A2(n8250), .ZN(n10881) );
  NOR2_X1 U9397 ( .A1(n10881), .A2(n8667), .ZN(n8200) );
  AOI211_X1 U9398 ( .C1(n9122), .C2(n10879), .A(n8201), .B(n8200), .ZN(n8202)
         );
  OAI211_X1 U9399 ( .C1(n10878), .C2(n8256), .A(n8203), .B(n8202), .ZN(
        P2_U3287) );
  INV_X1 U9400 ( .A(n8204), .ZN(n8227) );
  OAI222_X1 U9401 ( .A1(n8593), .A2(n8227), .B1(n8206), .B2(P2_U3152), .C1(
        n8205), .C2(n9696), .ZN(P2_U3334) );
  XNOR2_X1 U9402 ( .A(n8207), .B(n8208), .ZN(n8213) );
  AND2_X1 U9403 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10674) );
  OAI22_X1 U9404 ( .A1(n9798), .A2(n8428), .B1(n9799), .B2(n8209), .ZN(n8210)
         );
  AOI211_X1 U9405 ( .C1(n9750), .C2(n10100), .A(n10674), .B(n8210), .ZN(n8212)
         );
  NAND2_X1 U9406 ( .A1(n10564), .A2(n9803), .ZN(n8211) );
  OAI211_X1 U9407 ( .C1(n8213), .C2(n9805), .A(n8212), .B(n8211), .ZN(P1_U3234) );
  OAI21_X1 U9408 ( .B1(n8216), .B2(n8418), .A(n8402), .ZN(n8217) );
  INV_X1 U9409 ( .A(n8217), .ZN(n8225) );
  INV_X1 U9410 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8218) );
  NAND2_X1 U9411 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8746) );
  OAI21_X1 U9412 ( .B1(n8929), .B2(n8218), .A(n8746), .ZN(n8219) );
  AOI21_X1 U9413 ( .B1(n8959), .B2(n8394), .A(n8219), .ZN(n8224) );
  AOI21_X1 U9414 ( .B1(n5864), .B2(n8221), .A(n8220), .ZN(n8393) );
  XNOR2_X1 U9415 ( .A(n8393), .B(n8401), .ZN(n8222) );
  NAND2_X1 U9416 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8222), .ZN(n8395) );
  OAI211_X1 U9417 ( .C1(n8222), .C2(P2_REG1_REG_15__SCAN_IN), .A(n8907), .B(
        n8395), .ZN(n8223) );
  OAI211_X1 U9418 ( .C1(n8225), .C2(n8961), .A(n8224), .B(n8223), .ZN(P2_U3260) );
  OAI222_X1 U9419 ( .A1(n8228), .A2(P1_U3084), .B1(n10596), .B2(n8227), .C1(
        n8226), .C2(n8813), .ZN(P1_U3329) );
  NAND2_X1 U9420 ( .A1(n8230), .A2(n8229), .ZN(n8232) );
  XNOR2_X1 U9421 ( .A(n8232), .B(n8231), .ZN(n8233) );
  NAND2_X1 U9422 ( .A1(n8233), .A2(n9756), .ZN(n8238) );
  NOR2_X1 U9423 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8234), .ZN(n10662) );
  INV_X1 U9424 ( .A(n10099), .ZN(n10928) );
  OAI22_X1 U9425 ( .A1(n9798), .A2(n10928), .B1(n9799), .B2(n8235), .ZN(n8236)
         );
  AOI211_X1 U9426 ( .C1(n9750), .C2(n10101), .A(n10662), .B(n8236), .ZN(n8237)
         );
  OAI211_X1 U9427 ( .C1(n10888), .C2(n9753), .A(n8238), .B(n8237), .ZN(
        P1_U3215) );
  OR2_X1 U9428 ( .A1(n8894), .A2(n10879), .ZN(n8265) );
  NAND2_X1 U9429 ( .A1(n8239), .A2(n8265), .ZN(n8240) );
  OR2_X1 U9430 ( .A1(n8240), .A2(n8264), .ZN(n8258) );
  NAND2_X1 U9431 ( .A1(n8240), .A2(n8264), .ZN(n8241) );
  NAND2_X1 U9432 ( .A1(n8258), .A2(n8241), .ZN(n10895) );
  AOI22_X1 U9433 ( .A1(n9139), .A2(n8892), .B1(n8894), .B2(n9137), .ZN(n8246)
         );
  NAND2_X1 U9434 ( .A1(n8273), .A2(n8242), .ZN(n8244) );
  NAND2_X1 U9435 ( .A1(n8244), .A2(n8264), .ZN(n8243) );
  OAI211_X1 U9436 ( .C1(n8244), .C2(n8264), .A(n8243), .B(n10798), .ZN(n8245)
         );
  OAI211_X1 U9437 ( .C1(n10895), .C2(n8247), .A(n8246), .B(n8245), .ZN(n10898)
         );
  NAND2_X1 U9438 ( .A1(n10898), .A2(n8422), .ZN(n8255) );
  OAI22_X1 U9439 ( .A1(n10815), .A2(n8249), .B1(n8248), .B2(n10809), .ZN(n8253) );
  INV_X1 U9440 ( .A(n8257), .ZN(n10896) );
  OR2_X1 U9441 ( .A1(n8250), .A2(n10896), .ZN(n8251) );
  NAND2_X1 U9442 ( .A1(n8280), .A2(n8251), .ZN(n10897) );
  NOR2_X1 U9443 ( .A1(n10897), .A2(n8667), .ZN(n8252) );
  AOI211_X1 U9444 ( .C1(n9122), .C2(n8257), .A(n8253), .B(n8252), .ZN(n8254)
         );
  OAI211_X1 U9445 ( .C1(n10895), .C2(n8256), .A(n8255), .B(n8254), .ZN(
        P2_U3286) );
  NAND2_X1 U9446 ( .A1(n8257), .A2(n8893), .ZN(n8259) );
  NAND2_X1 U9447 ( .A1(n8258), .A2(n8259), .ZN(n8271) );
  INV_X1 U9448 ( .A(n8276), .ZN(n8263) );
  OR2_X1 U9449 ( .A1(n8263), .A2(n8259), .ZN(n8262) );
  AND2_X1 U9450 ( .A1(n8260), .A2(n8262), .ZN(n8261) );
  NAND2_X1 U9451 ( .A1(n10870), .A2(n8261), .ZN(n8270) );
  INV_X1 U9452 ( .A(n8262), .ZN(n8268) );
  NOR2_X1 U9453 ( .A1(n8264), .A2(n8263), .ZN(n8266) );
  AND2_X1 U9454 ( .A1(n8266), .A2(n8265), .ZN(n8267) );
  OAI21_X1 U9455 ( .B1(n8271), .B2(n8276), .A(n8319), .ZN(n10908) );
  NAND2_X1 U9456 ( .A1(n8273), .A2(n8272), .ZN(n8275) );
  AND2_X1 U9457 ( .A1(n8275), .A2(n8274), .ZN(n8613) );
  XNOR2_X1 U9458 ( .A(n8613), .B(n8276), .ZN(n8277) );
  NAND2_X1 U9459 ( .A1(n8277), .A2(n10798), .ZN(n8279) );
  AOI22_X1 U9460 ( .A1(n9139), .A2(n8891), .B1(n8893), .B2(n9137), .ZN(n8278)
         );
  NAND2_X1 U9461 ( .A1(n8279), .A2(n8278), .ZN(n10909) );
  AOI21_X1 U9462 ( .B1(n8280), .B2(n10905), .A(n11000), .ZN(n8281) );
  NAND2_X1 U9463 ( .A1(n8281), .A2(n8604), .ZN(n10906) );
  NOR2_X1 U9464 ( .A1(n10906), .A2(n10812), .ZN(n8282) );
  OAI21_X1 U9465 ( .B1(n10909), .B2(n8282), .A(n8422), .ZN(n8286) );
  OAI22_X1 U9466 ( .A1(n10815), .A2(n7660), .B1(n8283), .B2(n10809), .ZN(n8284) );
  AOI21_X1 U9467 ( .B1(n9122), .B2(n10905), .A(n8284), .ZN(n8285) );
  OAI211_X1 U9468 ( .C1(n9146), .C2(n10908), .A(n8286), .B(n8285), .ZN(
        P2_U3285) );
  NAND2_X1 U9469 ( .A1(n8289), .A2(n8288), .ZN(n8290) );
  XNOR2_X1 U9470 ( .A(n8287), .B(n8290), .ZN(n8291) );
  NAND2_X1 U9471 ( .A1(n8291), .A2(n9756), .ZN(n8295) );
  OAI22_X1 U9472 ( .A1(n9800), .A2(n10928), .B1(n9799), .B2(n10941), .ZN(n8292) );
  AOI211_X1 U9473 ( .C1(n8454), .C2(n10097), .A(n8293), .B(n8292), .ZN(n8294)
         );
  OAI211_X1 U9474 ( .C1(n5350), .C2(n9753), .A(n8295), .B(n8294), .ZN(P1_U3222) );
  NOR3_X1 U9475 ( .A1(n8296), .A2(n8320), .A3(n8769), .ZN(n8297) );
  AOI21_X1 U9476 ( .B1(n8298), .B2(n10727), .A(n8297), .ZN(n8306) );
  NAND2_X1 U9477 ( .A1(n8729), .A2(n8299), .ZN(n8700) );
  INV_X1 U9478 ( .A(n8700), .ZN(n8710) );
  INV_X1 U9479 ( .A(n8609), .ZN(n10949) );
  INV_X1 U9480 ( .A(n10736), .ZN(n8750) );
  NOR2_X1 U9481 ( .A1(n10742), .A2(n8602), .ZN(n8302) );
  OAI21_X1 U9482 ( .B1(n8748), .B2(n8320), .A(n8300), .ZN(n8301) );
  AOI211_X1 U9483 ( .C1(n8750), .C2(n8890), .A(n8302), .B(n8301), .ZN(n8303)
         );
  OAI21_X1 U9484 ( .B1(n10949), .B2(n8856), .A(n8303), .ZN(n8304) );
  AOI21_X1 U9485 ( .B1(n8710), .B2(n10727), .A(n8304), .ZN(n8305) );
  OAI21_X1 U9486 ( .B1(n8307), .B2(n8306), .A(n8305), .ZN(P2_U3226) );
  INV_X1 U9487 ( .A(n8308), .ZN(n8311) );
  OAI222_X1 U9488 ( .A1(n9696), .A2(n8310), .B1(n8593), .B2(n8311), .C1(
        P2_U3152), .C2(n8309), .ZN(P2_U3333) );
  OAI222_X1 U9489 ( .A1(P1_U3084), .A2(n8312), .B1(n10596), .B2(n8311), .C1(
        n9361), .C2(n8813), .ZN(P1_U3328) );
  INV_X1 U9490 ( .A(n8387), .ZN(n8317) );
  AOI21_X1 U9491 ( .B1(n8315), .B2(n8314), .A(n8313), .ZN(n8316) );
  NOR2_X1 U9492 ( .A1(n8317), .A2(n8316), .ZN(n8318) );
  OAI222_X1 U9493 ( .A1(n9067), .A2(n8703), .B1(n8415), .B2(n8747), .C1(n9070), 
        .C2(n8318), .ZN(n10966) );
  INV_X1 U9494 ( .A(n10966), .ZN(n8329) );
  NOR2_X1 U9495 ( .A1(n8322), .A2(n8321), .ZN(n10963) );
  INV_X1 U9496 ( .A(n10963), .ZN(n8323) );
  NAND3_X1 U9497 ( .A1(n8323), .A2(n9114), .A3(n10968), .ZN(n8328) );
  OAI22_X1 U9498 ( .A1(n10815), .A2(n8324), .B1(n8706), .B2(n10809), .ZN(n8326) );
  OAI21_X1 U9499 ( .B1(n8605), .B2(n10964), .A(n8416), .ZN(n10965) );
  NOR2_X1 U9500 ( .A1(n10965), .A2(n8667), .ZN(n8325) );
  AOI211_X1 U9501 ( .C1(n9122), .C2(n8713), .A(n8326), .B(n8325), .ZN(n8327)
         );
  OAI211_X1 U9502 ( .C1(n8329), .C2(n10817), .A(n8328), .B(n8327), .ZN(
        P2_U3283) );
  XNOR2_X1 U9503 ( .A(n8331), .B(n8330), .ZN(n8332) );
  XNOR2_X1 U9504 ( .A(n8333), .B(n8332), .ZN(n8334) );
  NAND2_X1 U9505 ( .A1(n8334), .A2(n9756), .ZN(n8339) );
  OAI22_X1 U9506 ( .A1(n9800), .A2(n8428), .B1(n9799), .B2(n8437), .ZN(n8337)
         );
  OAI21_X1 U9507 ( .B1(n9798), .B2(n9830), .A(n8335), .ZN(n8336) );
  NOR2_X1 U9508 ( .A1(n8337), .A2(n8336), .ZN(n8338) );
  OAI211_X1 U9509 ( .C1(n5349), .C2(n9753), .A(n8339), .B(n8338), .ZN(P1_U3232) );
  NOR2_X1 U9510 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8376) );
  NOR2_X1 U9511 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8374) );
  NOR2_X1 U9512 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8372) );
  NOR2_X1 U9513 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8370) );
  NOR2_X1 U9514 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8368) );
  NOR2_X1 U9515 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8366) );
  NAND2_X1 U9516 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8364) );
  XOR2_X1 U9517 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10623) );
  NAND2_X1 U9518 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8362) );
  XOR2_X1 U9519 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10621) );
  NOR2_X1 U9520 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8346) );
  XNOR2_X1 U9521 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10612) );
  NAND2_X1 U9522 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8344) );
  XOR2_X1 U9523 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10610) );
  NAND2_X1 U9524 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8342) );
  XOR2_X1 U9525 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10608) );
  AOI21_X1 U9526 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10603) );
  NAND3_X1 U9527 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10605) );
  OAI21_X1 U9528 ( .B1(n10603), .B2(n8340), .A(n10605), .ZN(n10607) );
  NAND2_X1 U9529 ( .A1(n10608), .A2(n10607), .ZN(n8341) );
  NAND2_X1 U9530 ( .A1(n8342), .A2(n8341), .ZN(n10609) );
  NAND2_X1 U9531 ( .A1(n10610), .A2(n10609), .ZN(n8343) );
  NAND2_X1 U9532 ( .A1(n8344), .A2(n8343), .ZN(n10611) );
  NOR2_X1 U9533 ( .A1(n10612), .A2(n10611), .ZN(n8345) );
  NOR2_X1 U9534 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  NOR2_X1 U9535 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8347), .ZN(n10614) );
  AND2_X1 U9536 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8347), .ZN(n10613) );
  NOR2_X1 U9537 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10613), .ZN(n8348) );
  NOR2_X1 U9538 ( .A1(n10614), .A2(n8348), .ZN(n8349) );
  NAND2_X1 U9539 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n8349), .ZN(n8351) );
  XOR2_X1 U9540 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n8349), .Z(n10616) );
  NAND2_X1 U9541 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10616), .ZN(n8350) );
  NAND2_X1 U9542 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  NAND2_X1 U9543 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8352), .ZN(n8354) );
  XOR2_X1 U9544 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8352), .Z(n10617) );
  NAND2_X1 U9545 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10617), .ZN(n8353) );
  NAND2_X1 U9546 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  NAND2_X1 U9547 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8355), .ZN(n8357) );
  XOR2_X1 U9548 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n8355), .Z(n10618) );
  NAND2_X1 U9549 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10618), .ZN(n8356) );
  NAND2_X1 U9550 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  NAND2_X1 U9551 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n8358), .ZN(n8360) );
  XOR2_X1 U9552 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n8358), .Z(n10619) );
  NAND2_X1 U9553 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10619), .ZN(n8359) );
  NAND2_X1 U9554 ( .A1(n8360), .A2(n8359), .ZN(n10620) );
  NAND2_X1 U9555 ( .A1(n10621), .A2(n10620), .ZN(n8361) );
  NAND2_X1 U9556 ( .A1(n8362), .A2(n8361), .ZN(n10622) );
  NAND2_X1 U9557 ( .A1(n10623), .A2(n10622), .ZN(n8363) );
  NAND2_X1 U9558 ( .A1(n8364), .A2(n8363), .ZN(n10625) );
  XNOR2_X1 U9559 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10624) );
  NOR2_X1 U9560 ( .A1(n10625), .A2(n10624), .ZN(n8365) );
  NOR2_X1 U9561 ( .A1(n8366), .A2(n8365), .ZN(n10627) );
  XNOR2_X1 U9562 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10626) );
  NOR2_X1 U9563 ( .A1(n10627), .A2(n10626), .ZN(n8367) );
  NOR2_X1 U9564 ( .A1(n8368), .A2(n8367), .ZN(n10629) );
  XNOR2_X1 U9565 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10628) );
  NOR2_X1 U9566 ( .A1(n10629), .A2(n10628), .ZN(n8369) );
  NOR2_X1 U9567 ( .A1(n8370), .A2(n8369), .ZN(n10631) );
  XNOR2_X1 U9568 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10630) );
  NOR2_X1 U9569 ( .A1(n10631), .A2(n10630), .ZN(n8371) );
  NOR2_X1 U9570 ( .A1(n8372), .A2(n8371), .ZN(n10633) );
  XNOR2_X1 U9571 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10632) );
  NOR2_X1 U9572 ( .A1(n10633), .A2(n10632), .ZN(n8373) );
  NOR2_X1 U9573 ( .A1(n8374), .A2(n8373), .ZN(n10635) );
  XNOR2_X1 U9574 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10634) );
  NOR2_X1 U9575 ( .A1(n10635), .A2(n10634), .ZN(n8375) );
  NOR2_X1 U9576 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  AND2_X1 U9577 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8377), .ZN(n10636) );
  NOR2_X1 U9578 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10636), .ZN(n8378) );
  NOR2_X1 U9579 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8377), .ZN(n10637) );
  NOR2_X1 U9580 ( .A1(n8378), .A2(n10637), .ZN(n8380) );
  XNOR2_X1 U9581 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8379) );
  XNOR2_X1 U9582 ( .A(n8380), .B(n8379), .ZN(ADD_1071_U4) );
  AOI21_X1 U9583 ( .B1(n8382), .B2(n8381), .A(n5502), .ZN(n10980) );
  OAI22_X1 U9584 ( .A1(n10815), .A2(n8383), .B1(n8736), .B2(n10809), .ZN(n8385) );
  XNOR2_X1 U9585 ( .A(n8416), .B(n8744), .ZN(n10982) );
  NOR2_X1 U9586 ( .A1(n10982), .A2(n8667), .ZN(n8384) );
  AOI211_X1 U9587 ( .C1(n9122), .C2(n8744), .A(n8385), .B(n8384), .ZN(n8392)
         );
  NAND2_X1 U9588 ( .A1(n8387), .A2(n8386), .ZN(n8389) );
  XNOR2_X1 U9589 ( .A(n8389), .B(n8388), .ZN(n8390) );
  OAI222_X1 U9590 ( .A1(n9067), .A2(n8733), .B1(n8415), .B2(n8687), .C1(n8390), 
        .C2(n9070), .ZN(n10984) );
  NAND2_X1 U9591 ( .A1(n10984), .A2(n8422), .ZN(n8391) );
  OAI211_X1 U9592 ( .C1(n10980), .C2(n9146), .A(n8392), .B(n8391), .ZN(
        P2_U3282) );
  NAND2_X1 U9593 ( .A1(n8394), .A2(n8393), .ZN(n8396) );
  NAND2_X1 U9594 ( .A1(n8396), .A2(n8395), .ZN(n8398) );
  XNOR2_X1 U9595 ( .A(n8914), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8397) );
  NOR2_X1 U9596 ( .A1(n8398), .A2(n8397), .ZN(n8904) );
  AOI21_X1 U9597 ( .B1(n8398), .B2(n8397), .A(n8904), .ZN(n8410) );
  INV_X1 U9598 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U9599 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8686) );
  OAI21_X1 U9600 ( .B1(n8929), .B2(n8399), .A(n8686), .ZN(n8408) );
  NAND2_X1 U9601 ( .A1(n8401), .A2(n8400), .ZN(n8403) );
  NAND2_X1 U9602 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8914), .ZN(n8404) );
  OAI21_X1 U9603 ( .B1(n8914), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8404), .ZN(
        n8405) );
  NOR2_X1 U9604 ( .A1(n8406), .A2(n8405), .ZN(n8913) );
  AOI211_X1 U9605 ( .C1(n8406), .C2(n8405), .A(n8913), .B(n8961), .ZN(n8407)
         );
  AOI211_X1 U9606 ( .C1(n8959), .C2(n8914), .A(n8408), .B(n8407), .ZN(n8409)
         );
  OAI21_X1 U9607 ( .B1(n8410), .B2(n8957), .A(n8409), .ZN(P2_U3261) );
  INV_X1 U9608 ( .A(n8744), .ZN(n10981) );
  NAND2_X1 U9609 ( .A1(n10981), .A2(n8747), .ZN(n8411) );
  XNOR2_X1 U9610 ( .A(n8515), .B(n8514), .ZN(n11005) );
  INV_X1 U9611 ( .A(n11005), .ZN(n8424) );
  XNOR2_X1 U9612 ( .A(n8511), .B(n8510), .ZN(n8413) );
  OAI222_X1 U9613 ( .A1(n8415), .A2(n8414), .B1(n9067), .B2(n8747), .C1(n9070), 
        .C2(n8413), .ZN(n11003) );
  INV_X1 U9614 ( .A(n8760), .ZN(n10999) );
  OAI21_X1 U9615 ( .B1(n8417), .B2(n10999), .A(n8518), .ZN(n11001) );
  OAI22_X1 U9616 ( .A1(n10815), .A2(n8418), .B1(n8752), .B2(n10809), .ZN(n8419) );
  AOI21_X1 U9617 ( .B1(n8760), .B2(n9122), .A(n8419), .ZN(n8420) );
  OAI21_X1 U9618 ( .B1(n11001), .B2(n8667), .A(n8420), .ZN(n8421) );
  AOI21_X1 U9619 ( .B1(n11003), .B2(n8422), .A(n8421), .ZN(n8423) );
  OAI21_X1 U9620 ( .B1(n8424), .B2(n9146), .A(n8423), .ZN(P2_U3281) );
  NAND2_X1 U9621 ( .A1(n10564), .A2(n10099), .ZN(n8426) );
  NOR2_X1 U9622 ( .A1(n10564), .A2(n10099), .ZN(n8425) );
  NAND2_X1 U9623 ( .A1(n10917), .A2(n8428), .ZN(n9954) );
  NAND2_X1 U9624 ( .A1(n9952), .A2(n9954), .ZN(n10913) );
  NAND2_X1 U9625 ( .A1(n10917), .A2(n10098), .ZN(n8429) );
  OR2_X1 U9626 ( .A1(n8478), .A2(n10926), .ZN(n9953) );
  NAND2_X1 U9627 ( .A1(n8478), .A2(n10926), .ZN(n9832) );
  OAI21_X1 U9628 ( .B1(n5083), .B2(n10049), .A(n8488), .ZN(n10959) );
  INV_X1 U9629 ( .A(n10959), .ZN(n8444) );
  AND2_X1 U9630 ( .A1(n10564), .A2(n10928), .ZN(n9948) );
  NOR2_X1 U9631 ( .A1(n10913), .A2(n9948), .ZN(n8431) );
  INV_X1 U9632 ( .A(n8494), .ZN(n8432) );
  AOI21_X1 U9633 ( .B1(n10049), .B2(n8433), .A(n8432), .ZN(n8436) );
  NAND2_X1 U9634 ( .A1(n10959), .A2(n10426), .ZN(n8435) );
  AOI22_X1 U9635 ( .A1(n10768), .A2(n10098), .B1(n10096), .B2(n10769), .ZN(
        n8434) );
  OAI211_X1 U9636 ( .C1(n10554), .C2(n8436), .A(n8435), .B(n8434), .ZN(n10957)
         );
  NAND2_X1 U9637 ( .A1(n10957), .A2(n11019), .ZN(n8443) );
  OAI22_X1 U9638 ( .A1(n11019), .A2(n8438), .B1(n8437), .B2(n11014), .ZN(n8441) );
  NAND2_X1 U9639 ( .A1(n10919), .A2(n8478), .ZN(n8439) );
  NAND2_X1 U9640 ( .A1(n8473), .A2(n8439), .ZN(n10956) );
  NOR2_X1 U9641 ( .A1(n10956), .A2(n8588), .ZN(n8440) );
  AOI211_X1 U9642 ( .C1(n10413), .C2(n8478), .A(n8441), .B(n8440), .ZN(n8442)
         );
  OAI211_X1 U9643 ( .C1(n8444), .C2(n10938), .A(n8443), .B(n8442), .ZN(
        P1_U3278) );
  INV_X1 U9644 ( .A(n8445), .ZN(n8467) );
  OAI222_X1 U9645 ( .A1(n8593), .A2(n8467), .B1(n8447), .B2(P2_U3152), .C1(
        n8446), .C2(n9696), .ZN(P2_U3332) );
  XOR2_X1 U9646 ( .A(n8449), .B(n8448), .Z(n8450) );
  XNOR2_X1 U9647 ( .A(n8451), .B(n8450), .ZN(n8457) );
  OAI22_X1 U9648 ( .A1(n9800), .A2(n10926), .B1(n9799), .B2(n8471), .ZN(n8452)
         );
  AOI211_X1 U9649 ( .C1(n8454), .C2(n10095), .A(n8453), .B(n8452), .ZN(n8456)
         );
  NAND2_X1 U9650 ( .A1(n9831), .A2(n9803), .ZN(n8455) );
  OAI211_X1 U9651 ( .C1(n8457), .C2(n9805), .A(n8456), .B(n8455), .ZN(P1_U3213) );
  NAND2_X1 U9652 ( .A1(n7054), .A2(n8459), .ZN(n8460) );
  XNOR2_X1 U9653 ( .A(n8461), .B(n8460), .ZN(n8466) );
  NAND2_X1 U9654 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8910) );
  OAI21_X1 U9655 ( .B1(n10736), .B2(n8651), .A(n8910), .ZN(n8462) );
  AOI21_X1 U9656 ( .B1(n10731), .B2(n8887), .A(n8462), .ZN(n8463) );
  OAI21_X1 U9657 ( .B1(n8539), .B2(n10742), .A(n8463), .ZN(n8464) );
  AOI21_X1 U9658 ( .B1(n9223), .B2(n10733), .A(n8464), .ZN(n8465) );
  OAI21_X1 U9659 ( .B1(n8466), .B2(n8882), .A(n8465), .ZN(P2_U3230) );
  OAI222_X1 U9660 ( .A1(n8468), .A2(P1_U3084), .B1(n10596), .B2(n8467), .C1(
        n9580), .C2(n8813), .ZN(P1_U3327) );
  NAND2_X1 U9661 ( .A1(n8494), .A2(n9832), .ZN(n8469) );
  XOR2_X1 U9662 ( .A(n5078), .B(n8469), .Z(n8470) );
  AOI222_X1 U9663 ( .A1(n10097), .A2(n10768), .B1(n10095), .B2(n10769), .C1(
        n10930), .C2(n8470), .ZN(n10973) );
  OAI22_X1 U9664 ( .A1(n11019), .A2(n8472), .B1(n8471), .B2(n11014), .ZN(n8477) );
  INV_X1 U9665 ( .A(n9831), .ZN(n10974) );
  INV_X1 U9666 ( .A(n8473), .ZN(n8475) );
  INV_X1 U9667 ( .A(n8500), .ZN(n8474) );
  OAI211_X1 U9668 ( .C1(n10974), .C2(n8475), .A(n8474), .B(n11033), .ZN(n10972) );
  NOR2_X1 U9669 ( .A1(n10972), .A2(n10937), .ZN(n8476) );
  AOI211_X1 U9670 ( .C1(n10413), .C2(n9831), .A(n8477), .B(n8476), .ZN(n8481)
         );
  OR2_X1 U9671 ( .A1(n8478), .A2(n10097), .ZN(n8482) );
  NAND2_X1 U9672 ( .A1(n8488), .A2(n8482), .ZN(n8479) );
  XNOR2_X1 U9673 ( .A(n8479), .B(n5078), .ZN(n10976) );
  NAND2_X1 U9674 ( .A1(n10976), .A2(n10302), .ZN(n8480) );
  OAI211_X1 U9675 ( .C1(n10973), .C2(n10465), .A(n8481), .B(n8480), .ZN(
        P1_U3277) );
  OR2_X1 U9676 ( .A1(n9831), .A2(n10096), .ZN(n8484) );
  AND2_X1 U9677 ( .A1(n8482), .A2(n8484), .ZN(n8487) );
  NAND2_X1 U9678 ( .A1(n8569), .A2(n10555), .ZN(n9970) );
  INV_X1 U9679 ( .A(n10052), .ZN(n8483) );
  AND2_X1 U9680 ( .A1(n8487), .A2(n8483), .ZN(n8486) );
  INV_X1 U9681 ( .A(n8484), .ZN(n8485) );
  NAND2_X1 U9682 ( .A1(n8488), .A2(n8487), .ZN(n8490) );
  AND2_X1 U9683 ( .A1(n8490), .A2(n8489), .ZN(n8491) );
  NAND2_X1 U9684 ( .A1(n8491), .A2(n10052), .ZN(n8492) );
  NAND2_X1 U9685 ( .A1(n8570), .A2(n8492), .ZN(n10988) );
  INV_X1 U9686 ( .A(n9832), .ZN(n9961) );
  NOR2_X1 U9687 ( .A1(n5078), .A2(n9961), .ZN(n8493) );
  OR2_X1 U9688 ( .A1(n9831), .A2(n9830), .ZN(n9962) );
  NAND2_X1 U9689 ( .A1(n8495), .A2(n9962), .ZN(n8573) );
  XOR2_X1 U9690 ( .A(n10052), .B(n8573), .Z(n8497) );
  OAI22_X1 U9691 ( .A1(n10453), .A2(n10925), .B1(n9830), .B2(n10927), .ZN(
        n8496) );
  AOI21_X1 U9692 ( .B1(n8497), .B2(n10930), .A(n8496), .ZN(n8498) );
  OAI21_X1 U9693 ( .B1(n10988), .B2(n7857), .A(n8498), .ZN(n10992) );
  NAND2_X1 U9694 ( .A1(n10992), .A2(n11019), .ZN(n8505) );
  OAI22_X1 U9695 ( .A1(n11019), .A2(n8499), .B1(n8554), .B2(n11014), .ZN(n8503) );
  INV_X1 U9696 ( .A(n8569), .ZN(n10989) );
  NAND2_X1 U9697 ( .A1(n8500), .A2(n10989), .ZN(n10558) );
  OR2_X1 U9698 ( .A1(n8500), .A2(n10989), .ZN(n8501) );
  NAND2_X1 U9699 ( .A1(n10558), .A2(n8501), .ZN(n10991) );
  NOR2_X1 U9700 ( .A1(n10991), .A2(n8588), .ZN(n8502) );
  AOI211_X1 U9701 ( .C1(n10413), .C2(n8569), .A(n8503), .B(n8502), .ZN(n8504)
         );
  OAI211_X1 U9702 ( .C1(n10988), .C2(n10938), .A(n8505), .B(n8504), .ZN(
        P1_U3276) );
  INV_X1 U9703 ( .A(n8506), .ZN(n8777) );
  OAI222_X1 U9704 ( .A1(P1_U3084), .A2(n8508), .B1(n10596), .B2(n8777), .C1(
        n8507), .C2(n8813), .ZN(P1_U3326) );
  OAI21_X1 U9705 ( .B1(n8511), .B2(n8510), .A(n8509), .ZN(n8512) );
  XOR2_X1 U9706 ( .A(n8517), .B(n8512), .Z(n8513) );
  AOI222_X1 U9707 ( .A1(n10798), .A2(n8513), .B1(n9138), .B2(n8837), .C1(n8888), .C2(n9137), .ZN(n9231) );
  AOI21_X1 U9708 ( .B1(n8517), .B2(n8516), .A(n5086), .ZN(n9227) );
  NAND2_X1 U9709 ( .A1(n9227), .A2(n9114), .ZN(n8524) );
  AOI211_X1 U9710 ( .C1(n9229), .C2(n8518), .A(n11000), .B(n5077), .ZN(n9228)
         );
  INV_X1 U9711 ( .A(n9229), .ZN(n8519) );
  NOR2_X1 U9712 ( .A1(n8519), .A2(n9133), .ZN(n8522) );
  OAI22_X1 U9713 ( .A1(n10815), .A2(n8520), .B1(n8690), .B2(n10809), .ZN(n8521) );
  AOI211_X1 U9714 ( .C1(n9228), .C2(n9025), .A(n8522), .B(n8521), .ZN(n8523)
         );
  OAI211_X1 U9715 ( .C1(n10817), .C2(n9231), .A(n8524), .B(n8523), .ZN(
        P2_U3280) );
  NOR2_X1 U9716 ( .A1(n5275), .A2(n8526), .ZN(n8527) );
  XNOR2_X1 U9717 ( .A(n8528), .B(n8527), .ZN(n8533) );
  NAND2_X1 U9718 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8927) );
  OAI21_X1 U9719 ( .B1(n10736), .B2(n8652), .A(n8927), .ZN(n8529) );
  AOI21_X1 U9720 ( .B1(n10731), .B2(n9138), .A(n8529), .ZN(n8530) );
  OAI21_X1 U9721 ( .B1(n9129), .B2(n10742), .A(n8530), .ZN(n8531) );
  AOI21_X1 U9722 ( .B1(n9216), .B2(n10733), .A(n8531), .ZN(n8532) );
  OAI21_X1 U9723 ( .B1(n8533), .B2(n8882), .A(n8532), .ZN(P2_U3240) );
  XOR2_X1 U9724 ( .A(n8536), .B(n8534), .Z(n8535) );
  AOI222_X1 U9725 ( .A1(n10798), .A2(n8535), .B1(n9109), .B2(n8837), .C1(n8887), .C2(n9137), .ZN(n9225) );
  OAI21_X1 U9726 ( .B1(n8537), .B2(n8536), .A(n8650), .ZN(n9221) );
  NAND2_X1 U9727 ( .A1(n9221), .A2(n9114), .ZN(n8544) );
  XNOR2_X1 U9728 ( .A(n5077), .B(n8595), .ZN(n8538) );
  NOR2_X1 U9729 ( .A1(n8538), .A2(n11000), .ZN(n9222) );
  NOR2_X1 U9730 ( .A1(n8595), .A2(n9133), .ZN(n8542) );
  OAI22_X1 U9731 ( .A1(n10815), .A2(n8540), .B1(n8539), .B2(n10809), .ZN(n8541) );
  AOI211_X1 U9732 ( .C1(n9222), .C2(n9025), .A(n8542), .B(n8541), .ZN(n8543)
         );
  OAI211_X1 U9733 ( .C1(n10817), .C2(n9225), .A(n8544), .B(n8543), .ZN(
        P2_U3279) );
  INV_X1 U9734 ( .A(n8545), .ZN(n8568) );
  OAI222_X1 U9735 ( .A1(n9696), .A2(n8546), .B1(n8593), .B2(n8568), .C1(
        P2_U3152), .C2(n6364), .ZN(P2_U3330) );
  XNOR2_X1 U9736 ( .A(n8548), .B(n8547), .ZN(n8550) );
  INV_X1 U9737 ( .A(n8551), .ZN(n8549) );
  NAND2_X1 U9738 ( .A1(n8550), .A2(n8549), .ZN(n8553) );
  INV_X1 U9739 ( .A(n9738), .ZN(n8552) );
  AOI22_X1 U9740 ( .A1(n8553), .A2(n9739), .B1(n8552), .B2(n8551), .ZN(n8558)
         );
  OAI22_X1 U9741 ( .A1(n9800), .A2(n9830), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10184), .ZN(n8556) );
  OAI22_X1 U9742 ( .A1(n9798), .A2(n10453), .B1(n9799), .B2(n8554), .ZN(n8555)
         );
  AOI211_X1 U9743 ( .C1(n8569), .C2(n9803), .A(n8556), .B(n8555), .ZN(n8557)
         );
  OAI21_X1 U9744 ( .B1(n8558), .B2(n9805), .A(n8557), .ZN(P1_U3239) );
  NAND2_X1 U9745 ( .A1(n5041), .A2(n8559), .ZN(n8560) );
  XNOR2_X1 U9746 ( .A(n8561), .B(n8560), .ZN(n8566) );
  NAND2_X1 U9747 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8955) );
  OAI21_X1 U9748 ( .B1(n10736), .B2(n8653), .A(n8955), .ZN(n8562) );
  AOI21_X1 U9749 ( .B1(n10731), .B2(n9109), .A(n8562), .ZN(n8563) );
  OAI21_X1 U9750 ( .B1(n9115), .B2(n10742), .A(n8563), .ZN(n8564) );
  AOI21_X1 U9751 ( .B1(n9211), .B2(n10733), .A(n8564), .ZN(n8565) );
  OAI21_X1 U9752 ( .B1(n8566), .B2(n8882), .A(n8565), .ZN(P2_U3221) );
  OAI222_X1 U9753 ( .A1(P1_U3084), .A2(n6952), .B1(n10596), .B2(n8568), .C1(
        n8567), .C2(n8813), .ZN(P1_U3325) );
  NAND2_X1 U9754 ( .A1(n10557), .A2(n10453), .ZN(n9973) );
  NAND2_X1 U9755 ( .A1(n9972), .A2(n9973), .ZN(n10549) );
  NAND2_X1 U9756 ( .A1(n10550), .A2(n10549), .ZN(n10548) );
  NAND2_X1 U9757 ( .A1(n10557), .A2(n10094), .ZN(n8571) );
  NAND2_X1 U9758 ( .A1(n10543), .A2(n10556), .ZN(n9975) );
  OR2_X1 U9759 ( .A1(n10538), .A2(n10454), .ZN(n9980) );
  NAND2_X1 U9760 ( .A1(n10538), .A2(n10454), .ZN(n9979) );
  NAND2_X1 U9761 ( .A1(n9980), .A2(n9979), .ZN(n10054) );
  INV_X1 U9762 ( .A(n10054), .ZN(n9978) );
  NAND2_X1 U9763 ( .A1(n5087), .A2(n9978), .ZN(n8572) );
  AND2_X1 U9764 ( .A1(n8778), .A2(n8572), .ZN(n10536) );
  NAND2_X1 U9765 ( .A1(n8573), .A2(n10052), .ZN(n8574) );
  NAND2_X1 U9766 ( .A1(n8574), .A2(n9969), .ZN(n10552) );
  INV_X1 U9767 ( .A(n10549), .ZN(n10551) );
  NAND2_X1 U9768 ( .A1(n10552), .A2(n10551), .ZN(n8575) );
  NAND2_X1 U9769 ( .A1(n10452), .A2(n10457), .ZN(n8579) );
  INV_X1 U9770 ( .A(n8579), .ZN(n8576) );
  INV_X1 U9771 ( .A(n9976), .ZN(n8577) );
  OAI21_X1 U9772 ( .B1(n8576), .B2(n8577), .A(n10054), .ZN(n8580) );
  NOR2_X1 U9773 ( .A1(n10054), .A2(n8577), .ZN(n8578) );
  NAND2_X1 U9774 ( .A1(n8579), .A2(n8578), .ZN(n8800) );
  AOI21_X1 U9775 ( .B1(n8580), .B2(n8800), .A(n10554), .ZN(n8582) );
  OAI22_X1 U9776 ( .A1(n9790), .A2(n10925), .B1(n10556), .B2(n10927), .ZN(
        n8581) );
  AOI211_X1 U9777 ( .C1(n10536), .C2(n10426), .A(n8582), .B(n8581), .ZN(n10541) );
  OR2_X2 U9778 ( .A1(n10558), .A2(n10557), .ZN(n10559) );
  INV_X1 U9779 ( .A(n10538), .ZN(n8583) );
  NOR2_X1 U9780 ( .A1(n10461), .A2(n8583), .ZN(n8584) );
  OR2_X1 U9781 ( .A1(n10437), .A2(n8584), .ZN(n10537) );
  INV_X1 U9782 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8585) );
  OAI22_X1 U9783 ( .A1(n11019), .A2(n8585), .B1(n9789), .B2(n11014), .ZN(n8586) );
  AOI21_X1 U9784 ( .B1(n10538), .B2(n10413), .A(n8586), .ZN(n8587) );
  OAI21_X1 U9785 ( .B1(n10537), .B2(n8588), .A(n8587), .ZN(n8589) );
  AOI21_X1 U9786 ( .B1(n10536), .B2(n10433), .A(n8589), .ZN(n8590) );
  OAI21_X1 U9787 ( .B1(n10541), .B2(n10789), .A(n8590), .ZN(P1_U3273) );
  INV_X1 U9788 ( .A(n8791), .ZN(n8727) );
  OAI222_X1 U9789 ( .A1(n8593), .A2(n8727), .B1(n5031), .B2(P2_U3152), .C1(
        n8591), .C2(n9696), .ZN(P2_U3329) );
  INV_X1 U9790 ( .A(n9211), .ZN(n9118) );
  NAND2_X1 U9791 ( .A1(n9127), .A2(n9118), .ZN(n9117) );
  INV_X1 U9792 ( .A(n9178), .ZN(n9017) );
  INV_X1 U9793 ( .A(n9167), .ZN(n8987) );
  XOR2_X1 U9794 ( .A(n9148), .B(n8963), .Z(n9150) );
  INV_X1 U9795 ( .A(P2_B_REG_SCAN_IN), .ZN(n8596) );
  OR2_X1 U9796 ( .A1(n6363), .A2(n8596), .ZN(n8597) );
  NAND2_X1 U9797 ( .A1(n9139), .A2(n8597), .ZN(n8666) );
  NOR2_X1 U9798 ( .A1(n8598), .A2(n8666), .ZN(n9147) );
  INV_X1 U9799 ( .A(n9147), .ZN(n9153) );
  NOR2_X1 U9800 ( .A1(n9153), .A2(n10817), .ZN(n8966) );
  AOI21_X1 U9801 ( .B1(n10817), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8966), .ZN(
        n8600) );
  NAND2_X1 U9802 ( .A1(n9148), .A2(n9122), .ZN(n8599) );
  OAI211_X1 U9803 ( .C1(n9150), .C2(n8667), .A(n8600), .B(n8599), .ZN(P2_U3265) );
  AOI21_X1 U9804 ( .B1(n8614), .B2(n8601), .A(n5082), .ZN(n10948) );
  OAI22_X1 U9805 ( .A1(n10815), .A2(n8603), .B1(n8602), .B2(n10809), .ZN(n8608) );
  INV_X1 U9806 ( .A(n8604), .ZN(n8606) );
  OAI21_X1 U9807 ( .B1(n10949), .B2(n8606), .A(n5336), .ZN(n10950) );
  NOR2_X1 U9808 ( .A1(n10950), .A2(n8667), .ZN(n8607) );
  AOI211_X1 U9809 ( .C1(n9122), .C2(n8609), .A(n8608), .B(n8607), .ZN(n8620)
         );
  INV_X1 U9810 ( .A(n8610), .ZN(n8612) );
  OAI21_X1 U9811 ( .B1(n8613), .B2(n8612), .A(n8611), .ZN(n8615) );
  XNOR2_X1 U9812 ( .A(n8615), .B(n8614), .ZN(n8616) );
  NAND2_X1 U9813 ( .A1(n8616), .A2(n10798), .ZN(n8618) );
  AOI22_X1 U9814 ( .A1(n9139), .A2(n8890), .B1(n8892), .B2(n9137), .ZN(n8617)
         );
  NAND2_X1 U9815 ( .A1(n8618), .A2(n8617), .ZN(n10952) );
  NAND2_X1 U9816 ( .A1(n10952), .A2(n10815), .ZN(n8619) );
  OAI211_X1 U9817 ( .C1(n10948), .C2(n9146), .A(n8620), .B(n8619), .ZN(
        P2_U3284) );
  NAND2_X1 U9818 ( .A1(n6544), .A2(n9756), .ZN(n8632) );
  AOI21_X1 U9819 ( .B1(n8623), .B2(n8622), .A(n8621), .ZN(n8631) );
  AOI22_X1 U9820 ( .A1(n9750), .A2(n10105), .B1(n9803), .B2(n5207), .ZN(n8630)
         );
  INV_X1 U9821 ( .A(n9799), .ZN(n8627) );
  INV_X1 U9822 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8624) );
  NOR2_X1 U9823 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8624), .ZN(n10163) );
  NOR2_X1 U9824 ( .A1(n9798), .A2(n8625), .ZN(n8626) );
  AOI211_X1 U9825 ( .C1(n8628), .C2(n8627), .A(n10163), .B(n8626), .ZN(n8629)
         );
  OAI211_X1 U9826 ( .C1(n8632), .C2(n8631), .A(n8630), .B(n8629), .ZN(P1_U3228) );
  OAI222_X1 U9827 ( .A1(n6947), .A2(P1_U3084), .B1(n10596), .B2(n8634), .C1(
        n8633), .C2(n8813), .ZN(P1_U3332) );
  NAND2_X1 U9828 ( .A1(n8845), .A2(n8901), .ZN(n8635) );
  OAI21_X1 U9829 ( .B1(n8882), .B2(n8636), .A(n8635), .ZN(n8640) );
  INV_X1 U9830 ( .A(n8637), .ZN(n8638) );
  NAND3_X1 U9831 ( .A1(n8640), .A2(n8639), .A3(n8638), .ZN(n8646) );
  AOI22_X1 U9832 ( .A1(n8750), .A2(n8900), .B1(n10731), .B2(n8901), .ZN(n8645)
         );
  NAND2_X1 U9833 ( .A1(n10733), .A2(n8641), .ZN(n8644) );
  NAND2_X1 U9834 ( .A1(n8642), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8643) );
  AND4_X1 U9835 ( .A1(n8646), .A2(n8645), .A3(n8644), .A4(n8643), .ZN(n8647)
         );
  OAI21_X1 U9836 ( .B1(n8648), .B2(n8882), .A(n8647), .ZN(P2_U3239) );
  INV_X1 U9837 ( .A(n9216), .ZN(n9134) );
  NAND2_X1 U9838 ( .A1(n9113), .A2(n9112), .ZN(n9209) );
  INV_X1 U9839 ( .A(n9204), .ZN(n9099) );
  INV_X1 U9840 ( .A(n9087), .ZN(n8654) );
  INV_X1 U9841 ( .A(n9194), .ZN(n9066) );
  AOI21_X2 U9842 ( .B1(n9062), .B2(n9072), .A(n8656), .ZN(n9050) );
  INV_X1 U9843 ( .A(n9173), .ZN(n8999) );
  XNOR2_X1 U9844 ( .A(n8662), .B(n8661), .ZN(n9155) );
  INV_X1 U9845 ( .A(n9155), .ZN(n8673) );
  XNOR2_X1 U9846 ( .A(n8663), .B(n8661), .ZN(n8664) );
  OAI222_X1 U9847 ( .A1(n9067), .A2(n8817), .B1(n8666), .B2(n8665), .C1(n8664), 
        .C2(n9070), .ZN(n9159) );
  OAI21_X1 U9848 ( .B1(n9156), .B2(n8971), .A(n8964), .ZN(n9157) );
  NOR2_X1 U9849 ( .A1(n9157), .A2(n8667), .ZN(n8671) );
  AOI22_X1 U9850 ( .A1(n8668), .A2(n9130), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10817), .ZN(n8669) );
  OAI21_X1 U9851 ( .B1(n9156), .B2(n9133), .A(n8669), .ZN(n8670) );
  AOI211_X1 U9852 ( .C1(n9159), .C2(n10815), .A(n8671), .B(n8670), .ZN(n8672)
         );
  OAI21_X1 U9853 ( .B1(n8673), .B2(n9146), .A(n8672), .ZN(P2_U3267) );
  OAI21_X1 U9854 ( .B1(n8748), .B2(n8680), .A(n8674), .ZN(n8677) );
  OAI22_X1 U9855 ( .A1(n8856), .A2(n10838), .B1(n8675), .B2(n10742), .ZN(n8676) );
  AOI211_X1 U9856 ( .C1(n8750), .C2(n8896), .A(n8677), .B(n8676), .ZN(n8684)
         );
  INV_X1 U9857 ( .A(n8678), .ZN(n8682) );
  OAI22_X1 U9858 ( .A1(n8769), .A2(n8680), .B1(n8882), .B2(n8679), .ZN(n8681)
         );
  NAND3_X1 U9859 ( .A1(n8775), .A2(n8682), .A3(n8681), .ZN(n8683) );
  OAI211_X1 U9860 ( .C1(n8685), .C2(n8882), .A(n8684), .B(n8683), .ZN(P2_U3241) );
  OAI21_X1 U9861 ( .B1(n8748), .B2(n8687), .A(n8686), .ZN(n8688) );
  AOI21_X1 U9862 ( .B1(n8750), .B2(n9138), .A(n8688), .ZN(n8689) );
  OAI21_X1 U9863 ( .B1(n8690), .B2(n10742), .A(n8689), .ZN(n8696) );
  INV_X1 U9864 ( .A(n8762), .ZN(n8694) );
  AOI22_X1 U9865 ( .A1(n8691), .A2(n10727), .B1(n8845), .B2(n8888), .ZN(n8692)
         );
  NOR3_X1 U9866 ( .A1(n8694), .A2(n8693), .A3(n8692), .ZN(n8695) );
  AOI211_X1 U9867 ( .C1(n10733), .C2(n9229), .A(n8696), .B(n8695), .ZN(n8697)
         );
  OAI21_X1 U9868 ( .B1(n8698), .B2(n8882), .A(n8697), .ZN(P2_U3228) );
  NAND2_X1 U9869 ( .A1(n8700), .A2(n8699), .ZN(n8701) );
  NAND2_X1 U9870 ( .A1(n8701), .A2(n8709), .ZN(n8737) );
  OAI21_X1 U9871 ( .B1(n8748), .B2(n8703), .A(n8702), .ZN(n8704) );
  AOI21_X1 U9872 ( .B1(n8750), .B2(n8889), .A(n8704), .ZN(n8705) );
  OAI21_X1 U9873 ( .B1(n8706), .B2(n10742), .A(n8705), .ZN(n8712) );
  AOI22_X1 U9874 ( .A1(n8707), .A2(n10727), .B1(n8845), .B2(n8891), .ZN(n8708)
         );
  NOR3_X1 U9875 ( .A1(n8710), .A2(n8709), .A3(n8708), .ZN(n8711) );
  AOI211_X1 U9876 ( .C1(n10733), .C2(n8713), .A(n8712), .B(n8711), .ZN(n8714)
         );
  OAI21_X1 U9877 ( .B1(n8737), .B2(n8882), .A(n8714), .ZN(P2_U3236) );
  NAND2_X1 U9878 ( .A1(n9054), .A2(n10904), .ZN(n9191) );
  INV_X1 U9879 ( .A(n9191), .ZN(n8722) );
  INV_X1 U9880 ( .A(n9055), .ZN(n8718) );
  NAND2_X1 U9881 ( .A1(n8886), .A2(n8837), .ZN(n8716) );
  NAND2_X1 U9882 ( .A1(n9089), .A2(n9137), .ZN(n8715) );
  NAND2_X1 U9883 ( .A1(n8716), .A2(n8715), .ZN(n9047) );
  AOI22_X1 U9884 ( .A1(n9047), .A2(n8840), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8717) );
  OAI21_X1 U9885 ( .B1(n8718), .B2(n10742), .A(n8717), .ZN(n8721) );
  NOR3_X1 U9886 ( .A1(n8719), .A2(n9034), .A3(n8769), .ZN(n8720) );
  AOI211_X1 U9887 ( .C1(n8723), .C2(n8722), .A(n8721), .B(n8720), .ZN(n8724)
         );
  OAI21_X1 U9888 ( .B1(n8725), .B2(n8882), .A(n8724), .ZN(P2_U3218) );
  INV_X1 U9889 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8792) );
  OAI222_X1 U9890 ( .A1(n10596), .A2(n8727), .B1(n8726), .B2(P1_U3084), .C1(
        n8792), .C2(n8813), .ZN(P1_U3324) );
  NAND2_X1 U9891 ( .A1(n8729), .A2(n8728), .ZN(n8731) );
  AND2_X1 U9892 ( .A1(n8731), .A2(n8730), .ZN(n8753) );
  OAI21_X1 U9893 ( .B1(n8748), .B2(n8733), .A(n8732), .ZN(n8734) );
  AOI21_X1 U9894 ( .B1(n8750), .B2(n8888), .A(n8734), .ZN(n8735) );
  OAI21_X1 U9895 ( .B1(n8736), .B2(n10742), .A(n8735), .ZN(n8743) );
  INV_X1 U9896 ( .A(n8737), .ZN(n8741) );
  AOI22_X1 U9897 ( .A1(n8738), .A2(n10727), .B1(n8845), .B2(n8890), .ZN(n8739)
         );
  NOR3_X1 U9898 ( .A1(n8741), .A2(n8740), .A3(n8739), .ZN(n8742) );
  AOI211_X1 U9899 ( .C1(n10733), .C2(n8744), .A(n8743), .B(n8742), .ZN(n8745)
         );
  OAI21_X1 U9900 ( .B1(n8753), .B2(n8882), .A(n8745), .ZN(P2_U3217) );
  OAI21_X1 U9901 ( .B1(n8748), .B2(n8747), .A(n8746), .ZN(n8749) );
  AOI21_X1 U9902 ( .B1(n8750), .B2(n8887), .A(n8749), .ZN(n8751) );
  OAI21_X1 U9903 ( .B1(n8752), .B2(n10742), .A(n8751), .ZN(n8759) );
  INV_X1 U9904 ( .A(n8753), .ZN(n8757) );
  AOI22_X1 U9905 ( .A1(n8754), .A2(n10727), .B1(n8845), .B2(n8889), .ZN(n8755)
         );
  NOR3_X1 U9906 ( .A1(n8757), .A2(n8756), .A3(n8755), .ZN(n8758) );
  AOI211_X1 U9907 ( .C1(n10733), .C2(n8760), .A(n8759), .B(n8758), .ZN(n8761)
         );
  OAI21_X1 U9908 ( .B1(n8762), .B2(n8882), .A(n8761), .ZN(P2_U3243) );
  NOR2_X1 U9909 ( .A1(n10742), .A2(n10808), .ZN(n8767) );
  NAND2_X1 U9910 ( .A1(n8897), .A2(n8837), .ZN(n8764) );
  NAND2_X1 U9911 ( .A1(n8899), .A2(n9137), .ZN(n8763) );
  AND2_X1 U9912 ( .A1(n8764), .A2(n8763), .ZN(n10800) );
  OAI22_X1 U9913 ( .A1(n8765), .A2(n10800), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9543), .ZN(n8766) );
  AOI211_X1 U9914 ( .C1(n10733), .C2(n10806), .A(n8767), .B(n8766), .ZN(n8774)
         );
  OAI22_X1 U9915 ( .A1(n8769), .A2(n10737), .B1(n8882), .B2(n8768), .ZN(n8770)
         );
  NAND3_X1 U9916 ( .A1(n8772), .A2(n8771), .A3(n8770), .ZN(n8773) );
  OAI211_X1 U9917 ( .C1(n8775), .C2(n8882), .A(n8774), .B(n8773), .ZN(P2_U3229) );
  OAI222_X1 U9918 ( .A1(n9699), .A2(n8777), .B1(n6363), .B2(P2_U3152), .C1(
        n8776), .C2(n9696), .ZN(P2_U3331) );
  OR2_X1 U9919 ( .A1(n10532), .A2(n10421), .ZN(n8779) );
  NAND2_X1 U9920 ( .A1(n10532), .A2(n10421), .ZN(n8780) );
  NAND2_X1 U9921 ( .A1(n8781), .A2(n8780), .ZN(n10417) );
  XNOR2_X1 U9922 ( .A(n10526), .B(n10447), .ZN(n9986) );
  NAND2_X1 U9923 ( .A1(n10518), .A2(n10385), .ZN(n9988) );
  AND2_X1 U9924 ( .A1(n10515), .A2(n10404), .ZN(n8782) );
  NAND2_X1 U9925 ( .A1(n10508), .A2(n10387), .ZN(n9999) );
  NAND2_X1 U9926 ( .A1(n10351), .A2(n9999), .ZN(n10056) );
  NAND2_X1 U9927 ( .A1(n10367), .A2(n10056), .ZN(n8784) );
  INV_X1 U9928 ( .A(n10387), .ZN(n10357) );
  OR2_X1 U9929 ( .A1(n10508), .A2(n10357), .ZN(n8783) );
  NOR2_X1 U9930 ( .A1(n10348), .A2(n10378), .ZN(n8786) );
  NAND2_X1 U9931 ( .A1(n10348), .A2(n10378), .ZN(n8785) );
  NAND2_X1 U9932 ( .A1(n10500), .A2(n10321), .ZN(n10007) );
  NAND2_X1 U9933 ( .A1(n10313), .A2(n8788), .ZN(n10301) );
  NAND2_X1 U9934 ( .A1(n10488), .A2(n10322), .ZN(n9920) );
  NAND2_X1 U9935 ( .A1(n10301), .A2(n10300), .ZN(n10299) );
  OR2_X1 U9936 ( .A1(n10488), .A2(n10092), .ZN(n8789) );
  NAND2_X1 U9937 ( .A1(n10299), .A2(n8789), .ZN(n10279) );
  NAND2_X1 U9938 ( .A1(n10481), .A2(n8790), .ZN(n10015) );
  NOR2_X1 U9939 ( .A1(n10279), .A2(n10282), .ZN(n10281) );
  NAND2_X1 U9940 ( .A1(n8791), .A2(n9807), .ZN(n8794) );
  OR2_X1 U9941 ( .A1(n9822), .A2(n8792), .ZN(n8793) );
  OR2_X2 U9942 ( .A1(n10303), .A2(n10481), .ZN(n10291) );
  NOR2_X2 U9943 ( .A1(n10476), .A2(n10291), .ZN(n10272) );
  AOI21_X1 U9944 ( .B1(n10476), .B2(n10291), .A(n10272), .ZN(n10477) );
  INV_X1 U9945 ( .A(n10476), .ZN(n8799) );
  INV_X1 U9946 ( .A(n8796), .ZN(n8797) );
  AOI22_X1 U9947 ( .A1(n10465), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8797), .B2(
        n10463), .ZN(n8798) );
  OAI21_X1 U9948 ( .B1(n8799), .B2(n11012), .A(n8798), .ZN(n8812) );
  NAND2_X1 U9949 ( .A1(n8800), .A2(n9979), .ZN(n10444) );
  OR2_X1 U9950 ( .A1(n10532), .A2(n9790), .ZN(n9983) );
  NAND2_X1 U9951 ( .A1(n10532), .A2(n9790), .ZN(n9984) );
  NAND2_X1 U9952 ( .A1(n10444), .A2(n10445), .ZN(n10443) );
  INV_X1 U9953 ( .A(n9986), .ZN(n10419) );
  INV_X1 U9954 ( .A(n10447), .ZN(n9827) );
  OR2_X1 U9955 ( .A1(n10526), .A2(n9827), .ZN(n9862) );
  OR2_X1 U9956 ( .A1(n10515), .A2(n9722), .ZN(n9995) );
  NAND2_X1 U9957 ( .A1(n10384), .A2(n9995), .ZN(n8801) );
  NAND2_X1 U9958 ( .A1(n10515), .A2(n9722), .ZN(n9996) );
  NAND2_X1 U9959 ( .A1(n8801), .A2(n9996), .ZN(n10376) );
  INV_X1 U9960 ( .A(n9999), .ZN(n8802) );
  INV_X1 U9961 ( .A(n10378), .ZN(n10342) );
  OR2_X1 U9962 ( .A1(n10348), .A2(n10342), .ZN(n10004) );
  NAND2_X1 U9963 ( .A1(n10348), .A2(n10342), .ZN(n10005) );
  INV_X1 U9964 ( .A(n10008), .ZN(n10317) );
  NOR2_X1 U9965 ( .A1(n10316), .A2(n10317), .ZN(n8804) );
  INV_X1 U9966 ( .A(n10296), .ZN(n9875) );
  NOR2_X1 U9967 ( .A1(n10300), .A2(n9875), .ZN(n8805) );
  INV_X1 U9968 ( .A(n10282), .ZN(n10059) );
  OAI21_X1 U9969 ( .B1(n10283), .B2(n10059), .A(n9825), .ZN(n8806) );
  XOR2_X1 U9970 ( .A(n10062), .B(n8806), .Z(n8811) );
  INV_X1 U9971 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U9972 ( .A1(n6644), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U9973 ( .A1(n5033), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8807) );
  OAI211_X1 U9974 ( .C1(n9813), .C2(n8809), .A(n8808), .B(n8807), .ZN(n10091)
         );
  NAND2_X1 U9975 ( .A1(n10640), .A2(P1_B_REG_SCAN_IN), .ZN(n8810) );
  AND2_X1 U9976 ( .A1(n10769), .A2(n8810), .ZN(n10265) );
  INV_X1 U9977 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9821) );
  OAI222_X1 U9978 ( .A1(n10596), .A2(n9820), .B1(n6405), .B2(P1_U3084), .C1(
        n9821), .C2(n8813), .ZN(P1_U3323) );
  XNOR2_X1 U9979 ( .A(n8815), .B(n8814), .ZN(n8821) );
  NOR2_X1 U9980 ( .A1(n8984), .A2(n10742), .ZN(n8819) );
  AOI22_X1 U9981 ( .A1(n8991), .A2(n10731), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8816) );
  OAI21_X1 U9982 ( .B1(n8817), .B2(n10736), .A(n8816), .ZN(n8818) );
  AOI211_X1 U9983 ( .C1(n9167), .C2(n10733), .A(n8819), .B(n8818), .ZN(n8820)
         );
  OAI21_X1 U9984 ( .B1(n8821), .B2(n8882), .A(n8820), .ZN(P2_U3216) );
  XNOR2_X1 U9985 ( .A(n8823), .B(n8822), .ZN(n8830) );
  AOI22_X1 U9986 ( .A1(n10731), .A2(n9110), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8826) );
  INV_X1 U9987 ( .A(n10742), .ZN(n8876) );
  INV_X1 U9988 ( .A(n8824), .ZN(n9084) );
  NAND2_X1 U9989 ( .A1(n8876), .A2(n9084), .ZN(n8825) );
  OAI211_X1 U9990 ( .C1(n8827), .C2(n10736), .A(n8826), .B(n8825), .ZN(n8828)
         );
  AOI21_X1 U9991 ( .B1(n9199), .B2(n10733), .A(n8828), .ZN(n8829) );
  OAI21_X1 U9992 ( .B1(n8830), .B2(n8882), .A(n8829), .ZN(P2_U3225) );
  NAND2_X1 U9993 ( .A1(n8832), .A2(n8831), .ZN(n8836) );
  INV_X1 U9994 ( .A(n8833), .ZN(n8834) );
  AOI21_X1 U9995 ( .B1(n8836), .B2(n8835), .A(n8834), .ZN(n8844) );
  NAND2_X1 U9996 ( .A1(n8991), .A2(n8837), .ZN(n8839) );
  NAND2_X1 U9997 ( .A1(n8886), .A2(n9137), .ZN(n8838) );
  NAND2_X1 U9998 ( .A1(n8839), .A2(n8838), .ZN(n9021) );
  AOI22_X1 U9999 ( .A1(n9021), .A2(n8840), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8841) );
  OAI21_X1 U10000 ( .B1(n9014), .B2(n10742), .A(n8841), .ZN(n8842) );
  AOI21_X1 U10001 ( .B1(n9178), .B2(n10733), .A(n8842), .ZN(n8843) );
  OAI21_X1 U10002 ( .B1(n8844), .B2(n8882), .A(n8843), .ZN(P2_U3227) );
  INV_X1 U10003 ( .A(n9182), .ZN(n9033) );
  NAND2_X1 U10004 ( .A1(n8886), .A2(n8845), .ZN(n8849) );
  OR2_X1 U10005 ( .A1(n8846), .A2(n8882), .ZN(n8848) );
  MUX2_X1 U10006 ( .A(n8849), .B(n8848), .S(n8847), .Z(n8855) );
  NOR2_X1 U10007 ( .A1(n10742), .A2(n9030), .ZN(n8853) );
  OAI22_X1 U10008 ( .A1(n8851), .A2(n10736), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8850), .ZN(n8852) );
  AOI211_X1 U10009 ( .C1(n10731), .C2(n9075), .A(n8853), .B(n8852), .ZN(n8854)
         );
  OAI211_X1 U10010 ( .C1(n9033), .C2(n8856), .A(n8855), .B(n8854), .ZN(
        P2_U3231) );
  XNOR2_X1 U10011 ( .A(n8858), .B(n8857), .ZN(n8864) );
  AOI22_X1 U10012 ( .A1(n10731), .A2(n9140), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3152), .ZN(n8861) );
  INV_X1 U10013 ( .A(n8859), .ZN(n9097) );
  NAND2_X1 U10014 ( .A1(n8876), .A2(n9097), .ZN(n8860) );
  OAI211_X1 U10015 ( .C1(n9068), .C2(n10736), .A(n8861), .B(n8860), .ZN(n8862)
         );
  AOI21_X1 U10016 ( .B1(n9204), .B2(n10733), .A(n8862), .ZN(n8863) );
  OAI21_X1 U10017 ( .B1(n8864), .B2(n8882), .A(n8863), .ZN(P2_U3235) );
  INV_X1 U10018 ( .A(n8865), .ZN(n8866) );
  AOI21_X1 U10019 ( .B1(n8868), .B2(n8867), .A(n8866), .ZN(n8873) );
  AOI22_X1 U10020 ( .A1(n10731), .A2(n9102), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3152), .ZN(n8870) );
  NAND2_X1 U10021 ( .A1(n8876), .A2(n9064), .ZN(n8869) );
  OAI211_X1 U10022 ( .C1(n9034), .C2(n10736), .A(n8870), .B(n8869), .ZN(n8871)
         );
  AOI21_X1 U10023 ( .B1(n9194), .B2(n10733), .A(n8871), .ZN(n8872) );
  OAI21_X1 U10024 ( .B1(n8873), .B2(n8882), .A(n8872), .ZN(P2_U3237) );
  XNOR2_X1 U10025 ( .A(n8875), .B(n8874), .ZN(n8883) );
  AOI22_X1 U10026 ( .A1(n9040), .A2(n10731), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3152), .ZN(n8878) );
  NAND2_X1 U10027 ( .A1(n9003), .A2(n8876), .ZN(n8877) );
  OAI211_X1 U10028 ( .C1(n8879), .C2(n10736), .A(n8878), .B(n8877), .ZN(n8880)
         );
  AOI21_X1 U10029 ( .B1(n9173), .B2(n10733), .A(n8880), .ZN(n8881) );
  OAI21_X1 U10030 ( .B1(n8883), .B2(n8882), .A(n8881), .ZN(P2_U3242) );
  MUX2_X1 U10031 ( .A(n8884), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8902), .Z(
        P2_U3583) );
  INV_X1 U10032 ( .A(n8885), .ZN(n8976) );
  MUX2_X1 U10033 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8976), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10034 ( .A(n8992), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8902), .Z(
        P2_U3580) );
  MUX2_X1 U10035 ( .A(n9000), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8902), .Z(
        P2_U3579) );
  MUX2_X1 U10036 ( .A(n8991), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8902), .Z(
        P2_U3578) );
  MUX2_X1 U10037 ( .A(n9040), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8902), .Z(
        P2_U3577) );
  MUX2_X1 U10038 ( .A(n8886), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8902), .Z(
        P2_U3576) );
  MUX2_X1 U10039 ( .A(n9075), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8902), .Z(
        P2_U3575) );
  MUX2_X1 U10040 ( .A(n9089), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8902), .Z(
        P2_U3574) );
  MUX2_X1 U10041 ( .A(n9102), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8902), .Z(
        P2_U3573) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9110), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10043 ( .A(n9140), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8902), .Z(
        P2_U3571) );
  MUX2_X1 U10044 ( .A(n9109), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8902), .Z(
        P2_U3570) );
  MUX2_X1 U10045 ( .A(n9138), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8902), .Z(
        P2_U3569) );
  MUX2_X1 U10046 ( .A(n8887), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8902), .Z(
        P2_U3568) );
  MUX2_X1 U10047 ( .A(n8888), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8902), .Z(
        P2_U3567) );
  MUX2_X1 U10048 ( .A(n8889), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8902), .Z(
        P2_U3566) );
  MUX2_X1 U10049 ( .A(n8890), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8902), .Z(
        P2_U3565) );
  MUX2_X1 U10050 ( .A(n8891), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8902), .Z(
        P2_U3564) );
  MUX2_X1 U10051 ( .A(n8892), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8902), .Z(
        P2_U3563) );
  MUX2_X1 U10052 ( .A(n8893), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8902), .Z(
        P2_U3562) );
  MUX2_X1 U10053 ( .A(n8894), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8902), .Z(
        P2_U3561) );
  MUX2_X1 U10054 ( .A(n8895), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8902), .Z(
        P2_U3560) );
  MUX2_X1 U10055 ( .A(n8896), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8902), .Z(
        P2_U3559) );
  MUX2_X1 U10056 ( .A(n8897), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8902), .Z(
        P2_U3558) );
  MUX2_X1 U10057 ( .A(n8898), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8902), .Z(
        P2_U3557) );
  MUX2_X1 U10058 ( .A(n8899), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8902), .Z(
        P2_U3556) );
  MUX2_X1 U10059 ( .A(n8900), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8902), .Z(
        P2_U3555) );
  MUX2_X1 U10060 ( .A(n10730), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8902), .Z(
        P2_U3554) );
  MUX2_X1 U10061 ( .A(n8901), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8902), .Z(
        P2_U3553) );
  MUX2_X1 U10062 ( .A(n8903), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8902), .Z(
        P2_U3552) );
  INV_X1 U10063 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8912) );
  XNOR2_X1 U10064 ( .A(n8932), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8909) );
  INV_X1 U10065 ( .A(n8914), .ZN(n8906) );
  AOI21_X1 U10066 ( .B1(n8906), .B2(n8905), .A(n8904), .ZN(n8908) );
  NAND2_X1 U10067 ( .A1(n8909), .A2(n8908), .ZN(n8930) );
  OAI211_X1 U10068 ( .C1(n8909), .C2(n8908), .A(n8907), .B(n8930), .ZN(n8911)
         );
  OAI211_X1 U10069 ( .C1(n8929), .C2(n8912), .A(n8911), .B(n8910), .ZN(n8919)
         );
  AOI21_X1 U10070 ( .B1(n8914), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8913), .ZN(
        n8917) );
  NAND2_X1 U10071 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n8924), .ZN(n8915) );
  OAI21_X1 U10072 ( .B1(n8924), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8915), .ZN(
        n8916) );
  AOI211_X1 U10073 ( .C1(n8917), .C2(n8916), .A(n8923), .B(n8961), .ZN(n8918)
         );
  AOI211_X1 U10074 ( .C1(n8959), .C2(n8924), .A(n8919), .B(n8918), .ZN(n8920)
         );
  INV_X1 U10075 ( .A(n8920), .ZN(P2_U3262) );
  OR2_X1 U10076 ( .A1(n8939), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U10077 ( .A1(n8939), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U10078 ( .A1(n8922), .A2(n8921), .ZN(n8926) );
  AOI21_X1 U10079 ( .B1(n8926), .B2(n8925), .A(n8942), .ZN(n8941) );
  INV_X1 U10080 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8928) );
  OAI21_X1 U10081 ( .B1(n8929), .B2(n8928), .A(n8927), .ZN(n8938) );
  OAI21_X1 U10082 ( .B1(n8932), .B2(n8931), .A(n8930), .ZN(n8935) );
  INV_X1 U10083 ( .A(n8939), .ZN(n8943) );
  NAND2_X1 U10084 ( .A1(n8943), .A2(n8933), .ZN(n8947) );
  OAI21_X1 U10085 ( .B1(n8943), .B2(n8933), .A(n8947), .ZN(n8934) );
  NOR2_X1 U10086 ( .A1(n8934), .A2(n8935), .ZN(n8949) );
  AOI21_X1 U10087 ( .B1(n8935), .B2(n8934), .A(n8949), .ZN(n8936) );
  NOR2_X1 U10088 ( .A1(n8957), .A2(n8936), .ZN(n8937) );
  AOI211_X1 U10089 ( .C1(n8959), .C2(n8939), .A(n8938), .B(n8937), .ZN(n8940)
         );
  OAI21_X1 U10090 ( .B1(n8941), .B2(n8961), .A(n8940), .ZN(P2_U3263) );
  MUX2_X1 U10091 ( .A(n9116), .B(P2_REG2_REG_19__SCAN_IN), .S(n10812), .Z(
        n8946) );
  AOI21_X1 U10092 ( .B1(n8944), .B2(n8943), .A(n8942), .ZN(n8945) );
  XOR2_X1 U10093 ( .A(n8946), .B(n8945), .Z(n8962) );
  INV_X1 U10094 ( .A(n8947), .ZN(n8948) );
  NOR2_X1 U10095 ( .A1(n8949), .A2(n8948), .ZN(n8952) );
  XNOR2_X1 U10096 ( .A(n10812), .B(n8950), .ZN(n8951) );
  XNOR2_X1 U10097 ( .A(n8952), .B(n8951), .ZN(n8956) );
  NAND2_X1 U10098 ( .A1(n8953), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8954) );
  OAI211_X1 U10099 ( .C1(n8957), .C2(n8956), .A(n8955), .B(n8954), .ZN(n8958)
         );
  AOI21_X1 U10100 ( .B1(n10812), .B2(n8959), .A(n8958), .ZN(n8960) );
  OAI21_X1 U10101 ( .B1(n8962), .B2(n8961), .A(n8960), .ZN(P2_U3264) );
  INV_X1 U10102 ( .A(n8963), .ZN(n9152) );
  NAND2_X1 U10103 ( .A1(n8965), .A2(n8964), .ZN(n9151) );
  NAND3_X1 U10104 ( .A1(n9152), .A2(n9144), .A3(n9151), .ZN(n8968) );
  AOI21_X1 U10105 ( .B1(n10817), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8966), .ZN(
        n8967) );
  OAI211_X1 U10106 ( .C1(n5338), .C2(n9133), .A(n8968), .B(n8967), .ZN(
        P2_U3266) );
  XNOR2_X1 U10107 ( .A(n8970), .B(n8969), .ZN(n9166) );
  AOI21_X1 U10108 ( .B1(n9162), .B2(n8981), .A(n8971), .ZN(n9163) );
  AOI22_X1 U10109 ( .A1(n8972), .A2(n9130), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10817), .ZN(n8973) );
  OAI21_X1 U10110 ( .B1(n5342), .B2(n9133), .A(n8973), .ZN(n8978) );
  AOI211_X1 U10111 ( .C1(n9144), .C2(n9163), .A(n8978), .B(n8977), .ZN(n8979)
         );
  OAI21_X1 U10112 ( .B1(n9166), .B2(n9146), .A(n8979), .ZN(P2_U3268) );
  XOR2_X1 U10113 ( .A(n8989), .B(n8980), .Z(n9171) );
  INV_X1 U10114 ( .A(n9002), .ZN(n8983) );
  INV_X1 U10115 ( .A(n8981), .ZN(n8982) );
  AOI21_X1 U10116 ( .B1(n9167), .B2(n8983), .A(n8982), .ZN(n9168) );
  INV_X1 U10117 ( .A(n8984), .ZN(n8985) );
  AOI22_X1 U10118 ( .A1(n8985), .A2(n9130), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10817), .ZN(n8986) );
  OAI21_X1 U10119 ( .B1(n8987), .B2(n9133), .A(n8986), .ZN(n8996) );
  OAI211_X1 U10120 ( .C1(n8990), .C2(n8989), .A(n8988), .B(n10798), .ZN(n8994)
         );
  AOI22_X1 U10121 ( .A1(n8992), .A2(n9139), .B1(n9137), .B2(n8991), .ZN(n8993)
         );
  NOR2_X1 U10122 ( .A1(n9170), .A2(n10817), .ZN(n8995) );
  AOI211_X1 U10123 ( .C1(n9144), .C2(n9168), .A(n8996), .B(n8995), .ZN(n8997)
         );
  OAI21_X1 U10124 ( .B1(n9171), .B2(n9146), .A(n8997), .ZN(P2_U3269) );
  XNOR2_X1 U10125 ( .A(n8998), .B(n5493), .ZN(n9176) );
  NOR2_X1 U10126 ( .A1(n8999), .A2(n9133), .ZN(n9007) );
  XNOR2_X1 U10127 ( .A(n5046), .B(n5493), .ZN(n9001) );
  AOI222_X1 U10128 ( .A1(n10798), .A2(n9001), .B1(n9000), .B2(n9139), .C1(
        n9040), .C2(n9137), .ZN(n9175) );
  AOI211_X1 U10129 ( .C1(n9173), .C2(n9011), .A(n11000), .B(n9002), .ZN(n9172)
         );
  AOI22_X1 U10130 ( .A1(n9172), .A2(n9004), .B1(n9130), .B2(n9003), .ZN(n9005)
         );
  AOI21_X1 U10131 ( .B1(n9175), .B2(n9005), .A(n10817), .ZN(n9006) );
  AOI211_X1 U10132 ( .C1(n10817), .C2(P2_REG2_REG_26__SCAN_IN), .A(n9007), .B(
        n9006), .ZN(n9008) );
  OAI21_X1 U10133 ( .B1(n9176), .B2(n9146), .A(n9008), .ZN(P2_U3270) );
  XOR2_X1 U10134 ( .A(n9019), .B(n9009), .Z(n9181) );
  INV_X1 U10135 ( .A(n9010), .ZN(n9013) );
  INV_X1 U10136 ( .A(n9011), .ZN(n9012) );
  AOI211_X1 U10137 ( .C1(n9178), .C2(n9013), .A(n11000), .B(n9012), .ZN(n9177)
         );
  INV_X1 U10138 ( .A(n9014), .ZN(n9015) );
  AOI22_X1 U10139 ( .A1(n9015), .A2(n9130), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10817), .ZN(n9016) );
  OAI21_X1 U10140 ( .B1(n9017), .B2(n9133), .A(n9016), .ZN(n9024) );
  AOI211_X1 U10141 ( .C1(n9020), .C2(n9019), .A(n9070), .B(n9018), .ZN(n9022)
         );
  NOR2_X1 U10142 ( .A1(n9022), .A2(n9021), .ZN(n9180) );
  NOR2_X1 U10143 ( .A1(n9180), .A2(n10817), .ZN(n9023) );
  AOI211_X1 U10144 ( .C1(n9177), .C2(n9025), .A(n9024), .B(n9023), .ZN(n9026)
         );
  OAI21_X1 U10145 ( .B1(n9181), .B2(n9146), .A(n9026), .ZN(P2_U3271) );
  INV_X1 U10146 ( .A(n9027), .ZN(n9028) );
  AOI21_X1 U10147 ( .B1(n5269), .B2(n9029), .A(n9028), .ZN(n9186) );
  XOR2_X1 U10148 ( .A(n9182), .B(n9051), .Z(n9183) );
  INV_X1 U10149 ( .A(n9030), .ZN(n9031) );
  AOI22_X1 U10150 ( .A1(n9031), .A2(n9130), .B1(n10817), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n9032) );
  OAI21_X1 U10151 ( .B1(n9033), .B2(n9133), .A(n9032), .ZN(n9042) );
  NOR2_X1 U10152 ( .A1(n9034), .A2(n9067), .ZN(n9039) );
  AOI211_X1 U10153 ( .C1(n9037), .C2(n9036), .A(n9070), .B(n9035), .ZN(n9038)
         );
  AOI211_X1 U10154 ( .C1(n9139), .C2(n9040), .A(n9039), .B(n9038), .ZN(n9185)
         );
  NOR2_X1 U10155 ( .A1(n9185), .A2(n10817), .ZN(n9041) );
  AOI211_X1 U10156 ( .C1(n9183), .C2(n9144), .A(n9042), .B(n9041), .ZN(n9043)
         );
  OAI21_X1 U10157 ( .B1(n9186), .B2(n9146), .A(n9043), .ZN(P2_U3272) );
  OAI21_X1 U10158 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9048) );
  AOI21_X1 U10159 ( .B1(n9048), .B2(n10798), .A(n9047), .ZN(n9192) );
  OR2_X1 U10160 ( .A1(n9050), .A2(n9049), .ZN(n9188) );
  NAND3_X1 U10161 ( .A1(n9188), .A2(n9187), .A3(n9114), .ZN(n9060) );
  INV_X1 U10162 ( .A(n9063), .ZN(n9053) );
  INV_X1 U10163 ( .A(n9051), .ZN(n9052) );
  AOI21_X1 U10164 ( .B1(n9054), .B2(n9053), .A(n9052), .ZN(n9189) );
  AOI22_X1 U10165 ( .A1(n10817), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9055), 
        .B2(n9130), .ZN(n9056) );
  OAI21_X1 U10166 ( .B1(n9057), .B2(n9133), .A(n9056), .ZN(n9058) );
  AOI21_X1 U10167 ( .B1(n9189), .B2(n9144), .A(n9058), .ZN(n9059) );
  OAI211_X1 U10168 ( .C1(n10817), .C2(n9192), .A(n9060), .B(n9059), .ZN(
        P2_U3273) );
  XNOR2_X1 U10169 ( .A(n9062), .B(n9061), .ZN(n9198) );
  AOI21_X1 U10170 ( .B1(n9194), .B2(n9082), .A(n9063), .ZN(n9195) );
  AOI22_X1 U10171 ( .A1(n10817), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9064), 
        .B2(n9130), .ZN(n9065) );
  OAI21_X1 U10172 ( .B1(n9066), .B2(n9133), .A(n9065), .ZN(n9077) );
  NOR2_X1 U10173 ( .A1(n9068), .A2(n9067), .ZN(n9074) );
  AOI211_X1 U10174 ( .C1(n9072), .C2(n9071), .A(n9070), .B(n9069), .ZN(n9073)
         );
  AOI211_X1 U10175 ( .C1(n9139), .C2(n9075), .A(n9074), .B(n9073), .ZN(n9197)
         );
  NOR2_X1 U10176 ( .A1(n9197), .A2(n10817), .ZN(n9076) );
  AOI211_X1 U10177 ( .C1(n9195), .C2(n9144), .A(n9077), .B(n9076), .ZN(n9078)
         );
  OAI21_X1 U10178 ( .B1(n9198), .B2(n9146), .A(n9078), .ZN(P2_U3274) );
  INV_X1 U10179 ( .A(n9079), .ZN(n9080) );
  AOI21_X1 U10180 ( .B1(n9087), .B2(n9081), .A(n9080), .ZN(n9203) );
  INV_X1 U10181 ( .A(n9096), .ZN(n9083) );
  AOI21_X1 U10182 ( .B1(n9199), .B2(n9083), .A(n5332), .ZN(n9200) );
  AOI22_X1 U10183 ( .A1(n10817), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9084), 
        .B2(n9130), .ZN(n9085) );
  OAI21_X1 U10184 ( .B1(n9086), .B2(n9133), .A(n9085), .ZN(n9092) );
  XNOR2_X1 U10185 ( .A(n9088), .B(n9087), .ZN(n9090) );
  AOI222_X1 U10186 ( .A1(n10798), .A2(n9090), .B1(n9089), .B2(n9139), .C1(
        n9110), .C2(n9137), .ZN(n9202) );
  NOR2_X1 U10187 ( .A1(n9202), .A2(n10817), .ZN(n9091) );
  AOI211_X1 U10188 ( .C1(n9200), .C2(n9144), .A(n9092), .B(n9091), .ZN(n9093)
         );
  OAI21_X1 U10189 ( .B1(n9203), .B2(n9146), .A(n9093), .ZN(P2_U3275) );
  OAI21_X1 U10190 ( .B1(n9095), .B2(n9100), .A(n9094), .ZN(n9208) );
  AOI21_X1 U10191 ( .B1(n9204), .B2(n9117), .A(n9096), .ZN(n9205) );
  AOI22_X1 U10192 ( .A1(n10817), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9097), 
        .B2(n9130), .ZN(n9098) );
  OAI21_X1 U10193 ( .B1(n9099), .B2(n9133), .A(n9098), .ZN(n9105) );
  XNOR2_X1 U10194 ( .A(n9101), .B(n9100), .ZN(n9103) );
  AOI222_X1 U10195 ( .A1(n10798), .A2(n9103), .B1(n9102), .B2(n9139), .C1(
        n9140), .C2(n9137), .ZN(n9207) );
  NOR2_X1 U10196 ( .A1(n9207), .A2(n10817), .ZN(n9104) );
  AOI211_X1 U10197 ( .C1(n9205), .C2(n9144), .A(n9105), .B(n9104), .ZN(n9106)
         );
  OAI21_X1 U10198 ( .B1(n9208), .B2(n9146), .A(n9106), .ZN(P2_U3276) );
  XNOR2_X1 U10199 ( .A(n9108), .B(n9107), .ZN(n9111) );
  AOI222_X1 U10200 ( .A1(n10798), .A2(n9111), .B1(n9110), .B2(n9139), .C1(
        n9109), .C2(n9137), .ZN(n9214) );
  OR2_X1 U10201 ( .A1(n9113), .A2(n9112), .ZN(n9210) );
  NAND3_X1 U10202 ( .A1(n9210), .A2(n9209), .A3(n9114), .ZN(n9124) );
  OAI22_X1 U10203 ( .A1(n10815), .A2(n9116), .B1(n9115), .B2(n10809), .ZN(
        n9121) );
  OAI211_X1 U10204 ( .C1(n9127), .C2(n9118), .A(n9117), .B(n10803), .ZN(n9213)
         );
  NOR2_X1 U10205 ( .A1(n9213), .A2(n9119), .ZN(n9120) );
  AOI211_X1 U10206 ( .C1(n9122), .C2(n9211), .A(n9121), .B(n9120), .ZN(n9123)
         );
  OAI211_X1 U10207 ( .C1(n10817), .C2(n9214), .A(n9124), .B(n9123), .ZN(
        P2_U3277) );
  XNOR2_X1 U10208 ( .A(n9126), .B(n9125), .ZN(n9220) );
  AOI21_X1 U10209 ( .B1(n9216), .B2(n9128), .A(n9127), .ZN(n9217) );
  INV_X1 U10210 ( .A(n9129), .ZN(n9131) );
  AOI22_X1 U10211 ( .A1(n10817), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9131), 
        .B2(n9130), .ZN(n9132) );
  OAI21_X1 U10212 ( .B1(n9134), .B2(n9133), .A(n9132), .ZN(n9143) );
  XNOR2_X1 U10213 ( .A(n9136), .B(n9135), .ZN(n9141) );
  AOI222_X1 U10214 ( .A1(n10798), .A2(n9141), .B1(n9140), .B2(n9139), .C1(
        n9138), .C2(n9137), .ZN(n9219) );
  NOR2_X1 U10215 ( .A1(n9219), .A2(n10817), .ZN(n9142) );
  AOI211_X1 U10216 ( .C1(n9217), .C2(n9144), .A(n9143), .B(n9142), .ZN(n9145)
         );
  OAI21_X1 U10217 ( .B1(n9220), .B2(n9146), .A(n9145), .ZN(P2_U3278) );
  AOI21_X1 U10218 ( .B1(n9148), .B2(n10904), .A(n9147), .ZN(n9149) );
  OAI21_X1 U10219 ( .B1(n9150), .B2(n11000), .A(n9149), .ZN(n9233) );
  MUX2_X1 U10220 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9233), .S(n11007), .Z(
        P2_U3551) );
  NAND3_X1 U10221 ( .A1(n9152), .A2(n10803), .A3(n9151), .ZN(n9154) );
  OAI211_X1 U10222 ( .C1(n5338), .C2(n10998), .A(n9154), .B(n9153), .ZN(n9234)
         );
  MUX2_X1 U10223 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9234), .S(n11007), .Z(
        P2_U3550) );
  NAND2_X1 U10224 ( .A1(n9155), .A2(n11004), .ZN(n9161) );
  OAI22_X1 U10225 ( .A1(n9157), .A2(n11000), .B1(n9156), .B2(n10998), .ZN(
        n9158) );
  NOR2_X1 U10226 ( .A1(n9159), .A2(n9158), .ZN(n9160) );
  NAND2_X1 U10227 ( .A1(n9161), .A2(n9160), .ZN(n9235) );
  MUX2_X1 U10228 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9235), .S(n11007), .Z(
        P2_U3549) );
  AOI22_X1 U10229 ( .A1(n9163), .A2(n10803), .B1(n10904), .B2(n9162), .ZN(
        n9164) );
  OAI211_X1 U10230 ( .C1(n9166), .C2(n10962), .A(n9165), .B(n9164), .ZN(n9236)
         );
  MUX2_X1 U10231 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9236), .S(n11007), .Z(
        P2_U3548) );
  AOI22_X1 U10232 ( .A1(n9168), .A2(n10803), .B1(n10904), .B2(n9167), .ZN(
        n9169) );
  OAI211_X1 U10233 ( .C1(n9171), .C2(n10962), .A(n9170), .B(n9169), .ZN(n9237)
         );
  MUX2_X1 U10234 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9237), .S(n11007), .Z(
        P2_U3547) );
  AOI21_X1 U10235 ( .B1(n10904), .B2(n9173), .A(n9172), .ZN(n9174) );
  OAI211_X1 U10236 ( .C1(n9176), .C2(n10962), .A(n9175), .B(n9174), .ZN(n9238)
         );
  MUX2_X1 U10237 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9238), .S(n11007), .Z(
        P2_U3546) );
  AOI21_X1 U10238 ( .B1(n10904), .B2(n9178), .A(n9177), .ZN(n9179) );
  OAI211_X1 U10239 ( .C1(n9181), .C2(n10962), .A(n9180), .B(n9179), .ZN(n9239)
         );
  MUX2_X1 U10240 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9239), .S(n11007), .Z(
        P2_U3545) );
  AOI22_X1 U10241 ( .A1(n9183), .A2(n10803), .B1(n10904), .B2(n9182), .ZN(
        n9184) );
  OAI211_X1 U10242 ( .C1(n9186), .C2(n10962), .A(n9185), .B(n9184), .ZN(n9240)
         );
  MUX2_X1 U10243 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9240), .S(n11007), .Z(
        P2_U3544) );
  NAND3_X1 U10244 ( .A1(n9188), .A2(n9187), .A3(n11004), .ZN(n9193) );
  NAND2_X1 U10245 ( .A1(n9189), .A2(n10803), .ZN(n9190) );
  NAND4_X1 U10246 ( .A1(n9193), .A2(n9192), .A3(n9191), .A4(n9190), .ZN(n9241)
         );
  MUX2_X1 U10247 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9241), .S(n11007), .Z(
        P2_U3543) );
  AOI22_X1 U10248 ( .A1(n9195), .A2(n10803), .B1(n10904), .B2(n9194), .ZN(
        n9196) );
  OAI211_X1 U10249 ( .C1(n9198), .C2(n10962), .A(n9197), .B(n9196), .ZN(n9242)
         );
  MUX2_X1 U10250 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9242), .S(n11007), .Z(
        P2_U3542) );
  AOI22_X1 U10251 ( .A1(n9200), .A2(n10803), .B1(n10904), .B2(n9199), .ZN(
        n9201) );
  OAI211_X1 U10252 ( .C1(n9203), .C2(n10962), .A(n9202), .B(n9201), .ZN(n9243)
         );
  MUX2_X1 U10253 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9243), .S(n11007), .Z(
        P2_U3541) );
  AOI22_X1 U10254 ( .A1(n9205), .A2(n10803), .B1(n10904), .B2(n9204), .ZN(
        n9206) );
  OAI211_X1 U10255 ( .C1(n9208), .C2(n10962), .A(n9207), .B(n9206), .ZN(n9244)
         );
  MUX2_X1 U10256 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9244), .S(n11007), .Z(
        P2_U3540) );
  NAND3_X1 U10257 ( .A1(n9210), .A2(n9209), .A3(n11004), .ZN(n9215) );
  NAND2_X1 U10258 ( .A1(n9211), .A2(n10904), .ZN(n9212) );
  NAND4_X1 U10259 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n9245)
         );
  MUX2_X1 U10260 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9245), .S(n11007), .Z(
        P2_U3539) );
  AOI22_X1 U10261 ( .A1(n9217), .A2(n10803), .B1(n10904), .B2(n9216), .ZN(
        n9218) );
  OAI211_X1 U10262 ( .C1(n9220), .C2(n10962), .A(n9219), .B(n9218), .ZN(n9246)
         );
  MUX2_X1 U10263 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9246), .S(n11007), .Z(
        P2_U3538) );
  INV_X1 U10264 ( .A(n9221), .ZN(n9226) );
  AOI21_X1 U10265 ( .B1(n10904), .B2(n9223), .A(n9222), .ZN(n9224) );
  OAI211_X1 U10266 ( .C1(n9226), .C2(n10962), .A(n9225), .B(n9224), .ZN(n9247)
         );
  MUX2_X1 U10267 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9247), .S(n11007), .Z(
        P2_U3537) );
  INV_X1 U10268 ( .A(n9227), .ZN(n9232) );
  AOI21_X1 U10269 ( .B1(n10904), .B2(n9229), .A(n9228), .ZN(n9230) );
  OAI211_X1 U10270 ( .C1(n9232), .C2(n10962), .A(n9231), .B(n9230), .ZN(n9248)
         );
  MUX2_X1 U10271 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9248), .S(n11007), .Z(
        P2_U3536) );
  MUX2_X1 U10272 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9233), .S(n11011), .Z(
        P2_U3519) );
  MUX2_X1 U10273 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9234), .S(n11011), .Z(
        P2_U3518) );
  MUX2_X1 U10274 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9235), .S(n11011), .Z(
        P2_U3517) );
  MUX2_X1 U10275 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9236), .S(n11011), .Z(
        P2_U3516) );
  MUX2_X1 U10276 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9237), .S(n11011), .Z(
        P2_U3515) );
  MUX2_X1 U10277 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9238), .S(n11011), .Z(
        P2_U3514) );
  MUX2_X1 U10278 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9239), .S(n11011), .Z(
        P2_U3513) );
  MUX2_X1 U10279 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9240), .S(n11011), .Z(
        P2_U3512) );
  MUX2_X1 U10280 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9241), .S(n11011), .Z(
        P2_U3511) );
  MUX2_X1 U10281 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9242), .S(n11011), .Z(
        P2_U3510) );
  MUX2_X1 U10282 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9243), .S(n11011), .Z(
        P2_U3509) );
  MUX2_X1 U10283 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9244), .S(n11011), .Z(
        P2_U3508) );
  MUX2_X1 U10284 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9245), .S(n11011), .Z(
        P2_U3507) );
  MUX2_X1 U10285 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9246), .S(n11011), .Z(
        P2_U3505) );
  MUX2_X1 U10286 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9247), .S(n11011), .Z(
        P2_U3502) );
  MUX2_X1 U10287 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9248), .S(n11011), .Z(
        P2_U3499) );
  NAND2_X1 U10288 ( .A1(n10602), .A2(P2_D_REG_29__SCAN_IN), .ZN(n9689) );
  XOR2_X1 U10289 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n9250) );
  XNOR2_X1 U10290 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n9249)
         );
  NAND2_X1 U10291 ( .A1(n9250), .A2(n9249), .ZN(n9353) );
  INV_X1 U10292 ( .A(n9353), .ZN(n9360) );
  XOR2_X1 U10293 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .Z(n9359) );
  XNOR2_X1 U10294 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .ZN(n9358)
         );
  XNOR2_X1 U10295 ( .A(SI_31_), .B(keyinput_1), .ZN(n9253) );
  XNOR2_X1 U10296 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n9252) );
  XNOR2_X1 U10297 ( .A(SI_30_), .B(keyinput_2), .ZN(n9251) );
  NOR3_X1 U10298 ( .A1(n9253), .A2(n9252), .A3(n9251), .ZN(n9257) );
  XNOR2_X1 U10299 ( .A(n9471), .B(keyinput_3), .ZN(n9256) );
  XNOR2_X1 U10300 ( .A(n9469), .B(keyinput_7), .ZN(n9255) );
  XNOR2_X1 U10301 ( .A(SI_23_), .B(keyinput_9), .ZN(n9254) );
  NOR4_X1 U10302 ( .A1(n9257), .A2(n9256), .A3(n9255), .A4(n9254), .ZN(n9266)
         );
  XNOR2_X1 U10303 ( .A(n9463), .B(keyinput_5), .ZN(n9263) );
  XNOR2_X1 U10304 ( .A(n9258), .B(keyinput_4), .ZN(n9262) );
  XNOR2_X1 U10305 ( .A(n9259), .B(keyinput_6), .ZN(n9261) );
  XNOR2_X1 U10306 ( .A(SI_24_), .B(keyinput_8), .ZN(n9260) );
  NOR4_X1 U10307 ( .A1(n9263), .A2(n9262), .A3(n9261), .A4(n9260), .ZN(n9265)
         );
  XNOR2_X1 U10308 ( .A(SI_22_), .B(keyinput_10), .ZN(n9264) );
  AOI21_X1 U10309 ( .B1(n9266), .B2(n9265), .A(n9264), .ZN(n9275) );
  XOR2_X1 U10310 ( .A(SI_18_), .B(keyinput_14), .Z(n9274) );
  XNOR2_X1 U10311 ( .A(n9267), .B(keyinput_11), .ZN(n9273) );
  XNOR2_X1 U10312 ( .A(n9268), .B(keyinput_13), .ZN(n9271) );
  XNOR2_X1 U10313 ( .A(SI_17_), .B(keyinput_15), .ZN(n9270) );
  XNOR2_X1 U10314 ( .A(SI_20_), .B(keyinput_12), .ZN(n9269) );
  NAND3_X1 U10315 ( .A1(n9271), .A2(n9270), .A3(n9269), .ZN(n9272) );
  NOR4_X1 U10316 ( .A1(n9275), .A2(n9274), .A3(n9273), .A4(n9272), .ZN(n9278)
         );
  XOR2_X1 U10317 ( .A(SI_15_), .B(keyinput_17), .Z(n9277) );
  XNOR2_X1 U10318 ( .A(SI_16_), .B(keyinput_16), .ZN(n9276) );
  NOR3_X1 U10319 ( .A1(n9278), .A2(n9277), .A3(n9276), .ZN(n9281) );
  XNOR2_X1 U10320 ( .A(n9484), .B(keyinput_18), .ZN(n9280) );
  XNOR2_X1 U10321 ( .A(SI_13_), .B(keyinput_19), .ZN(n9279) );
  OAI21_X1 U10322 ( .B1(n9281), .B2(n9280), .A(n9279), .ZN(n9288) );
  XNOR2_X1 U10323 ( .A(SI_12_), .B(keyinput_20), .ZN(n9287) );
  XNOR2_X1 U10324 ( .A(SI_10_), .B(keyinput_22), .ZN(n9285) );
  XNOR2_X1 U10325 ( .A(SI_11_), .B(keyinput_21), .ZN(n9284) );
  XNOR2_X1 U10326 ( .A(SI_9_), .B(keyinput_23), .ZN(n9283) );
  XNOR2_X1 U10327 ( .A(SI_8_), .B(keyinput_24), .ZN(n9282) );
  NAND4_X1 U10328 ( .A1(n9285), .A2(n9284), .A3(n9283), .A4(n9282), .ZN(n9286)
         );
  AOI21_X1 U10329 ( .B1(n9288), .B2(n9287), .A(n9286), .ZN(n9291) );
  XNOR2_X1 U10330 ( .A(SI_7_), .B(keyinput_25), .ZN(n9290) );
  XNOR2_X1 U10331 ( .A(n9499), .B(keyinput_26), .ZN(n9289) );
  OAI21_X1 U10332 ( .B1(n9291), .B2(n9290), .A(n9289), .ZN(n9294) );
  XNOR2_X1 U10333 ( .A(n9504), .B(keyinput_28), .ZN(n9293) );
  XNOR2_X1 U10334 ( .A(n9503), .B(keyinput_27), .ZN(n9292) );
  NAND3_X1 U10335 ( .A1(n9294), .A2(n9293), .A3(n9292), .ZN(n9298) );
  XNOR2_X1 U10336 ( .A(n9510), .B(keyinput_31), .ZN(n9297) );
  XNOR2_X1 U10337 ( .A(SI_3_), .B(keyinput_29), .ZN(n9296) );
  XNOR2_X1 U10338 ( .A(SI_2_), .B(keyinput_30), .ZN(n9295) );
  NAND4_X1 U10339 ( .A1(n9298), .A2(n9297), .A3(n9296), .A4(n9295), .ZN(n9302)
         );
  XOR2_X1 U10340 ( .A(SI_0_), .B(keyinput_32), .Z(n9301) );
  XNOR2_X1 U10341 ( .A(n5400), .B(keyinput_33), .ZN(n9300) );
  XNOR2_X1 U10342 ( .A(P2_U3152), .B(keyinput_34), .ZN(n9299) );
  AOI211_X1 U10343 ( .C1(n9302), .C2(n9301), .A(n9300), .B(n9299), .ZN(n9307)
         );
  XNOR2_X1 U10344 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n9306) );
  XNOR2_X1 U10345 ( .A(n9303), .B(keyinput_36), .ZN(n9305) );
  XNOR2_X1 U10346 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n9304)
         );
  OAI211_X1 U10347 ( .C1(n9307), .C2(n9306), .A(n9305), .B(n9304), .ZN(n9310)
         );
  XOR2_X1 U10348 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .Z(n9309) );
  XNOR2_X1 U10349 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n9308)
         );
  AOI21_X1 U10350 ( .B1(n9310), .B2(n9309), .A(n9308), .ZN(n9317) );
  XOR2_X1 U10351 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .Z(n9316) );
  XOR2_X1 U10352 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n9314) );
  XNOR2_X1 U10353 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n9313) );
  XNOR2_X1 U10354 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_41), .ZN(n9312)
         );
  XNOR2_X1 U10355 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n9311)
         );
  NOR4_X1 U10356 ( .A1(n9314), .A2(n9313), .A3(n9312), .A4(n9311), .ZN(n9315)
         );
  OAI21_X1 U10357 ( .B1(n9317), .B2(n9316), .A(n9315), .ZN(n9321) );
  XNOR2_X1 U10358 ( .A(n9318), .B(keyinput_45), .ZN(n9320) );
  XNOR2_X1 U10359 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n9319)
         );
  AOI21_X1 U10360 ( .B1(n9321), .B2(n9320), .A(n9319), .ZN(n9326) );
  XNOR2_X1 U10361 ( .A(n9322), .B(keyinput_47), .ZN(n9325) );
  XNOR2_X1 U10362 ( .A(n9323), .B(keyinput_48), .ZN(n9324) );
  OAI21_X1 U10363 ( .B1(n9326), .B2(n9325), .A(n9324), .ZN(n9333) );
  XNOR2_X1 U10364 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n9332) );
  XNOR2_X1 U10365 ( .A(n9327), .B(keyinput_50), .ZN(n9330) );
  XNOR2_X1 U10366 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n9329) );
  XNOR2_X1 U10367 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n9328)
         );
  NAND3_X1 U10368 ( .A1(n9330), .A2(n9329), .A3(n9328), .ZN(n9331) );
  AOI21_X1 U10369 ( .B1(n9333), .B2(n9332), .A(n9331), .ZN(n9336) );
  XNOR2_X1 U10370 ( .A(n9552), .B(keyinput_53), .ZN(n9335) );
  XOR2_X1 U10371 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n9334) );
  OAI21_X1 U10372 ( .B1(n9336), .B2(n9335), .A(n9334), .ZN(n9343) );
  XNOR2_X1 U10373 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n9342)
         );
  XNOR2_X1 U10374 ( .A(n9337), .B(keyinput_56), .ZN(n9340) );
  XNOR2_X1 U10375 ( .A(n9557), .B(keyinput_57), .ZN(n9339) );
  XNOR2_X1 U10376 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n9338)
         );
  NAND3_X1 U10377 ( .A1(n9340), .A2(n9339), .A3(n9338), .ZN(n9341) );
  AOI21_X1 U10378 ( .B1(n9343), .B2(n9342), .A(n9341), .ZN(n9349) );
  XNOR2_X1 U10379 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n9348) );
  XNOR2_X1 U10380 ( .A(n9564), .B(keyinput_61), .ZN(n9346) );
  XNOR2_X1 U10381 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n9345)
         );
  XNOR2_X1 U10382 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n9344)
         );
  NOR3_X1 U10383 ( .A1(n9346), .A2(n9345), .A3(n9344), .ZN(n9347) );
  OAI21_X1 U10384 ( .B1(n9349), .B2(n9348), .A(n9347), .ZN(n9352) );
  XNOR2_X1 U10385 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_63), .ZN(n9351)
         );
  XNOR2_X1 U10386 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .ZN(n9350) );
  NAND3_X1 U10387 ( .A1(n9352), .A2(n9351), .A3(n9350), .ZN(n9356) );
  XNOR2_X1 U10388 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .ZN(n9355)
         );
  XNOR2_X1 U10389 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .ZN(n9354)
         );
  AOI211_X1 U10390 ( .C1(n9356), .C2(n9355), .A(n9354), .B(n9353), .ZN(n9357)
         );
  AOI211_X1 U10391 ( .C1(n9360), .C2(n9359), .A(n9358), .B(n9357), .ZN(n9364)
         );
  XNOR2_X1 U10392 ( .A(n9361), .B(keyinput_71), .ZN(n9363) );
  XNOR2_X1 U10393 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .ZN(n9362)
         );
  NOR3_X1 U10394 ( .A1(n9364), .A2(n9363), .A3(n9362), .ZN(n9375) );
  XNOR2_X1 U10395 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n9366)
         );
  XNOR2_X1 U10396 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n9365)
         );
  NOR2_X1 U10397 ( .A1(n9366), .A2(n9365), .ZN(n9371) );
  XNOR2_X1 U10398 ( .A(n9367), .B(keyinput_73), .ZN(n9370) );
  XNOR2_X1 U10399 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .ZN(n9369)
         );
  XNOR2_X1 U10400 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n9368)
         );
  NAND4_X1 U10401 ( .A1(n9371), .A2(n9370), .A3(n9369), .A4(n9368), .ZN(n9374)
         );
  XOR2_X1 U10402 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .Z(n9373) );
  XNOR2_X1 U10403 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n9372)
         );
  OAI211_X1 U10404 ( .C1(n9375), .C2(n9374), .A(n9373), .B(n9372), .ZN(n9378)
         );
  XNOR2_X1 U10405 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n9377)
         );
  XNOR2_X1 U10406 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .ZN(n9376)
         );
  NAND3_X1 U10407 ( .A1(n9378), .A2(n9377), .A3(n9376), .ZN(n9381) );
  XNOR2_X1 U10408 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n9380)
         );
  XNOR2_X1 U10409 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n9379)
         );
  NAND3_X1 U10410 ( .A1(n9381), .A2(n9380), .A3(n9379), .ZN(n9390) );
  XNOR2_X1 U10411 ( .A(n9382), .B(keyinput_84), .ZN(n9389) );
  XOR2_X1 U10412 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .Z(n9387) );
  XNOR2_X1 U10413 ( .A(n9383), .B(keyinput_87), .ZN(n9386) );
  XNOR2_X1 U10414 ( .A(n9384), .B(keyinput_86), .ZN(n9385) );
  NAND3_X1 U10415 ( .A1(n9387), .A2(n9386), .A3(n9385), .ZN(n9388) );
  AOI21_X1 U10416 ( .B1(n9390), .B2(n9389), .A(n9388), .ZN(n9393) );
  XNOR2_X1 U10417 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n9392)
         );
  XNOR2_X1 U10418 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n9391)
         );
  OAI21_X1 U10419 ( .B1(n9393), .B2(n9392), .A(n9391), .ZN(n9396) );
  XNOR2_X1 U10420 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n9395)
         );
  XNOR2_X1 U10421 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_91), .ZN(n9394) );
  AOI21_X1 U10422 ( .B1(n9396), .B2(n9395), .A(n9394), .ZN(n9400) );
  XNOR2_X1 U10423 ( .A(n9620), .B(keyinput_93), .ZN(n9399) );
  XNOR2_X1 U10424 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_94), .ZN(n9398) );
  XNOR2_X1 U10425 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_92), .ZN(n9397) );
  NOR4_X1 U10426 ( .A1(n9400), .A2(n9399), .A3(n9398), .A4(n9397), .ZN(n9403)
         );
  XNOR2_X1 U10427 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .ZN(n9402) );
  XNOR2_X1 U10428 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_95), .ZN(n9401) );
  NOR3_X1 U10429 ( .A1(n9403), .A2(n9402), .A3(n9401), .ZN(n9408) );
  XNOR2_X1 U10430 ( .A(n9404), .B(keyinput_97), .ZN(n9407) );
  XNOR2_X1 U10431 ( .A(n9629), .B(keyinput_98), .ZN(n9406) );
  XNOR2_X1 U10432 ( .A(n9630), .B(keyinput_99), .ZN(n9405) );
  OAI211_X1 U10433 ( .C1(n9408), .C2(n9407), .A(n9406), .B(n9405), .ZN(n9411)
         );
  XNOR2_X1 U10434 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_100), .ZN(n9410) );
  XNOR2_X1 U10435 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_101), .ZN(n9409) );
  NAND3_X1 U10436 ( .A1(n9411), .A2(n9410), .A3(n9409), .ZN(n9419) );
  XNOR2_X1 U10437 ( .A(n9638), .B(keyinput_102), .ZN(n9418) );
  XNOR2_X1 U10438 ( .A(n9412), .B(keyinput_104), .ZN(n9416) );
  XNOR2_X1 U10439 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_105), .ZN(n9415) );
  XNOR2_X1 U10440 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_103), .ZN(n9414) );
  XNOR2_X1 U10441 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_106), .ZN(n9413) );
  NAND4_X1 U10442 ( .A1(n9416), .A2(n9415), .A3(n9414), .A4(n9413), .ZN(n9417)
         );
  AOI21_X1 U10443 ( .B1(n9419), .B2(n9418), .A(n9417), .ZN(n9422) );
  XNOR2_X1 U10444 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_107), .ZN(n9421) );
  XNOR2_X1 U10445 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_108), .ZN(n9420) );
  OAI21_X1 U10446 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9425) );
  XNOR2_X1 U10447 ( .A(n5547), .B(keyinput_110), .ZN(n9424) );
  XNOR2_X1 U10448 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_109), .ZN(n9423) );
  NAND3_X1 U10449 ( .A1(n9425), .A2(n9424), .A3(n9423), .ZN(n9430) );
  XNOR2_X1 U10450 ( .A(n9657), .B(keyinput_111), .ZN(n9429) );
  XNOR2_X1 U10451 ( .A(n9426), .B(keyinput_112), .ZN(n9428) );
  XNOR2_X1 U10452 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_113), .ZN(n9427) );
  AOI211_X1 U10453 ( .C1(n9430), .C2(n9429), .A(n9428), .B(n9427), .ZN(n9435)
         );
  XNOR2_X1 U10454 ( .A(n9431), .B(keyinput_114), .ZN(n9434) );
  XOR2_X1 U10455 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_116), .Z(n9433) );
  XOR2_X1 U10456 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_115), .Z(n9432) );
  OAI211_X1 U10457 ( .C1(n9435), .C2(n9434), .A(n9433), .B(n9432), .ZN(n9442)
         );
  XOR2_X1 U10458 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_117), .Z(n9441) );
  XNOR2_X1 U10459 ( .A(n9669), .B(keyinput_119), .ZN(n9438) );
  XNOR2_X1 U10460 ( .A(n9673), .B(keyinput_118), .ZN(n9437) );
  XNOR2_X1 U10461 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_121), .ZN(n9436) );
  NOR3_X1 U10462 ( .A1(n9438), .A2(n9437), .A3(n9436), .ZN(n9440) );
  XNOR2_X1 U10463 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_120), .ZN(n9439) );
  NAND4_X1 U10464 ( .A1(n9442), .A2(n9441), .A3(n9440), .A4(n9439), .ZN(n9445)
         );
  XOR2_X1 U10465 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .Z(n9444) );
  XNOR2_X1 U10466 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_123), .ZN(n9443) );
  AOI21_X1 U10467 ( .B1(n9445), .B2(n9444), .A(n9443), .ZN(n9449) );
  XNOR2_X1 U10468 ( .A(n9446), .B(keyinput_124), .ZN(n9448) );
  INV_X1 U10469 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10599) );
  XNOR2_X1 U10470 ( .A(n10599), .B(keyinput_125), .ZN(n9447) );
  OAI21_X1 U10471 ( .B1(n9449), .B2(n9448), .A(n9447), .ZN(n9452) );
  XOR2_X1 U10472 ( .A(keyinput_127), .B(P1_D_REG_4__SCAN_IN), .Z(n9451) );
  XOR2_X1 U10473 ( .A(keyinput_126), .B(P1_D_REG_3__SCAN_IN), .Z(n9450) );
  NAND3_X1 U10474 ( .A1(n9452), .A2(n9451), .A3(n9450), .ZN(n9687) );
  XOR2_X1 U10475 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_254), .Z(n9686) );
  XOR2_X1 U10476 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_255), .Z(n9685) );
  XNOR2_X1 U10477 ( .A(n9453), .B(keyinput_140), .ZN(n9459) );
  XNOR2_X1 U10478 ( .A(SI_17_), .B(keyinput_143), .ZN(n9455) );
  XNOR2_X1 U10479 ( .A(SI_21_), .B(keyinput_139), .ZN(n9454) );
  NAND2_X1 U10480 ( .A1(n9455), .A2(n9454), .ZN(n9458) );
  XNOR2_X1 U10481 ( .A(SI_19_), .B(keyinput_141), .ZN(n9457) );
  XNOR2_X1 U10482 ( .A(SI_18_), .B(keyinput_142), .ZN(n9456) );
  NOR4_X1 U10483 ( .A1(n9459), .A2(n9458), .A3(n9457), .A4(n9456), .ZN(n9483)
         );
  XOR2_X1 U10484 ( .A(SI_31_), .B(keyinput_129), .Z(n9462) );
  XOR2_X1 U10485 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n9461) );
  XOR2_X1 U10486 ( .A(SI_30_), .B(keyinput_130), .Z(n9460) );
  NAND3_X1 U10487 ( .A1(n9462), .A2(n9461), .A3(n9460), .ZN(n9467) );
  XNOR2_X1 U10488 ( .A(n9463), .B(keyinput_133), .ZN(n9466) );
  XNOR2_X1 U10489 ( .A(SI_26_), .B(keyinput_134), .ZN(n9465) );
  XNOR2_X1 U10490 ( .A(SI_28_), .B(keyinput_132), .ZN(n9464) );
  NAND4_X1 U10491 ( .A1(n9467), .A2(n9466), .A3(n9465), .A4(n9464), .ZN(n9479)
         );
  XNOR2_X1 U10492 ( .A(n9468), .B(keyinput_137), .ZN(n9475) );
  XNOR2_X1 U10493 ( .A(n9469), .B(keyinput_135), .ZN(n9474) );
  XNOR2_X1 U10494 ( .A(n9470), .B(keyinput_136), .ZN(n9473) );
  XNOR2_X1 U10495 ( .A(n9471), .B(keyinput_131), .ZN(n9472) );
  NAND4_X1 U10496 ( .A1(n9475), .A2(n9474), .A3(n9473), .A4(n9472), .ZN(n9478)
         );
  XNOR2_X1 U10497 ( .A(n9476), .B(keyinput_138), .ZN(n9477) );
  OAI21_X1 U10498 ( .B1(n9479), .B2(n9478), .A(n9477), .ZN(n9482) );
  XOR2_X1 U10499 ( .A(SI_15_), .B(keyinput_145), .Z(n9481) );
  XNOR2_X1 U10500 ( .A(SI_16_), .B(keyinput_144), .ZN(n9480) );
  AOI211_X1 U10501 ( .C1(n9483), .C2(n9482), .A(n9481), .B(n9480), .ZN(n9488)
         );
  XNOR2_X1 U10502 ( .A(n9484), .B(keyinput_146), .ZN(n9487) );
  XNOR2_X1 U10503 ( .A(n9485), .B(keyinput_147), .ZN(n9486) );
  OAI21_X1 U10504 ( .B1(n9488), .B2(n9487), .A(n9486), .ZN(n9497) );
  XNOR2_X1 U10505 ( .A(n9489), .B(keyinput_148), .ZN(n9496) );
  XNOR2_X1 U10506 ( .A(n9490), .B(keyinput_151), .ZN(n9494) );
  XNOR2_X1 U10507 ( .A(SI_8_), .B(keyinput_152), .ZN(n9493) );
  XNOR2_X1 U10508 ( .A(SI_11_), .B(keyinput_149), .ZN(n9492) );
  XNOR2_X1 U10509 ( .A(SI_10_), .B(keyinput_150), .ZN(n9491) );
  NAND4_X1 U10510 ( .A1(n9494), .A2(n9493), .A3(n9492), .A4(n9491), .ZN(n9495)
         );
  AOI21_X1 U10511 ( .B1(n9497), .B2(n9496), .A(n9495), .ZN(n9502) );
  XNOR2_X1 U10512 ( .A(n9498), .B(keyinput_153), .ZN(n9501) );
  XNOR2_X1 U10513 ( .A(n9499), .B(keyinput_154), .ZN(n9500) );
  OAI21_X1 U10514 ( .B1(n9502), .B2(n9501), .A(n9500), .ZN(n9507) );
  XNOR2_X1 U10515 ( .A(n9503), .B(keyinput_155), .ZN(n9506) );
  XNOR2_X1 U10516 ( .A(n9504), .B(keyinput_156), .ZN(n9505) );
  NAND3_X1 U10517 ( .A1(n9507), .A2(n9506), .A3(n9505), .ZN(n9514) );
  XNOR2_X1 U10518 ( .A(n9508), .B(keyinput_158), .ZN(n9513) );
  XNOR2_X1 U10519 ( .A(n9509), .B(keyinput_157), .ZN(n9512) );
  XNOR2_X1 U10520 ( .A(n9510), .B(keyinput_159), .ZN(n9511) );
  NAND4_X1 U10521 ( .A1(n9514), .A2(n9513), .A3(n9512), .A4(n9511), .ZN(n9519)
         );
  XOR2_X1 U10522 ( .A(SI_0_), .B(keyinput_160), .Z(n9518) );
  XNOR2_X1 U10523 ( .A(P2_U3152), .B(keyinput_162), .ZN(n9517) );
  XNOR2_X1 U10524 ( .A(n5400), .B(keyinput_161), .ZN(n9516) );
  AOI211_X1 U10525 ( .C1(n9519), .C2(n9518), .A(n9517), .B(n9516), .ZN(n9524)
         );
  XNOR2_X1 U10526 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n9523)
         );
  XNOR2_X1 U10527 ( .A(n9520), .B(keyinput_165), .ZN(n9522) );
  XNOR2_X1 U10528 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n9521)
         );
  OAI211_X1 U10529 ( .C1(n9524), .C2(n9523), .A(n9522), .B(n9521), .ZN(n9527)
         );
  XOR2_X1 U10530 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .Z(n9526) );
  XNOR2_X1 U10531 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n9525)
         );
  AOI21_X1 U10532 ( .B1(n9527), .B2(n9526), .A(n9525), .ZN(n9535) );
  XOR2_X1 U10533 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .Z(n9534) );
  XOR2_X1 U10534 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .Z(n9532) );
  XNOR2_X1 U10535 ( .A(n9528), .B(keyinput_171), .ZN(n9531) );
  XNOR2_X1 U10536 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n9530)
         );
  XNOR2_X1 U10537 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n9529)
         );
  NOR4_X1 U10538 ( .A1(n9532), .A2(n9531), .A3(n9530), .A4(n9529), .ZN(n9533)
         );
  OAI21_X1 U10539 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9539) );
  XNOR2_X1 U10540 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n9538)
         );
  XNOR2_X1 U10541 ( .A(n9536), .B(keyinput_174), .ZN(n9537) );
  AOI21_X1 U10542 ( .B1(n9539), .B2(n9538), .A(n9537), .ZN(n9542) );
  XNOR2_X1 U10543 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n9541)
         );
  XNOR2_X1 U10544 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n9540)
         );
  OAI21_X1 U10545 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(n9551) );
  XNOR2_X1 U10546 ( .A(n9543), .B(keyinput_177), .ZN(n9550) );
  INV_X1 U10547 ( .A(keyinput_180), .ZN(n9548) );
  XNOR2_X1 U10548 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n9547)
         );
  INV_X1 U10549 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9544) );
  OAI22_X1 U10550 ( .A1(n9544), .A2(keyinput_180), .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_179), .ZN(n9545) );
  AOI21_X1 U10551 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_179), .A(n9545), 
        .ZN(n9546) );
  OAI211_X1 U10552 ( .C1(P2_REG3_REG_4__SCAN_IN), .C2(n9548), .A(n9547), .B(
        n9546), .ZN(n9549) );
  AOI21_X1 U10553 ( .B1(n9551), .B2(n9550), .A(n9549), .ZN(n9555) );
  XNOR2_X1 U10554 ( .A(n9552), .B(keyinput_181), .ZN(n9554) );
  XOR2_X1 U10555 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .Z(n9553) );
  OAI21_X1 U10556 ( .B1(n9555), .B2(n9554), .A(n9553), .ZN(n9563) );
  XNOR2_X1 U10557 ( .A(n9556), .B(keyinput_183), .ZN(n9562) );
  XNOR2_X1 U10558 ( .A(n9557), .B(keyinput_185), .ZN(n9560) );
  XNOR2_X1 U10559 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n9559)
         );
  XNOR2_X1 U10560 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n9558)
         );
  NAND3_X1 U10561 ( .A1(n9560), .A2(n9559), .A3(n9558), .ZN(n9561) );
  AOI21_X1 U10562 ( .B1(n9563), .B2(n9562), .A(n9561), .ZN(n9571) );
  XNOR2_X1 U10563 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .ZN(n9570)
         );
  XNOR2_X1 U10564 ( .A(n9564), .B(keyinput_189), .ZN(n9568) );
  XNOR2_X1 U10565 ( .A(n9565), .B(keyinput_190), .ZN(n9567) );
  XNOR2_X1 U10566 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n9566)
         );
  NOR3_X1 U10567 ( .A1(n9568), .A2(n9567), .A3(n9566), .ZN(n9569) );
  OAI21_X1 U10568 ( .B1(n9571), .B2(n9570), .A(n9569), .ZN(n9574) );
  XOR2_X1 U10569 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .Z(n9573) );
  XNOR2_X1 U10570 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n9572)
         );
  NAND3_X1 U10571 ( .A1(n9574), .A2(n9573), .A3(n9572), .ZN(n9579) );
  XNOR2_X1 U10572 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n9578)
         );
  XOR2_X1 U10573 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .Z(n9577)
         );
  XNOR2_X1 U10574 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .ZN(n9576)
         );
  XNOR2_X1 U10575 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n9575)
         );
  NAND2_X1 U10576 ( .A1(n9576), .A2(n9575), .ZN(n9582) );
  AOI211_X1 U10577 ( .C1(n9579), .C2(n9578), .A(n9577), .B(n9582), .ZN(n9587)
         );
  XOR2_X1 U10578 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .Z(n9583)
         );
  XNOR2_X1 U10579 ( .A(n9580), .B(keyinput_198), .ZN(n9581) );
  OAI21_X1 U10580 ( .B1(n9583), .B2(n9582), .A(n9581), .ZN(n9586) );
  XNOR2_X1 U10581 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n9585)
         );
  XNOR2_X1 U10582 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n9584)
         );
  OAI211_X1 U10583 ( .C1(n9587), .C2(n9586), .A(n9585), .B(n9584), .ZN(n9599)
         );
  XNOR2_X1 U10584 ( .A(n9588), .B(keyinput_202), .ZN(n9591) );
  XNOR2_X1 U10585 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .ZN(n9590)
         );
  XNOR2_X1 U10586 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .ZN(n9589)
         );
  NAND3_X1 U10587 ( .A1(n9591), .A2(n9590), .A3(n9589), .ZN(n9595) );
  XNOR2_X1 U10588 ( .A(n9592), .B(keyinput_204), .ZN(n9594) );
  XNOR2_X1 U10589 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .ZN(n9593)
         );
  NOR3_X1 U10590 ( .A1(n9595), .A2(n9594), .A3(n9593), .ZN(n9598) );
  XOR2_X1 U10591 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .Z(n9597)
         );
  XNOR2_X1 U10592 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n9596)
         );
  AOI211_X1 U10593 ( .C1(n9599), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9607)
         );
  XOR2_X1 U10594 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .Z(n9602)
         );
  XNOR2_X1 U10595 ( .A(n9600), .B(keyinput_208), .ZN(n9601) );
  NAND2_X1 U10596 ( .A1(n9602), .A2(n9601), .ZN(n9606) );
  XNOR2_X1 U10597 ( .A(n9603), .B(keyinput_211), .ZN(n9605) );
  XNOR2_X1 U10598 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .ZN(n9604)
         );
  OAI211_X1 U10599 ( .C1(n9607), .C2(n9606), .A(n9605), .B(n9604), .ZN(n9613)
         );
  XNOR2_X1 U10600 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n9612)
         );
  XOR2_X1 U10601 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .Z(n9610)
         );
  XNOR2_X1 U10602 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .ZN(n9609)
         );
  XNOR2_X1 U10603 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n9608)
         );
  NAND3_X1 U10604 ( .A1(n9610), .A2(n9609), .A3(n9608), .ZN(n9611) );
  AOI21_X1 U10605 ( .B1(n9613), .B2(n9612), .A(n9611), .ZN(n9616) );
  XNOR2_X1 U10606 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .ZN(n9615)
         );
  XNOR2_X1 U10607 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .ZN(n9614)
         );
  OAI21_X1 U10608 ( .B1(n9616), .B2(n9615), .A(n9614), .ZN(n9619) );
  XNOR2_X1 U10609 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_218), .ZN(n9618)
         );
  XOR2_X1 U10610 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_219), .Z(n9617) );
  AOI21_X1 U10611 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(n9624) );
  XNOR2_X1 U10612 ( .A(n6370), .B(keyinput_222), .ZN(n9623) );
  XNOR2_X1 U10613 ( .A(n9620), .B(keyinput_221), .ZN(n9622) );
  XNOR2_X1 U10614 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_220), .ZN(n9621) );
  NOR4_X1 U10615 ( .A1(n9624), .A2(n9623), .A3(n9622), .A4(n9621), .ZN(n9628)
         );
  XNOR2_X1 U10616 ( .A(n9625), .B(keyinput_223), .ZN(n9627) );
  XNOR2_X1 U10617 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_224), .ZN(n9626) );
  NOR3_X1 U10618 ( .A1(n9628), .A2(n9627), .A3(n9626), .ZN(n9634) );
  XNOR2_X1 U10619 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_225), .ZN(n9633) );
  XNOR2_X1 U10620 ( .A(n9629), .B(keyinput_226), .ZN(n9632) );
  XNOR2_X1 U10621 ( .A(n9630), .B(keyinput_227), .ZN(n9631) );
  OAI211_X1 U10622 ( .C1(n9634), .C2(n9633), .A(n9632), .B(n9631), .ZN(n9637)
         );
  XNOR2_X1 U10623 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_228), .ZN(n9636) );
  XNOR2_X1 U10624 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_229), .ZN(n9635) );
  NAND3_X1 U10625 ( .A1(n9637), .A2(n9636), .A3(n9635), .ZN(n9647) );
  XNOR2_X1 U10626 ( .A(n9638), .B(keyinput_230), .ZN(n9646) );
  XOR2_X1 U10627 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_234), .Z(n9644) );
  XNOR2_X1 U10628 ( .A(n9639), .B(keyinput_231), .ZN(n9643) );
  XNOR2_X1 U10629 ( .A(n9640), .B(keyinput_233), .ZN(n9642) );
  XNOR2_X1 U10630 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_232), .ZN(n9641) );
  NAND4_X1 U10631 ( .A1(n9644), .A2(n9643), .A3(n9642), .A4(n9641), .ZN(n9645)
         );
  AOI21_X1 U10632 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n9652) );
  XNOR2_X1 U10633 ( .A(n9648), .B(keyinput_235), .ZN(n9651) );
  XNOR2_X1 U10634 ( .A(n9649), .B(keyinput_236), .ZN(n9650) );
  OAI21_X1 U10635 ( .B1(n9652), .B2(n9651), .A(n9650), .ZN(n9656) );
  XNOR2_X1 U10636 ( .A(n9653), .B(keyinput_237), .ZN(n9655) );
  XNOR2_X1 U10637 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_238), .ZN(n9654) );
  NAND3_X1 U10638 ( .A1(n9656), .A2(n9655), .A3(n9654), .ZN(n9661) );
  XNOR2_X1 U10639 ( .A(n9657), .B(keyinput_239), .ZN(n9660) );
  XNOR2_X1 U10640 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_240), .ZN(n9659) );
  XNOR2_X1 U10641 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_241), .ZN(n9658) );
  AOI211_X1 U10642 ( .C1(n9661), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9665)
         );
  XNOR2_X1 U10643 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_242), .ZN(n9664) );
  XOR2_X1 U10644 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_243), .Z(n9663) );
  XOR2_X1 U10645 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_244), .Z(n9662) );
  OAI211_X1 U10646 ( .C1(n9665), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9677)
         );
  INV_X1 U10647 ( .A(keyinput_248), .ZN(n9672) );
  AOI22_X1 U10648 ( .A1(n9668), .A2(keyinput_249), .B1(n9666), .B2(
        keyinput_248), .ZN(n9667) );
  OAI21_X1 U10649 ( .B1(n9668), .B2(keyinput_249), .A(n9667), .ZN(n9671) );
  XNOR2_X1 U10650 ( .A(n9669), .B(keyinput_247), .ZN(n9670) );
  AOI211_X1 U10651 ( .C1(P1_IR_REG_29__SCAN_IN), .C2(n9672), .A(n9671), .B(
        n9670), .ZN(n9676) );
  XOR2_X1 U10652 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_245), .Z(n9675) );
  XNOR2_X1 U10653 ( .A(n9673), .B(keyinput_246), .ZN(n9674) );
  NAND4_X1 U10654 ( .A1(n9677), .A2(n9676), .A3(n9675), .A4(n9674), .ZN(n9680)
         );
  XNOR2_X1 U10655 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_250), .ZN(n9679) );
  XNOR2_X1 U10656 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_251), .ZN(n9678) );
  AOI21_X1 U10657 ( .B1(n9680), .B2(n9679), .A(n9678), .ZN(n9683) );
  XNOR2_X1 U10658 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_252), .ZN(n9682) );
  XNOR2_X1 U10659 ( .A(n10599), .B(keyinput_253), .ZN(n9681) );
  OAI21_X1 U10660 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n9684) );
  NAND4_X1 U10661 ( .A1(n9687), .A2(n9686), .A3(n9685), .A4(n9684), .ZN(n9688)
         );
  XOR2_X1 U10662 ( .A(n9689), .B(n9688), .Z(P2_U3299) );
  INV_X1 U10663 ( .A(n9808), .ZN(n10597) );
  INV_X1 U10664 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9691) );
  NAND3_X1 U10665 ( .A1(n9691), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9693) );
  OAI22_X1 U10666 ( .A1(n9690), .A2(n9693), .B1(n9692), .B2(n9696), .ZN(n9694)
         );
  INV_X1 U10667 ( .A(n9694), .ZN(n9695) );
  OAI21_X1 U10668 ( .B1(n10597), .B2(n9699), .A(n9695), .ZN(P2_U3327) );
  OAI222_X1 U10669 ( .A1(n9699), .A2(n9820), .B1(n9698), .B2(P2_U3152), .C1(
        n9697), .C2(n9696), .ZN(P2_U3328) );
  MUX2_X1 U10670 ( .A(n9700), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10671 ( .A1(n5047), .A2(n9701), .ZN(n9703) );
  XNOR2_X1 U10672 ( .A(n9703), .B(n9702), .ZN(n9708) );
  OAI22_X1 U10673 ( .A1(n9798), .A2(n10342), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9704), .ZN(n9706) );
  OAI22_X1 U10674 ( .A1(n9800), .A2(n9722), .B1(n9799), .B2(n10371), .ZN(n9705) );
  AOI211_X1 U10675 ( .C1(n10508), .C2(n9803), .A(n9706), .B(n9705), .ZN(n9707)
         );
  OAI21_X1 U10676 ( .B1(n9708), .B2(n9805), .A(n9707), .ZN(P1_U3214) );
  OAI21_X1 U10677 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9712) );
  NAND2_X1 U10678 ( .A1(n9712), .A2(n9756), .ZN(n9717) );
  NOR2_X1 U10679 ( .A1(n9713), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10258) );
  INV_X1 U10680 ( .A(n10440), .ZN(n9714) );
  OAI22_X1 U10681 ( .A1(n9798), .A2(n9827), .B1(n9799), .B2(n9714), .ZN(n9715)
         );
  AOI211_X1 U10682 ( .C1(n9750), .C2(n10446), .A(n10258), .B(n9715), .ZN(n9716) );
  OAI211_X1 U10683 ( .C1(n10442), .C2(n9753), .A(n9717), .B(n9716), .ZN(
        P1_U3217) );
  NOR2_X1 U10684 ( .A1(n9718), .A2(n5097), .ZN(n9719) );
  XNOR2_X1 U10685 ( .A(n9720), .B(n9719), .ZN(n9727) );
  INV_X1 U10686 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9721) );
  OAI22_X1 U10687 ( .A1(n9798), .A2(n9722), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9721), .ZN(n9725) );
  INV_X1 U10688 ( .A(n9723), .ZN(n10410) );
  OAI22_X1 U10689 ( .A1(n9800), .A2(n9827), .B1(n9799), .B2(n10410), .ZN(n9724) );
  AOI211_X1 U10690 ( .C1(n10518), .C2(n9803), .A(n9725), .B(n9724), .ZN(n9726)
         );
  OAI21_X1 U10691 ( .B1(n9727), .B2(n9805), .A(n9726), .ZN(P1_U3221) );
  XNOR2_X1 U10692 ( .A(n9729), .B(n9728), .ZN(n9730) );
  XNOR2_X1 U10693 ( .A(n9731), .B(n9730), .ZN(n9736) );
  OAI22_X1 U10694 ( .A1(n9798), .A2(n10344), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9732), .ZN(n9734) );
  OAI22_X1 U10695 ( .A1(n9800), .A2(n10342), .B1(n9799), .B2(n10336), .ZN(
        n9733) );
  AOI211_X1 U10696 ( .C1(n10500), .C2(n9803), .A(n9734), .B(n9733), .ZN(n9735)
         );
  OAI21_X1 U10697 ( .B1(n9736), .B2(n9805), .A(n9735), .ZN(P1_U3223) );
  INV_X1 U10698 ( .A(n10557), .ZN(n11013) );
  NOR2_X1 U10699 ( .A1(n11013), .A2(n11029), .ZN(n10561) );
  INV_X1 U10700 ( .A(n10561), .ZN(n9744) );
  AOI21_X1 U10701 ( .B1(n9739), .B2(n9738), .A(n9737), .ZN(n9740) );
  OAI21_X1 U10702 ( .B1(n5537), .B2(n9740), .A(n9756), .ZN(n9743) );
  AND2_X1 U10703 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10203) );
  OAI22_X1 U10704 ( .A1(n9798), .A2(n10556), .B1(n9799), .B2(n11015), .ZN(
        n9741) );
  AOI211_X1 U10705 ( .C1(n9750), .C2(n10095), .A(n10203), .B(n9741), .ZN(n9742) );
  OAI211_X1 U10706 ( .C1(n9764), .C2(n9744), .A(n9743), .B(n9742), .ZN(
        P1_U3224) );
  INV_X1 U10707 ( .A(n10543), .ZN(n10467) );
  OAI21_X1 U10708 ( .B1(n9747), .B2(n9745), .A(n9746), .ZN(n9748) );
  NAND2_X1 U10709 ( .A1(n9748), .A2(n9756), .ZN(n9752) );
  AND2_X1 U10710 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10213) );
  OAI22_X1 U10711 ( .A1(n9798), .A2(n10454), .B1(n9799), .B2(n10462), .ZN(
        n9749) );
  AOI211_X1 U10712 ( .C1(n9750), .C2(n10094), .A(n10213), .B(n9749), .ZN(n9751) );
  OAI211_X1 U10713 ( .C1(n10467), .C2(n9753), .A(n9752), .B(n9751), .ZN(
        P1_U3226) );
  NAND2_X1 U10714 ( .A1(n10348), .A2(n10827), .ZN(n10504) );
  XNOR2_X1 U10715 ( .A(n9755), .B(n9754), .ZN(n9757) );
  NAND2_X1 U10716 ( .A1(n9757), .A2(n9756), .ZN(n9763) );
  INV_X1 U10717 ( .A(n10362), .ZN(n9758) );
  OAI22_X1 U10718 ( .A1(n10387), .A2(n9800), .B1(n9799), .B2(n9758), .ZN(n9761) );
  INV_X1 U10719 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9759) );
  OAI22_X1 U10720 ( .A1(n9798), .A2(n10321), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9759), .ZN(n9760) );
  NOR2_X1 U10721 ( .A1(n9761), .A2(n9760), .ZN(n9762) );
  OAI211_X1 U10722 ( .C1(n9764), .C2(n10504), .A(n9763), .B(n9762), .ZN(
        P1_U3227) );
  INV_X1 U10723 ( .A(n9765), .ZN(n9767) );
  NAND2_X1 U10724 ( .A1(n9767), .A2(n9766), .ZN(n9768) );
  XNOR2_X1 U10725 ( .A(n9769), .B(n9768), .ZN(n9775) );
  INV_X1 U10726 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9770) );
  OAI22_X1 U10727 ( .A1(n9800), .A2(n9790), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9770), .ZN(n9773) );
  OAI22_X1 U10728 ( .A1(n9798), .A2(n10385), .B1(n9799), .B2(n9771), .ZN(n9772) );
  AOI211_X1 U10729 ( .C1(n10526), .C2(n9803), .A(n9773), .B(n9772), .ZN(n9774)
         );
  OAI21_X1 U10730 ( .B1(n9775), .B2(n9805), .A(n9774), .ZN(P1_U3231) );
  NAND2_X1 U10731 ( .A1(n5080), .A2(n9776), .ZN(n9777) );
  XNOR2_X1 U10732 ( .A(n9778), .B(n9777), .ZN(n9783) );
  INV_X1 U10733 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9779) );
  OAI22_X1 U10734 ( .A1(n9798), .A2(n10387), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9779), .ZN(n9781) );
  OAI22_X1 U10735 ( .A1(n9800), .A2(n10385), .B1(n9799), .B2(n10390), .ZN(
        n9780) );
  AOI211_X1 U10736 ( .C1(n10515), .C2(n9803), .A(n9781), .B(n9780), .ZN(n9782)
         );
  OAI21_X1 U10737 ( .B1(n9783), .B2(n9805), .A(n9782), .ZN(P1_U3233) );
  AOI21_X1 U10738 ( .B1(n9786), .B2(n9788), .A(n9785), .ZN(n9787) );
  AOI21_X1 U10739 ( .B1(n5210), .B2(n9788), .A(n9787), .ZN(n9794) );
  NAND2_X1 U10740 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10243)
         );
  OAI21_X1 U10741 ( .B1(n9800), .B2(n10556), .A(n10243), .ZN(n9792) );
  OAI22_X1 U10742 ( .A1(n9798), .A2(n9790), .B1(n9799), .B2(n9789), .ZN(n9791)
         );
  AOI211_X1 U10743 ( .C1(n10538), .C2(n9803), .A(n9792), .B(n9791), .ZN(n9793)
         );
  OAI21_X1 U10744 ( .B1(n9794), .B2(n9805), .A(n9793), .ZN(P1_U3236) );
  XNOR2_X1 U10745 ( .A(n9796), .B(n9795), .ZN(n9806) );
  INV_X1 U10746 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9797) );
  OAI22_X1 U10747 ( .A1(n9798), .A2(n10322), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9797), .ZN(n9802) );
  OAI22_X1 U10748 ( .A1(n9800), .A2(n10321), .B1(n9799), .B2(n10327), .ZN(
        n9801) );
  AOI211_X1 U10749 ( .C1(n10493), .C2(n9803), .A(n9802), .B(n9801), .ZN(n9804)
         );
  OAI21_X1 U10750 ( .B1(n9806), .B2(n9805), .A(n9804), .ZN(P1_U3238) );
  NAND2_X1 U10751 ( .A1(n9808), .A2(n9807), .ZN(n9811) );
  INV_X1 U10752 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9809) );
  OR2_X1 U10753 ( .A1(n9822), .A2(n9809), .ZN(n9810) );
  NAND2_X1 U10754 ( .A1(n5033), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9818) );
  INV_X1 U10755 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9812) );
  OR2_X1 U10756 ( .A1(n9813), .A2(n9812), .ZN(n9817) );
  INV_X1 U10757 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9814) );
  OR2_X1 U10758 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  AND3_X1 U10759 ( .A1(n9818), .A2(n9817), .A3(n9816), .ZN(n10267) );
  NAND2_X1 U10760 ( .A1(n10473), .A2(n10267), .ZN(n10029) );
  OR2_X1 U10761 ( .A1(n9822), .A2(n9821), .ZN(n9823) );
  NAND2_X1 U10762 ( .A1(n11030), .A2(n10091), .ZN(n9913) );
  NAND2_X1 U10763 ( .A1(n10029), .A2(n9913), .ZN(n10064) );
  INV_X1 U10764 ( .A(n10064), .ZN(n9882) );
  INV_X1 U10765 ( .A(n9825), .ZN(n9826) );
  OR2_X1 U10766 ( .A1(n9918), .A2(n9826), .ZN(n10027) );
  AND2_X1 U10767 ( .A1(n10007), .A2(n10005), .ZN(n9872) );
  NAND4_X1 U10768 ( .A1(n9999), .A2(n9979), .A3(n9973), .A4(n9975), .ZN(n9829)
         );
  NAND3_X1 U10769 ( .A1(n9863), .A2(n9827), .A3(n10526), .ZN(n9828) );
  AND2_X1 U10770 ( .A1(n9828), .A2(n9988), .ZN(n9990) );
  NAND3_X1 U10771 ( .A1(n9990), .A2(n9996), .A3(n9984), .ZN(n9883) );
  OR2_X1 U10772 ( .A1(n9829), .A2(n9883), .ZN(n9869) );
  INV_X1 U10773 ( .A(n9869), .ZN(n9852) );
  NAND2_X1 U10774 ( .A1(n9831), .A2(n9830), .ZN(n9963) );
  NAND2_X1 U10775 ( .A1(n9970), .A2(n9963), .ZN(n9858) );
  INV_X1 U10776 ( .A(n9858), .ZN(n9899) );
  NAND2_X1 U10777 ( .A1(n9832), .A2(n9954), .ZN(n9855) );
  INV_X1 U10778 ( .A(n9945), .ZN(n9833) );
  INV_X1 U10779 ( .A(n9948), .ZN(n10921) );
  OAI211_X1 U10780 ( .C1(n9833), .C2(n9942), .A(n10921), .B(n9944), .ZN(n9834)
         );
  NOR2_X1 U10781 ( .A1(n9855), .A2(n9834), .ZN(n9898) );
  NAND2_X1 U10782 ( .A1(n6469), .A2(n9835), .ZN(n9838) );
  NAND2_X1 U10783 ( .A1(n10107), .A2(n9836), .ZN(n9837) );
  NAND3_X1 U10784 ( .A1(n9838), .A2(n9837), .A3(n9916), .ZN(n9840) );
  NAND2_X1 U10785 ( .A1(n9840), .A2(n9839), .ZN(n9842) );
  OAI211_X1 U10786 ( .C1(n9843), .C2(n9842), .A(n9885), .B(n9841), .ZN(n9846)
         );
  INV_X1 U10787 ( .A(n9844), .ZN(n9892) );
  NAND3_X1 U10788 ( .A1(n9846), .A2(n9892), .A3(n9845), .ZN(n9850) );
  INV_X1 U10789 ( .A(n9933), .ZN(n9847) );
  NOR2_X1 U10790 ( .A1(n9848), .A2(n9847), .ZN(n9849) );
  NAND2_X1 U10791 ( .A1(n9928), .A2(n9937), .ZN(n9895) );
  AOI21_X1 U10792 ( .B1(n9850), .B2(n9849), .A(n9895), .ZN(n9851) );
  NAND4_X1 U10793 ( .A1(n9852), .A2(n9899), .A3(n9898), .A4(n9851), .ZN(n9874)
         );
  NAND3_X1 U10794 ( .A1(n9945), .A2(n9938), .A3(n9941), .ZN(n9857) );
  NOR2_X1 U10795 ( .A1(n10564), .A2(n10928), .ZN(n9947) );
  INV_X1 U10796 ( .A(n9947), .ZN(n9853) );
  AND2_X1 U10797 ( .A1(n9952), .A2(n9853), .ZN(n9854) );
  OAI211_X1 U10798 ( .C1(n9855), .C2(n9854), .A(n9962), .B(n9953), .ZN(n9856)
         );
  AOI21_X1 U10799 ( .B1(n9898), .B2(n9857), .A(n9856), .ZN(n9859) );
  OAI211_X1 U10800 ( .C1(n9859), .C2(n9858), .A(n9969), .B(n9972), .ZN(n9860)
         );
  INV_X1 U10801 ( .A(n9860), .ZN(n9870) );
  NAND2_X1 U10802 ( .A1(n9980), .A2(n9976), .ZN(n9861) );
  NAND2_X1 U10803 ( .A1(n9861), .A2(n9979), .ZN(n9866) );
  INV_X1 U10804 ( .A(n9983), .ZN(n9864) );
  NAND2_X1 U10805 ( .A1(n9863), .A2(n9862), .ZN(n9989) );
  OAI211_X1 U10806 ( .C1(n9864), .C2(n9989), .A(n9990), .B(n9996), .ZN(n9865)
         );
  OAI211_X1 U10807 ( .C1(n9883), .C2(n9866), .A(n9995), .B(n9865), .ZN(n9867)
         );
  NAND2_X1 U10808 ( .A1(n9867), .A2(n9999), .ZN(n9868) );
  OAI211_X1 U10809 ( .C1(n9870), .C2(n9869), .A(n10001), .B(n9868), .ZN(n9871)
         );
  NAND2_X1 U10810 ( .A1(n9872), .A2(n9871), .ZN(n9873) );
  AND3_X1 U10811 ( .A1(n9921), .A2(n9873), .A3(n10008), .ZN(n9904) );
  OAI21_X1 U10812 ( .B1(n5391), .B2(n9874), .A(n9904), .ZN(n9876) );
  NAND2_X1 U10813 ( .A1(n9919), .A2(n9875), .ZN(n9907) );
  OAI21_X1 U10814 ( .B1(n9876), .B2(n10300), .A(n9907), .ZN(n9878) );
  AND2_X1 U10815 ( .A1(n10015), .A2(n9920), .ZN(n9908) );
  INV_X1 U10816 ( .A(n9908), .ZN(n9877) );
  NOR2_X1 U10817 ( .A1(n9878), .A2(n9877), .ZN(n9880) );
  INV_X1 U10818 ( .A(n10091), .ZN(n9879) );
  NAND2_X1 U10819 ( .A1(n10275), .A2(n9879), .ZN(n10060) );
  INV_X1 U10820 ( .A(n9910), .ZN(n10025) );
  OAI211_X1 U10821 ( .C1(n10027), .C2(n9880), .A(n10060), .B(n10025), .ZN(
        n9881) );
  INV_X1 U10822 ( .A(n10473), .ZN(n10271) );
  INV_X1 U10823 ( .A(n10267), .ZN(n10090) );
  AOI21_X1 U10824 ( .B1(n9882), .B2(n9881), .A(n10031), .ZN(n10079) );
  NOR2_X1 U10825 ( .A1(n10079), .A2(n10260), .ZN(n10078) );
  INV_X1 U10826 ( .A(n10027), .ZN(n9912) );
  INV_X1 U10827 ( .A(n9883), .ZN(n9903) );
  INV_X1 U10828 ( .A(n9975), .ZN(n9901) );
  NAND3_X1 U10829 ( .A1(n9886), .A2(n9885), .A3(n9884), .ZN(n9893) );
  NAND2_X1 U10830 ( .A1(n9888), .A2(n9887), .ZN(n9890) );
  NAND3_X1 U10831 ( .A1(n9890), .A2(n9889), .A3(n9923), .ZN(n9891) );
  NAND3_X1 U10832 ( .A1(n9893), .A2(n9892), .A3(n9891), .ZN(n9896) );
  AND2_X1 U10833 ( .A1(n9933), .A2(n9894), .ZN(n9927) );
  AOI21_X1 U10834 ( .B1(n9896), .B2(n9927), .A(n9895), .ZN(n9897) );
  NAND4_X1 U10835 ( .A1(n9973), .A2(n9899), .A3(n9898), .A4(n9897), .ZN(n9900)
         );
  NOR2_X1 U10836 ( .A1(n9901), .A2(n9900), .ZN(n9902) );
  NAND4_X1 U10837 ( .A1(n9903), .A2(n9902), .A3(n9979), .A4(n9999), .ZN(n9905)
         );
  OAI211_X1 U10838 ( .C1(n5391), .C2(n9905), .A(n9904), .B(n9919), .ZN(n9906)
         );
  NAND3_X1 U10839 ( .A1(n9908), .A2(n9907), .A3(n9906), .ZN(n9911) );
  NAND2_X1 U10840 ( .A1(n10275), .A2(n10267), .ZN(n9909) );
  NAND2_X1 U10841 ( .A1(n10060), .A2(n9909), .ZN(n10030) );
  AOI211_X1 U10842 ( .C1(n9912), .C2(n9911), .A(n9910), .B(n10030), .ZN(n9917)
         );
  INV_X1 U10843 ( .A(n9913), .ZN(n9914) );
  NAND2_X1 U10844 ( .A1(n9914), .A2(n10090), .ZN(n9915) );
  NAND2_X1 U10845 ( .A1(n10029), .A2(n9915), .ZN(n10021) );
  INV_X1 U10846 ( .A(n10031), .ZN(n10063) );
  AND2_X1 U10847 ( .A1(n10063), .A2(n9916), .ZN(n10070) );
  OAI21_X1 U10848 ( .B1(n9917), .B2(n10021), .A(n10070), .ZN(n10067) );
  NAND2_X1 U10849 ( .A1(n10064), .A2(n10473), .ZN(n10019) );
  NOR2_X1 U10850 ( .A1(n9918), .A2(n10024), .ZN(n10017) );
  INV_X1 U10851 ( .A(n10024), .ZN(n10020) );
  MUX2_X1 U10852 ( .A(n9920), .B(n9919), .S(n10020), .Z(n10014) );
  INV_X1 U10853 ( .A(n10300), .ZN(n10012) );
  MUX2_X1 U10854 ( .A(n10296), .B(n9921), .S(n10024), .Z(n10011) );
  INV_X1 U10855 ( .A(n9922), .ZN(n9924) );
  NAND2_X1 U10856 ( .A1(n9931), .A2(n9927), .ZN(n9929) );
  NAND2_X1 U10857 ( .A1(n9929), .A2(n9928), .ZN(n9936) );
  AOI21_X1 U10858 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(n9935) );
  MUX2_X1 U10859 ( .A(n9938), .B(n9937), .S(n10024), .Z(n9939) );
  MUX2_X1 U10860 ( .A(n9942), .B(n9941), .S(n10024), .Z(n9943) );
  MUX2_X1 U10861 ( .A(n9945), .B(n9944), .S(n10024), .Z(n9946) );
  MUX2_X1 U10862 ( .A(n9948), .B(n9947), .S(n10024), .Z(n9949) );
  NOR2_X1 U10863 ( .A1(n10913), .A2(n9949), .ZN(n9950) );
  NAND2_X1 U10864 ( .A1(n9951), .A2(n9950), .ZN(n9955) );
  AOI21_X1 U10865 ( .B1(n9955), .B2(n9952), .A(n9961), .ZN(n9957) );
  INV_X1 U10866 ( .A(n9953), .ZN(n9959) );
  AOI21_X1 U10867 ( .B1(n9955), .B2(n9954), .A(n9959), .ZN(n9956) );
  MUX2_X1 U10868 ( .A(n9957), .B(n9956), .S(n10024), .Z(n9958) );
  NAND2_X1 U10869 ( .A1(n9963), .A2(n9959), .ZN(n9960) );
  NAND2_X1 U10870 ( .A1(n9960), .A2(n9962), .ZN(n9966) );
  NAND2_X1 U10871 ( .A1(n9962), .A2(n9961), .ZN(n9964) );
  NAND2_X1 U10872 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  MUX2_X1 U10873 ( .A(n9966), .B(n9965), .S(n10024), .Z(n9967) );
  INV_X1 U10874 ( .A(n9967), .ZN(n9968) );
  MUX2_X1 U10875 ( .A(n9970), .B(n9969), .S(n10024), .Z(n9971) );
  MUX2_X1 U10876 ( .A(n9973), .B(n9972), .S(n10024), .Z(n9974) );
  MUX2_X1 U10877 ( .A(n9976), .B(n9975), .S(n10024), .Z(n9977) );
  MUX2_X1 U10878 ( .A(n9980), .B(n9979), .S(n10020), .Z(n9981) );
  INV_X1 U10879 ( .A(n10445), .ZN(n10436) );
  AOI21_X1 U10880 ( .B1(n9982), .B2(n9981), .A(n10436), .ZN(n9994) );
  INV_X1 U10881 ( .A(n10399), .ZN(n9987) );
  MUX2_X1 U10882 ( .A(n9984), .B(n9983), .S(n10024), .Z(n9985) );
  NAND3_X1 U10883 ( .A1(n9987), .A2(n9986), .A3(n9985), .ZN(n9993) );
  AND2_X1 U10884 ( .A1(n9995), .A2(n9996), .ZN(n10034) );
  NAND2_X1 U10885 ( .A1(n9989), .A2(n9988), .ZN(n9991) );
  MUX2_X1 U10886 ( .A(n9991), .B(n9990), .S(n10024), .Z(n9992) );
  OAI211_X1 U10887 ( .C1(n9994), .C2(n9993), .A(n10034), .B(n9992), .ZN(n9998)
         );
  INV_X1 U10888 ( .A(n10056), .ZN(n10375) );
  MUX2_X1 U10889 ( .A(n9996), .B(n9995), .S(n10024), .Z(n9997) );
  NAND3_X1 U10890 ( .A1(n9998), .A2(n10375), .A3(n9997), .ZN(n10003) );
  AND2_X1 U10891 ( .A1(n10005), .A2(n9999), .ZN(n10000) );
  MUX2_X1 U10892 ( .A(n10001), .B(n10000), .S(n10024), .Z(n10002) );
  MUX2_X1 U10893 ( .A(n10005), .B(n10004), .S(n10024), .Z(n10006) );
  INV_X1 U10894 ( .A(n10316), .ZN(n10010) );
  MUX2_X1 U10895 ( .A(n10008), .B(n10007), .S(n10024), .Z(n10009) );
  NAND3_X1 U10896 ( .A1(n10282), .A2(n10014), .A3(n10013), .ZN(n10023) );
  NAND3_X1 U10897 ( .A1(n10025), .A2(n10015), .A3(n10023), .ZN(n10016) );
  AOI21_X1 U10898 ( .B1(n10017), .B2(n10016), .A(n10030), .ZN(n10018) );
  NAND2_X1 U10899 ( .A1(n10021), .A2(n10020), .ZN(n10022) );
  INV_X1 U10900 ( .A(n10023), .ZN(n10026) );
  OAI211_X1 U10901 ( .C1(n10027), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10028) );
  OAI21_X1 U10902 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(n10032) );
  NOR4_X1 U10903 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10041) );
  NAND4_X1 U10904 ( .A1(n10041), .A2(n10040), .A3(n10765), .A4(n10039), .ZN(
        n10045) );
  NOR4_X1 U10905 ( .A1(n10045), .A2(n10044), .A3(n10043), .A4(n10042), .ZN(
        n10048) );
  INV_X1 U10906 ( .A(n10913), .ZN(n10923) );
  NAND4_X1 U10907 ( .A1(n10048), .A2(n10047), .A3(n10923), .A4(n10046), .ZN(
        n10050) );
  NOR3_X1 U10908 ( .A1(n10050), .A2(n5078), .A3(n10049), .ZN(n10051) );
  NAND4_X1 U10909 ( .A1(n10457), .A2(n10551), .A3(n10052), .A4(n10051), .ZN(
        n10053) );
  OR4_X1 U10910 ( .A1(n10399), .A2(n10436), .A3(n10054), .A4(n10053), .ZN(
        n10055) );
  NOR4_X1 U10911 ( .A1(n10056), .A2(n10383), .A3(n10419), .A4(n10055), .ZN(
        n10057) );
  XNOR2_X1 U10912 ( .A(n10348), .B(n10378), .ZN(n10353) );
  NAND3_X1 U10913 ( .A1(n10341), .A2(n10057), .A3(n10353), .ZN(n10058) );
  NOR4_X1 U10914 ( .A1(n10059), .A2(n10300), .A3(n10316), .A4(n10058), .ZN(
        n10061) );
  NAND4_X1 U10915 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n10065) );
  OAI21_X1 U10916 ( .B1(n10065), .B2(n10064), .A(n6947), .ZN(n10068) );
  MUX2_X1 U10917 ( .A(n10067), .B(n10066), .S(n10785), .Z(n10075) );
  INV_X1 U10918 ( .A(n10068), .ZN(n10069) );
  NAND2_X1 U10919 ( .A1(n10069), .A2(n10260), .ZN(n10074) );
  INV_X1 U10920 ( .A(n10070), .ZN(n10071) );
  NOR3_X1 U10921 ( .A1(n10072), .A2(n10086), .A3(n10071), .ZN(n10073) );
  AOI21_X1 U10922 ( .B1(n10075), .B2(n10074), .A(n10073), .ZN(n10077) );
  MUX2_X1 U10923 ( .A(n10078), .B(n10077), .S(n10076), .Z(n10089) );
  INV_X1 U10924 ( .A(n10079), .ZN(n10082) );
  OAI21_X1 U10925 ( .B1(n10082), .B2(n10081), .A(n10080), .ZN(n10088) );
  NAND4_X1 U10926 ( .A1(n10768), .A2(n10588), .A3(n10083), .A4(n10640), .ZN(
        n10084) );
  OAI211_X1 U10927 ( .C1(n10086), .C2(n10085), .A(n10084), .B(P1_B_REG_SCAN_IN), .ZN(n10087) );
  OAI21_X1 U10928 ( .B1(n10089), .B2(n10088), .A(n10087), .ZN(P1_U3240) );
  MUX2_X1 U10929 ( .A(n10090), .B(P1_DATAO_REG_31__SCAN_IN), .S(n10106), .Z(
        P1_U3586) );
  MUX2_X1 U10930 ( .A(n10091), .B(P1_DATAO_REG_30__SCAN_IN), .S(n10106), .Z(
        P1_U3585) );
  MUX2_X1 U10931 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10297), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10932 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10092), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10933 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10298), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10934 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10358), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10935 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10378), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10936 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10357), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10937 ( .A(n10404), .B(P1_DATAO_REG_22__SCAN_IN), .S(n10106), .Z(
        P1_U3577) );
  MUX2_X1 U10938 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10422), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10939 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10447), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10940 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10421), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10941 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10446), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10942 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10093), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10943 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10094), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10944 ( .A(n10095), .B(P1_DATAO_REG_15__SCAN_IN), .S(n10106), .Z(
        P1_U3570) );
  MUX2_X1 U10945 ( .A(n10096), .B(P1_DATAO_REG_14__SCAN_IN), .S(n10106), .Z(
        P1_U3569) );
  MUX2_X1 U10946 ( .A(n10097), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10106), .Z(
        P1_U3568) );
  MUX2_X1 U10947 ( .A(n10098), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10106), .Z(
        P1_U3567) );
  MUX2_X1 U10948 ( .A(n10099), .B(P1_DATAO_REG_11__SCAN_IN), .S(n10106), .Z(
        P1_U3566) );
  MUX2_X1 U10949 ( .A(n10100), .B(P1_DATAO_REG_10__SCAN_IN), .S(n10106), .Z(
        P1_U3565) );
  MUX2_X1 U10950 ( .A(n10101), .B(P1_DATAO_REG_9__SCAN_IN), .S(n10106), .Z(
        P1_U3564) );
  MUX2_X1 U10951 ( .A(n10102), .B(P1_DATAO_REG_8__SCAN_IN), .S(n10106), .Z(
        P1_U3563) );
  MUX2_X1 U10952 ( .A(n10103), .B(P1_DATAO_REG_7__SCAN_IN), .S(n10106), .Z(
        P1_U3562) );
  MUX2_X1 U10953 ( .A(n10770), .B(P1_DATAO_REG_6__SCAN_IN), .S(n10106), .Z(
        P1_U3561) );
  MUX2_X1 U10954 ( .A(n10104), .B(P1_DATAO_REG_5__SCAN_IN), .S(n10106), .Z(
        P1_U3560) );
  MUX2_X1 U10955 ( .A(n7834), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10106), .Z(
        P1_U3559) );
  MUX2_X1 U10956 ( .A(n10105), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10106), .Z(
        P1_U3558) );
  MUX2_X1 U10957 ( .A(n7832), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10106), .Z(
        P1_U3557) );
  MUX2_X1 U10958 ( .A(n10107), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10106), .Z(
        P1_U3556) );
  MUX2_X1 U10959 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6469), .S(P1_U4006), .Z(
        P1_U3555) );
  AOI211_X1 U10960 ( .C1(n10121), .C2(n10109), .A(n10108), .B(n10657), .ZN(
        n10110) );
  AOI21_X1 U10961 ( .B1(n10672), .B2(n10111), .A(n10110), .ZN(n10118) );
  AOI22_X1 U10962 ( .A1(n10667), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .ZN(n10117) );
  NAND2_X1 U10963 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10114) );
  AOI21_X1 U10964 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(n10115) );
  NAND2_X1 U10965 ( .A1(n10689), .A2(n10115), .ZN(n10116) );
  NAND3_X1 U10966 ( .A1(n10118), .A2(n10117), .A3(n10116), .ZN(P1_U3242) );
  AOI21_X1 U10967 ( .B1(n10640), .B2(n10119), .A(n6952), .ZN(n10639) );
  NOR2_X1 U10968 ( .A1(n10120), .A2(n6952), .ZN(n10123) );
  NOR2_X1 U10969 ( .A1(n6952), .A2(n10121), .ZN(n10122) );
  MUX2_X1 U10970 ( .A(n10123), .B(n10122), .S(n10640), .Z(n10124) );
  INV_X1 U10971 ( .A(n10124), .ZN(n10125) );
  OAI211_X1 U10972 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10639), .A(n10125), .B(
        P1_U4006), .ZN(n10167) );
  AOI211_X1 U10973 ( .C1(n10128), .C2(n10127), .A(n10126), .B(n10657), .ZN(
        n10129) );
  AOI21_X1 U10974 ( .B1(n10672), .B2(n10130), .A(n10129), .ZN(n10139) );
  AOI21_X1 U10975 ( .B1(n10133), .B2(n10132), .A(n10131), .ZN(n10137) );
  INV_X1 U10976 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10135) );
  OAI22_X1 U10977 ( .A1(n10679), .A2(n10135), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10134), .ZN(n10136) );
  AOI21_X1 U10978 ( .B1(n10689), .B2(n10137), .A(n10136), .ZN(n10138) );
  NAND3_X1 U10979 ( .A1(n10167), .A2(n10139), .A3(n10138), .ZN(P1_U3243) );
  AOI211_X1 U10980 ( .C1(n10142), .C2(n10141), .A(n10140), .B(n10657), .ZN(
        n10143) );
  AOI21_X1 U10981 ( .B1(n10672), .B2(n10144), .A(n10143), .ZN(n10151) );
  AOI21_X1 U10982 ( .B1(n10667), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n10145), .ZN(
        n10150) );
  OAI211_X1 U10983 ( .C1(n10148), .C2(n10147), .A(n10689), .B(n10146), .ZN(
        n10149) );
  NAND3_X1 U10984 ( .A1(n10151), .A2(n10150), .A3(n10149), .ZN(P1_U3244) );
  OAI21_X1 U10985 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(n10156) );
  AOI22_X1 U10986 ( .A1(n10690), .A2(n10156), .B1(n10672), .B2(n10155), .ZN(
        n10166) );
  INV_X1 U10987 ( .A(n10157), .ZN(n10160) );
  OAI21_X1 U10988 ( .B1(n10160), .B2(n10159), .A(n10158), .ZN(n10164) );
  INV_X1 U10989 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10161) );
  NOR2_X1 U10990 ( .A1(n10679), .A2(n10161), .ZN(n10162) );
  AOI211_X1 U10991 ( .C1(n10689), .C2(n10164), .A(n10163), .B(n10162), .ZN(
        n10165) );
  NAND3_X1 U10992 ( .A1(n10167), .A2(n10166), .A3(n10165), .ZN(P1_U3245) );
  OAI21_X1 U10993 ( .B1(n10170), .B2(n10169), .A(n10168), .ZN(n10171) );
  NAND2_X1 U10994 ( .A1(n10171), .A2(n10689), .ZN(n10180) );
  AOI21_X1 U10995 ( .B1(n10667), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n10172), .ZN(
        n10179) );
  AOI211_X1 U10996 ( .C1(n10175), .C2(n10174), .A(n10173), .B(n10657), .ZN(
        n10176) );
  AOI21_X1 U10997 ( .B1(n10672), .B2(n10177), .A(n10176), .ZN(n10178) );
  NAND3_X1 U10998 ( .A1(n10180), .A2(n10179), .A3(n10178), .ZN(P1_U3250) );
  INV_X1 U10999 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10187) );
  AOI21_X1 U11000 ( .B1(n10182), .B2(n8171), .A(n10181), .ZN(n10204) );
  XNOR2_X1 U11001 ( .A(n10194), .B(n10204), .ZN(n10183) );
  NAND2_X1 U11002 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10183), .ZN(n10206) );
  OAI211_X1 U11003 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n10183), .A(n10689), 
        .B(n10206), .ZN(n10186) );
  OR2_X1 U11004 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10184), .ZN(n10185) );
  OAI211_X1 U11005 ( .C1(n10187), .C2(n10679), .A(n10186), .B(n10185), .ZN(
        n10192) );
  AOI211_X1 U11006 ( .C1(n10190), .C2(n8499), .A(n10196), .B(n10657), .ZN(
        n10191) );
  AOI211_X1 U11007 ( .C1(n10672), .C2(n10205), .A(n10192), .B(n10191), .ZN(
        n10193) );
  INV_X1 U11008 ( .A(n10193), .ZN(P1_U3256) );
  NAND2_X1 U11009 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10222), .ZN(n10197) );
  OAI21_X1 U11010 ( .B1(n10222), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10197), 
        .ZN(n10198) );
  NOR2_X1 U11011 ( .A1(n10199), .A2(n10198), .ZN(n10216) );
  AOI211_X1 U11012 ( .C1(n10199), .C2(n10198), .A(n10216), .B(n10657), .ZN(
        n10200) );
  INV_X1 U11013 ( .A(n10200), .ZN(n10212) );
  INV_X1 U11014 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10201) );
  NOR2_X1 U11015 ( .A1(n10679), .A2(n10201), .ZN(n10202) );
  AOI211_X1 U11016 ( .C1(n10222), .C2(n10672), .A(n10203), .B(n10202), .ZN(
        n10211) );
  NAND2_X1 U11017 ( .A1(n10205), .A2(n10204), .ZN(n10207) );
  NAND2_X1 U11018 ( .A1(n10207), .A2(n10206), .ZN(n10209) );
  XOR2_X1 U11019 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10222), .Z(n10208) );
  NAND2_X1 U11020 ( .A1(n10208), .A2(n10209), .ZN(n10223) );
  OAI211_X1 U11021 ( .C1(n10209), .C2(n10208), .A(n10689), .B(n10223), .ZN(
        n10210) );
  NAND3_X1 U11022 ( .A1(n10212), .A2(n10211), .A3(n10210), .ZN(P1_U3257) );
  INV_X1 U11023 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10215) );
  INV_X1 U11024 ( .A(n10213), .ZN(n10214) );
  OAI21_X1 U11025 ( .B1(n10679), .B2(n10215), .A(n10214), .ZN(n10221) );
  AOI21_X1 U11026 ( .B1(n10222), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10216), 
        .ZN(n10219) );
  NAND2_X1 U11027 ( .A1(n10238), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10217) );
  OAI21_X1 U11028 ( .B1(n10238), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10217), 
        .ZN(n10218) );
  NOR2_X1 U11029 ( .A1(n10219), .A2(n10218), .ZN(n10237) );
  AOI211_X1 U11030 ( .C1(n10219), .C2(n10218), .A(n10237), .B(n10657), .ZN(
        n10220) );
  AOI211_X1 U11031 ( .C1(n10672), .C2(n10238), .A(n10221), .B(n10220), .ZN(
        n10229) );
  INV_X1 U11032 ( .A(n10238), .ZN(n10234) );
  XNOR2_X1 U11033 ( .A(n10234), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10227) );
  INV_X1 U11034 ( .A(n10222), .ZN(n10225) );
  OAI21_X1 U11035 ( .B1(n10225), .B2(n10224), .A(n10223), .ZN(n10226) );
  NAND2_X1 U11036 ( .A1(n10227), .A2(n10226), .ZN(n10232) );
  OAI211_X1 U11037 ( .C1(n10227), .C2(n10226), .A(n10689), .B(n10232), .ZN(
        n10228) );
  NAND2_X1 U11038 ( .A1(n10229), .A2(n10228), .ZN(P1_U3258) );
  INV_X1 U11039 ( .A(n10255), .ZN(n10231) );
  NAND2_X1 U11040 ( .A1(n10231), .A2(n10230), .ZN(n10251) );
  OAI21_X1 U11041 ( .B1(n10231), .B2(n10230), .A(n10251), .ZN(n10236) );
  OAI21_X1 U11042 ( .B1(n10234), .B2(n10233), .A(n10232), .ZN(n10235) );
  NOR2_X1 U11043 ( .A1(n10235), .A2(n10236), .ZN(n10249) );
  AOI21_X1 U11044 ( .B1(n10236), .B2(n10235), .A(n10249), .ZN(n10248) );
  AOI21_X1 U11045 ( .B1(n10238), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10237), 
        .ZN(n10241) );
  MUX2_X1 U11046 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n8585), .S(n10255), .Z(
        n10239) );
  INV_X1 U11047 ( .A(n10239), .ZN(n10240) );
  NOR2_X1 U11048 ( .A1(n10241), .A2(n10240), .ZN(n10254) );
  AOI211_X1 U11049 ( .C1(n10241), .C2(n10240), .A(n10254), .B(n10657), .ZN(
        n10242) );
  INV_X1 U11050 ( .A(n10242), .ZN(n10247) );
  INV_X1 U11051 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10244) );
  OAI21_X1 U11052 ( .B1(n10679), .B2(n10244), .A(n10243), .ZN(n10245) );
  AOI21_X1 U11053 ( .B1(n10255), .B2(n10672), .A(n10245), .ZN(n10246) );
  OAI211_X1 U11054 ( .C1(n10248), .C2(n10264), .A(n10247), .B(n10246), .ZN(
        P1_U3259) );
  INV_X1 U11055 ( .A(n10249), .ZN(n10250) );
  NAND2_X1 U11056 ( .A1(n10251), .A2(n10250), .ZN(n10253) );
  XNOR2_X1 U11057 ( .A(n10785), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10252) );
  XNOR2_X1 U11058 ( .A(n10253), .B(n10252), .ZN(n10263) );
  INV_X1 U11059 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10256) );
  MUX2_X1 U11060 ( .A(n10256), .B(P1_REG2_REG_19__SCAN_IN), .S(n10260), .Z(
        n10257) );
  INV_X1 U11061 ( .A(n10672), .ZN(n10261) );
  AOI21_X1 U11062 ( .B1(n10667), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n10258), 
        .ZN(n10259) );
  OAI21_X1 U11063 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(n10262) );
  XNOR2_X1 U11064 ( .A(n10273), .B(n10473), .ZN(n10472) );
  NAND2_X1 U11065 ( .A1(n10472), .A2(n10470), .ZN(n10270) );
  INV_X1 U11066 ( .A(n10265), .ZN(n10266) );
  NOR2_X1 U11067 ( .A1(n10267), .A2(n10266), .ZN(n11032) );
  INV_X1 U11068 ( .A(n11032), .ZN(n10268) );
  NOR2_X1 U11069 ( .A1(n10268), .A2(n10465), .ZN(n10276) );
  AOI21_X1 U11070 ( .B1(n10789), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10276), 
        .ZN(n10269) );
  OAI211_X1 U11071 ( .C1(n10271), .C2(n11012), .A(n10270), .B(n10269), .ZN(
        P1_U3261) );
  INV_X1 U11072 ( .A(n10272), .ZN(n10274) );
  NAND2_X1 U11073 ( .A1(n11034), .A2(n10470), .ZN(n10278) );
  AOI21_X1 U11074 ( .B1(n10789), .B2(P1_REG2_REG_30__SCAN_IN), .A(n10276), 
        .ZN(n10277) );
  OAI211_X1 U11075 ( .C1(n11030), .C2(n11012), .A(n10278), .B(n10277), .ZN(
        P1_U3262) );
  AND2_X1 U11076 ( .A1(n10279), .A2(n10282), .ZN(n10280) );
  XNOR2_X1 U11077 ( .A(n10283), .B(n10282), .ZN(n10286) );
  OAI22_X1 U11078 ( .A1(n10284), .A2(n10925), .B1(n10322), .B2(n10927), .ZN(
        n10285) );
  OAI22_X1 U11079 ( .A1(n11019), .A2(n10288), .B1(n10287), .B2(n11014), .ZN(
        n10289) );
  AOI21_X1 U11080 ( .B1(n10481), .B2(n10413), .A(n10289), .ZN(n10293) );
  NAND2_X1 U11081 ( .A1(n10303), .A2(n10481), .ZN(n10290) );
  NAND2_X1 U11082 ( .A1(n10482), .A2(n10470), .ZN(n10292) );
  OAI211_X1 U11083 ( .C1(n10484), .C2(n10789), .A(n10293), .B(n10292), .ZN(
        n10294) );
  INV_X1 U11084 ( .A(n10294), .ZN(n10295) );
  OAI21_X1 U11085 ( .B1(n10485), .B2(n11021), .A(n10295), .ZN(P1_U3263) );
  OAI21_X1 U11086 ( .B1(n10301), .B2(n10300), .A(n10299), .ZN(n10486) );
  NAND2_X1 U11087 ( .A1(n10486), .A2(n10302), .ZN(n10312) );
  INV_X1 U11088 ( .A(n10325), .ZN(n10305) );
  INV_X1 U11089 ( .A(n10303), .ZN(n10304) );
  AOI211_X1 U11090 ( .C1(n10488), .C2(n10305), .A(n10990), .B(n10304), .ZN(
        n10487) );
  NOR2_X1 U11091 ( .A1(n10306), .A2(n11012), .ZN(n10310) );
  OAI22_X1 U11092 ( .A1(n11019), .A2(n10308), .B1(n10307), .B2(n11014), .ZN(
        n10309) );
  AOI211_X1 U11093 ( .C1(n10487), .C2(n11023), .A(n10310), .B(n10309), .ZN(
        n10311) );
  OAI211_X1 U11094 ( .C1(n10789), .C2(n10490), .A(n10312), .B(n10311), .ZN(
        P1_U3264) );
  INV_X1 U11095 ( .A(n10315), .ZN(n10318) );
  OAI21_X1 U11096 ( .B1(n10318), .B2(n10317), .A(n10316), .ZN(n10320) );
  AOI21_X1 U11097 ( .B1(n10320), .B2(n10319), .A(n10554), .ZN(n10324) );
  OAI22_X1 U11098 ( .A1(n10322), .A2(n10925), .B1(n10321), .B2(n10927), .ZN(
        n10323) );
  AOI211_X1 U11099 ( .C1(n10492), .C2(n10426), .A(n10324), .B(n10323), .ZN(
        n10496) );
  AOI21_X1 U11100 ( .B1(n10493), .B2(n10334), .A(n10325), .ZN(n10494) );
  INV_X1 U11101 ( .A(n10493), .ZN(n10326) );
  NOR2_X1 U11102 ( .A1(n10326), .A2(n11012), .ZN(n10330) );
  OAI22_X1 U11103 ( .A1(n11019), .A2(n10328), .B1(n10327), .B2(n11014), .ZN(
        n10329) );
  AOI211_X1 U11104 ( .C1(n10494), .C2(n10470), .A(n10330), .B(n10329), .ZN(
        n10332) );
  NAND2_X1 U11105 ( .A1(n10492), .A2(n10433), .ZN(n10331) );
  OAI211_X1 U11106 ( .C1(n10496), .C2(n10789), .A(n10332), .B(n10331), .ZN(
        P1_U3265) );
  XOR2_X1 U11107 ( .A(n10341), .B(n10333), .Z(n10502) );
  INV_X1 U11108 ( .A(n10334), .ZN(n10335) );
  AOI211_X1 U11109 ( .C1(n10500), .C2(n10349), .A(n10990), .B(n10335), .ZN(
        n10499) );
  NOR2_X1 U11110 ( .A1(n5343), .A2(n11012), .ZN(n10339) );
  OAI22_X1 U11111 ( .A1(n11019), .A2(n10337), .B1(n10336), .B2(n11014), .ZN(
        n10338) );
  AOI211_X1 U11112 ( .C1(n10499), .C2(n11023), .A(n10339), .B(n10338), .ZN(
        n10346) );
  XOR2_X1 U11113 ( .A(n10341), .B(n10340), .Z(n10343) );
  OAI222_X1 U11114 ( .A1(n10925), .A2(n10344), .B1(n10343), .B2(n10554), .C1(
        n10927), .C2(n10342), .ZN(n10498) );
  NAND2_X1 U11115 ( .A1(n10498), .A2(n11019), .ZN(n10345) );
  OAI211_X1 U11116 ( .C1(n10502), .C2(n11021), .A(n10346), .B(n10345), .ZN(
        P1_U3266) );
  XNOR2_X1 U11117 ( .A(n10347), .B(n10353), .ZN(n10507) );
  AOI22_X1 U11118 ( .A1(n10348), .A2(n10413), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10465), .ZN(n10366) );
  AOI21_X1 U11119 ( .B1(n10368), .B2(n10348), .A(n10990), .ZN(n10350) );
  NAND2_X1 U11120 ( .A1(n10350), .A2(n10349), .ZN(n10503) );
  NAND2_X1 U11121 ( .A1(n10352), .A2(n10351), .ZN(n10355) );
  INV_X1 U11122 ( .A(n10353), .ZN(n10354) );
  XNOR2_X1 U11123 ( .A(n10355), .B(n10354), .ZN(n10356) );
  NAND2_X1 U11124 ( .A1(n10356), .A2(n10930), .ZN(n10506) );
  NAND2_X1 U11125 ( .A1(n10357), .A2(n10768), .ZN(n10360) );
  NAND2_X1 U11126 ( .A1(n10358), .A2(n10769), .ZN(n10359) );
  AND2_X1 U11127 ( .A1(n10360), .A2(n10359), .ZN(n10505) );
  INV_X1 U11128 ( .A(n10505), .ZN(n10361) );
  AOI21_X1 U11129 ( .B1(n10362), .B2(n10463), .A(n10361), .ZN(n10363) );
  OAI211_X1 U11130 ( .C1(n10785), .C2(n10503), .A(n10506), .B(n10363), .ZN(
        n10364) );
  NAND2_X1 U11131 ( .A1(n10364), .A2(n11019), .ZN(n10365) );
  OAI211_X1 U11132 ( .C1(n10507), .C2(n11021), .A(n10366), .B(n10365), .ZN(
        P1_U3267) );
  XNOR2_X1 U11133 ( .A(n10367), .B(n10375), .ZN(n10512) );
  INV_X1 U11134 ( .A(n10388), .ZN(n10370) );
  INV_X1 U11135 ( .A(n10368), .ZN(n10369) );
  AOI21_X1 U11136 ( .B1(n10508), .B2(n10370), .A(n10369), .ZN(n10509) );
  INV_X1 U11137 ( .A(n10371), .ZN(n10372) );
  AOI22_X1 U11138 ( .A1(n10465), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10372), 
        .B2(n10463), .ZN(n10373) );
  OAI21_X1 U11139 ( .B1(n10374), .B2(n11012), .A(n10373), .ZN(n10380) );
  XNOR2_X1 U11140 ( .A(n10376), .B(n10375), .ZN(n10377) );
  AOI222_X1 U11141 ( .A1(n10404), .A2(n10768), .B1(n10378), .B2(n10769), .C1(
        n10930), .C2(n10377), .ZN(n10511) );
  NOR2_X1 U11142 ( .A1(n10511), .A2(n10465), .ZN(n10379) );
  AOI211_X1 U11143 ( .C1(n10509), .C2(n10470), .A(n10380), .B(n10379), .ZN(
        n10381) );
  OAI21_X1 U11144 ( .B1(n10512), .B2(n11021), .A(n10381), .ZN(P1_U3268) );
  XNOR2_X1 U11145 ( .A(n10382), .B(n10383), .ZN(n10517) );
  XNOR2_X1 U11146 ( .A(n10384), .B(n10383), .ZN(n10386) );
  OAI222_X1 U11147 ( .A1(n10925), .A2(n10387), .B1(n10386), .B2(n10554), .C1(
        n10927), .C2(n10385), .ZN(n10513) );
  INV_X1 U11148 ( .A(n10409), .ZN(n10389) );
  AOI211_X1 U11149 ( .C1(n10515), .C2(n10389), .A(n10990), .B(n10388), .ZN(
        n10514) );
  NAND2_X1 U11150 ( .A1(n10514), .A2(n11023), .ZN(n10393) );
  INV_X1 U11151 ( .A(n10390), .ZN(n10391) );
  AOI22_X1 U11152 ( .A1(n10465), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10391), 
        .B2(n10463), .ZN(n10392) );
  OAI211_X1 U11153 ( .C1(n10394), .C2(n11012), .A(n10393), .B(n10392), .ZN(
        n10395) );
  AOI21_X1 U11154 ( .B1(n10513), .B2(n11019), .A(n10395), .ZN(n10396) );
  OAI21_X1 U11155 ( .B1(n10517), .B2(n11021), .A(n10396), .ZN(P1_U3269) );
  OAI21_X1 U11156 ( .B1(n10398), .B2(n10399), .A(n10397), .ZN(n10524) );
  NAND2_X1 U11157 ( .A1(n10400), .A2(n10399), .ZN(n10401) );
  NAND2_X1 U11158 ( .A1(n10402), .A2(n10401), .ZN(n10403) );
  NAND2_X1 U11159 ( .A1(n10403), .A2(n10930), .ZN(n10406) );
  AOI22_X1 U11160 ( .A1(n10768), .A2(n10447), .B1(n10404), .B2(n10769), .ZN(
        n10405) );
  NAND2_X1 U11161 ( .A1(n10406), .A2(n10405), .ZN(n10522) );
  NAND2_X1 U11162 ( .A1(n10427), .A2(n10518), .ZN(n10407) );
  NAND2_X1 U11163 ( .A1(n10407), .A2(n11033), .ZN(n10408) );
  OR2_X1 U11164 ( .A1(n10409), .A2(n10408), .ZN(n10520) );
  OAI22_X1 U11165 ( .A1(n11019), .A2(n10411), .B1(n10410), .B2(n11014), .ZN(
        n10412) );
  AOI21_X1 U11166 ( .B1(n10518), .B2(n10413), .A(n10412), .ZN(n10414) );
  OAI21_X1 U11167 ( .B1(n10520), .B2(n10937), .A(n10414), .ZN(n10415) );
  AOI21_X1 U11168 ( .B1(n10522), .B2(n11019), .A(n10415), .ZN(n10416) );
  OAI21_X1 U11169 ( .B1(n10524), .B2(n11021), .A(n10416), .ZN(P1_U3270) );
  INV_X1 U11170 ( .A(n10417), .ZN(n10418) );
  OAI21_X1 U11171 ( .B1(n10418), .B2(n10419), .A(n5429), .ZN(n10525) );
  XNOR2_X1 U11172 ( .A(n10420), .B(n10419), .ZN(n10424) );
  AOI22_X1 U11173 ( .A1(n10422), .A2(n10769), .B1(n10768), .B2(n10421), .ZN(
        n10423) );
  OAI21_X1 U11174 ( .B1(n10424), .B2(n10554), .A(n10423), .ZN(n10425) );
  AOI21_X1 U11175 ( .B1(n10525), .B2(n10426), .A(n10425), .ZN(n10529) );
  INV_X1 U11176 ( .A(n10526), .ZN(n10431) );
  AOI21_X1 U11177 ( .B1(n10526), .B2(n10438), .A(n5351), .ZN(n10527) );
  NAND2_X1 U11178 ( .A1(n10527), .A2(n10470), .ZN(n10430) );
  AOI22_X1 U11179 ( .A1(n10465), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10428), 
        .B2(n10463), .ZN(n10429) );
  OAI211_X1 U11180 ( .C1(n10431), .C2(n11012), .A(n10430), .B(n10429), .ZN(
        n10432) );
  AOI21_X1 U11181 ( .B1(n10525), .B2(n10433), .A(n10432), .ZN(n10434) );
  OAI21_X1 U11182 ( .B1(n10529), .B2(n10789), .A(n10434), .ZN(P1_U3271) );
  XNOR2_X1 U11183 ( .A(n10435), .B(n10436), .ZN(n10535) );
  INV_X1 U11184 ( .A(n10437), .ZN(n10439) );
  AOI211_X1 U11185 ( .C1(n10532), .C2(n10439), .A(n10990), .B(n5352), .ZN(
        n10531) );
  AOI22_X1 U11186 ( .A1(n10465), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10440), 
        .B2(n10463), .ZN(n10441) );
  OAI21_X1 U11187 ( .B1(n10442), .B2(n11012), .A(n10441), .ZN(n10450) );
  OAI21_X1 U11188 ( .B1(n10445), .B2(n10444), .A(n10443), .ZN(n10448) );
  AOI222_X1 U11189 ( .A1(n10930), .A2(n10448), .B1(n10447), .B2(n10769), .C1(
        n10446), .C2(n10768), .ZN(n10534) );
  NOR2_X1 U11190 ( .A1(n10534), .A2(n10465), .ZN(n10449) );
  AOI211_X1 U11191 ( .C1(n10531), .C2(n11023), .A(n10450), .B(n10449), .ZN(
        n10451) );
  OAI21_X1 U11192 ( .B1(n10535), .B2(n11021), .A(n10451), .ZN(P1_U3272) );
  XOR2_X1 U11193 ( .A(n10457), .B(n10452), .Z(n10460) );
  OAI22_X1 U11194 ( .A1(n10454), .A2(n10925), .B1(n10453), .B2(n10927), .ZN(
        n10459) );
  AOI21_X1 U11195 ( .B1(n10457), .B2(n10456), .A(n10455), .ZN(n10547) );
  NOR2_X1 U11196 ( .A1(n10547), .A2(n7857), .ZN(n10458) );
  AOI211_X1 U11197 ( .C1(n10930), .C2(n10460), .A(n10459), .B(n10458), .ZN(
        n10546) );
  AOI21_X1 U11198 ( .B1(n10543), .B2(n10559), .A(n10461), .ZN(n10544) );
  INV_X1 U11199 ( .A(n10462), .ZN(n10464) );
  AOI22_X1 U11200 ( .A1(n10465), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10464), 
        .B2(n10463), .ZN(n10466) );
  OAI21_X1 U11201 ( .B1(n10467), .B2(n11012), .A(n10466), .ZN(n10469) );
  NOR2_X1 U11202 ( .A1(n10547), .A2(n10938), .ZN(n10468) );
  AOI211_X1 U11203 ( .C1(n10544), .C2(n10470), .A(n10469), .B(n10468), .ZN(
        n10471) );
  OAI21_X1 U11204 ( .B1(n10546), .B2(n10465), .A(n10471), .ZN(P1_U3274) );
  NAND2_X1 U11205 ( .A1(n10472), .A2(n11033), .ZN(n10475) );
  AOI21_X1 U11206 ( .B1(n10473), .B2(n10827), .A(n11032), .ZN(n10474) );
  NAND2_X1 U11207 ( .A1(n10475), .A2(n10474), .ZN(n10569) );
  MUX2_X1 U11208 ( .A(n10569), .B(P1_REG1_REG_31__SCAN_IN), .S(n11035), .Z(
        P1_U3554) );
  AND2_X1 U11209 ( .A1(n7857), .A2(n10718), .ZN(n10832) );
  AOI22_X1 U11210 ( .A1(n10477), .A2(n11033), .B1(n10827), .B2(n10476), .ZN(
        n10478) );
  OAI211_X1 U11211 ( .C1(n10480), .C2(n10832), .A(n10479), .B(n10478), .ZN(
        n10570) );
  MUX2_X1 U11212 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10570), .S(n11036), .Z(
        P1_U3552) );
  AOI22_X1 U11213 ( .A1(n10482), .A2(n11033), .B1(n10827), .B2(n10481), .ZN(
        n10483) );
  OAI211_X1 U11214 ( .C1(n10485), .C2(n10832), .A(n10484), .B(n10483), .ZN(
        n10571) );
  MUX2_X1 U11215 ( .A(n10571), .B(P1_REG1_REG_28__SCAN_IN), .S(n11035), .Z(
        P1_U3551) );
  INV_X1 U11216 ( .A(n10486), .ZN(n10491) );
  AOI21_X1 U11217 ( .B1(n10827), .B2(n10488), .A(n10487), .ZN(n10489) );
  OAI211_X1 U11218 ( .C1(n10491), .C2(n10832), .A(n10490), .B(n10489), .ZN(
        n10572) );
  MUX2_X1 U11219 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10572), .S(n11036), .Z(
        P1_U3550) );
  INV_X1 U11220 ( .A(n10492), .ZN(n10497) );
  AOI22_X1 U11221 ( .A1(n10494), .A2(n11033), .B1(n10827), .B2(n10493), .ZN(
        n10495) );
  OAI211_X1 U11222 ( .C1(n10497), .C2(n10718), .A(n10496), .B(n10495), .ZN(
        n10573) );
  MUX2_X1 U11223 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10573), .S(n11036), .Z(
        P1_U3549) );
  AOI211_X1 U11224 ( .C1(n10827), .C2(n10500), .A(n10499), .B(n10498), .ZN(
        n10501) );
  OAI21_X1 U11225 ( .B1(n10502), .B2(n10832), .A(n10501), .ZN(n10574) );
  MUX2_X1 U11226 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10574), .S(n11036), .Z(
        P1_U3548) );
  OAI21_X1 U11227 ( .B1(n10507), .B2(n10832), .A(n5048), .ZN(n10575) );
  MUX2_X1 U11228 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10575), .S(n11036), .Z(
        P1_U3547) );
  AOI22_X1 U11229 ( .A1(n10509), .A2(n11033), .B1(n10827), .B2(n10508), .ZN(
        n10510) );
  OAI211_X1 U11230 ( .C1(n10512), .C2(n10832), .A(n10511), .B(n10510), .ZN(
        n10576) );
  MUX2_X1 U11231 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10576), .S(n11036), .Z(
        P1_U3546) );
  AOI211_X1 U11232 ( .C1(n10827), .C2(n10515), .A(n10514), .B(n10513), .ZN(
        n10516) );
  OAI21_X1 U11233 ( .B1(n10517), .B2(n10832), .A(n10516), .ZN(n10577) );
  MUX2_X1 U11234 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10577), .S(n11036), .Z(
        P1_U3545) );
  NAND2_X1 U11235 ( .A1(n10518), .A2(n10827), .ZN(n10519) );
  NAND2_X1 U11236 ( .A1(n10520), .A2(n10519), .ZN(n10521) );
  NOR2_X1 U11237 ( .A1(n10522), .A2(n10521), .ZN(n10523) );
  OAI21_X1 U11238 ( .B1(n10524), .B2(n10832), .A(n10523), .ZN(n10578) );
  MUX2_X1 U11239 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10578), .S(n11036), .Z(
        P1_U3544) );
  INV_X1 U11240 ( .A(n10525), .ZN(n10530) );
  AOI22_X1 U11241 ( .A1(n10527), .A2(n11033), .B1(n10827), .B2(n10526), .ZN(
        n10528) );
  OAI211_X1 U11242 ( .C1(n10530), .C2(n10718), .A(n10529), .B(n10528), .ZN(
        n10579) );
  MUX2_X1 U11243 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10579), .S(n11036), .Z(
        P1_U3543) );
  AOI21_X1 U11244 ( .B1(n10827), .B2(n10532), .A(n10531), .ZN(n10533) );
  OAI211_X1 U11245 ( .C1(n10535), .C2(n10832), .A(n10534), .B(n10533), .ZN(
        n10580) );
  MUX2_X1 U11246 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10580), .S(n11036), .Z(
        P1_U3542) );
  INV_X1 U11247 ( .A(n10536), .ZN(n10542) );
  INV_X1 U11248 ( .A(n10537), .ZN(n10539) );
  AOI22_X1 U11249 ( .A1(n10539), .A2(n11033), .B1(n10827), .B2(n10538), .ZN(
        n10540) );
  OAI211_X1 U11250 ( .C1(n10718), .C2(n10542), .A(n10541), .B(n10540), .ZN(
        n10581) );
  MUX2_X1 U11251 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10581), .S(n11036), .Z(
        P1_U3541) );
  AOI22_X1 U11252 ( .A1(n10544), .A2(n11033), .B1(n10827), .B2(n10543), .ZN(
        n10545) );
  OAI211_X1 U11253 ( .C1(n10547), .C2(n10718), .A(n10546), .B(n10545), .ZN(
        n10582) );
  MUX2_X1 U11254 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10582), .S(n11036), .Z(
        P1_U3540) );
  OAI21_X1 U11255 ( .B1(n10550), .B2(n10549), .A(n10548), .ZN(n11022) );
  XNOR2_X1 U11256 ( .A(n10552), .B(n10551), .ZN(n10553) );
  OAI222_X1 U11257 ( .A1(n10925), .A2(n10556), .B1(n10927), .B2(n10555), .C1(
        n10554), .C2(n10553), .ZN(n11020) );
  AOI21_X1 U11258 ( .B1(n10558), .B2(n10557), .A(n10990), .ZN(n10560) );
  AND2_X1 U11259 ( .A1(n10560), .A2(n10559), .ZN(n11024) );
  NOR3_X1 U11260 ( .A1(n11020), .A2(n10561), .A3(n11024), .ZN(n10562) );
  OAI21_X1 U11261 ( .B1(n11022), .B2(n10832), .A(n10562), .ZN(n10583) );
  MUX2_X1 U11262 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10583), .S(n11036), .Z(
        P1_U3539) );
  INV_X1 U11263 ( .A(n10563), .ZN(n10568) );
  AOI22_X1 U11264 ( .A1(n10565), .A2(n11033), .B1(n10827), .B2(n10564), .ZN(
        n10566) );
  OAI211_X1 U11265 ( .C1(n10718), .C2(n10568), .A(n10567), .B(n10566), .ZN(
        n10584) );
  MUX2_X1 U11266 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10584), .S(n11036), .Z(
        P1_U3534) );
  MUX2_X1 U11267 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10569), .S(n11040), .Z(
        P1_U3522) );
  MUX2_X1 U11268 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10570), .S(n11040), .Z(
        P1_U3520) );
  MUX2_X1 U11269 ( .A(n10571), .B(P1_REG0_REG_28__SCAN_IN), .S(n11037), .Z(
        P1_U3519) );
  MUX2_X1 U11270 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10572), .S(n11040), .Z(
        P1_U3518) );
  MUX2_X1 U11271 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10573), .S(n11040), .Z(
        P1_U3517) );
  MUX2_X1 U11272 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10574), .S(n11040), .Z(
        P1_U3516) );
  MUX2_X1 U11273 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10575), .S(n11040), .Z(
        P1_U3515) );
  MUX2_X1 U11274 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10576), .S(n11040), .Z(
        P1_U3514) );
  MUX2_X1 U11275 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10577), .S(n11040), .Z(
        P1_U3513) );
  MUX2_X1 U11276 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10578), .S(n11040), .Z(
        P1_U3512) );
  MUX2_X1 U11277 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10579), .S(n11040), .Z(
        P1_U3511) );
  MUX2_X1 U11278 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10580), .S(n11040), .Z(
        P1_U3510) );
  MUX2_X1 U11279 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10581), .S(n11040), .Z(
        P1_U3508) );
  MUX2_X1 U11280 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10582), .S(n11040), .Z(
        P1_U3505) );
  MUX2_X1 U11281 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10583), .S(n11040), .Z(
        P1_U3502) );
  MUX2_X1 U11282 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10584), .S(n11040), .Z(
        P1_U3487) );
  MUX2_X1 U11283 ( .A(n10586), .B(P1_D_REG_1__SCAN_IN), .S(n10585), .Z(
        P1_U3441) );
  INV_X1 U11284 ( .A(n10587), .ZN(n10589) );
  AND2_X1 U11285 ( .A1(n10589), .A2(n10588), .ZN(n10600) );
  MUX2_X1 U11286 ( .A(P1_D_REG_0__SCAN_IN), .B(n10590), .S(n10600), .Z(
        P1_U3440) );
  INV_X1 U11287 ( .A(n10591), .ZN(n10592) );
  NOR4_X1 U11288 ( .A1(n10592), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n6577), .ZN(n10593) );
  AOI21_X1 U11289 ( .B1(n10594), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10593), 
        .ZN(n10595) );
  OAI21_X1 U11290 ( .B1(n10597), .B2(n10596), .A(n10595), .ZN(P1_U3322) );
  MUX2_X1 U11291 ( .A(n10598), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11292 ( .A1(n10600), .A2(n10599), .ZN(P1_U3321) );
  AND2_X1 U11293 ( .A1(n10601), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U11294 ( .A1(n10601), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  AND2_X1 U11295 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10601), .ZN(P1_U3318) );
  AND2_X1 U11296 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10601), .ZN(P1_U3317) );
  AND2_X1 U11297 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10601), .ZN(P1_U3316) );
  AND2_X1 U11298 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10601), .ZN(P1_U3315) );
  AND2_X1 U11299 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10601), .ZN(P1_U3314) );
  AND2_X1 U11300 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10601), .ZN(P1_U3313) );
  AND2_X1 U11301 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10601), .ZN(P1_U3312) );
  AND2_X1 U11302 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10601), .ZN(P1_U3311) );
  AND2_X1 U11303 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10601), .ZN(P1_U3310) );
  AND2_X1 U11304 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10601), .ZN(P1_U3309) );
  AND2_X1 U11305 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10601), .ZN(P1_U3308) );
  AND2_X1 U11306 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10601), .ZN(P1_U3307) );
  AND2_X1 U11307 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10601), .ZN(P1_U3306) );
  AND2_X1 U11308 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10601), .ZN(P1_U3305) );
  AND2_X1 U11309 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10601), .ZN(P1_U3304) );
  AND2_X1 U11310 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10601), .ZN(P1_U3303) );
  AND2_X1 U11311 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10601), .ZN(P1_U3302) );
  AND2_X1 U11312 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10601), .ZN(P1_U3301) );
  AND2_X1 U11313 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10601), .ZN(P1_U3300) );
  AND2_X1 U11314 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10601), .ZN(P1_U3299) );
  AND2_X1 U11315 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10601), .ZN(P1_U3298) );
  AND2_X1 U11316 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10601), .ZN(P1_U3297) );
  AND2_X1 U11317 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10601), .ZN(P1_U3296) );
  AND2_X1 U11318 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10601), .ZN(P1_U3295) );
  AND2_X1 U11319 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10601), .ZN(P1_U3294) );
  AND2_X1 U11320 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10601), .ZN(P1_U3293) );
  AND2_X1 U11321 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10601), .ZN(P1_U3292) );
  AND2_X1 U11322 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10602), .ZN(P2_U3326) );
  AND2_X1 U11323 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10602), .ZN(P2_U3325) );
  AND2_X1 U11324 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10602), .ZN(P2_U3324) );
  AND2_X1 U11325 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10602), .ZN(P2_U3323) );
  AND2_X1 U11326 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10602), .ZN(P2_U3322) );
  AND2_X1 U11327 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10602), .ZN(P2_U3321) );
  AND2_X1 U11328 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10602), .ZN(P2_U3320) );
  AND2_X1 U11329 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10602), .ZN(P2_U3319) );
  AND2_X1 U11330 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10602), .ZN(P2_U3318) );
  AND2_X1 U11331 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10602), .ZN(P2_U3317) );
  AND2_X1 U11332 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10602), .ZN(P2_U3316) );
  AND2_X1 U11333 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10602), .ZN(P2_U3315) );
  AND2_X1 U11334 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10602), .ZN(P2_U3314) );
  AND2_X1 U11335 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10602), .ZN(P2_U3313) );
  AND2_X1 U11336 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10602), .ZN(P2_U3312) );
  AND2_X1 U11337 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10602), .ZN(P2_U3311) );
  AND2_X1 U11338 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10602), .ZN(P2_U3310) );
  AND2_X1 U11339 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10602), .ZN(P2_U3309) );
  AND2_X1 U11340 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10602), .ZN(P2_U3308) );
  AND2_X1 U11341 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10602), .ZN(P2_U3307) );
  AND2_X1 U11342 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10602), .ZN(P2_U3306) );
  AND2_X1 U11343 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10602), .ZN(P2_U3305) );
  AND2_X1 U11344 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10602), .ZN(P2_U3304) );
  AND2_X1 U11345 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10602), .ZN(P2_U3303) );
  AND2_X1 U11346 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10602), .ZN(P2_U3302) );
  AND2_X1 U11347 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10602), .ZN(P2_U3301) );
  AND2_X1 U11348 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10602), .ZN(P2_U3300) );
  AND2_X1 U11349 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10602), .ZN(P2_U3298) );
  AND2_X1 U11350 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10602), .ZN(P2_U3297) );
  XOR2_X1 U11351 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11352 ( .A(n10603), .ZN(n10604) );
  NAND2_X1 U11353 ( .A1(n10605), .A2(n10604), .ZN(n10606) );
  XNOR2_X1 U11354 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10606), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11355 ( .A(n10608), .B(n10607), .Z(ADD_1071_U54) );
  XOR2_X1 U11356 ( .A(n10610), .B(n10609), .Z(ADD_1071_U53) );
  XNOR2_X1 U11357 ( .A(n10612), .B(n10611), .ZN(ADD_1071_U52) );
  NOR2_X1 U11358 ( .A1(n10614), .A2(n10613), .ZN(n10615) );
  XOR2_X1 U11359 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10615), .Z(ADD_1071_U51) );
  XOR2_X1 U11360 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10616), .Z(ADD_1071_U50) );
  XOR2_X1 U11361 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10617), .Z(ADD_1071_U49) );
  XOR2_X1 U11362 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10618), .Z(ADD_1071_U48) );
  XOR2_X1 U11363 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10619), .Z(ADD_1071_U47) );
  XOR2_X1 U11364 ( .A(n10621), .B(n10620), .Z(ADD_1071_U63) );
  XOR2_X1 U11365 ( .A(n10623), .B(n10622), .Z(ADD_1071_U62) );
  XNOR2_X1 U11366 ( .A(n10625), .B(n10624), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11367 ( .A(n10627), .B(n10626), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11368 ( .A(n10629), .B(n10628), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11369 ( .A(n10631), .B(n10630), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11370 ( .A(n10633), .B(n10632), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11371 ( .A(n10635), .B(n10634), .ZN(ADD_1071_U56) );
  NOR2_X1 U11372 ( .A1(n10637), .A2(n10636), .ZN(n10638) );
  XOR2_X1 U11373 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10638), .Z(ADD_1071_U55)
         );
  OAI21_X1 U11374 ( .B1(n10640), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10639), .ZN(
        n10641) );
  XOR2_X1 U11375 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10641), .Z(n10644) );
  AOI22_X1 U11376 ( .A1(n10667), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10642) );
  OAI21_X1 U11377 ( .B1(n10644), .B2(n10643), .A(n10642), .ZN(P1_U3241) );
  AOI211_X1 U11378 ( .C1(n10647), .C2(n10646), .A(n10645), .B(n10657), .ZN(
        n10648) );
  AOI211_X1 U11379 ( .C1(n10672), .C2(n10650), .A(n10649), .B(n10648), .ZN(
        n10656) );
  AOI21_X1 U11380 ( .B1(n10653), .B2(n10652), .A(n10651), .ZN(n10654) );
  AOI22_X1 U11381 ( .A1(n10654), .A2(n10689), .B1(n10667), .B2(
        P1_ADDR_REG_6__SCAN_IN), .ZN(n10655) );
  NAND2_X1 U11382 ( .A1(n10656), .A2(n10655), .ZN(P1_U3247) );
  AOI211_X1 U11383 ( .C1(n10660), .C2(n10659), .A(n10658), .B(n10657), .ZN(
        n10661) );
  AOI211_X1 U11384 ( .C1(n10663), .C2(n10672), .A(n10662), .B(n10661), .ZN(
        n10670) );
  OAI21_X1 U11385 ( .B1(n10666), .B2(n10665), .A(n10664), .ZN(n10668) );
  AOI22_X1 U11386 ( .A1(n10668), .A2(n10689), .B1(n10667), .B2(
        P1_ADDR_REG_10__SCAN_IN), .ZN(n10669) );
  NAND2_X1 U11387 ( .A1(n10670), .A2(n10669), .ZN(P1_U3251) );
  INV_X1 U11388 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10671) );
  NOR2_X1 U11389 ( .A1(n10671), .A2(n10686), .ZN(n10673) );
  AOI21_X1 U11390 ( .B1(n10689), .B2(n10673), .A(n10672), .ZN(n10695) );
  INV_X1 U11391 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10678) );
  INV_X1 U11392 ( .A(n10674), .ZN(n10677) );
  NAND3_X1 U11393 ( .A1(n10675), .A2(n10682), .A3(n5159), .ZN(n10676) );
  OAI211_X1 U11394 ( .C1(n10679), .C2(n10678), .A(n10677), .B(n10676), .ZN(
        n10680) );
  INV_X1 U11395 ( .A(n10680), .ZN(n10693) );
  AOI211_X1 U11396 ( .C1(n10684), .C2(n10683), .A(n10682), .B(n10681), .ZN(
        n10691) );
  AOI21_X1 U11397 ( .B1(n10687), .B2(n10686), .A(n10685), .ZN(n10688) );
  AOI22_X1 U11398 ( .A1(n10691), .A2(n10690), .B1(n10689), .B2(n10688), .ZN(
        n10692) );
  OAI211_X1 U11399 ( .C1(n10695), .C2(n10694), .A(n10693), .B(n10692), .ZN(
        P1_U3252) );
  XNOR2_X1 U11400 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11401 ( .A(n10696), .ZN(n10697) );
  OAI211_X1 U11402 ( .C1(n10699), .C2(n10718), .A(n10698), .B(n10697), .ZN(
        n10700) );
  NOR2_X1 U11403 ( .A1(n10701), .A2(n10700), .ZN(n10704) );
  AOI22_X1 U11404 ( .A1(n11036), .A2(n10704), .B1(n10702), .B2(n11035), .ZN(
        P1_U3524) );
  INV_X1 U11405 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U11406 ( .A1(n11040), .A2(n10704), .B1(n10703), .B2(n11037), .ZN(
        P1_U3457) );
  INV_X1 U11407 ( .A(n10832), .ZN(n10977) );
  OAI21_X1 U11408 ( .B1(n10706), .B2(n10990), .A(n10705), .ZN(n10708) );
  AOI211_X1 U11409 ( .C1(n10977), .C2(n10709), .A(n10708), .B(n10707), .ZN(
        n10712) );
  AOI22_X1 U11410 ( .A1(n11036), .A2(n10712), .B1(n10710), .B2(n11035), .ZN(
        P1_U3525) );
  INV_X1 U11411 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U11412 ( .A1(n11040), .A2(n10712), .B1(n10711), .B2(n11037), .ZN(
        P1_U3460) );
  OAI22_X1 U11413 ( .A1(n10713), .A2(n11000), .B1(n7609), .B2(n10998), .ZN(
        n10715) );
  AOI211_X1 U11414 ( .C1(n10901), .C2(n10716), .A(n10715), .B(n10714), .ZN(
        n10717) );
  AOI22_X1 U11415 ( .A1(n11007), .A2(n10717), .B1(n7306), .B2(n11006), .ZN(
        P2_U3522) );
  AOI22_X1 U11416 ( .A1(n11011), .A2(n10717), .B1(n5609), .B2(n11008), .ZN(
        P2_U3457) );
  INV_X1 U11417 ( .A(n10718), .ZN(n10995) );
  OAI22_X1 U11418 ( .A1(n10720), .A2(n10990), .B1(n10719), .B2(n11029), .ZN(
        n10721) );
  AOI21_X1 U11419 ( .B1(n10722), .B2(n10995), .A(n10721), .ZN(n10723) );
  AND2_X1 U11420 ( .A1(n10724), .A2(n10723), .ZN(n10726) );
  AOI22_X1 U11421 ( .A1(n11036), .A2(n10726), .B1(n7246), .B2(n11035), .ZN(
        P1_U3526) );
  INV_X1 U11422 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U11423 ( .A1(n11040), .A2(n10726), .B1(n10725), .B2(n11037), .ZN(
        P1_U3463) );
  OAI211_X1 U11424 ( .C1(n10729), .C2(n5099), .A(n10728), .B(n10727), .ZN(
        n10740) );
  AOI22_X1 U11425 ( .A1(n10731), .A2(n10730), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10735) );
  NAND2_X1 U11426 ( .A1(n10733), .A2(n10732), .ZN(n10734) );
  OAI211_X1 U11427 ( .C1(n10737), .C2(n10736), .A(n10735), .B(n10734), .ZN(
        n10738) );
  INV_X1 U11428 ( .A(n10738), .ZN(n10739) );
  AND2_X1 U11429 ( .A1(n10740), .A2(n10739), .ZN(n10741) );
  OAI21_X1 U11430 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n10742), .A(n10741), .ZN(
        P2_U3220) );
  OAI22_X1 U11431 ( .A1(n10744), .A2(n10990), .B1(n10743), .B2(n11029), .ZN(
        n10745) );
  AOI21_X1 U11432 ( .B1(n10746), .B2(n10977), .A(n10745), .ZN(n10747) );
  AND2_X1 U11433 ( .A1(n10748), .A2(n10747), .ZN(n10751) );
  INV_X1 U11434 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U11435 ( .A1(n11036), .A2(n10751), .B1(n10749), .B2(n11035), .ZN(
        P1_U3527) );
  INV_X1 U11436 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U11437 ( .A1(n11040), .A2(n10751), .B1(n10750), .B2(n11037), .ZN(
        P1_U3466) );
  OAI22_X1 U11438 ( .A1(n10753), .A2(n11000), .B1(n10752), .B2(n10998), .ZN(
        n10755) );
  AOI211_X1 U11439 ( .C1(n11004), .C2(n10756), .A(n10755), .B(n10754), .ZN(
        n10757) );
  AOI22_X1 U11440 ( .A1(n11007), .A2(n10757), .B1(n7407), .B2(n11006), .ZN(
        P2_U3524) );
  AOI22_X1 U11441 ( .A1(n11011), .A2(n10757), .B1(n5639), .B2(n11008), .ZN(
        P2_U3463) );
  NAND2_X1 U11442 ( .A1(n7904), .A2(n10765), .ZN(n10758) );
  AND2_X1 U11443 ( .A1(n10759), .A2(n10758), .ZN(n10777) );
  NAND2_X1 U11444 ( .A1(n10760), .A2(n10781), .ZN(n10761) );
  NAND2_X1 U11445 ( .A1(n10761), .A2(n11033), .ZN(n10763) );
  OR2_X1 U11446 ( .A1(n10763), .A2(n10762), .ZN(n10784) );
  OAI21_X1 U11447 ( .B1(n10764), .B2(n11029), .A(n10784), .ZN(n10773) );
  XNOR2_X1 U11448 ( .A(n10766), .B(n10765), .ZN(n10767) );
  NAND2_X1 U11449 ( .A1(n10767), .A2(n10930), .ZN(n10772) );
  AOI22_X1 U11450 ( .A1(n10770), .A2(n10769), .B1(n10768), .B2(n7834), .ZN(
        n10771) );
  NAND2_X1 U11451 ( .A1(n10772), .A2(n10771), .ZN(n10786) );
  AOI211_X1 U11452 ( .C1(n10777), .C2(n10977), .A(n10773), .B(n10786), .ZN(
        n10775) );
  AOI22_X1 U11453 ( .A1(n11036), .A2(n10775), .B1(n6532), .B2(n11035), .ZN(
        P1_U3528) );
  INV_X1 U11454 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U11455 ( .A1(n11040), .A2(n10775), .B1(n10774), .B2(n11037), .ZN(
        P1_U3469) );
  NAND2_X1 U11456 ( .A1(n10777), .A2(n10776), .ZN(n10783) );
  NOR2_X1 U11457 ( .A1(n11014), .A2(n10778), .ZN(n10779) );
  AOI21_X1 U11458 ( .B1(n10781), .B2(n10780), .A(n10779), .ZN(n10782) );
  OAI211_X1 U11459 ( .C1(n10785), .C2(n10784), .A(n10783), .B(n10782), .ZN(
        n10787) );
  NOR2_X1 U11460 ( .A1(n10787), .A2(n10786), .ZN(n10788) );
  AOI22_X1 U11461 ( .A1(n10789), .A2(n6530), .B1(n10788), .B2(n11019), .ZN(
        P1_U3286) );
  NAND2_X1 U11462 ( .A1(n10791), .A2(n10790), .ZN(n10792) );
  XNOR2_X1 U11463 ( .A(n10793), .B(n10792), .ZN(n10818) );
  AND2_X1 U11464 ( .A1(n10818), .A2(n10794), .ZN(n10814) );
  OAI21_X1 U11465 ( .B1(n10797), .B2(n10796), .A(n10795), .ZN(n10799) );
  NAND2_X1 U11466 ( .A1(n10799), .A2(n10798), .ZN(n10801) );
  NAND2_X1 U11467 ( .A1(n10801), .A2(n10800), .ZN(n10822) );
  XNOR2_X1 U11468 ( .A(n10802), .B(n10820), .ZN(n10804) );
  NAND2_X1 U11469 ( .A1(n10804), .A2(n10803), .ZN(n10819) );
  NAND2_X1 U11470 ( .A1(n10806), .A2(n10805), .ZN(n10807) );
  OAI21_X1 U11471 ( .B1(n10809), .B2(n10808), .A(n10807), .ZN(n10810) );
  INV_X1 U11472 ( .A(n10810), .ZN(n10811) );
  OAI21_X1 U11473 ( .B1(n10819), .B2(n10812), .A(n10811), .ZN(n10813) );
  NOR3_X1 U11474 ( .A1(n10814), .A2(n10822), .A3(n10813), .ZN(n10816) );
  AOI22_X1 U11475 ( .A1(n10817), .A2(n5659), .B1(n10816), .B2(n10815), .ZN(
        P2_U3291) );
  AND2_X1 U11476 ( .A1(n10818), .A2(n11004), .ZN(n10823) );
  OAI21_X1 U11477 ( .B1(n10820), .B2(n10998), .A(n10819), .ZN(n10821) );
  NOR3_X1 U11478 ( .A1(n10823), .A2(n10822), .A3(n10821), .ZN(n10825) );
  AOI22_X1 U11479 ( .A1(n11007), .A2(n10825), .B1(n7408), .B2(n11006), .ZN(
        P2_U3525) );
  INV_X1 U11480 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U11481 ( .A1(n11011), .A2(n10825), .B1(n10824), .B2(n11008), .ZN(
        P2_U3466) );
  AOI22_X1 U11482 ( .A1(n10828), .A2(n11033), .B1(n10827), .B2(n10826), .ZN(
        n10829) );
  OAI211_X1 U11483 ( .C1(n10832), .C2(n10831), .A(n10830), .B(n10829), .ZN(
        n10833) );
  INV_X1 U11484 ( .A(n10833), .ZN(n10835) );
  AOI22_X1 U11485 ( .A1(n11036), .A2(n10835), .B1(n6550), .B2(n11035), .ZN(
        P1_U3529) );
  INV_X1 U11486 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U11487 ( .A1(n11040), .A2(n10835), .B1(n10834), .B2(n11037), .ZN(
        P1_U3472) );
  AND3_X1 U11488 ( .A1(n10837), .A2(n11004), .A3(n10836), .ZN(n10842) );
  OAI22_X1 U11489 ( .A1(n10839), .A2(n11000), .B1(n10838), .B2(n10998), .ZN(
        n10840) );
  NOR3_X1 U11490 ( .A1(n10842), .A2(n10841), .A3(n10840), .ZN(n10844) );
  AOI22_X1 U11491 ( .A1(n11007), .A2(n10844), .B1(n7436), .B2(n11006), .ZN(
        P2_U3526) );
  INV_X1 U11492 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U11493 ( .A1(n11011), .A2(n10844), .B1(n10843), .B2(n11008), .ZN(
        P2_U3469) );
  OAI21_X1 U11494 ( .B1(n10846), .B2(n11029), .A(n10845), .ZN(n10847) );
  AOI21_X1 U11495 ( .B1(n10848), .B2(n10995), .A(n10847), .ZN(n10849) );
  AND2_X1 U11496 ( .A1(n10850), .A2(n10849), .ZN(n10852) );
  AOI22_X1 U11497 ( .A1(n11036), .A2(n10852), .B1(n7271), .B2(n11035), .ZN(
        P1_U3530) );
  INV_X1 U11498 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U11499 ( .A1(n11040), .A2(n10852), .B1(n10851), .B2(n11037), .ZN(
        P1_U3475) );
  OAI22_X1 U11500 ( .A1(n10854), .A2(n11000), .B1(n10853), .B2(n10998), .ZN(
        n10856) );
  AOI211_X1 U11501 ( .C1(n11004), .C2(n10857), .A(n10856), .B(n10855), .ZN(
        n10859) );
  AOI22_X1 U11502 ( .A1(n11007), .A2(n10859), .B1(n7439), .B2(n11006), .ZN(
        P2_U3527) );
  INV_X1 U11503 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U11504 ( .A1(n11011), .A2(n10859), .B1(n10858), .B2(n11008), .ZN(
        P2_U3472) );
  INV_X1 U11505 ( .A(n10860), .ZN(n10865) );
  OAI22_X1 U11506 ( .A1(n10862), .A2(n10990), .B1(n10861), .B2(n11029), .ZN(
        n10864) );
  AOI211_X1 U11507 ( .C1(n10995), .C2(n10865), .A(n10864), .B(n10863), .ZN(
        n10867) );
  AOI22_X1 U11508 ( .A1(n11036), .A2(n10867), .B1(n6585), .B2(n11035), .ZN(
        P1_U3531) );
  INV_X1 U11509 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U11510 ( .A1(n11040), .A2(n10867), .B1(n10866), .B2(n11037), .ZN(
        P1_U3478) );
  INV_X1 U11511 ( .A(n10868), .ZN(n10873) );
  NAND3_X1 U11512 ( .A1(n10870), .A2(n11004), .A3(n10869), .ZN(n10872) );
  OAI211_X1 U11513 ( .C1(n10873), .C2(n10998), .A(n10872), .B(n10871), .ZN(
        n10874) );
  NOR2_X1 U11514 ( .A1(n10875), .A2(n10874), .ZN(n10877) );
  AOI22_X1 U11515 ( .A1(n11007), .A2(n10877), .B1(n7440), .B2(n11006), .ZN(
        P2_U3528) );
  INV_X1 U11516 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U11517 ( .A1(n11011), .A2(n10877), .B1(n10876), .B2(n11008), .ZN(
        P2_U3475) );
  INV_X1 U11518 ( .A(n10878), .ZN(n10884) );
  INV_X1 U11519 ( .A(n10879), .ZN(n10880) );
  OAI22_X1 U11520 ( .A1(n10881), .A2(n11000), .B1(n10880), .B2(n10998), .ZN(
        n10883) );
  AOI211_X1 U11521 ( .C1(n10901), .C2(n10884), .A(n10883), .B(n10882), .ZN(
        n10886) );
  AOI22_X1 U11522 ( .A1(n11007), .A2(n10886), .B1(n7470), .B2(n11006), .ZN(
        P2_U3529) );
  INV_X1 U11523 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U11524 ( .A1(n11011), .A2(n10886), .B1(n10885), .B2(n11008), .ZN(
        P2_U3478) );
  OAI21_X1 U11525 ( .B1(n10888), .B2(n11029), .A(n10887), .ZN(n10889) );
  AOI21_X1 U11526 ( .B1(n10890), .B2(n10995), .A(n10889), .ZN(n10891) );
  AND2_X1 U11527 ( .A1(n10892), .A2(n10891), .ZN(n10894) );
  AOI22_X1 U11528 ( .A1(n11036), .A2(n10894), .B1(n6624), .B2(n11035), .ZN(
        P1_U3533) );
  INV_X1 U11529 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U11530 ( .A1(n11040), .A2(n10894), .B1(n10893), .B2(n11037), .ZN(
        P1_U3484) );
  INV_X1 U11531 ( .A(n10895), .ZN(n10900) );
  OAI22_X1 U11532 ( .A1(n10897), .A2(n11000), .B1(n10896), .B2(n10998), .ZN(
        n10899) );
  AOI211_X1 U11533 ( .C1(n10901), .C2(n10900), .A(n10899), .B(n10898), .ZN(
        n10903) );
  AOI22_X1 U11534 ( .A1(n11007), .A2(n10903), .B1(n7530), .B2(n11006), .ZN(
        P2_U3530) );
  INV_X1 U11535 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U11536 ( .A1(n11011), .A2(n10903), .B1(n10902), .B2(n11008), .ZN(
        P2_U3481) );
  NAND2_X1 U11537 ( .A1(n10905), .A2(n10904), .ZN(n10907) );
  OAI211_X1 U11538 ( .C1(n10908), .C2(n10962), .A(n10907), .B(n10906), .ZN(
        n10910) );
  NOR2_X1 U11539 ( .A1(n10910), .A2(n10909), .ZN(n10912) );
  AOI22_X1 U11540 ( .A1(n11007), .A2(n10912), .B1(n7555), .B2(n11006), .ZN(
        P2_U3531) );
  INV_X1 U11541 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U11542 ( .A1(n11011), .A2(n10912), .B1(n10911), .B2(n11008), .ZN(
        P2_U3484) );
  OR2_X1 U11543 ( .A1(n10914), .A2(n10913), .ZN(n10915) );
  NAND2_X1 U11544 ( .A1(n10916), .A2(n10915), .ZN(n10939) );
  INV_X1 U11545 ( .A(n10939), .ZN(n10934) );
  AOI21_X1 U11546 ( .B1(n10918), .B2(n10917), .A(n10990), .ZN(n10920) );
  NAND2_X1 U11547 ( .A1(n10920), .A2(n10919), .ZN(n10936) );
  OAI21_X1 U11548 ( .B1(n5350), .B2(n11029), .A(n10936), .ZN(n10933) );
  NAND2_X1 U11549 ( .A1(n10922), .A2(n10921), .ZN(n10924) );
  XNOR2_X1 U11550 ( .A(n10924), .B(n10923), .ZN(n10931) );
  OAI22_X1 U11551 ( .A1(n10928), .A2(n10927), .B1(n10926), .B2(n10925), .ZN(
        n10929) );
  AOI21_X1 U11552 ( .B1(n10931), .B2(n10930), .A(n10929), .ZN(n10932) );
  OAI21_X1 U11553 ( .B1(n10939), .B2(n7857), .A(n10932), .ZN(n10945) );
  AOI211_X1 U11554 ( .C1(n10995), .C2(n10934), .A(n10933), .B(n10945), .ZN(
        n10935) );
  AOI22_X1 U11555 ( .A1(n11036), .A2(n10935), .B1(n7675), .B2(n11035), .ZN(
        P1_U3535) );
  AOI22_X1 U11556 ( .A1(n11040), .A2(n10935), .B1(n6662), .B2(n11037), .ZN(
        P1_U3490) );
  OAI22_X1 U11557 ( .A1(n10939), .A2(n10938), .B1(n10937), .B2(n10936), .ZN(
        n10940) );
  INV_X1 U11558 ( .A(n10940), .ZN(n10947) );
  NOR2_X1 U11559 ( .A1(n5350), .A2(n11012), .ZN(n10944) );
  INV_X1 U11560 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10942) );
  OAI22_X1 U11561 ( .A1(n11019), .A2(n10942), .B1(n10941), .B2(n11014), .ZN(
        n10943) );
  AOI211_X1 U11562 ( .C1(n10945), .C2(n11019), .A(n10944), .B(n10943), .ZN(
        n10946) );
  NAND2_X1 U11563 ( .A1(n10947), .A2(n10946), .ZN(P1_U3279) );
  INV_X1 U11564 ( .A(n10948), .ZN(n10953) );
  OAI22_X1 U11565 ( .A1(n10950), .A2(n11000), .B1(n10949), .B2(n10998), .ZN(
        n10951) );
  AOI211_X1 U11566 ( .C1(n10953), .C2(n11004), .A(n10952), .B(n10951), .ZN(
        n10955) );
  AOI22_X1 U11567 ( .A1(n11007), .A2(n10955), .B1(n5786), .B2(n11006), .ZN(
        P2_U3532) );
  INV_X1 U11568 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U11569 ( .A1(n11011), .A2(n10955), .B1(n10954), .B2(n11008), .ZN(
        P2_U3487) );
  OAI22_X1 U11570 ( .A1(n10956), .A2(n10990), .B1(n5349), .B2(n11029), .ZN(
        n10958) );
  AOI211_X1 U11571 ( .C1(n10995), .C2(n10959), .A(n10958), .B(n10957), .ZN(
        n10961) );
  AOI22_X1 U11572 ( .A1(n11036), .A2(n10961), .B1(n7863), .B2(n11035), .ZN(
        P1_U3536) );
  INV_X1 U11573 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U11574 ( .A1(n11040), .A2(n10961), .B1(n10960), .B2(n11037), .ZN(
        P1_U3493) );
  NOR2_X1 U11575 ( .A1(n10963), .A2(n10962), .ZN(n10969) );
  OAI22_X1 U11576 ( .A1(n10965), .A2(n11000), .B1(n10964), .B2(n10998), .ZN(
        n10967) );
  AOI211_X1 U11577 ( .C1(n10969), .C2(n10968), .A(n10967), .B(n10966), .ZN(
        n10971) );
  AOI22_X1 U11578 ( .A1(n11007), .A2(n10971), .B1(n5849), .B2(n11006), .ZN(
        P2_U3533) );
  INV_X1 U11579 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U11580 ( .A1(n11011), .A2(n10971), .B1(n10970), .B2(n11008), .ZN(
        P2_U3490) );
  OAI211_X1 U11581 ( .C1(n10974), .C2(n11029), .A(n10973), .B(n10972), .ZN(
        n10975) );
  AOI21_X1 U11582 ( .B1(n10977), .B2(n10976), .A(n10975), .ZN(n10979) );
  AOI22_X1 U11583 ( .A1(n11036), .A2(n10979), .B1(n8171), .B2(n11035), .ZN(
        P1_U3537) );
  INV_X1 U11584 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U11585 ( .A1(n11040), .A2(n10979), .B1(n10978), .B2(n11037), .ZN(
        P1_U3496) );
  INV_X1 U11586 ( .A(n10980), .ZN(n10985) );
  OAI22_X1 U11587 ( .A1(n10982), .A2(n11000), .B1(n10981), .B2(n10998), .ZN(
        n10983) );
  AOI211_X1 U11588 ( .C1(n10985), .C2(n11004), .A(n10984), .B(n10983), .ZN(
        n10987) );
  AOI22_X1 U11589 ( .A1(n11007), .A2(n10987), .B1(n5864), .B2(n11006), .ZN(
        P2_U3534) );
  INV_X1 U11590 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U11591 ( .A1(n11011), .A2(n10987), .B1(n10986), .B2(n11008), .ZN(
        P2_U3493) );
  INV_X1 U11592 ( .A(n10988), .ZN(n10994) );
  OAI22_X1 U11593 ( .A1(n10991), .A2(n10990), .B1(n10989), .B2(n11029), .ZN(
        n10993) );
  AOI211_X1 U11594 ( .C1(n10995), .C2(n10994), .A(n10993), .B(n10992), .ZN(
        n10997) );
  AOI22_X1 U11595 ( .A1(n11036), .A2(n10997), .B1(n6721), .B2(n11035), .ZN(
        P1_U3538) );
  INV_X1 U11596 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U11597 ( .A1(n11040), .A2(n10997), .B1(n10996), .B2(n11037), .ZN(
        P1_U3499) );
  OAI22_X1 U11598 ( .A1(n11001), .A2(n11000), .B1(n10999), .B2(n10998), .ZN(
        n11002) );
  AOI211_X1 U11599 ( .C1(n11005), .C2(n11004), .A(n11003), .B(n11002), .ZN(
        n11010) );
  AOI22_X1 U11600 ( .A1(n11007), .A2(n11010), .B1(n5883), .B2(n11006), .ZN(
        P2_U3535) );
  INV_X1 U11601 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U11602 ( .A1(n11011), .A2(n11010), .B1(n11009), .B2(n11008), .ZN(
        P2_U3496) );
  NOR2_X1 U11603 ( .A1(n11013), .A2(n11012), .ZN(n11018) );
  INV_X1 U11604 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11016) );
  OAI22_X1 U11605 ( .A1(n11019), .A2(n11016), .B1(n11015), .B2(n11014), .ZN(
        n11017) );
  AOI211_X1 U11606 ( .C1(n11020), .C2(n11019), .A(n11018), .B(n11017), .ZN(
        n11028) );
  OR2_X1 U11607 ( .A1(n11022), .A2(n11021), .ZN(n11026) );
  NAND2_X1 U11608 ( .A1(n11024), .A2(n11023), .ZN(n11025) );
  AND2_X1 U11609 ( .A1(n11026), .A2(n11025), .ZN(n11027) );
  NAND2_X1 U11610 ( .A1(n11028), .A2(n11027), .ZN(P1_U3275) );
  NOR2_X1 U11611 ( .A1(n11030), .A2(n11029), .ZN(n11031) );
  AOI22_X1 U11612 ( .A1(n11036), .A2(n11039), .B1(n8809), .B2(n11035), .ZN(
        P1_U3553) );
  INV_X1 U11613 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U11614 ( .A1(n11040), .A2(n11039), .B1(n11038), .B2(n11037), .ZN(
        P1_U3521) );
  XNOR2_X1 U11615 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X2 U5099 ( .A(n5957), .ZN(n5637) );
  CLKBUF_X1 U5101 ( .A(n6484), .Z(n6920) );
  CLKBUF_X2 U5113 ( .A(n8592), .Z(n5031) );
endmodule

