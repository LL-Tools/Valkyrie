

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567;

  XNOR2_X1 U2247 ( .A(n2583), .B(IR_REG_24__SCAN_IN), .ZN(n2593) );
  INV_X2 U2248 ( .A(n3324), .ZN(n3358) );
  XNOR2_X1 U2249 ( .A(n2236), .B(n2235), .ZN(n2241) );
  XNOR2_X1 U2250 ( .A(n2531), .B(IR_REG_22__SCAN_IN), .ZN(n3701) );
  OR2_X2 U2251 ( .A1(n3443), .A2(n3440), .ZN(n2198) );
  AND2_X4 U2252 ( .A1(n2237), .A2(n2241), .ZN(n2258) );
  NAND2_X2 U2253 ( .A1(n2593), .A2(n2592), .ZN(n2805) );
  AND2_X2 U2254 ( .A1(n2252), .A2(n2251), .ZN(n2647) );
  OR2_X2 U2255 ( .A1(n3139), .A2(n3246), .ZN(n3229) );
  BUF_X2 U2256 ( .A(n3338), .Z(n3353) );
  NAND2_X1 U2257 ( .A1(n4276), .A2(n4330), .ZN(n4029) );
  INV_X1 U2258 ( .A(n3614), .ZN(n3625) );
  XNOR2_X1 U2259 ( .A(n2530), .B(n2529), .ZN(n3694) );
  INV_X2 U2260 ( .A(n2254), .ZN(n3538) );
  INV_X2 U2261 ( .A(n2647), .ZN(n2522) );
  AND2_X1 U2262 ( .A1(n2226), .A2(n2222), .ZN(n2214) );
  NOR2_X1 U2263 ( .A1(n2225), .A2(n2224), .ZN(n2226) );
  NOR2_X1 U2264 ( .A1(n2231), .A2(IR_REG_25__SCAN_IN), .ZN(n2122) );
  AND3_X1 U2265 ( .A1(n2060), .A2(n2200), .A3(n2215), .ZN(n2304) );
  NOR2_X1 U2266 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2215)
         );
  INV_X1 U2267 ( .A(IR_REG_15__SCAN_IN), .ZN(n2420) );
  INV_X1 U2268 ( .A(IR_REG_14__SCAN_IN), .ZN(n2417) );
  NOR2_X1 U2269 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2200)
         );
  INV_X1 U2270 ( .A(IR_REG_13__SCAN_IN), .ZN(n2397) );
  INV_X1 U2271 ( .A(IR_REG_16__SCAN_IN), .ZN(n4225) );
  NOR2_X1 U2272 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2222)
         );
  NOR2_X2 U2273 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2060)
         );
  INV_X1 U2274 ( .A(IR_REG_11__SCAN_IN), .ZN(n2394) );
  INV_X1 U2275 ( .A(IR_REG_10__SCAN_IN), .ZN(n2393) );
  INV_X1 U2276 ( .A(IR_REG_12__SCAN_IN), .ZN(n2392) );
  INV_X1 U2277 ( .A(n2779), .ZN(n2005) );
  AND2_X4 U2278 ( .A1(n2805), .A2(n2932), .ZN(n2779) );
  NOR2_X2 U2279 ( .A1(n2083), .A2(n3117), .ZN(n3196) );
  OAI21_X2 U2280 ( .B1(n2579), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2651) );
  NOR2_X4 U2281 ( .A1(n3229), .A2(n3266), .ZN(n4047) );
  INV_X2 U2282 ( .A(n2647), .ZN(n2006) );
  OAI21_X1 U2283 ( .B1(n2134), .B2(n2133), .A(n2039), .ZN(n2132) );
  AND4_X1 U2284 ( .A1(n2317), .A2(n2122), .A3(n2214), .A4(n2232), .ZN(n2566)
         );
  NOR2_X1 U2285 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2232)
         );
  NAND2_X1 U2286 ( .A1(n3870), .A2(n2614), .ZN(n2152) );
  NAND2_X1 U2287 ( .A1(n3855), .A2(n3876), .ZN(n2153) );
  NAND2_X1 U2288 ( .A1(n2125), .A2(n2123), .ZN(n3939) );
  INV_X1 U2289 ( .A(n2124), .ZN(n2123) );
  AOI21_X1 U2290 ( .B1(n3582), .B2(n2129), .A(n3581), .ZN(n2124) );
  NAND2_X1 U2291 ( .A1(n3625), .A2(n3694), .ZN(n2725) );
  INV_X1 U2292 ( .A(IR_REG_23__SCAN_IN), .ZN(n2595) );
  OAI21_X1 U2293 ( .B1(n2581), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2594) );
  NOR2_X1 U2294 ( .A1(n2523), .A2(n2218), .ZN(n2524) );
  OR2_X1 U2295 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2218)
         );
  INV_X1 U2296 ( .A(IR_REG_2__SCAN_IN), .ZN(n2270) );
  INV_X1 U2297 ( .A(n2060), .ZN(n2255) );
  AOI21_X1 U2298 ( .B1(n2194), .B2(n2193), .A(n2035), .ZN(n2192) );
  NOR2_X1 U2299 ( .A1(n2196), .A2(n2195), .ZN(n2193) );
  INV_X1 U2300 ( .A(n3378), .ZN(n2194) );
  AND2_X1 U2301 ( .A1(n4328), .A2(n2630), .ZN(n2592) );
  NAND2_X1 U2302 ( .A1(n2109), .A2(n2108), .ZN(n2107) );
  INV_X1 U2303 ( .A(n2712), .ZN(n2108) );
  OR2_X1 U2304 ( .A1(n4353), .A2(n2168), .ZN(n2166) );
  NAND2_X1 U2305 ( .A1(n2169), .A2(REG1_REG_8__SCAN_IN), .ZN(n2168) );
  OAI21_X1 U2306 ( .B1(n4400), .B2(n3739), .A(n3738), .ZN(n3740) );
  OR2_X1 U2307 ( .A1(n4398), .A2(REG2_REG_13__SCAN_IN), .ZN(n3738) );
  OR2_X1 U2308 ( .A1(n4420), .A2(n4421), .ZN(n2158) );
  AOI22_X1 U2309 ( .A1(n4038), .A2(n2423), .B1(n3275), .B2(n3455), .ZN(n4019)
         );
  OAI21_X1 U2310 ( .B1(n3085), .B2(n2357), .A(n2356), .ZN(n3115) );
  AND2_X1 U2311 ( .A1(n2565), .A2(n3614), .ZN(n4276) );
  NAND2_X1 U2312 ( .A1(n2805), .A2(n4485), .ZN(n2740) );
  INV_X1 U2313 ( .A(IR_REG_6__SCAN_IN), .ZN(n2221) );
  AND2_X1 U2314 ( .A1(n2210), .A2(n3385), .ZN(n2207) );
  OAI21_X1 U2315 ( .B1(n2208), .B2(n2206), .A(n2046), .ZN(n2205) );
  INV_X1 U2316 ( .A(n3385), .ZN(n2206) );
  INV_X1 U2317 ( .A(IR_REG_27__SCAN_IN), .ZN(n2248) );
  INV_X1 U2318 ( .A(n2220), .ZN(n2182) );
  OAI21_X1 U2319 ( .B1(REG1_REG_7__SCAN_IN), .B2(n2882), .A(n2079), .ZN(n2883)
         );
  NAND2_X1 U2320 ( .A1(n2080), .A2(n2888), .ZN(n2079) );
  NAND2_X1 U2321 ( .A1(n2882), .A2(REG1_REG_7__SCAN_IN), .ZN(n2080) );
  INV_X1 U2322 ( .A(n4364), .ZN(n2169) );
  NOR2_X1 U2323 ( .A1(n4372), .A2(n2064), .ZN(n3754) );
  AND2_X1 U2324 ( .A1(n4498), .A2(REG1_REG_11__SCAN_IN), .ZN(n2064) );
  INV_X1 U2325 ( .A(n3587), .ZN(n2142) );
  OR2_X1 U2326 ( .A1(n2459), .A2(n3488), .ZN(n2463) );
  NOR2_X1 U2327 ( .A1(n2128), .A2(n3990), .ZN(n2127) );
  INV_X1 U2328 ( .A(n2216), .ZN(n2128) );
  INV_X1 U2329 ( .A(n2308), .ZN(n2119) );
  AND2_X1 U2330 ( .A1(n3701), .A2(n3625), .ZN(n2728) );
  NOR2_X1 U2331 ( .A1(n2433), .A2(n4046), .ZN(n2084) );
  OR2_X1 U2332 ( .A1(n4010), .A2(n4023), .ZN(n2447) );
  INV_X1 U2333 ( .A(IR_REG_18__SCAN_IN), .ZN(n2456) );
  INV_X1 U2334 ( .A(IR_REG_3__SCAN_IN), .ZN(n2280) );
  NAND2_X1 U2335 ( .A1(n3097), .A2(n3096), .ZN(n2203) );
  AND2_X1 U2336 ( .A1(n2187), .A2(n2192), .ZN(n2186) );
  NAND2_X1 U2337 ( .A1(n2010), .A2(n2199), .ZN(n2190) );
  NAND2_X1 U2338 ( .A1(n2836), .A2(n2835), .ZN(n2202) );
  NAND2_X1 U2339 ( .A1(n3301), .A2(n3300), .ZN(n3302) );
  INV_X1 U2340 ( .A(n3410), .ZN(n3301) );
  NAND2_X1 U2341 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2309) );
  NAND2_X1 U2342 ( .A1(n2828), .A2(n2664), .ZN(n2689) );
  AOI21_X1 U2343 ( .B1(n2681), .B2(REG2_REG_3__SCAN_IN), .A(n2219), .ZN(n2683)
         );
  NAND2_X1 U2344 ( .A1(n4342), .A2(n2711), .ZN(n2109) );
  OAI211_X1 U2345 ( .C1(n2854), .C2(n2068), .A(n2067), .B(n2021), .ZN(n2703)
         );
  NAND2_X1 U2346 ( .A1(n2071), .A2(REG1_REG_4__SCAN_IN), .ZN(n2068) );
  NAND2_X1 U2347 ( .A1(n2155), .A2(n2071), .ZN(n2067) );
  NAND2_X1 U2348 ( .A1(n2884), .A2(n2169), .ZN(n2167) );
  XNOR2_X1 U2349 ( .A(n3732), .B(n2077), .ZN(n2893) );
  XNOR2_X1 U2350 ( .A(n3754), .B(n2093), .ZN(n4384) );
  NAND2_X1 U2351 ( .A1(n2159), .A2(n2063), .ZN(n4393) );
  NAND2_X1 U2352 ( .A1(n3755), .A2(n2163), .ZN(n2159) );
  OR2_X1 U2353 ( .A1(n4384), .A2(n2160), .ZN(n2063) );
  NAND2_X1 U2354 ( .A1(n2163), .A2(REG1_REG_12__SCAN_IN), .ZN(n2160) );
  OR2_X1 U2355 ( .A1(n4384), .A2(n4385), .ZN(n2162) );
  NAND2_X1 U2356 ( .A1(n4377), .A2(n3735), .ZN(n3736) );
  INV_X1 U2357 ( .A(n2156), .ZN(n3760) );
  NAND2_X1 U2358 ( .A1(n3762), .A2(n3763), .ZN(n3768) );
  OR2_X1 U2359 ( .A1(n4443), .A2(n4444), .ZN(n2066) );
  NOR2_X1 U2360 ( .A1(n2099), .A2(n2098), .ZN(n2097) );
  INV_X1 U2361 ( .A(n3746), .ZN(n2098) );
  INV_X1 U2362 ( .A(n2101), .ZN(n2099) );
  OR2_X1 U2363 ( .A1(n3802), .A2(n3801), .ZN(n4062) );
  OAI22_X1 U2364 ( .A1(n2139), .A2(n2515), .B1(n3518), .B2(n3823), .ZN(n3798)
         );
  NOR2_X1 U2365 ( .A1(n3836), .A2(n3811), .ZN(n2515) );
  NAND2_X1 U2366 ( .A1(n2147), .A2(n2152), .ZN(n2144) );
  NAND2_X1 U2367 ( .A1(n2149), .A2(n2152), .ZN(n2145) );
  AND2_X1 U2368 ( .A1(n2153), .A2(n2486), .ZN(n2150) );
  NAND2_X1 U2369 ( .A1(n3972), .A2(n3974), .ZN(n2129) );
  NAND2_X1 U2370 ( .A1(n2448), .A2(n2127), .ZN(n2130) );
  AND2_X1 U2371 ( .A1(n3962), .A2(n3963), .ZN(n3990) );
  NAND2_X1 U2372 ( .A1(n4047), .A2(n2084), .ZN(n4030) );
  OAI21_X1 U2373 ( .B1(n2546), .B2(n2057), .A(n2055), .ZN(n4020) );
  INV_X1 U2374 ( .A(n2056), .ZN(n2055) );
  OAI21_X1 U2375 ( .B1(n2011), .B2(n2057), .A(n4021), .ZN(n2056) );
  INV_X1 U2376 ( .A(n3548), .ZN(n2057) );
  NAND2_X1 U2377 ( .A1(n2546), .A2(n2011), .ZN(n4039) );
  AND4_X1 U2378 ( .A1(n2416), .A2(n2415), .A3(n2414), .A4(n2413), .ZN(n3455)
         );
  AOI21_X1 U2379 ( .B1(n2135), .B2(n2366), .A(n2019), .ZN(n2134) );
  INV_X1 U2380 ( .A(n3186), .ZN(n3590) );
  NAND2_X1 U2381 ( .A1(n3191), .A2(n3117), .ZN(n2138) );
  NOR2_X1 U2382 ( .A1(n2136), .A2(n3590), .ZN(n2135) );
  INV_X1 U2383 ( .A(n2138), .ZN(n2136) );
  OAI21_X1 U2384 ( .B1(n3086), .B2(n3646), .A(n3644), .ZN(n3116) );
  OR2_X1 U2385 ( .A1(n2330), .A2(n2329), .ZN(n2346) );
  OR2_X1 U2386 ( .A1(n2343), .A2(n2342), .ZN(n2344) );
  NAND2_X1 U2387 ( .A1(n2951), .A2(n2297), .ZN(n2980) );
  NAND2_X1 U2388 ( .A1(n2564), .A2(n2563), .ZN(n4040) );
  NAND2_X1 U2389 ( .A1(n2532), .A2(n3780), .ZN(n4270) );
  NAND2_X1 U2390 ( .A1(n3813), .A2(n3364), .ZN(n3802) );
  NAND2_X1 U2391 ( .A1(n3976), .A2(n3953), .ZN(n3952) );
  NAND2_X1 U2392 ( .A1(n4276), .A2(n3694), .ZN(n4548) );
  AND2_X1 U2393 ( .A1(n2594), .A2(n2582), .ZN(n2583) );
  INV_X1 U2394 ( .A(IR_REG_19__SCAN_IN), .ZN(n2526) );
  AND2_X1 U2395 ( .A1(n2431), .A2(n2422), .ZN(n3759) );
  NOR2_X1 U2396 ( .A1(n2401), .A2(n2418), .ZN(n4398) );
  XNOR2_X1 U2397 ( .A(n2271), .B(n2270), .ZN(n2824) );
  AOI21_X1 U2398 ( .B1(n2023), .B2(n2913), .A(n2177), .ZN(n2176) );
  NAND2_X1 U2399 ( .A1(n2877), .A2(n2876), .ZN(n2902) );
  AND2_X1 U2400 ( .A1(n2738), .A2(n4476), .ZN(n3517) );
  NAND4_X1 U2401 ( .A1(n2492), .A2(n2491), .A3(n2490), .A4(n2489), .ZN(n3895)
         );
  NAND4_X1 U2402 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n3869)
         );
  INV_X1 U2403 ( .A(n3455), .ZN(n4025) );
  NAND2_X1 U2404 ( .A1(n2240), .A2(n2113), .ZN(n2112) );
  OR2_X1 U2405 ( .A1(n2254), .A2(n2253), .ZN(n2111) );
  NAND2_X1 U2406 ( .A1(n2265), .A2(REG3_REG_1__SCAN_IN), .ZN(n2114) );
  XNOR2_X1 U2407 ( .A(n2668), .B(REG1_REG_1__SCAN_IN), .ZN(n3722) );
  XNOR2_X1 U2408 ( .A(n2683), .B(n2682), .ZN(n2853) );
  XNOR2_X1 U2409 ( .A(n2703), .B(n4505), .ZN(n4349) );
  NAND2_X1 U2410 ( .A1(n4349), .A2(REG1_REG_6__SCAN_IN), .ZN(n4348) );
  NOR2_X1 U2411 ( .A1(n2076), .A2(n4331), .ZN(n2075) );
  INV_X1 U2412 ( .A(n2164), .ZN(n2076) );
  AND3_X1 U2413 ( .A1(n3750), .A2(n2074), .A3(REG1_REG_10__SCAN_IN), .ZN(n3751) );
  XNOR2_X1 U2414 ( .A(n3736), .B(n2093), .ZN(n4390) );
  NAND2_X1 U2415 ( .A1(n4390), .A2(REG2_REG_12__SCAN_IN), .ZN(n4389) );
  AOI21_X1 U2416 ( .B1(n4450), .B2(n4449), .A(n2049), .ZN(n2171) );
  INV_X1 U2417 ( .A(n2066), .ZN(n4442) );
  NAND2_X1 U2418 ( .A1(n2174), .A2(n4435), .ZN(n2173) );
  NAND2_X1 U2419 ( .A1(n4443), .A2(n4444), .ZN(n2174) );
  NAND2_X1 U2420 ( .A1(n3773), .A2(n2102), .ZN(n4446) );
  INV_X1 U2421 ( .A(n4476), .ZN(n4453) );
  NOR2_X1 U2422 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2062)
         );
  AND2_X1 U2423 ( .A1(n3220), .A2(n2543), .ZN(n3617) );
  INV_X1 U2424 ( .A(n2385), .ZN(n2133) );
  NOR2_X1 U2425 ( .A1(n3280), .A2(n3279), .ZN(n3451) );
  AOI21_X1 U2426 ( .B1(n2702), .B2(REG2_REG_5__SCAN_IN), .A(n2708), .ZN(n2710)
         );
  INV_X1 U2427 ( .A(n4394), .ZN(n2163) );
  NOR2_X1 U2428 ( .A1(n4393), .A2(n2044), .ZN(n3756) );
  NAND2_X1 U2429 ( .A1(n2158), .A2(n2157), .ZN(n2156) );
  NAND2_X1 U2430 ( .A1(n3759), .A2(REG1_REG_15__SCAN_IN), .ZN(n2157) );
  NAND2_X1 U2431 ( .A1(n4449), .A2(REG2_REG_18__SCAN_IN), .ZN(n2101) );
  OR2_X1 U2432 ( .A1(n3961), .A2(n3885), .ZN(n3941) );
  NAND2_X1 U2433 ( .A1(n2061), .A2(n3883), .ZN(n3961) );
  INV_X1 U2434 ( .A(n4008), .ZN(n2061) );
  OR2_X1 U2435 ( .A1(n2273), .A2(n2774), .ZN(n3627) );
  OR2_X1 U2436 ( .A1(n3194), .A2(n3140), .ZN(n3139) );
  NAND2_X1 U2437 ( .A1(n3058), .A2(n2009), .ZN(n2083) );
  NOR2_X1 U2438 ( .A1(n3040), .A2(n2916), .ZN(n2082) );
  INV_X1 U2439 ( .A(n2231), .ZN(n2121) );
  NAND2_X1 U2440 ( .A1(n2317), .A2(n2214), .ZN(n2435) );
  OR2_X1 U2441 ( .A1(n2396), .A2(n2395), .ZN(n2400) );
  NOR2_X1 U2442 ( .A1(n2901), .A2(n2178), .ZN(n2177) );
  NOR2_X1 U2443 ( .A1(n3513), .A2(n2197), .ZN(n2196) );
  INV_X1 U2444 ( .A(n3441), .ZN(n2197) );
  NAND2_X1 U2445 ( .A1(n3264), .A2(n2209), .ZN(n2208) );
  INV_X1 U2446 ( .A(n3262), .ZN(n2209) );
  NAND2_X1 U2447 ( .A1(n3262), .A2(n3265), .ZN(n2210) );
  OR2_X1 U2448 ( .A1(n2449), .A2(n3413), .ZN(n2459) );
  INV_X1 U2449 ( .A(n3357), .ZN(n3348) );
  AND2_X1 U2450 ( .A1(n2487), .A2(REG3_REG_24__SCAN_IN), .ZN(n2495) );
  NOR2_X1 U2451 ( .A1(n2386), .A2(n3243), .ZN(n2402) );
  INV_X1 U2452 ( .A(n2179), .ZN(n3493) );
  AOI21_X1 U2453 ( .B1(n2007), .B2(n3483), .A(n3428), .ZN(n2180) );
  NAND2_X1 U2454 ( .A1(n2007), .A2(n2182), .ZN(n2181) );
  NAND2_X1 U2455 ( .A1(n2781), .A2(n2780), .ZN(n2782) );
  NAND2_X1 U2456 ( .A1(n2442), .A2(REG3_REG_18__SCAN_IN), .ZN(n2449) );
  AND2_X1 U2457 ( .A1(n2495), .A2(REG3_REG_25__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U2458 ( .A1(n2237), .A2(n2635), .ZN(n2254) );
  AND2_X1 U2459 ( .A1(n2241), .A2(REG2_REG_1__SCAN_IN), .ZN(n2113) );
  NAND2_X1 U2460 ( .A1(n2258), .A2(REG0_REG_1__SCAN_IN), .ZN(n2110) );
  NAND2_X1 U2461 ( .A1(n2823), .A2(n2822), .ZN(n2821) );
  XNOR2_X1 U2462 ( .A(n2680), .B(n2671), .ZN(n2681) );
  INV_X1 U2463 ( .A(n2694), .ZN(n2071) );
  INV_X1 U2464 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2091) );
  INV_X1 U2465 ( .A(n2279), .ZN(n2201) );
  XNOR2_X1 U2466 ( .A(n2883), .B(n4362), .ZN(n4353) );
  NAND2_X1 U2467 ( .A1(n2107), .A2(n2032), .ZN(n2889) );
  NOR2_X1 U2468 ( .A1(n4353), .A2(n4354), .ZN(n4352) );
  NOR2_X1 U2469 ( .A1(n2165), .A2(n2040), .ZN(n2164) );
  INV_X1 U2470 ( .A(n2167), .ZN(n2165) );
  NAND2_X1 U2471 ( .A1(n4367), .A2(n2892), .ZN(n3732) );
  INV_X1 U2472 ( .A(n4493), .ZN(n3757) );
  XNOR2_X1 U2473 ( .A(n2156), .B(n4490), .ZN(n4433) );
  NAND2_X1 U2474 ( .A1(n3768), .A2(n2048), .ZN(n4443) );
  NOR2_X1 U2475 ( .A1(n4447), .A2(n2103), .ZN(n2100) );
  NAND2_X1 U2476 ( .A1(n2095), .A2(n2101), .ZN(n2094) );
  INV_X1 U2477 ( .A(n2100), .ZN(n2095) );
  NOR2_X1 U2478 ( .A1(n4062), .A2(n4065), .ZN(n4061) );
  NOR2_X1 U2479 ( .A1(n2509), .A2(n4179), .ZN(n2516) );
  OR2_X1 U2480 ( .A1(n2145), .A2(n2016), .ZN(n2143) );
  INV_X1 U2481 ( .A(n2141), .ZN(n2140) );
  OAI21_X1 U2482 ( .B1(n2144), .B2(n2016), .A(n2142), .ZN(n2141) );
  INV_X1 U2483 ( .A(n3895), .ZN(n3855) );
  AOI21_X1 U2484 ( .B1(n3924), .B2(n3923), .A(n3889), .ZN(n3909) );
  NAND2_X1 U2485 ( .A1(n3947), .A2(n3932), .ZN(n2469) );
  NOR2_X1 U2486 ( .A1(n3947), .A2(n3932), .ZN(n2470) );
  OR2_X1 U2487 ( .A1(n3952), .A2(n2613), .ZN(n3931) );
  AND2_X1 U2488 ( .A1(n2440), .A2(REG3_REG_17__SCAN_IN), .ZN(n2442) );
  NAND2_X1 U2489 ( .A1(n4020), .A2(n3551), .ZN(n4008) );
  INV_X1 U2490 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U2491 ( .A1(n4019), .A2(n4018), .ZN(n4017) );
  INV_X1 U2492 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3528) );
  OR2_X1 U2493 ( .A1(n3266), .A2(n3707), .ZN(n2410) );
  INV_X1 U2494 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2375) );
  NAND2_X1 U2495 ( .A1(n3116), .A2(n3661), .ZN(n2541) );
  AND4_X1 U2496 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n3244)
         );
  NAND2_X1 U2497 ( .A1(n2540), .A2(n3652), .ZN(n3086) );
  OAI21_X1 U2498 ( .B1(n2980), .B2(n2020), .A(n2115), .ZN(n2320) );
  INV_X1 U2499 ( .A(n2116), .ZN(n2115) );
  INV_X1 U2500 ( .A(n3651), .ZN(n2058) );
  OR2_X1 U2501 ( .A1(n2957), .A2(n2850), .ZN(n2977) );
  NAND2_X1 U2502 ( .A1(n3627), .A2(n3630), .ZN(n3598) );
  OR2_X1 U2503 ( .A1(n2804), .A2(n2740), .ZN(n2928) );
  INV_X1 U2504 ( .A(n3607), .ZN(n4065) );
  AND2_X1 U2505 ( .A1(n2087), .A2(n2086), .ZN(n4070) );
  INV_X1 U2506 ( .A(n3793), .ZN(n2086) );
  NAND2_X1 U2507 ( .A1(n2088), .A2(n4040), .ZN(n2087) );
  OR2_X1 U2508 ( .A1(n3804), .A2(n3803), .ZN(n2089) );
  NAND2_X1 U2509 ( .A1(n2085), .A2(n3841), .ZN(n3840) );
  NAND2_X1 U2510 ( .A1(n3899), .A2(n3876), .ZN(n3875) );
  NAND2_X1 U2511 ( .A1(n2522), .A2(DATAI_23_), .ZN(n3901) );
  NOR2_X1 U2512 ( .A1(n3931), .A2(n3917), .ZN(n3916) );
  AND2_X1 U2513 ( .A1(n3916), .A2(n3901), .ZN(n3899) );
  AND2_X1 U2514 ( .A1(n4003), .A2(n2612), .ZN(n3976) );
  NAND2_X1 U2515 ( .A1(n2448), .A2(n2216), .ZN(n3989) );
  NAND2_X1 U2516 ( .A1(n4047), .A2(n3275), .ZN(n4032) );
  NAND2_X1 U2517 ( .A1(n3196), .A2(n3195), .ZN(n3194) );
  INV_X1 U2518 ( .A(n3032), .ZN(n3040) );
  NAND2_X1 U2519 ( .A1(n3058), .A2(n2082), .ZN(n3090) );
  NAND2_X1 U2520 ( .A1(n3058), .A2(n2991), .ZN(n3039) );
  NOR2_X1 U2521 ( .A1(n2977), .A2(n2976), .ZN(n3056) );
  AND2_X1 U2522 ( .A1(n3056), .A2(n3055), .ZN(n3058) );
  NAND2_X1 U2523 ( .A1(n2980), .A2(n2308), .ZN(n2120) );
  NOR2_X1 U2524 ( .A1(n3017), .A2(n2793), .ZN(n2943) );
  INV_X1 U2525 ( .A(n4548), .ZN(n4545) );
  NAND2_X1 U2526 ( .A1(n2525), .A2(n2581), .ZN(n3614) );
  NAND2_X1 U2527 ( .A1(n2213), .A2(n2211), .ZN(n2525) );
  NAND2_X1 U2528 ( .A1(n2212), .A2(IR_REG_31__SCAN_IN), .ZN(n2211) );
  INV_X1 U2529 ( .A(IR_REG_20__SCAN_IN), .ZN(n2529) );
  OR2_X1 U2530 ( .A1(n2353), .A2(IR_REG_9__SCAN_IN), .ZN(n2396) );
  INV_X1 U2531 ( .A(IR_REG_7__SCAN_IN), .ZN(n2327) );
  AND2_X1 U2532 ( .A1(n2292), .A2(n2282), .ZN(n2688) );
  OAI211_X1 U2533 ( .C1(IR_REG_31__SCAN_IN), .C2(IR_REG_1__SCAN_IN), .A(n2154), 
        .B(n2255), .ZN(n2668) );
  NAND2_X1 U2534 ( .A1(n2022), .A2(IR_REG_1__SCAN_IN), .ZN(n2154) );
  NAND2_X1 U2535 ( .A1(n2191), .A2(n3512), .ZN(n3379) );
  NAND2_X1 U2536 ( .A1(n2198), .A2(n2196), .ZN(n2191) );
  NAND2_X1 U2537 ( .A1(n2204), .A2(n2208), .ZN(n3387) );
  NAND2_X1 U2538 ( .A1(n3263), .A2(n2210), .ZN(n2204) );
  INV_X1 U2539 ( .A(n3106), .ZN(n3107) );
  NAND2_X1 U2540 ( .A1(n2203), .A2(n3101), .ZN(n3105) );
  INV_X1 U2541 ( .A(n2936), .ZN(n2942) );
  INV_X1 U2542 ( .A(n2192), .ZN(n2185) );
  NAND2_X1 U2543 ( .A1(n2189), .A2(n3362), .ZN(n2188) );
  INV_X1 U2544 ( .A(n2190), .ZN(n2189) );
  INV_X1 U2545 ( .A(n3140), .ZN(n3172) );
  NAND2_X1 U2546 ( .A1(n2006), .A2(DATAI_25_), .ZN(n3857) );
  INV_X1 U2547 ( .A(n2875), .ZN(n2976) );
  CLKBUF_X1 U2548 ( .A(n3460), .Z(n3465) );
  NAND2_X1 U2549 ( .A1(n2006), .A2(DATAI_24_), .ZN(n3876) );
  INV_X1 U2550 ( .A(n2845), .ZN(n2846) );
  NAND2_X1 U2551 ( .A1(n2202), .A2(n2840), .ZN(n2844) );
  INV_X1 U2552 ( .A(n2958), .ZN(n2850) );
  AND4_X1 U2553 ( .A1(n2335), .A2(n2334), .A3(n2333), .A4(n2332), .ZN(n3081)
         );
  INV_X1 U2554 ( .A(n4277), .ZN(n3601) );
  NAND2_X1 U2555 ( .A1(n2522), .A2(DATAI_20_), .ZN(n3953) );
  CLKBUF_X1 U2556 ( .A(n3405), .Z(n3506) );
  AND4_X1 U2557 ( .A1(n2301), .A2(n2300), .A3(n2299), .A4(n2298), .ZN(n3048)
         );
  NAND2_X1 U2558 ( .A1(n2902), .A2(n2901), .ZN(n2915) );
  NAND2_X1 U2559 ( .A1(n2198), .A2(n3441), .ZN(n3515) );
  INV_X1 U2560 ( .A(n3517), .ZN(n3532) );
  OR2_X1 U2561 ( .A1(n2811), .A2(n2810), .ZN(n3533) );
  NAND4_X1 U2562 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(n3820)
         );
  NAND4_X1 U2563 ( .A1(n2514), .A2(n2513), .A3(n2512), .A4(n2511), .ZN(n3836)
         );
  NAND4_X1 U2564 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n3852)
         );
  NAND4_X1 U2565 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n3870)
         );
  OAI211_X1 U2566 ( .C1(n3487), .C2(n2468), .A(n2462), .B(n2461), .ZN(n3969)
         );
  INV_X1 U2567 ( .A(n3081), .ZN(n3712) );
  NAND4_X1 U2568 ( .A1(n2291), .A2(n2290), .A3(n2289), .A4(n2288), .ZN(n3717)
         );
  NAND3_X1 U2569 ( .A1(n2263), .A2(n2262), .A3(n2261), .ZN(n3720) );
  NAND2_X1 U2570 ( .A1(n3538), .A2(REG1_REG_0__SCAN_IN), .ZN(n2261) );
  INV_X1 U2571 ( .A(U4043), .ZN(n3719) );
  AND2_X1 U2572 ( .A1(n2650), .A2(n2649), .ZN(n2666) );
  NAND2_X1 U2573 ( .A1(n2663), .A2(n2662), .ZN(n2828) );
  XNOR2_X1 U2574 ( .A(n2689), .B(n2671), .ZN(n2687) );
  INV_X1 U2575 ( .A(n2072), .ZN(n2695) );
  INV_X1 U2576 ( .A(n2090), .ZN(n2686) );
  OAI21_X1 U2577 ( .B1(n2853), .B2(n2091), .A(n2092), .ZN(n2090) );
  INV_X1 U2578 ( .A(n2107), .ZN(n2887) );
  INV_X1 U2579 ( .A(n2109), .ZN(n2713) );
  NAND2_X1 U2580 ( .A1(n4348), .A2(n2704), .ZN(n2882) );
  XNOR2_X1 U2581 ( .A(n4362), .B(n2889), .ZN(n4359) );
  NAND2_X1 U2582 ( .A1(n2166), .A2(n2167), .ZN(n4363) );
  NOR2_X1 U2583 ( .A1(n3751), .A2(n3752), .ZN(n4374) );
  INV_X1 U2584 ( .A(n2162), .ZN(n4383) );
  INV_X1 U2585 ( .A(n3755), .ZN(n2161) );
  NAND2_X1 U2586 ( .A1(n4389), .A2(n3737), .ZN(n4400) );
  XNOR2_X1 U2587 ( .A(n3740), .B(n3757), .ZN(n4408) );
  NOR2_X1 U2588 ( .A1(n4408), .A2(n4409), .ZN(n4407) );
  OAI21_X1 U2589 ( .B1(n4408), .B2(n2105), .A(n2104), .ZN(n4415) );
  NAND2_X1 U2590 ( .A1(n2106), .A2(REG2_REG_14__SCAN_IN), .ZN(n2105) );
  NAND2_X1 U2591 ( .A1(n3741), .A2(n2106), .ZN(n2104) );
  INV_X1 U2592 ( .A(n4416), .ZN(n2106) );
  INV_X1 U2593 ( .A(n2158), .ZN(n4419) );
  AND2_X1 U2594 ( .A1(n2066), .A2(n2065), .ZN(n3771) );
  NAND2_X1 U2595 ( .A1(n4449), .A2(REG1_REG_18__SCAN_IN), .ZN(n2065) );
  NAND2_X1 U2596 ( .A1(n2096), .A2(n2094), .ZN(n3777) );
  OAI21_X1 U2597 ( .B1(n3882), .B2(n2145), .A(n2144), .ZN(n3829) );
  INV_X1 U2598 ( .A(n2146), .ZN(n3847) );
  AOI21_X1 U2599 ( .B1(n3882), .B2(n2150), .A(n2148), .ZN(n2146) );
  NAND2_X1 U2600 ( .A1(n3882), .A2(n2486), .ZN(n2151) );
  NAND2_X1 U2601 ( .A1(n3897), .A2(n2033), .ZN(n4087) );
  NAND2_X1 U2602 ( .A1(n3926), .A2(n4024), .ZN(n2054) );
  AND2_X1 U2603 ( .A1(n2130), .A2(n2129), .ZN(n3959) );
  NAND2_X1 U2604 ( .A1(n4039), .A2(n3548), .ZN(n4022) );
  NAND2_X1 U2605 ( .A1(n2131), .A2(n2134), .ZN(n3138) );
  NAND2_X1 U2606 ( .A1(n3115), .A2(n2135), .ZN(n2131) );
  NAND2_X1 U2607 ( .A1(n2137), .A2(n2138), .ZN(n3188) );
  OR2_X1 U2608 ( .A1(n3115), .A2(n2366), .ZN(n2137) );
  AND2_X1 U2609 ( .A1(n4470), .A2(n2982), .ZN(n3999) );
  OR2_X1 U2610 ( .A1(n2740), .A2(n2737), .ZN(n4476) );
  NOR2_X1 U2611 ( .A1(n4463), .A2(n2981), .ZN(n4466) );
  NOR2_X1 U2612 ( .A1(n4087), .A2(n2053), .ZN(n4300) );
  NOR2_X1 U2613 ( .A1(n2008), .A2(n4540), .ZN(n2053) );
  AND2_X2 U2614 ( .A1(n2610), .A2(n2618), .ZN(n4555) );
  AND2_X1 U2615 ( .A1(n2588), .A2(n2589), .ZN(n2645) );
  NAND2_X1 U2616 ( .A1(n2641), .A2(IR_REG_31__SCAN_IN), .ZN(n2233) );
  INV_X1 U2617 ( .A(n2241), .ZN(n2635) );
  XNOR2_X1 U2618 ( .A(n2586), .B(IR_REG_26__SCAN_IN), .ZN(n2630) );
  INV_X1 U2619 ( .A(n2579), .ZN(n2585) );
  CLKBUF_X1 U2620 ( .A(n2593), .Z(n4329) );
  AND2_X1 U2621 ( .A1(n2806), .A2(STATE_REG_SCAN_IN), .ZN(n4485) );
  XNOR2_X1 U2622 ( .A(n2527), .B(n2526), .ZN(n3780) );
  XNOR2_X1 U2623 ( .A(n2382), .B(IR_REG_11__SCAN_IN), .ZN(n4498) );
  INV_X1 U2624 ( .A(IR_REG_4__SCAN_IN), .ZN(n2293) );
  NAND2_X1 U2625 ( .A1(n3750), .A2(n2074), .ZN(n2885) );
  OR2_X1 U2626 ( .A1(n2173), .A2(n4442), .ZN(n2172) );
  OAI21_X1 U2627 ( .B1(n4451), .B2(n4452), .A(n2171), .ZN(n2170) );
  OAI21_X1 U2628 ( .B1(n4300), .B2(n4564), .A(n2050), .ZN(U3541) );
  AND2_X1 U2629 ( .A1(n2052), .A2(n2051), .ZN(n2050) );
  OR2_X1 U2630 ( .A1(n4567), .A2(n4191), .ZN(n2051) );
  OR2_X1 U2631 ( .A1(n4303), .A2(n4268), .ZN(n2052) );
  OR2_X1 U2632 ( .A1(n3373), .A2(n4325), .ZN(n2616) );
  NOR2_X1 U2633 ( .A1(n3308), .A2(n2220), .ZN(n3429) );
  NOR2_X1 U2634 ( .A1(n3430), .A2(n3427), .ZN(n2007) );
  XNOR2_X1 U2635 ( .A(n3892), .B(n3882), .ZN(n2008) );
  NAND2_X1 U2636 ( .A1(n2201), .A2(n2215), .ZN(n2302) );
  AND2_X1 U2637 ( .A1(n2082), .A2(n2081), .ZN(n2009) );
  INV_X1 U2638 ( .A(IR_REG_28__SCAN_IN), .ZN(n2567) );
  NOR2_X1 U2639 ( .A1(n3378), .A2(n2195), .ZN(n2010) );
  AND2_X1 U2640 ( .A1(n2043), .A2(n3546), .ZN(n2011) );
  INV_X1 U2641 ( .A(n2914), .ZN(n2178) );
  NAND2_X1 U2642 ( .A1(n2317), .A2(n2222), .ZN(n2353) );
  AND2_X1 U2643 ( .A1(n3714), .A2(n2909), .ZN(n2012) );
  NAND2_X1 U2644 ( .A1(n3869), .A2(n2485), .ZN(n2013) );
  XNOR2_X1 U2645 ( .A(n2233), .B(IR_REG_30__SCAN_IN), .ZN(n2240) );
  NAND4_X1 U2646 ( .A1(n2269), .A2(n2268), .A3(n2267), .A4(n2266), .ZN(n2273)
         );
  OR2_X1 U2647 ( .A1(n2913), .A2(n2914), .ZN(n2014) );
  NAND4_X1 U2648 ( .A1(n2111), .A2(n2114), .A3(n2110), .A4(n2112), .ZN(n4273)
         );
  INV_X1 U2649 ( .A(n4273), .ZN(n2257) );
  AND3_X1 U2650 ( .A1(n2317), .A2(n2214), .A3(n2121), .ZN(n2015) );
  AND2_X1 U2651 ( .A1(n3852), .A2(n2615), .ZN(n2016) );
  NOR2_X1 U2652 ( .A1(n3429), .A2(n3483), .ZN(n2017) );
  NOR2_X1 U2653 ( .A1(n4448), .A2(n2170), .ZN(n2018) );
  AND2_X1 U2654 ( .A1(n3173), .A2(n3195), .ZN(n2019) );
  OR2_X1 U2655 ( .A1(n2012), .A2(n2217), .ZN(n2020) );
  NAND2_X1 U2656 ( .A1(n2702), .A2(REG1_REG_5__SCAN_IN), .ZN(n2021) );
  INV_X1 U2657 ( .A(IR_REG_29__SCAN_IN), .ZN(n2235) );
  AND2_X1 U2658 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2022)
         );
  NAND2_X1 U2659 ( .A1(n2901), .A2(n2178), .ZN(n2023) );
  OAI21_X1 U2660 ( .B1(n2148), .B2(n2150), .A(n2502), .ZN(n2147) );
  INV_X1 U2661 ( .A(n2149), .ZN(n2148) );
  NAND2_X1 U2662 ( .A1(n2024), .A2(n2153), .ZN(n2149) );
  NAND2_X1 U2663 ( .A1(n2494), .A2(n2013), .ZN(n2024) );
  AND2_X1 U2664 ( .A1(n2135), .A2(n2385), .ZN(n2025) );
  AND2_X1 U2665 ( .A1(n2151), .A2(n2013), .ZN(n2026) );
  AND2_X1 U2666 ( .A1(n2014), .A2(n2876), .ZN(n2027) );
  INV_X1 U2667 ( .A(n2139), .ZN(n3809) );
  OAI21_X1 U2668 ( .B1(n3882), .B2(n2143), .A(n2140), .ZN(n2139) );
  AND2_X1 U2669 ( .A1(n3773), .A2(n2100), .ZN(n2028) );
  AND2_X1 U2670 ( .A1(n2846), .A2(n2840), .ZN(n2029) );
  AND2_X1 U2671 ( .A1(n3107), .A2(n3101), .ZN(n2030) );
  OR2_X1 U2672 ( .A1(n2685), .A2(n2091), .ZN(n2031) );
  INV_X1 U2673 ( .A(IR_REG_21__SCAN_IN), .ZN(n2212) );
  INV_X1 U2674 ( .A(n3440), .ZN(n2199) );
  OR2_X1 U2675 ( .A1(n2888), .A2(n2990), .ZN(n2032) );
  INV_X1 U2676 ( .A(n3091), .ZN(n2081) );
  INV_X1 U2677 ( .A(n3512), .ZN(n2195) );
  INV_X1 U2678 ( .A(n4046), .ZN(n3275) );
  INV_X1 U2679 ( .A(n3467), .ZN(n4010) );
  AND2_X1 U2680 ( .A1(n3896), .A2(n2054), .ZN(n2033) );
  NOR2_X1 U2681 ( .A1(n4407), .A2(n3741), .ZN(n2034) );
  AND2_X1 U2682 ( .A1(n3355), .A2(n3354), .ZN(n2035) );
  INV_X1 U2683 ( .A(n2085), .ZN(n3856) );
  NOR2_X1 U2684 ( .A1(n3875), .A2(n2614), .ZN(n2085) );
  INV_X1 U2685 ( .A(n4041), .ZN(n4014) );
  AND2_X1 U2686 ( .A1(n2137), .A2(n2135), .ZN(n2036) );
  AND2_X1 U2687 ( .A1(n2546), .A2(n3546), .ZN(n2037) );
  AND2_X1 U2688 ( .A1(n2162), .A2(n2161), .ZN(n2038) );
  NAND2_X1 U2689 ( .A1(n3244), .A2(n3172), .ZN(n2039) );
  AND2_X1 U2690 ( .A1(n2886), .A2(REG1_REG_9__SCAN_IN), .ZN(n2040) );
  INV_X1 U2691 ( .A(n3581), .ZN(n2126) );
  AND2_X1 U2692 ( .A1(n2084), .A2(n3467), .ZN(n2041) );
  AND2_X1 U2693 ( .A1(n2127), .A2(n2126), .ZN(n2042) );
  NAND2_X2 U2694 ( .A1(n2931), .A2(n4476), .ZN(n4470) );
  AND2_X1 U2695 ( .A1(n3549), .A2(n3548), .ZN(n2043) );
  INV_X1 U2696 ( .A(n3753), .ZN(n2093) );
  INV_X1 U2697 ( .A(n3932), .ZN(n2613) );
  NAND2_X1 U2698 ( .A1(n2295), .A2(DATAI_21_), .ZN(n3932) );
  NAND2_X1 U2699 ( .A1(n2120), .A2(n2118), .ZN(n3047) );
  NAND2_X1 U2700 ( .A1(n2175), .A2(n2176), .ZN(n2999) );
  AND2_X1 U2701 ( .A1(n4398), .A2(REG1_REG_13__SCAN_IN), .ZN(n2044) );
  NOR2_X1 U2702 ( .A1(n4352), .A2(n2884), .ZN(n2045) );
  AND2_X2 U2703 ( .A1(n2618), .A2(n2930), .ZN(n4567) );
  AND2_X1 U2704 ( .A1(n2666), .A2(n2665), .ZN(n4435) );
  INV_X1 U2705 ( .A(n4024), .ZN(n4044) );
  INV_X1 U2706 ( .A(n2693), .ZN(n2155) );
  NAND2_X1 U2707 ( .A1(n4270), .A2(n4549), .ZN(n4533) );
  INV_X1 U2708 ( .A(n4533), .ZN(n4540) );
  NAND2_X1 U2709 ( .A1(n3274), .A2(n3273), .ZN(n2046) );
  AND3_X1 U2710 ( .A1(n2070), .A2(n2071), .A3(n2069), .ZN(n2047) );
  OR2_X1 U2711 ( .A1(n3774), .A2(REG1_REG_17__SCAN_IN), .ZN(n2048) );
  INV_X1 U2712 ( .A(n2103), .ZN(n2102) );
  NOR2_X1 U2713 ( .A1(n3774), .A2(REG2_REG_17__SCAN_IN), .ZN(n2103) );
  AND2_X1 U2714 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n2049) );
  INV_X1 U2715 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2073) );
  OAI21_X1 U2716 ( .B1(n2986), .B2(n2539), .A(n3648), .ZN(n3031) );
  OAI21_X2 U2717 ( .B1(n2059), .B2(n2058), .A(n3639), .ZN(n2986) );
  INV_X1 U2718 ( .A(n3049), .ZN(n2059) );
  NAND2_X1 U2719 ( .A1(n2060), .A2(n2270), .ZN(n2279) );
  NAND2_X1 U2720 ( .A1(IR_REG_31__SCAN_IN), .A2(n2255), .ZN(n2271) );
  OAI21_X2 U2721 ( .B1(n3941), .B2(n3888), .A(n3887), .ZN(n3924) );
  NAND2_X1 U2722 ( .A1(n2566), .A2(n2567), .ZN(n2234) );
  NAND2_X1 U2723 ( .A1(n2566), .A2(n2062), .ZN(n2641) );
  OAI21_X1 U2724 ( .B1(n2952), .B2(n2537), .A(n3636), .ZN(n2971) );
  NAND2_X1 U2725 ( .A1(n2933), .A2(n3632), .ZN(n2952) );
  NAND2_X1 U2726 ( .A1(n2934), .A2(n2935), .ZN(n2933) );
  NAND2_X1 U2727 ( .A1(n2687), .A2(REG1_REG_3__SCAN_IN), .ZN(n2691) );
  NOR2_X1 U2728 ( .A1(n4404), .A2(n3758), .ZN(n4420) );
  OAI21_X1 U2729 ( .B1(n2854), .B2(n2073), .A(n2693), .ZN(n2072) );
  NAND2_X1 U2730 ( .A1(n2693), .A2(n2073), .ZN(n2069) );
  NAND2_X1 U2731 ( .A1(n2854), .A2(n2693), .ZN(n2070) );
  NAND2_X1 U2732 ( .A1(n2166), .A2(n2164), .ZN(n2078) );
  NAND2_X1 U2733 ( .A1(n2075), .A2(n2166), .ZN(n2074) );
  NAND2_X1 U2734 ( .A1(n2078), .A2(n4331), .ZN(n3750) );
  INV_X1 U2735 ( .A(n4331), .ZN(n2077) );
  INV_X1 U2736 ( .A(n2083), .ZN(n3126) );
  AND2_X2 U2737 ( .A1(n4047), .A2(n2041), .ZN(n4003) );
  NOR2_X2 U2738 ( .A1(n3840), .A2(n3811), .ZN(n3813) );
  OAI211_X1 U2739 ( .C1(n4069), .C2(n4548), .A(n4070), .B(n4071), .ZN(n4285)
         );
  XNOR2_X1 U2740 ( .A(n3788), .B(n3606), .ZN(n2088) );
  NAND2_X1 U2741 ( .A1(n4062), .A2(n2089), .ZN(n4069) );
  NAND3_X1 U2742 ( .A1(n2214), .A2(n2317), .A3(n2122), .ZN(n2579) );
  AND2_X2 U2743 ( .A1(n2304), .A2(n2221), .ZN(n2317) );
  OAI22_X1 U2744 ( .A1(n2685), .A2(n2092), .B1(n2853), .B2(n2031), .ZN(n2708)
         );
  NAND2_X1 U2745 ( .A1(n2684), .A2(n2856), .ZN(n2092) );
  NAND2_X1 U2746 ( .A1(n3745), .A2(n2097), .ZN(n2096) );
  NAND2_X1 U2747 ( .A1(n3745), .A2(n3746), .ZN(n3773) );
  AOI21_X1 U2748 ( .B1(n3759), .B2(REG2_REG_15__SCAN_IN), .A(n4415), .ZN(n3743) );
  AOI21_X1 U2749 ( .B1(n3782), .B2(n4437), .A(n3781), .ZN(n3783) );
  NAND2_X1 U2750 ( .A1(n2172), .A2(n2018), .ZN(U3258) );
  NAND2_X1 U2751 ( .A1(n2250), .A2(n2249), .ZN(n2252) );
  AND2_X2 U2752 ( .A1(n2240), .A2(n2241), .ZN(n2497) );
  OAI21_X1 U2753 ( .B1(n2117), .B2(n2012), .A(n2319), .ZN(n2116) );
  NAND2_X1 U2754 ( .A1(n2118), .A2(n2119), .ZN(n2117) );
  INV_X1 U2755 ( .A(n2217), .ZN(n2118) );
  NAND2_X1 U2756 ( .A1(n2448), .A2(n2042), .ZN(n2125) );
  INV_X1 U2757 ( .A(n2130), .ZN(n3988) );
  AOI21_X1 U2758 ( .B1(n3115), .B2(n2025), .A(n2132), .ZN(n3219) );
  NAND2_X1 U2759 ( .A1(n2877), .A2(n2027), .ZN(n2175) );
  OAI21_X1 U2760 ( .B1(n3308), .B2(n2181), .A(n2180), .ZN(n2179) );
  OAI211_X1 U2761 ( .C1(n3443), .C2(n2188), .A(n2184), .B(n2183), .ZN(n3369)
         );
  NAND2_X1 U2762 ( .A1(n3443), .A2(n2186), .ZN(n2183) );
  AOI22_X1 U2763 ( .A1(n2186), .A2(n2190), .B1(n2185), .B2(n3362), .ZN(n2184)
         );
  INV_X1 U2764 ( .A(n3362), .ZN(n2187) );
  NAND2_X1 U2765 ( .A1(n2202), .A2(n2029), .ZN(n2873) );
  NAND2_X1 U2766 ( .A1(n2203), .A2(n2030), .ZN(n3148) );
  AOI21_X1 U2767 ( .B1(n3263), .B2(n2207), .A(n2205), .ZN(n3280) );
  OAI21_X1 U2768 ( .B1(n2524), .B2(n2640), .A(IR_REG_21__SCAN_IN), .ZN(n2213)
         );
  CLKBUF_X1 U2769 ( .A(n3450), .Z(n3523) );
  CLKBUF_X1 U2770 ( .A(n3451), .Z(n3525) );
  OR2_X1 U2771 ( .A1(n3352), .A2(n2727), .ZN(n2734) );
  INV_X1 U2772 ( .A(n4028), .ZN(n2433) );
  OR2_X1 U2773 ( .A1(n3985), .A2(n3467), .ZN(n2216) );
  AND2_X1 U2774 ( .A1(n3715), .A2(n2976), .ZN(n2217) );
  INV_X1 U2775 ( .A(n2707), .ZN(n2702) );
  NAND2_X1 U2776 ( .A1(n2006), .A2(DATAI_22_), .ZN(n3910) );
  INV_X1 U2777 ( .A(n3910), .ZN(n3917) );
  INV_X1 U2778 ( .A(n4505), .ZN(n2709) );
  INV_X1 U2779 ( .A(IR_REG_31__SCAN_IN), .ZN(n2640) );
  AND2_X1 U2780 ( .A1(n2680), .A2(n2688), .ZN(n2219) );
  AND2_X1 U2781 ( .A1(n2355), .A2(n2396), .ZN(n2886) );
  OR2_X1 U2782 ( .A1(n3307), .A2(n3409), .ZN(n2220) );
  INV_X1 U2783 ( .A(IR_REG_9__SCAN_IN), .ZN(n2223) );
  AND2_X1 U2784 ( .A1(n3887), .A2(n3674), .ZN(n2552) );
  AND2_X1 U2785 ( .A1(n3584), .A2(n3864), .ZN(n3681) );
  AND2_X1 U2786 ( .A1(n2556), .A2(n2555), .ZN(n3553) );
  NAND2_X1 U2787 ( .A1(n3503), .A2(n3406), .ZN(n3300) );
  OR2_X1 U2788 ( .A1(n2651), .A2(n2248), .ZN(n2249) );
  NAND2_X1 U2789 ( .A1(n2886), .A2(REG2_REG_9__SCAN_IN), .ZN(n2892) );
  NAND2_X1 U2790 ( .A1(n4041), .A2(n2433), .ZN(n2434) );
  INV_X1 U2791 ( .A(IR_REG_17__SCAN_IN), .ZN(n2436) );
  INV_X1 U2792 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2358) );
  INV_X2 U2793 ( .A(n3338), .ZN(n3356) );
  INV_X1 U2794 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2329) );
  INV_X1 U2795 ( .A(n2791), .ZN(n2787) );
  NOR2_X1 U2796 ( .A1(n2463), .A2(n3434), .ZN(n2472) );
  INV_X1 U2797 ( .A(n2688), .ZN(n2671) );
  NAND2_X1 U2798 ( .A1(n2503), .A2(REG3_REG_26__SCAN_IN), .ZN(n2509) );
  NAND2_X1 U2799 ( .A1(n3926), .A2(n3917), .ZN(n2478) );
  INV_X1 U2800 ( .A(n3946), .ZN(n4272) );
  INV_X1 U2801 ( .A(n3810), .ZN(n3818) );
  INV_X1 U2802 ( .A(n3388), .ZN(n3266) );
  INV_X1 U2803 ( .A(n2909), .ZN(n3055) );
  OR2_X1 U2804 ( .A1(n2396), .A2(IR_REG_10__SCAN_IN), .ZN(n2373) );
  AND2_X1 U2805 ( .A1(n2479), .A2(REG3_REG_23__SCAN_IN), .ZN(n2487) );
  NOR2_X1 U2806 ( .A1(n2359), .A2(n2358), .ZN(n2367) );
  XNOR2_X1 U2807 ( .A(n2782), .B(n3324), .ZN(n2783) );
  OR2_X1 U2808 ( .A1(n2376), .A2(n2375), .ZN(n2386) );
  NOR2_X1 U2809 ( .A1(n2425), .A2(n2424), .ZN(n2440) );
  INV_X1 U2810 ( .A(n3869), .ZN(n3911) );
  AND2_X1 U2811 ( .A1(REG3_REG_22__SCAN_IN), .A2(n2472), .ZN(n2479) );
  OR2_X1 U2812 ( .A1(n2411), .A2(n3528), .ZN(n2425) );
  INV_X1 U2813 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4231) );
  INV_X1 U2814 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3243) );
  OR2_X1 U2815 ( .A1(n3820), .A2(n3364), .ZN(n3785) );
  INV_X1 U2816 ( .A(n3870), .ZN(n3839) );
  INV_X1 U2817 ( .A(n3926), .ZN(n3898) );
  AOI21_X1 U2818 ( .B1(n3939), .B2(n3578), .A(n3580), .ZN(n3922) );
  INV_X1 U2819 ( .A(n4023), .ZN(n3985) );
  INV_X1 U2820 ( .A(n3780), .ZN(n3769) );
  OR3_X1 U2821 ( .A1(n2930), .A2(n2929), .A3(n2928), .ZN(n2931) );
  INV_X1 U2822 ( .A(n2723), .ZN(n2606) );
  INV_X1 U2823 ( .A(n3841), .ZN(n2615) );
  OR2_X1 U2824 ( .A1(n3701), .A2(n4467), .ZN(n4549) );
  NOR2_X1 U2825 ( .A1(n2400), .A2(IR_REG_13__SCAN_IN), .ZN(n2418) );
  INV_X1 U2826 ( .A(n3973), .ZN(n3415) );
  INV_X1 U2827 ( .A(n3023), .ZN(n3419) );
  OR2_X1 U2828 ( .A1(n2346), .A2(n4231), .ZN(n2359) );
  INV_X1 U2829 ( .A(n3974), .ZN(n3991) );
  NOR2_X1 U2830 ( .A1(n2309), .A2(n2238), .ZN(n2321) );
  AND2_X1 U2831 ( .A1(n2260), .A2(n2259), .ZN(n2262) );
  AND2_X1 U2832 ( .A1(n2666), .A2(n4335), .ZN(n4450) );
  AND2_X1 U2833 ( .A1(n2666), .A2(n3698), .ZN(n4437) );
  AND2_X1 U2834 ( .A1(n2516), .A2(REG3_REG_28__SCAN_IN), .ZN(n3795) );
  AND2_X1 U2835 ( .A1(n2728), .A2(n2735), .ZN(n4024) );
  AOI21_X1 U2836 ( .B1(n2606), .B2(n4132), .A(n2645), .ZN(n2930) );
  INV_X1 U2837 ( .A(n3117), .ZN(n3125) );
  AND3_X1 U2838 ( .A1(n2609), .A2(n2608), .A3(n2607), .ZN(n2618) );
  NAND2_X1 U2839 ( .A1(n2587), .A2(n2630), .ZN(n2723) );
  XNOR2_X1 U2840 ( .A(n2594), .B(n2595), .ZN(n2806) );
  AND2_X1 U2841 ( .A1(n2650), .A2(n2648), .ZN(n4427) );
  INV_X1 U2842 ( .A(n3533), .ZN(n3114) );
  OR3_X1 U2843 ( .A1(n2741), .A2(n2740), .A3(n2739), .ZN(n3536) );
  OAI211_X1 U2844 ( .C1(n3433), .C2(n2468), .A(n2467), .B(n2466), .ZN(n3706)
         );
  INV_X1 U2845 ( .A(n3244), .ZN(n3709) );
  OR2_X1 U2846 ( .A1(n2623), .A2(n2805), .ZN(n3716) );
  INV_X1 U2847 ( .A(n4502), .ZN(n4362) );
  INV_X1 U2848 ( .A(n4498), .ZN(n4382) );
  INV_X1 U2849 ( .A(n4435), .ZN(n4441) );
  INV_X1 U2850 ( .A(n3999), .ZN(n4054) );
  INV_X1 U2851 ( .A(n4458), .ZN(n4050) );
  OR2_X1 U2852 ( .A1(n3373), .A2(n4268), .ZN(n2621) );
  NAND2_X1 U2853 ( .A1(n4567), .A2(n4545), .ZN(n4268) );
  INV_X1 U2854 ( .A(n4567), .ZN(n4564) );
  NAND2_X1 U2855 ( .A1(n4555), .A2(n4545), .ZN(n4325) );
  INV_X1 U2856 ( .A(n4555), .ZN(n4553) );
  INV_X1 U2857 ( .A(n4484), .ZN(n4483) );
  NAND2_X1 U2858 ( .A1(n2723), .A2(n2644), .ZN(n4484) );
  INV_X1 U2859 ( .A(n2886), .ZN(n4501) );
  INV_X1 U2860 ( .A(n3716), .ZN(U4043) );
  NAND4_X1 U2861 ( .A1(n2397), .A2(n2417), .A3(n2393), .A4(n2420), .ZN(n2225)
         );
  NAND4_X1 U2862 ( .A1(n2392), .A2(n4225), .A3(n2394), .A4(n2223), .ZN(n2224)
         );
  NOR2_X1 U2863 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2230)
         );
  NOR2_X1 U2864 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2229)
         );
  NOR2_X1 U2865 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2228)
         );
  NOR2_X1 U2866 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2227)
         );
  NAND4_X1 U2867 ( .A1(n2230), .A2(n2229), .A3(n2228), .A4(n2227), .ZN(n2231)
         );
  INV_X1 U2868 ( .A(n2240), .ZN(n2237) );
  NAND2_X1 U2869 ( .A1(n2234), .A2(IR_REG_31__SCAN_IN), .ZN(n2236) );
  NAND2_X1 U2870 ( .A1(n3538), .A2(REG1_REG_18__SCAN_IN), .ZN(n2245) );
  NAND2_X1 U2871 ( .A1(n2258), .A2(REG0_REG_18__SCAN_IN), .ZN(n2244) );
  AND2_X4 U2872 ( .A1(n2240), .A2(n2635), .ZN(n2265) );
  NAND2_X1 U2873 ( .A1(REG3_REG_5__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2238) );
  NAND2_X1 U2874 ( .A1(n2321), .A2(REG3_REG_7__SCAN_IN), .ZN(n2330) );
  NAND2_X1 U2875 ( .A1(n2367), .A2(REG3_REG_11__SCAN_IN), .ZN(n2376) );
  NAND2_X1 U2876 ( .A1(n2402), .A2(REG3_REG_14__SCAN_IN), .ZN(n2411) );
  OR2_X1 U2877 ( .A1(n2442), .A2(REG3_REG_18__SCAN_IN), .ZN(n2239) );
  AND2_X1 U2878 ( .A1(n2449), .A2(n2239), .ZN(n3994) );
  NAND2_X1 U2879 ( .A1(n2265), .A2(n3994), .ZN(n2243) );
  NAND2_X1 U2880 ( .A1(n2497), .A2(REG2_REG_18__SCAN_IN), .ZN(n2242) );
  NAND4_X1 U2881 ( .A1(n2245), .A2(n2244), .A3(n2243), .A4(n2242), .ZN(n4011)
         );
  INV_X1 U2882 ( .A(n4011), .ZN(n3972) );
  INV_X1 U2883 ( .A(n2435), .ZN(n2246) );
  NAND2_X1 U2884 ( .A1(n2246), .A2(n2436), .ZN(n2455) );
  NAND2_X1 U2885 ( .A1(n2455), .A2(IR_REG_31__SCAN_IN), .ZN(n2247) );
  XNOR2_X1 U2886 ( .A(n2247), .B(IR_REG_18__SCAN_IN), .ZN(n4449) );
  INV_X1 U2887 ( .A(n4449), .ZN(n4488) );
  INV_X1 U2888 ( .A(DATAI_18_), .ZN(n4487) );
  NAND2_X1 U2889 ( .A1(n2651), .A2(n2567), .ZN(n2250) );
  NAND2_X1 U2890 ( .A1(n2567), .A2(IR_REG_27__SCAN_IN), .ZN(n2251) );
  MUX2_X1 U2891 ( .A(n4488), .B(n4487), .S(n2295), .Z(n3974) );
  INV_X1 U2892 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2253) );
  INV_X1 U2893 ( .A(DATAI_1_), .ZN(n2256) );
  INV_X1 U2894 ( .A(n2647), .ZN(n2295) );
  MUX2_X1 U2895 ( .A(n2668), .B(n2256), .S(n2006), .Z(n3023) );
  NAND2_X1 U2896 ( .A1(n2257), .A2(n3419), .ZN(n2534) );
  NAND2_X1 U2897 ( .A1(n4273), .A2(n3023), .ZN(n3623) );
  NAND2_X1 U2898 ( .A1(n2534), .A2(n3623), .ZN(n2533) );
  NAND2_X1 U2899 ( .A1(n2497), .A2(REG2_REG_0__SCAN_IN), .ZN(n2263) );
  NAND2_X1 U2900 ( .A1(n2258), .A2(REG0_REG_0__SCAN_IN), .ZN(n2260) );
  NAND2_X1 U2901 ( .A1(n2265), .A2(REG3_REG_0__SCAN_IN), .ZN(n2259) );
  MUX2_X1 U2902 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(n2647), .Z(n4277) );
  AND2_X1 U2903 ( .A1(n3720), .A2(n4277), .ZN(n3018) );
  AND2_X1 U2904 ( .A1(n4273), .A2(n3419), .ZN(n2264) );
  AOI21_X1 U2905 ( .B1(n2533), .B2(n3018), .A(n2264), .ZN(n2754) );
  NAND2_X1 U2906 ( .A1(n2265), .A2(REG3_REG_2__SCAN_IN), .ZN(n2269) );
  NAND2_X1 U2907 ( .A1(n2258), .A2(REG0_REG_2__SCAN_IN), .ZN(n2268) );
  NAND2_X1 U2908 ( .A1(n2497), .A2(REG2_REG_2__SCAN_IN), .ZN(n2267) );
  NAND2_X1 U2909 ( .A1(n3538), .A2(REG1_REG_2__SCAN_IN), .ZN(n2266) );
  INV_X1 U2910 ( .A(DATAI_2_), .ZN(n2272) );
  MUX2_X1 U2911 ( .A(n2824), .B(n2272), .S(n2295), .Z(n2774) );
  NAND2_X1 U2912 ( .A1(n2273), .A2(n2774), .ZN(n3630) );
  NAND2_X1 U2913 ( .A1(n2754), .A2(n3598), .ZN(n2756) );
  INV_X1 U2914 ( .A(n2273), .ZN(n2938) );
  NAND2_X1 U2915 ( .A1(n2938), .A2(n2774), .ZN(n2274) );
  NAND2_X1 U2916 ( .A1(n2756), .A2(n2274), .ZN(n2927) );
  NAND2_X1 U2917 ( .A1(n3538), .A2(REG1_REG_3__SCAN_IN), .ZN(n2278) );
  INV_X1 U2918 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2286) );
  NAND2_X1 U2919 ( .A1(n2265), .A2(n2286), .ZN(n2277) );
  NAND2_X1 U2920 ( .A1(n2258), .A2(REG0_REG_3__SCAN_IN), .ZN(n2276) );
  NAND2_X1 U2921 ( .A1(n2497), .A2(REG2_REG_3__SCAN_IN), .ZN(n2275) );
  NAND4_X1 U2922 ( .A1(n2278), .A2(n2277), .A3(n2276), .A4(n2275), .ZN(n3718)
         );
  NAND2_X1 U2923 ( .A1(n2279), .A2(IR_REG_31__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2924 ( .A1(n2281), .A2(n2280), .ZN(n2292) );
  OR2_X1 U2925 ( .A1(n2281), .A2(n2280), .ZN(n2282) );
  MUX2_X1 U2926 ( .A(n2688), .B(DATAI_3_), .S(n2522), .Z(n2936) );
  NAND2_X1 U2927 ( .A1(n3718), .A2(n2936), .ZN(n2283) );
  NAND2_X1 U2928 ( .A1(n2927), .A2(n2283), .ZN(n2285) );
  INV_X1 U2929 ( .A(n3718), .ZN(n2848) );
  NAND2_X1 U2930 ( .A1(n2848), .A2(n2942), .ZN(n2284) );
  NAND2_X1 U2931 ( .A1(n2285), .A2(n2284), .ZN(n2948) );
  INV_X1 U2932 ( .A(n2948), .ZN(n2296) );
  NAND2_X1 U2933 ( .A1(n2497), .A2(REG2_REG_4__SCAN_IN), .ZN(n2291) );
  NAND2_X1 U2934 ( .A1(n3538), .A2(REG1_REG_4__SCAN_IN), .ZN(n2290) );
  INV_X1 U2935 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4220) );
  NAND2_X1 U2936 ( .A1(n2286), .A2(n4220), .ZN(n2287) );
  AND2_X1 U2937 ( .A1(n2287), .A2(n2309), .ZN(n2834) );
  NAND2_X1 U2938 ( .A1(n2265), .A2(n2834), .ZN(n2289) );
  NAND2_X1 U2939 ( .A1(n2258), .A2(REG0_REG_4__SCAN_IN), .ZN(n2288) );
  NAND2_X1 U2940 ( .A1(n2292), .A2(IR_REG_31__SCAN_IN), .ZN(n2294) );
  XNOR2_X1 U2941 ( .A(n2294), .B(n2293), .ZN(n2682) );
  INV_X1 U2942 ( .A(DATAI_4_), .ZN(n2624) );
  MUX2_X1 U2943 ( .A(n2682), .B(n2624), .S(n2522), .Z(n2958) );
  OR2_X1 U2944 ( .A1(n3717), .A2(n2958), .ZN(n3633) );
  NAND2_X1 U2945 ( .A1(n3717), .A2(n2958), .ZN(n3636) );
  NAND2_X1 U2946 ( .A1(n3633), .A2(n3636), .ZN(n2949) );
  NAND2_X1 U2947 ( .A1(n2296), .A2(n2949), .ZN(n2951) );
  NAND2_X1 U2948 ( .A1(n3717), .A2(n2850), .ZN(n2297) );
  NAND2_X1 U2949 ( .A1(n3538), .A2(REG1_REG_5__SCAN_IN), .ZN(n2301) );
  NAND2_X1 U2950 ( .A1(n2258), .A2(REG0_REG_5__SCAN_IN), .ZN(n2300) );
  XNOR2_X1 U2951 ( .A(n2309), .B(REG3_REG_5__SCAN_IN), .ZN(n2869) );
  NAND2_X1 U2952 ( .A1(n2265), .A2(n2869), .ZN(n2299) );
  NAND2_X1 U2953 ( .A1(n2497), .A2(REG2_REG_5__SCAN_IN), .ZN(n2298) );
  NAND2_X1 U2954 ( .A1(n2302), .A2(IR_REG_31__SCAN_IN), .ZN(n2303) );
  MUX2_X1 U2955 ( .A(IR_REG_31__SCAN_IN), .B(n2303), .S(IR_REG_5__SCAN_IN), 
        .Z(n2306) );
  INV_X1 U2956 ( .A(n2304), .ZN(n2305) );
  NAND2_X1 U2957 ( .A1(n2306), .A2(n2305), .ZN(n2707) );
  INV_X1 U2958 ( .A(DATAI_5_), .ZN(n2307) );
  MUX2_X1 U2959 ( .A(n2707), .B(n2307), .S(n2522), .Z(n2875) );
  NAND2_X1 U2960 ( .A1(n3048), .A2(n2875), .ZN(n2308) );
  INV_X1 U2961 ( .A(n3048), .ZN(n3715) );
  NAND2_X1 U2962 ( .A1(n2497), .A2(REG2_REG_6__SCAN_IN), .ZN(n2315) );
  NAND2_X1 U2963 ( .A1(n3538), .A2(REG1_REG_6__SCAN_IN), .ZN(n2314) );
  INV_X1 U2964 ( .A(n2309), .ZN(n2310) );
  AOI21_X1 U2965 ( .B1(n2310), .B2(REG3_REG_5__SCAN_IN), .A(
        REG3_REG_6__SCAN_IN), .ZN(n2311) );
  OR2_X1 U2966 ( .A1(n2311), .A2(n2321), .ZN(n2912) );
  INV_X1 U2967 ( .A(n2912), .ZN(n4454) );
  NAND2_X1 U2968 ( .A1(n2265), .A2(n4454), .ZN(n2313) );
  NAND2_X1 U2969 ( .A1(n2258), .A2(REG0_REG_6__SCAN_IN), .ZN(n2312) );
  NAND4_X1 U2970 ( .A1(n2315), .A2(n2314), .A3(n2313), .A4(n2312), .ZN(n3714)
         );
  NOR2_X1 U2971 ( .A1(n2304), .A2(n2640), .ZN(n2316) );
  MUX2_X1 U2972 ( .A(n2640), .B(n2316), .S(IR_REG_6__SCAN_IN), .Z(n2318) );
  OR2_X1 U2973 ( .A1(n2318), .A2(n2317), .ZN(n4505) );
  MUX2_X1 U2974 ( .A(n2709), .B(DATAI_6_), .S(n2522), .Z(n2909) );
  INV_X1 U2975 ( .A(n3714), .ZN(n2922) );
  NAND2_X1 U2976 ( .A1(n2922), .A2(n3055), .ZN(n2319) );
  INV_X1 U2977 ( .A(n2320), .ZN(n2995) );
  NAND2_X1 U2978 ( .A1(n2497), .A2(REG2_REG_7__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U2979 ( .A1(n3538), .A2(REG1_REG_7__SCAN_IN), .ZN(n2325) );
  OR2_X1 U2980 ( .A1(n2321), .A2(REG3_REG_7__SCAN_IN), .ZN(n2322) );
  AND2_X1 U2981 ( .A1(n2330), .A2(n2322), .ZN(n2994) );
  NAND2_X1 U2982 ( .A1(n2265), .A2(n2994), .ZN(n2324) );
  NAND2_X1 U2983 ( .A1(n2258), .A2(REG0_REG_7__SCAN_IN), .ZN(n2323) );
  NAND4_X1 U2984 ( .A1(n2326), .A2(n2325), .A3(n2324), .A4(n2323), .ZN(n3713)
         );
  OR2_X1 U2985 ( .A1(n2317), .A2(n2640), .ZN(n2328) );
  NAND2_X1 U2986 ( .A1(n2328), .A2(n2327), .ZN(n2336) );
  OAI21_X1 U2987 ( .B1(n2328), .B2(n2327), .A(n2336), .ZN(n2888) );
  INV_X1 U2988 ( .A(DATAI_7_), .ZN(n4177) );
  MUX2_X1 U2989 ( .A(n2888), .B(n4177), .S(n2522), .Z(n2991) );
  OR2_X1 U2990 ( .A1(n3713), .A2(n2991), .ZN(n2538) );
  NAND2_X1 U2991 ( .A1(n3713), .A2(n2991), .ZN(n3648) );
  NAND2_X1 U2992 ( .A1(n2538), .A2(n3648), .ZN(n3638) );
  NAND2_X1 U2993 ( .A1(n3538), .A2(REG1_REG_8__SCAN_IN), .ZN(n2335) );
  NAND2_X1 U2994 ( .A1(n2258), .A2(REG0_REG_8__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U2995 ( .A1(n2330), .A2(n2329), .ZN(n2331) );
  AND2_X1 U2996 ( .A1(n2346), .A2(n2331), .ZN(n3041) );
  NAND2_X1 U2997 ( .A1(n2265), .A2(n3041), .ZN(n2333) );
  NAND2_X1 U2998 ( .A1(n2497), .A2(REG2_REG_8__SCAN_IN), .ZN(n2332) );
  NAND2_X1 U2999 ( .A1(n2336), .A2(IR_REG_31__SCAN_IN), .ZN(n2337) );
  XNOR2_X1 U3000 ( .A(n2337), .B(IR_REG_8__SCAN_IN), .ZN(n4502) );
  INV_X1 U3001 ( .A(DATAI_8_), .ZN(n2338) );
  MUX2_X1 U3002 ( .A(n4362), .B(n2338), .S(n2522), .Z(n3032) );
  NAND2_X1 U3003 ( .A1(n3081), .A2(n3032), .ZN(n2340) );
  AND2_X1 U3004 ( .A1(n3638), .A2(n2340), .ZN(n2339) );
  NAND2_X1 U3005 ( .A1(n2995), .A2(n2339), .ZN(n2345) );
  INV_X1 U3006 ( .A(n2340), .ZN(n2343) );
  INV_X1 U3007 ( .A(n2991), .ZN(n2916) );
  NAND2_X1 U3008 ( .A1(n3713), .A2(n2916), .ZN(n3036) );
  NAND2_X1 U3009 ( .A1(n3712), .A2(n3040), .ZN(n2341) );
  AND2_X1 U3010 ( .A1(n3036), .A2(n2341), .ZN(n2342) );
  NAND2_X1 U3011 ( .A1(n2345), .A2(n2344), .ZN(n3085) );
  NAND2_X1 U3012 ( .A1(n2497), .A2(REG2_REG_9__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U3013 ( .A1(n3538), .A2(REG1_REG_9__SCAN_IN), .ZN(n2351) );
  NAND2_X1 U3014 ( .A1(n2346), .A2(n4231), .ZN(n2347) );
  NAND2_X1 U3015 ( .A1(n2359), .A2(n2347), .ZN(n3092) );
  INV_X1 U3016 ( .A(n3092), .ZN(n2348) );
  NAND2_X1 U3017 ( .A1(n2265), .A2(n2348), .ZN(n2350) );
  NAND2_X1 U3018 ( .A1(n2258), .A2(REG0_REG_9__SCAN_IN), .ZN(n2349) );
  NAND4_X1 U3019 ( .A1(n2352), .A2(n2351), .A3(n2350), .A4(n2349), .ZN(n3711)
         );
  NAND2_X1 U3020 ( .A1(n2353), .A2(IR_REG_31__SCAN_IN), .ZN(n2354) );
  MUX2_X1 U3021 ( .A(IR_REG_31__SCAN_IN), .B(n2354), .S(IR_REG_9__SCAN_IN), 
        .Z(n2355) );
  MUX2_X1 U3022 ( .A(n2886), .B(DATAI_9_), .S(n2522), .Z(n3091) );
  AND2_X1 U3023 ( .A1(n3711), .A2(n3091), .ZN(n2357) );
  OR2_X1 U3024 ( .A1(n3711), .A2(n3091), .ZN(n2356) );
  NAND2_X1 U3025 ( .A1(n3538), .A2(REG1_REG_10__SCAN_IN), .ZN(n2364) );
  NAND2_X1 U3026 ( .A1(n2258), .A2(REG0_REG_10__SCAN_IN), .ZN(n2363) );
  AND2_X1 U3027 ( .A1(n2359), .A2(n2358), .ZN(n2360) );
  NOR2_X1 U3028 ( .A1(n2367), .A2(n2360), .ZN(n3127) );
  NAND2_X1 U3029 ( .A1(n2265), .A2(n3127), .ZN(n2362) );
  NAND2_X1 U3030 ( .A1(n2497), .A2(REG2_REG_10__SCAN_IN), .ZN(n2361) );
  NAND4_X1 U3031 ( .A1(n2364), .A2(n2363), .A3(n2362), .A4(n2361), .ZN(n3191)
         );
  NAND2_X1 U3032 ( .A1(n2396), .A2(IR_REG_31__SCAN_IN), .ZN(n2365) );
  XNOR2_X1 U3033 ( .A(n2365), .B(IR_REG_10__SCAN_IN), .ZN(n4331) );
  MUX2_X1 U3034 ( .A(n4331), .B(DATAI_10_), .S(n2522), .Z(n3117) );
  NOR2_X1 U3035 ( .A1(n3191), .A2(n3117), .ZN(n2366) );
  INV_X1 U3036 ( .A(n3191), .ZN(n3154) );
  NAND2_X1 U3037 ( .A1(n3538), .A2(REG1_REG_11__SCAN_IN), .ZN(n2372) );
  NAND2_X1 U3038 ( .A1(n2258), .A2(REG0_REG_11__SCAN_IN), .ZN(n2371) );
  OR2_X1 U3039 ( .A1(n2367), .A2(REG3_REG_11__SCAN_IN), .ZN(n2368) );
  AND2_X1 U3040 ( .A1(n2368), .A2(n2376), .ZN(n3197) );
  NAND2_X1 U3041 ( .A1(n2265), .A2(n3197), .ZN(n2370) );
  NAND2_X1 U3042 ( .A1(n2497), .A2(REG2_REG_11__SCAN_IN), .ZN(n2369) );
  NAND4_X1 U3043 ( .A1(n2372), .A2(n2371), .A3(n2370), .A4(n2369), .ZN(n3710)
         );
  NAND2_X1 U3044 ( .A1(n2373), .A2(IR_REG_31__SCAN_IN), .ZN(n2382) );
  INV_X1 U3045 ( .A(DATAI_11_), .ZN(n2374) );
  MUX2_X1 U3046 ( .A(n4382), .B(n2374), .S(n2522), .Z(n3195) );
  OR2_X1 U3047 ( .A1(n3710), .A2(n3195), .ZN(n3621) );
  NAND2_X1 U3048 ( .A1(n3710), .A2(n3195), .ZN(n3660) );
  NAND2_X1 U3049 ( .A1(n3621), .A2(n3660), .ZN(n3186) );
  INV_X1 U3050 ( .A(n3710), .ZN(n3173) );
  NAND2_X1 U3051 ( .A1(n2497), .A2(REG2_REG_12__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3052 ( .A1(n3538), .A2(REG1_REG_12__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U3053 ( .A1(n2376), .A2(n2375), .ZN(n2377) );
  AND2_X1 U3054 ( .A1(n2386), .A2(n2377), .ZN(n3176) );
  NAND2_X1 U3055 ( .A1(n2265), .A2(n3176), .ZN(n2379) );
  NAND2_X1 U3056 ( .A1(n2258), .A2(REG0_REG_12__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3057 ( .A1(n2382), .A2(n2394), .ZN(n2383) );
  NAND2_X1 U3058 ( .A1(n2383), .A2(IR_REG_31__SCAN_IN), .ZN(n2384) );
  XNOR2_X1 U3059 ( .A(n2384), .B(IR_REG_12__SCAN_IN), .ZN(n3753) );
  MUX2_X1 U3060 ( .A(n3753), .B(DATAI_12_), .S(n2522), .Z(n3140) );
  NAND2_X1 U3061 ( .A1(n3709), .A2(n3140), .ZN(n2385) );
  NAND2_X1 U3062 ( .A1(n2497), .A2(REG2_REG_13__SCAN_IN), .ZN(n2391) );
  NAND2_X1 U3063 ( .A1(n3538), .A2(REG1_REG_13__SCAN_IN), .ZN(n2390) );
  AND2_X1 U3064 ( .A1(n2386), .A2(n3243), .ZN(n2387) );
  NOR2_X1 U3065 ( .A1(n2402), .A2(n2387), .ZN(n3247) );
  NAND2_X1 U3066 ( .A1(n2265), .A2(n3247), .ZN(n2389) );
  NAND2_X1 U3067 ( .A1(n2258), .A2(REG0_REG_13__SCAN_IN), .ZN(n2388) );
  NAND4_X1 U3068 ( .A1(n2391), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n3708)
         );
  NAND3_X1 U3069 ( .A1(n2394), .A2(n2393), .A3(n2392), .ZN(n2395) );
  NAND2_X1 U3070 ( .A1(n2400), .A2(IR_REG_31__SCAN_IN), .ZN(n2398) );
  MUX2_X1 U3071 ( .A(n2398), .B(IR_REG_31__SCAN_IN), .S(n2397), .Z(n2399) );
  INV_X1 U3072 ( .A(n2399), .ZN(n2401) );
  MUX2_X1 U3073 ( .A(n4398), .B(DATAI_13_), .S(n2006), .Z(n3246) );
  OR2_X1 U3074 ( .A1(n3708), .A2(n3246), .ZN(n3217) );
  AND2_X1 U3075 ( .A1(n3708), .A2(n3246), .ZN(n3216) );
  AOI21_X1 U3076 ( .B1(n3219), .B2(n3217), .A(n3216), .ZN(n3207) );
  NAND2_X1 U3077 ( .A1(n2497), .A2(REG2_REG_14__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U3078 ( .A1(n3538), .A2(REG1_REG_14__SCAN_IN), .ZN(n2406) );
  OR2_X1 U3079 ( .A1(n2402), .A2(REG3_REG_14__SCAN_IN), .ZN(n2403) );
  AND2_X1 U3080 ( .A1(n2411), .A2(n2403), .ZN(n3392) );
  NAND2_X1 U3081 ( .A1(n2265), .A2(n3392), .ZN(n2405) );
  NAND2_X1 U3082 ( .A1(n2258), .A2(REG0_REG_14__SCAN_IN), .ZN(n2404) );
  NAND4_X1 U3083 ( .A1(n2407), .A2(n2406), .A3(n2405), .A4(n2404), .ZN(n3707)
         );
  OR2_X1 U3084 ( .A1(n2418), .A2(n2640), .ZN(n2408) );
  XNOR2_X1 U3085 ( .A(n2408), .B(IR_REG_14__SCAN_IN), .ZN(n4493) );
  INV_X1 U3086 ( .A(DATAI_14_), .ZN(n2409) );
  MUX2_X1 U3087 ( .A(n3757), .B(n2409), .S(n2522), .Z(n3388) );
  OR2_X1 U3088 ( .A1(n3707), .A2(n3388), .ZN(n3546) );
  NAND2_X1 U3089 ( .A1(n3707), .A2(n3388), .ZN(n3547) );
  NAND2_X1 U3090 ( .A1(n3546), .A2(n3547), .ZN(n3209) );
  NAND2_X1 U3091 ( .A1(n3207), .A2(n3209), .ZN(n3208) );
  NAND2_X1 U3092 ( .A1(n3208), .A2(n2410), .ZN(n4038) );
  NAND2_X1 U3093 ( .A1(n2497), .A2(REG2_REG_15__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U3094 ( .A1(n3538), .A2(REG1_REG_15__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3095 ( .A1(n2411), .A2(n3528), .ZN(n2412) );
  AND2_X1 U3096 ( .A1(n2425), .A2(n2412), .ZN(n4048) );
  NAND2_X1 U3097 ( .A1(n2265), .A2(n4048), .ZN(n2414) );
  NAND2_X1 U3098 ( .A1(n2258), .A2(REG0_REG_15__SCAN_IN), .ZN(n2413) );
  NAND2_X1 U3099 ( .A1(n2418), .A2(n2417), .ZN(n2419) );
  NAND2_X1 U3100 ( .A1(n2419), .A2(IR_REG_31__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U3101 ( .A1(n2421), .A2(n2420), .ZN(n2431) );
  OR2_X1 U3102 ( .A1(n2421), .A2(n2420), .ZN(n2422) );
  MUX2_X1 U3103 ( .A(n3759), .B(DATAI_15_), .S(n2522), .Z(n4046) );
  NAND2_X1 U3104 ( .A1(n4025), .A2(n4046), .ZN(n2423) );
  NAND2_X1 U3105 ( .A1(n2497), .A2(REG2_REG_16__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3106 ( .A1(n3538), .A2(REG1_REG_16__SCAN_IN), .ZN(n2429) );
  AND2_X1 U3107 ( .A1(n2425), .A2(n2424), .ZN(n2426) );
  NOR2_X1 U3108 ( .A1(n2440), .A2(n2426), .ZN(n4033) );
  NAND2_X1 U3109 ( .A1(n2265), .A2(n4033), .ZN(n2428) );
  NAND2_X1 U3110 ( .A1(n2258), .A2(REG0_REG_16__SCAN_IN), .ZN(n2427) );
  NAND4_X1 U3111 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .ZN(n4041)
         );
  NAND2_X1 U3112 ( .A1(n2431), .A2(IR_REG_31__SCAN_IN), .ZN(n2432) );
  XNOR2_X1 U3113 ( .A(n2432), .B(n4225), .ZN(n4490) );
  INV_X1 U3114 ( .A(DATAI_16_), .ZN(n4489) );
  MUX2_X1 U3115 ( .A(n4490), .B(n4489), .S(n2006), .Z(n4028) );
  OR2_X1 U3116 ( .A1(n4041), .A2(n4028), .ZN(n3669) );
  NAND2_X1 U3117 ( .A1(n4041), .A2(n4028), .ZN(n3551) );
  NAND2_X1 U3118 ( .A1(n3669), .A2(n3551), .ZN(n4018) );
  NAND2_X1 U3119 ( .A1(n4017), .A2(n2434), .ZN(n4002) );
  NAND2_X1 U3120 ( .A1(n2435), .A2(IR_REG_31__SCAN_IN), .ZN(n2437) );
  MUX2_X1 U3121 ( .A(n2437), .B(IR_REG_31__SCAN_IN), .S(n2436), .Z(n2438) );
  NAND2_X1 U3122 ( .A1(n2438), .A2(n2455), .ZN(n3749) );
  INV_X1 U3123 ( .A(DATAI_17_), .ZN(n2439) );
  MUX2_X1 U3124 ( .A(n3749), .B(n2439), .S(n2006), .Z(n3467) );
  NAND2_X1 U3125 ( .A1(n3538), .A2(REG1_REG_17__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3126 ( .A1(n2258), .A2(REG0_REG_17__SCAN_IN), .ZN(n2445) );
  NOR2_X1 U3127 ( .A1(n2440), .A2(REG3_REG_17__SCAN_IN), .ZN(n2441) );
  OR2_X1 U3128 ( .A1(n2442), .A2(n2441), .ZN(n4004) );
  INV_X1 U3129 ( .A(n4004), .ZN(n3470) );
  NAND2_X1 U3130 ( .A1(n2265), .A2(n3470), .ZN(n2444) );
  NAND2_X1 U3131 ( .A1(n2497), .A2(REG2_REG_17__SCAN_IN), .ZN(n2443) );
  NAND4_X1 U3132 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n4023)
         );
  NAND2_X1 U3133 ( .A1(n4002), .A2(n2447), .ZN(n2448) );
  OR2_X1 U3134 ( .A1(n4011), .A2(n3974), .ZN(n3962) );
  NAND2_X1 U3135 ( .A1(n4011), .A2(n3974), .ZN(n3963) );
  INV_X1 U3136 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3413) );
  NAND2_X1 U3137 ( .A1(n2449), .A2(n3413), .ZN(n2450) );
  AND2_X1 U3138 ( .A1(n2459), .A2(n2450), .ZN(n3977) );
  NAND2_X1 U3139 ( .A1(n3977), .A2(n2265), .ZN(n2454) );
  NAND2_X1 U3140 ( .A1(n3538), .A2(REG1_REG_19__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U3141 ( .A1(n2258), .A2(REG0_REG_19__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3142 ( .A1(n2497), .A2(REG2_REG_19__SCAN_IN), .ZN(n2451) );
  NAND4_X1 U3143 ( .A1(n2454), .A2(n2453), .A3(n2452), .A4(n2451), .ZN(n3983)
         );
  INV_X1 U3144 ( .A(n2455), .ZN(n2457) );
  NAND2_X1 U3145 ( .A1(n2457), .A2(n2456), .ZN(n2523) );
  NAND2_X1 U3146 ( .A1(n2523), .A2(IR_REG_31__SCAN_IN), .ZN(n2527) );
  INV_X1 U3147 ( .A(DATAI_19_), .ZN(n2458) );
  MUX2_X1 U31480 ( .A(n3780), .B(n2458), .S(n2006), .Z(n3973) );
  OR2_X1 U31490 ( .A1(n3983), .A2(n3415), .ZN(n3582) );
  AND2_X1 U3150 ( .A1(n3983), .A2(n3415), .ZN(n3581) );
  INV_X1 U3151 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3488) );
  NAND2_X1 U3152 ( .A1(n2459), .A2(n3488), .ZN(n2460) );
  NAND2_X1 U3153 ( .A1(n2463), .A2(n2460), .ZN(n3487) );
  INV_X1 U3154 ( .A(n2265), .ZN(n2468) );
  AOI22_X1 U3155 ( .A1(n2497), .A2(REG2_REG_20__SCAN_IN), .B1(n2258), .B2(
        REG0_REG_20__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U3156 ( .A1(n3538), .A2(REG1_REG_20__SCAN_IN), .ZN(n2461) );
  INV_X1 U3157 ( .A(n3953), .ZN(n3944) );
  NAND2_X1 U3158 ( .A1(n3969), .A2(n3944), .ZN(n3578) );
  NOR2_X1 U3159 ( .A1(n3969), .A2(n3944), .ZN(n3580) );
  INV_X1 U3160 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3434) );
  NAND2_X1 U3161 ( .A1(n2463), .A2(n3434), .ZN(n2465) );
  INV_X1 U3162 ( .A(n2472), .ZN(n2464) );
  NAND2_X1 U3163 ( .A1(n2465), .A2(n2464), .ZN(n3433) );
  AOI22_X1 U3164 ( .A1(n2497), .A2(REG2_REG_21__SCAN_IN), .B1(n3538), .B2(
        REG1_REG_21__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U3165 ( .A1(n2258), .A2(REG0_REG_21__SCAN_IN), .ZN(n2466) );
  INV_X1 U3166 ( .A(n3706), .ZN(n3947) );
  OAI21_X1 U3167 ( .B1(n3922), .B2(n2470), .A(n2469), .ZN(n2471) );
  INV_X1 U3168 ( .A(n2471), .ZN(n3906) );
  NAND2_X1 U3169 ( .A1(n3538), .A2(REG1_REG_22__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U3170 ( .A1(n2258), .A2(REG0_REG_22__SCAN_IN), .ZN(n2476) );
  NOR2_X1 U3171 ( .A1(REG3_REG_22__SCAN_IN), .A2(n2472), .ZN(n2473) );
  NOR2_X1 U3172 ( .A1(n2479), .A2(n2473), .ZN(n3915) );
  NAND2_X1 U3173 ( .A1(n2265), .A2(n3915), .ZN(n2475) );
  NAND2_X1 U3174 ( .A1(n2497), .A2(REG2_REG_22__SCAN_IN), .ZN(n2474) );
  NAND4_X1 U3175 ( .A1(n2477), .A2(n2476), .A3(n2475), .A4(n2474), .ZN(n3926)
         );
  OR2_X1 U3176 ( .A1(n3926), .A2(n3910), .ZN(n3890) );
  NAND2_X1 U3177 ( .A1(n3926), .A2(n3910), .ZN(n2554) );
  NAND2_X1 U3178 ( .A1(n3890), .A2(n2554), .ZN(n3908) );
  NAND2_X1 U3179 ( .A1(n3906), .A2(n3908), .ZN(n3907) );
  NAND2_X1 U3180 ( .A1(n3907), .A2(n2478), .ZN(n3882) );
  NAND2_X1 U3181 ( .A1(n3538), .A2(REG1_REG_23__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3182 ( .A1(n2258), .A2(REG0_REG_23__SCAN_IN), .ZN(n2483) );
  NOR2_X1 U3183 ( .A1(n2479), .A2(REG3_REG_23__SCAN_IN), .ZN(n2480) );
  NOR2_X1 U3184 ( .A1(n2487), .A2(n2480), .ZN(n3902) );
  NAND2_X1 U3185 ( .A1(n2265), .A2(n3902), .ZN(n2482) );
  NAND2_X1 U3186 ( .A1(n2497), .A2(REG2_REG_23__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3187 ( .A1(n3911), .A2(n3901), .ZN(n2486) );
  INV_X1 U3188 ( .A(n3901), .ZN(n2485) );
  NAND2_X1 U3189 ( .A1(n2497), .A2(REG2_REG_24__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U3190 ( .A1(n3538), .A2(REG1_REG_24__SCAN_IN), .ZN(n2491) );
  NOR2_X1 U3191 ( .A1(n2487), .A2(REG3_REG_24__SCAN_IN), .ZN(n2488) );
  NOR2_X1 U3192 ( .A1(n2495), .A2(n2488), .ZN(n3877) );
  NAND2_X1 U3193 ( .A1(n2265), .A2(n3877), .ZN(n2490) );
  NAND2_X1 U3194 ( .A1(n2258), .A2(REG0_REG_24__SCAN_IN), .ZN(n2489) );
  INV_X1 U3195 ( .A(n3876), .ZN(n2493) );
  NAND2_X1 U3196 ( .A1(n3895), .A2(n2493), .ZN(n2494) );
  NAND2_X1 U3197 ( .A1(n3538), .A2(REG1_REG_25__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U3198 ( .A1(n2258), .A2(REG0_REG_25__SCAN_IN), .ZN(n2500) );
  NOR2_X1 U3199 ( .A1(n2495), .A2(REG3_REG_25__SCAN_IN), .ZN(n2496) );
  NOR2_X1 U3200 ( .A1(n2503), .A2(n2496), .ZN(n3859) );
  NAND2_X1 U3201 ( .A1(n2265), .A2(n3859), .ZN(n2499) );
  NAND2_X1 U3202 ( .A1(n2497), .A2(REG2_REG_25__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U3203 ( .A1(n3839), .A2(n3857), .ZN(n2502) );
  INV_X1 U3204 ( .A(n3857), .ZN(n2614) );
  NAND2_X1 U3205 ( .A1(n3538), .A2(REG1_REG_26__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3206 ( .A1(n2258), .A2(REG0_REG_26__SCAN_IN), .ZN(n2507) );
  OAI21_X1 U3207 ( .B1(n2503), .B2(REG3_REG_26__SCAN_IN), .A(n2509), .ZN(n2504) );
  INV_X1 U3208 ( .A(n2504), .ZN(n3842) );
  NAND2_X1 U3209 ( .A1(n2265), .A2(n3842), .ZN(n2506) );
  NAND2_X1 U32100 ( .A1(n2497), .A2(REG2_REG_26__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U32110 ( .A1(n2295), .A2(DATAI_26_), .ZN(n3841) );
  NOR2_X1 U32120 ( .A1(n3852), .A2(n2615), .ZN(n3587) );
  NAND2_X1 U32130 ( .A1(n3538), .A2(REG1_REG_27__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U32140 ( .A1(n2258), .A2(REG0_REG_27__SCAN_IN), .ZN(n2513) );
  INV_X1 U32150 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4179) );
  AND2_X1 U32160 ( .A1(n2509), .A2(n4179), .ZN(n2510) );
  NOR2_X1 U32170 ( .A1(n2516), .A2(n2510), .ZN(n3814) );
  NAND2_X1 U32180 ( .A1(n2265), .A2(n3814), .ZN(n2512) );
  NAND2_X1 U32190 ( .A1(n2497), .A2(REG2_REG_27__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U32200 ( .A1(n2006), .A2(DATAI_27_), .ZN(n3823) );
  INV_X1 U32210 ( .A(n3823), .ZN(n3811) );
  INV_X1 U32220 ( .A(n3836), .ZN(n3518) );
  NAND2_X1 U32230 ( .A1(n3538), .A2(REG1_REG_28__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U32240 ( .A1(n2258), .A2(REG0_REG_28__SCAN_IN), .ZN(n2520) );
  NOR2_X1 U32250 ( .A1(n2516), .A2(REG3_REG_28__SCAN_IN), .ZN(n2517) );
  NOR2_X1 U32260 ( .A1(n3795), .A2(n2517), .ZN(n3371) );
  NAND2_X1 U32270 ( .A1(n2265), .A2(n3371), .ZN(n2519) );
  NAND2_X1 U32280 ( .A1(n2497), .A2(REG2_REG_28__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U32290 ( .A1(n2522), .A2(DATAI_28_), .ZN(n3364) );
  NAND2_X1 U32300 ( .A1(n3820), .A2(n3364), .ZN(n3566) );
  NAND2_X1 U32310 ( .A1(n3785), .A2(n3566), .ZN(n3797) );
  XNOR2_X1 U32320 ( .A(n3798), .B(n3797), .ZN(n3377) );
  NAND2_X1 U32330 ( .A1(n2524), .A2(n2212), .ZN(n2581) );
  NAND2_X1 U32340 ( .A1(n2527), .A2(n2526), .ZN(n2528) );
  NAND2_X1 U32350 ( .A1(n2528), .A2(IR_REG_31__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U32360 ( .A1(n2581), .A2(IR_REG_31__SCAN_IN), .ZN(n2531) );
  XNOR2_X1 U32370 ( .A(n2725), .B(n3701), .ZN(n2532) );
  NAND2_X1 U32380 ( .A1(n3694), .A2(n3769), .ZN(n4467) );
  INV_X1 U32390 ( .A(n2533), .ZN(n3020) );
  NOR2_X1 U32400 ( .A1(n3720), .A2(n3601), .ZN(n3626) );
  NAND2_X1 U32410 ( .A1(n3020), .A2(n3626), .ZN(n3019) );
  NAND2_X1 U32420 ( .A1(n3019), .A2(n2534), .ZN(n2536) );
  INV_X1 U32430 ( .A(n3598), .ZN(n2535) );
  NAND2_X1 U32440 ( .A1(n2536), .A2(n2535), .ZN(n2758) );
  NAND2_X1 U32450 ( .A1(n2758), .A2(n3627), .ZN(n2934) );
  OR2_X1 U32460 ( .A1(n3718), .A2(n2942), .ZN(n3632) );
  NAND2_X1 U32470 ( .A1(n3718), .A2(n2942), .ZN(n3629) );
  NAND2_X1 U32480 ( .A1(n3632), .A2(n3629), .ZN(n3596) );
  INV_X1 U32490 ( .A(n3596), .ZN(n2935) );
  INV_X1 U32500 ( .A(n3633), .ZN(n2537) );
  AND2_X1 U32510 ( .A1(n3715), .A2(n2875), .ZN(n2970) );
  OR2_X1 U32520 ( .A1(n3715), .A2(n2875), .ZN(n3649) );
  OAI21_X1 U32530 ( .B1(n2971), .B2(n2970), .A(n3649), .ZN(n3049) );
  NAND2_X1 U32540 ( .A1(n3714), .A2(n3055), .ZN(n3651) );
  OR2_X1 U32550 ( .A1(n3714), .A2(n3055), .ZN(n3639) );
  INV_X1 U32560 ( .A(n2538), .ZN(n2539) );
  OR2_X1 U32570 ( .A1(n3712), .A2(n3032), .ZN(n3643) );
  NAND2_X1 U32580 ( .A1(n3031), .A2(n3643), .ZN(n2540) );
  NAND2_X1 U32590 ( .A1(n3712), .A2(n3032), .ZN(n3652) );
  AND2_X1 U32600 ( .A1(n3711), .A2(n2081), .ZN(n3646) );
  OR2_X1 U32610 ( .A1(n3711), .A2(n2081), .ZN(n3644) );
  NAND2_X1 U32620 ( .A1(n3191), .A2(n3125), .ZN(n3661) );
  OR2_X1 U32630 ( .A1(n3191), .A2(n3125), .ZN(n3655) );
  NAND2_X1 U32640 ( .A1(n2541), .A2(n3655), .ZN(n3187) );
  NAND2_X1 U32650 ( .A1(n3187), .A2(n3660), .ZN(n2542) );
  NAND2_X1 U32660 ( .A1(n2542), .A2(n3621), .ZN(n3222) );
  NAND2_X1 U32670 ( .A1(n3709), .A2(n3172), .ZN(n3220) );
  INV_X1 U32680 ( .A(n3246), .ZN(n3238) );
  NAND2_X1 U32690 ( .A1(n3708), .A2(n3238), .ZN(n2543) );
  NAND2_X1 U32700 ( .A1(n3222), .A2(n3617), .ZN(n2545) );
  NOR2_X1 U32710 ( .A1(n3709), .A2(n3172), .ZN(n3221) );
  NOR2_X1 U32720 ( .A1(n3708), .A2(n3238), .ZN(n2544) );
  AOI21_X1 U32730 ( .B1(n3617), .B2(n3221), .A(n2544), .ZN(n3620) );
  NAND2_X1 U32740 ( .A1(n2545), .A2(n3620), .ZN(n3550) );
  INV_X1 U32750 ( .A(n3209), .ZN(n3591) );
  NAND2_X1 U32760 ( .A1(n3550), .A2(n3591), .ZN(n2546) );
  OR2_X1 U32770 ( .A1(n4025), .A2(n3275), .ZN(n3549) );
  NAND2_X1 U32780 ( .A1(n4025), .A2(n3275), .ZN(n3548) );
  INV_X1 U32790 ( .A(n4018), .ZN(n4021) );
  NAND2_X1 U32800 ( .A1(n3983), .A2(n3973), .ZN(n2547) );
  AND2_X1 U32810 ( .A1(n2547), .A2(n3963), .ZN(n3884) );
  OR2_X1 U32820 ( .A1(n4023), .A2(n3467), .ZN(n3960) );
  NAND2_X1 U32830 ( .A1(n3962), .A2(n3960), .ZN(n2549) );
  NOR2_X1 U32840 ( .A1(n3983), .A2(n3973), .ZN(n2548) );
  AOI21_X1 U32850 ( .B1(n3884), .B2(n2549), .A(n2548), .ZN(n3940) );
  OR2_X1 U32860 ( .A1(n3969), .A2(n3953), .ZN(n2550) );
  NAND2_X1 U32870 ( .A1(n3940), .A2(n2550), .ZN(n2551) );
  NAND2_X1 U32880 ( .A1(n3969), .A2(n3953), .ZN(n3886) );
  NAND2_X1 U32890 ( .A1(n2551), .A2(n3886), .ZN(n3887) );
  OR2_X1 U32900 ( .A1(n3706), .A2(n3932), .ZN(n3577) );
  AND2_X1 U32910 ( .A1(n3577), .A2(n3890), .ZN(n3674) );
  NAND2_X1 U32920 ( .A1(n4008), .A2(n2552), .ZN(n2557) );
  INV_X1 U32930 ( .A(n2552), .ZN(n3554) );
  NAND2_X1 U32940 ( .A1(n4023), .A2(n3467), .ZN(n3883) );
  AND3_X1 U32950 ( .A1(n3884), .A2(n3886), .A3(n3883), .ZN(n3672) );
  OR2_X1 U32960 ( .A1(n3554), .A2(n3672), .ZN(n2556) );
  AND2_X1 U32970 ( .A1(n3706), .A2(n3932), .ZN(n3676) );
  NAND2_X1 U32980 ( .A1(n3869), .A2(n3901), .ZN(n2553) );
  NAND2_X1 U32990 ( .A1(n2554), .A2(n2553), .ZN(n3680) );
  AOI21_X1 U33000 ( .B1(n3676), .B2(n3890), .A(n3680), .ZN(n2555) );
  NAND2_X1 U33010 ( .A1(n2557), .A2(n3553), .ZN(n3865) );
  OR2_X1 U33020 ( .A1(n3895), .A2(n3876), .ZN(n3584) );
  OR2_X1 U33030 ( .A1(n3869), .A2(n3901), .ZN(n3864) );
  NAND2_X1 U33040 ( .A1(n3865), .A2(n3681), .ZN(n2558) );
  NAND2_X1 U33050 ( .A1(n3895), .A2(n3876), .ZN(n3583) );
  NAND2_X1 U33060 ( .A1(n2558), .A2(n3583), .ZN(n3849) );
  NAND2_X1 U33070 ( .A1(n3870), .A2(n3857), .ZN(n3604) );
  INV_X1 U33080 ( .A(n3604), .ZN(n2559) );
  OR2_X1 U33100 ( .A1(n3870), .A2(n3857), .ZN(n3830) );
  OR2_X1 U33110 ( .A1(n3852), .A2(n3841), .ZN(n2560) );
  NAND2_X1 U33120 ( .A1(n3830), .A2(n2560), .ZN(n3685) );
  INV_X1 U33130 ( .A(n3685), .ZN(n2561) );
  AND2_X1 U33140 ( .A1(n3852), .A2(n3841), .ZN(n3564) );
  AOI21_X2 U33150 ( .B1(n3831), .B2(n2561), .A(n3564), .ZN(n3819) );
  OR2_X1 U33160 ( .A1(n3836), .A2(n3823), .ZN(n2562) );
  NAND2_X1 U33170 ( .A1(n3836), .A2(n3823), .ZN(n3683) );
  NAND2_X1 U33180 ( .A1(n2562), .A2(n3683), .ZN(n3810) );
  INV_X1 U33190 ( .A(n2562), .ZN(n3559) );
  AOI21_X1 U33200 ( .B1(n3819), .B2(n3818), .A(n3559), .ZN(n3787) );
  XNOR2_X1 U33210 ( .A(n3787), .B(n3797), .ZN(n2576) );
  NAND2_X1 U33220 ( .A1(n3701), .A2(n3769), .ZN(n2564) );
  INV_X1 U33230 ( .A(n3694), .ZN(n4330) );
  NAND2_X1 U33240 ( .A1(n3625), .A2(n4330), .ZN(n2563) );
  INV_X1 U33250 ( .A(n3701), .ZN(n2565) );
  OR2_X1 U33260 ( .A1(n2566), .A2(n2640), .ZN(n2568) );
  XNOR2_X1 U33270 ( .A(n2568), .B(n2567), .ZN(n4335) );
  INV_X1 U33280 ( .A(n4335), .ZN(n2735) );
  NAND2_X1 U33290 ( .A1(n3836), .A2(n4024), .ZN(n2574) );
  NAND2_X1 U33300 ( .A1(n2497), .A2(REG2_REG_29__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U33310 ( .A1(n3538), .A2(REG1_REG_29__SCAN_IN), .ZN(n2571) );
  NAND2_X1 U33320 ( .A1(n2265), .A2(n3795), .ZN(n2570) );
  NAND2_X1 U33330 ( .A1(n2258), .A2(REG0_REG_29__SCAN_IN), .ZN(n2569) );
  NAND4_X1 U33340 ( .A1(n2572), .A2(n2571), .A3(n2570), .A4(n2569), .ZN(n3705)
         );
  NAND2_X1 U33350 ( .A1(n2728), .A2(n4335), .ZN(n3946) );
  NAND2_X1 U33360 ( .A1(n3705), .A2(n4272), .ZN(n2573) );
  OAI211_X1 U33370 ( .C1(n4029), .C2(n3364), .A(n2574), .B(n2573), .ZN(n2575)
         );
  AOI21_X1 U33380 ( .B1(n2576), .B2(n4040), .A(n2575), .ZN(n3370) );
  OAI21_X1 U33390 ( .B1(n3377), .B2(n4540), .A(n3370), .ZN(n2619) );
  NOR2_X1 U33400 ( .A1(n2015), .A2(n2640), .ZN(n2577) );
  MUX2_X1 U33410 ( .A(n2640), .B(n2577), .S(IR_REG_25__SCAN_IN), .Z(n2578) );
  INV_X1 U33420 ( .A(n2578), .ZN(n2580) );
  NAND2_X1 U33430 ( .A1(n2580), .A2(n2579), .ZN(n2591) );
  NAND2_X1 U33440 ( .A1(n2591), .A2(B_REG_SCAN_IN), .ZN(n2584) );
  OR2_X1 U33450 ( .A1(n2640), .A2(n2595), .ZN(n2582) );
  MUX2_X1 U33460 ( .A(n2584), .B(B_REG_SCAN_IN), .S(n4329), .Z(n2587) );
  OR2_X1 U33470 ( .A1(n2585), .A2(n2640), .ZN(n2586) );
  INV_X1 U33480 ( .A(D_REG_0__SCAN_IN), .ZN(n4132) );
  INV_X1 U33490 ( .A(n4329), .ZN(n2588) );
  INV_X1 U33500 ( .A(n2630), .ZN(n2589) );
  INV_X1 U33510 ( .A(n2930), .ZN(n2610) );
  NAND2_X1 U33520 ( .A1(n2589), .A2(n2591), .ZN(n2721) );
  OAI21_X1 U3353 ( .B1(n2723), .B2(D_REG_1__SCAN_IN), .A(n2721), .ZN(n2609) );
  NAND2_X1 U33540 ( .A1(n3694), .A2(n3780), .ZN(n2590) );
  AND2_X1 U3355 ( .A1(n2728), .A2(n2590), .ZN(n2804) );
  INV_X1 U3356 ( .A(n2591), .ZN(n4328) );
  NOR2_X1 U3357 ( .A1(n4549), .A2(n3625), .ZN(n2736) );
  NOR2_X1 U3358 ( .A1(n2928), .A2(n2736), .ZN(n2608) );
  NOR4_X1 U3359 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2599) );
  NOR4_X1 U3360 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2598) );
  NOR4_X1 U3361 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2597) );
  NOR4_X1 U3362 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2596) );
  AND4_X1 U3363 ( .A1(n2599), .A2(n2598), .A3(n2597), .A4(n2596), .ZN(n2605)
         );
  NOR2_X1 U3364 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_4__SCAN_IN), .ZN(n2603) );
  NOR4_X1 U3365 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2602) );
  NOR4_X1 U3366 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2601) );
  NOR4_X1 U3367 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2600) );
  AND4_X1 U3368 ( .A1(n2603), .A2(n2602), .A3(n2601), .A4(n2600), .ZN(n2604)
         );
  NAND2_X1 U3369 ( .A1(n2605), .A2(n2604), .ZN(n2720) );
  NAND2_X1 U3370 ( .A1(n2606), .A2(n2720), .ZN(n2607) );
  MUX2_X1 U3371 ( .A(REG0_REG_28__SCAN_IN), .B(n2619), .S(n4555), .Z(n2611) );
  INV_X1 U3372 ( .A(n2611), .ZN(n2617) );
  NAND2_X1 U3373 ( .A1(n3023), .A2(n3601), .ZN(n3017) );
  INV_X1 U3374 ( .A(n2774), .ZN(n2793) );
  NAND2_X1 U3375 ( .A1(n2943), .A2(n2942), .ZN(n2957) );
  NOR2_X1 U3376 ( .A1(n3415), .A2(n3991), .ZN(n2612) );
  OAI21_X1 U3377 ( .B1(n3813), .B2(n3364), .A(n3802), .ZN(n3373) );
  NAND2_X1 U3378 ( .A1(n2617), .A2(n2616), .ZN(U3514) );
  MUX2_X1 U3379 ( .A(REG1_REG_28__SCAN_IN), .B(n2619), .S(n4567), .Z(n2620) );
  INV_X1 U3380 ( .A(n2620), .ZN(n2622) );
  NAND2_X1 U3381 ( .A1(n2622), .A2(n2621), .ZN(U3546) );
  INV_X2 U3382 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3383 ( .A(n4485), .ZN(n2623) );
  MUX2_X1 U3384 ( .A(n2624), .B(n2682), .S(STATE_REG_SCAN_IN), .Z(n2625) );
  INV_X1 U3385 ( .A(n2625), .ZN(U3348) );
  INV_X1 U3386 ( .A(DATAI_3_), .ZN(n2626) );
  MUX2_X1 U3387 ( .A(n2671), .B(n2626), .S(U3149), .Z(n2627) );
  INV_X1 U3388 ( .A(n2627), .ZN(U3349) );
  MUX2_X1 U3389 ( .A(n2888), .B(n4177), .S(U3149), .Z(n2628) );
  INV_X1 U3390 ( .A(n2628), .ZN(U3345) );
  INV_X1 U3391 ( .A(n3749), .ZN(n3774) );
  NAND2_X1 U3392 ( .A1(n3774), .A2(STATE_REG_SCAN_IN), .ZN(n2629) );
  OAI21_X1 U3393 ( .B1(STATE_REG_SCAN_IN), .B2(n2439), .A(n2629), .ZN(U3335)
         );
  INV_X1 U3394 ( .A(DATAI_26_), .ZN(n4173) );
  NAND2_X1 U3395 ( .A1(n2630), .A2(STATE_REG_SCAN_IN), .ZN(n2631) );
  OAI21_X1 U3396 ( .B1(STATE_REG_SCAN_IN), .B2(n4173), .A(n2631), .ZN(U3326)
         );
  MUX2_X1 U3397 ( .A(n2458), .B(n3780), .S(STATE_REG_SCAN_IN), .Z(n2632) );
  INV_X1 U3398 ( .A(n2632), .ZN(U3333) );
  INV_X1 U3399 ( .A(DATAI_21_), .ZN(n2634) );
  NAND2_X1 U3400 ( .A1(n3625), .A2(STATE_REG_SCAN_IN), .ZN(n2633) );
  OAI21_X1 U3401 ( .B1(STATE_REG_SCAN_IN), .B2(n2634), .A(n2633), .ZN(U3331)
         );
  INV_X1 U3402 ( .A(DATAI_29_), .ZN(n2637) );
  NAND2_X1 U3403 ( .A1(n2635), .A2(STATE_REG_SCAN_IN), .ZN(n2636) );
  OAI21_X1 U3404 ( .B1(STATE_REG_SCAN_IN), .B2(n2637), .A(n2636), .ZN(U3323)
         );
  INV_X1 U3405 ( .A(DATAI_22_), .ZN(n2639) );
  NAND2_X1 U3406 ( .A1(n3701), .A2(STATE_REG_SCAN_IN), .ZN(n2638) );
  OAI21_X1 U3407 ( .B1(STATE_REG_SCAN_IN), .B2(n2639), .A(n2638), .ZN(U3330)
         );
  INV_X1 U3408 ( .A(DATAI_31_), .ZN(n2643) );
  OR4_X1 U3409 ( .A1(n2641), .A2(IR_REG_30__SCAN_IN), .A3(n2640), .A4(U3149), 
        .ZN(n2642) );
  OAI21_X1 U3410 ( .B1(STATE_REG_SCAN_IN), .B2(n2643), .A(n2642), .ZN(U3321)
         );
  INV_X1 U3411 ( .A(n2740), .ZN(n2644) );
  AOI22_X1 U3412 ( .A1(n4484), .A2(n4132), .B1(n2645), .B2(n4485), .ZN(U3458)
         );
  INV_X1 U3413 ( .A(D_REG_1__SCAN_IN), .ZN(n2719) );
  INV_X1 U3414 ( .A(n2721), .ZN(n2646) );
  AOI22_X1 U3415 ( .A1(n4484), .A2(n2719), .B1(n2646), .B2(n4485), .ZN(U3459)
         );
  OR2_X1 U3416 ( .A1(n2806), .A2(U3149), .ZN(n3703) );
  NAND2_X1 U3417 ( .A1(n2740), .A2(n3703), .ZN(n2650) );
  AOI21_X1 U3418 ( .B1(n2728), .B2(n2806), .A(n2647), .ZN(n2649) );
  INV_X1 U3419 ( .A(n2649), .ZN(n2648) );
  INV_X1 U3420 ( .A(n4427), .ZN(n4451) );
  INV_X1 U3421 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n2660) );
  XNOR2_X1 U3422 ( .A(n2651), .B(IR_REG_27__SCAN_IN), .ZN(n4327) );
  INV_X1 U3423 ( .A(n4327), .ZN(n2665) );
  INV_X1 U3424 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2745) );
  NAND3_X1 U3425 ( .A1(n4435), .A2(IR_REG_0__SCAN_IN), .A3(n2745), .ZN(n2659)
         );
  INV_X1 U3426 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2652) );
  AND2_X1 U3427 ( .A1(n4327), .A2(n2652), .ZN(n2653) );
  NOR2_X1 U3428 ( .A1(n4335), .A2(n2653), .ZN(n2816) );
  OAI21_X1 U3429 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4327), .A(n2816), .ZN(n2655)
         );
  INV_X1 U3430 ( .A(IR_REG_0__SCAN_IN), .ZN(n2654) );
  MUX2_X1 U3431 ( .A(n2816), .B(n2655), .S(n2654), .Z(n2656) );
  INV_X1 U3432 ( .A(n2656), .ZN(n2657) );
  AOI22_X1 U3433 ( .A1(n2666), .A2(n2657), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2658) );
  OAI211_X1 U3434 ( .C1(n4451), .C2(n2660), .A(n2659), .B(n2658), .ZN(U3240)
         );
  NOR2_X1 U3435 ( .A1(n4427), .A2(U4043), .ZN(U3148) );
  INV_X1 U3436 ( .A(n4450), .ZN(n4440) );
  AND2_X1 U3437 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3723)
         );
  NAND2_X1 U3438 ( .A1(n3722), .A2(n3723), .ZN(n3721) );
  INV_X1 U3439 ( .A(n2668), .ZN(n4333) );
  NAND2_X1 U3440 ( .A1(n4333), .A2(REG1_REG_1__SCAN_IN), .ZN(n2826) );
  NAND2_X1 U3441 ( .A1(n3721), .A2(n2826), .ZN(n2663) );
  INV_X1 U3442 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2661) );
  MUX2_X1 U3443 ( .A(n2661), .B(REG1_REG_2__SCAN_IN), .S(n2824), .Z(n2662) );
  INV_X1 U3444 ( .A(n2824), .ZN(n4332) );
  NAND2_X1 U3445 ( .A1(n4332), .A2(REG1_REG_2__SCAN_IN), .ZN(n2664) );
  XOR2_X1 U3446 ( .A(n2687), .B(REG1_REG_3__SCAN_IN), .Z(n2673) );
  NOR2_X1 U3447 ( .A1(n4335), .A2(n2665), .ZN(n3698) );
  INV_X1 U3448 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2667) );
  MUX2_X1 U3449 ( .A(n2667), .B(REG2_REG_2__SCAN_IN), .S(n2824), .Z(n2823) );
  XNOR2_X1 U3450 ( .A(n2668), .B(REG2_REG_1__SCAN_IN), .ZN(n3726) );
  AND2_X1 U3451 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2669)
         );
  NAND2_X1 U3452 ( .A1(n3726), .A2(n2669), .ZN(n3725) );
  NAND2_X1 U3453 ( .A1(n4333), .A2(REG2_REG_1__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U3454 ( .A1(n3725), .A2(n2670), .ZN(n2822) );
  OAI21_X1 U3455 ( .B1(n2667), .B2(n2824), .A(n2821), .ZN(n2680) );
  XNOR2_X1 U3456 ( .A(n2681), .B(n4122), .ZN(n2672) );
  AOI22_X1 U3457 ( .A1(n4435), .A2(n2673), .B1(n4437), .B2(n2672), .ZN(n2675)
         );
  AOI22_X1 U34580 ( .A1(n4427), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2674) );
  OAI211_X1 U34590 ( .C1(n2671), .C2(n4440), .A(n2675), .B(n2674), .ZN(U3243)
         );
  INV_X1 U3460 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4144) );
  NAND2_X1 U3461 ( .A1(U4043), .A2(n3983), .ZN(n2676) );
  OAI21_X1 U3462 ( .B1(U4043), .B2(n4144), .A(n2676), .ZN(U3569) );
  INV_X1 U3463 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4145) );
  NAND2_X1 U3464 ( .A1(U4043), .A2(n3191), .ZN(n2677) );
  OAI21_X1 U3465 ( .B1(U4043), .B2(n4145), .A(n2677), .ZN(U3560) );
  INV_X1 U3466 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4142) );
  NAND2_X1 U34670 ( .A1(U4043), .A2(n3926), .ZN(n2678) );
  OAI21_X1 U3468 ( .B1(U4043), .B2(n4142), .A(n2678), .ZN(U3572) );
  INV_X1 U34690 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4203) );
  NAND2_X1 U3470 ( .A1(U4043), .A2(n4273), .ZN(n2679) );
  OAI21_X1 U34710 ( .B1(U4043), .B2(n4203), .A(n2679), .ZN(U3551) );
  INV_X1 U3472 ( .A(n2682), .ZN(n2856) );
  INV_X1 U34730 ( .A(n2683), .ZN(n2684) );
  INV_X1 U3474 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4232) );
  MUX2_X1 U34750 ( .A(REG2_REG_5__SCAN_IN), .B(n4232), .S(n2707), .Z(n2685) );
  INV_X1 U3476 ( .A(n4437), .ZN(n4445) );
  AOI211_X1 U34770 ( .C1(n2686), .C2(n2685), .A(n2708), .B(n4445), .ZN(n2699)
         );
  NAND2_X1 U3478 ( .A1(n2689), .A2(n2688), .ZN(n2690) );
  NAND2_X1 U34790 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  XNOR2_X1 U3480 ( .A(n2692), .B(n2856), .ZN(n2854) );
  NAND2_X1 U34810 ( .A1(n2692), .A2(n2856), .ZN(n2693) );
  MUX2_X1 U3482 ( .A(REG1_REG_5__SCAN_IN), .B(n2701), .S(n2707), .Z(n2694) );
  AOI211_X1 U34830 ( .C1(n2695), .C2(n2694), .A(n2047), .B(n4441), .ZN(n2698)
         );
  AND2_X1 U3484 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2879) );
  AOI21_X1 U34850 ( .B1(n4427), .B2(ADDR_REG_5__SCAN_IN), .A(n2879), .ZN(n2696) );
  OAI21_X1 U3486 ( .B1(n4440), .B2(n2707), .A(n2696), .ZN(n2697) );
  OR3_X1 U34870 ( .A1(n2699), .A2(n2698), .A3(n2697), .ZN(U3245) );
  INV_X1 U3488 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2700) );
  MUX2_X1 U34890 ( .A(n2700), .B(REG1_REG_7__SCAN_IN), .S(n2888), .Z(n2706) );
  INV_X1 U3490 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U34910 ( .A1(n2709), .A2(n2703), .ZN(n2704) );
  OAI21_X1 U3492 ( .B1(n2706), .B2(n2882), .A(n4435), .ZN(n2705) );
  AOI21_X1 U34930 ( .B1(n2706), .B2(n2882), .A(n2705), .ZN(n2717) );
  OR2_X1 U3494 ( .A1(n2710), .A2(n4505), .ZN(n2711) );
  XNOR2_X1 U34950 ( .A(n2710), .B(n2709), .ZN(n4343) );
  NAND2_X1 U3496 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4343), .ZN(n4342) );
  INV_X1 U34970 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2990) );
  MUX2_X1 U3498 ( .A(REG2_REG_7__SCAN_IN), .B(n2990), .S(n2888), .Z(n2712) );
  AOI211_X1 U34990 ( .C1(n2713), .C2(n2712), .A(n4445), .B(n2887), .ZN(n2716)
         );
  INV_X1 U3500 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4180) );
  NOR2_X1 U35010 ( .A1(STATE_REG_SCAN_IN), .A2(n4180), .ZN(n2920) );
  AOI21_X1 U3502 ( .B1(n4427), .B2(ADDR_REG_7__SCAN_IN), .A(n2920), .ZN(n2714)
         );
  OAI21_X1 U35030 ( .B1(n4440), .B2(n2888), .A(n2714), .ZN(n2715) );
  OR3_X1 U3504 ( .A1(n2717), .A2(n2716), .A3(n2715), .ZN(U3247) );
  INV_X1 U35050 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4141) );
  NAND2_X1 U35060 ( .A1(U4043), .A2(n3870), .ZN(n2718) );
  OAI21_X1 U35070 ( .B1(U4043), .B2(n4141), .A(n2718), .ZN(U3575) );
  NOR2_X1 U35080 ( .A1(n2720), .A2(n2719), .ZN(n2722) );
  OAI21_X1 U35090 ( .B1(n2723), .B2(n2722), .A(n2721), .ZN(n2929) );
  INV_X1 U35100 ( .A(n2929), .ZN(n2724) );
  NAND2_X1 U35110 ( .A1(n2724), .A2(n2930), .ZN(n2741) );
  INV_X1 U35120 ( .A(n2725), .ZN(n2932) );
  INV_X4 U35130 ( .A(n2779), .ZN(n3352) );
  NAND2_X1 U35140 ( .A1(n3701), .A2(n3780), .ZN(n2772) );
  INV_X1 U35150 ( .A(n2772), .ZN(n2726) );
  NAND2_X1 U35160 ( .A1(n4485), .A2(n2726), .ZN(n2727) );
  INV_X1 U35170 ( .A(n2734), .ZN(n3699) );
  AND2_X1 U35180 ( .A1(n2741), .A2(n3699), .ZN(n2810) );
  INV_X1 U35190 ( .A(n2810), .ZN(n2733) );
  INV_X1 U35200 ( .A(n2928), .ZN(n2732) );
  INV_X1 U35210 ( .A(n2728), .ZN(n2730) );
  NAND2_X1 U35220 ( .A1(n4276), .A2(n3769), .ZN(n2729) );
  NAND3_X1 U35230 ( .A1(n4029), .A2(n2730), .A3(n2729), .ZN(n2739) );
  NAND2_X1 U35240 ( .A1(n2739), .A2(n4029), .ZN(n2731) );
  NAND2_X1 U35250 ( .A1(n2741), .A2(n2731), .ZN(n2809) );
  NAND3_X1 U35260 ( .A1(n2733), .A2(n2732), .A3(n2809), .ZN(n3420) );
  INV_X1 U35270 ( .A(n3420), .ZN(n2753) );
  INV_X1 U35280 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4475) );
  OR2_X1 U35290 ( .A1(n2741), .A2(n2734), .ZN(n2792) );
  OR2_X2 U35300 ( .A1(n2792), .A2(n2735), .ZN(n3529) );
  INV_X1 U35310 ( .A(n3529), .ZN(n3498) );
  OR3_X1 U35320 ( .A1(n2741), .A2(n4029), .A3(n2740), .ZN(n2738) );
  INV_X1 U35330 ( .A(n2736), .ZN(n2737) );
  AND2_X4 U35340 ( .A1(n2805), .A2(n2725), .ZN(n3357) );
  NAND2_X2 U35350 ( .A1(n3357), .A2(n4548), .ZN(n3338) );
  NAND2_X1 U35360 ( .A1(n3356), .A2(n3720), .ZN(n2744) );
  INV_X1 U35370 ( .A(n2805), .ZN(n2742) );
  AOI22_X1 U35380 ( .A1(n2779), .A2(n4277), .B1(n2742), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2743) );
  NAND2_X1 U35390 ( .A1(n2744), .A2(n2743), .ZN(n2750) );
  NAND2_X1 U35400 ( .A1(n3720), .A2(n2779), .ZN(n2748) );
  NAND2_X1 U35410 ( .A1(n3357), .A2(n4277), .ZN(n2775) );
  OR2_X1 U35420 ( .A1(n2805), .A2(n2745), .ZN(n2746) );
  AND2_X1 U35430 ( .A1(n2775), .A2(n2746), .ZN(n2747) );
  NAND2_X1 U35440 ( .A1(n2748), .A2(n2747), .ZN(n2749) );
  NAND2_X1 U35450 ( .A1(n2750), .A2(n2749), .ZN(n2778) );
  OAI21_X1 U35460 ( .B1(n2750), .B2(n2749), .A(n2778), .ZN(n2820) );
  OAI22_X1 U35470 ( .A1(n3517), .A2(n3601), .B1(n3536), .B2(n2820), .ZN(n2751)
         );
  AOI21_X1 U35480 ( .B1(n3498), .B2(n4273), .A(n2751), .ZN(n2752) );
  OAI21_X1 U35490 ( .B1(n2753), .B2(n4475), .A(n2752), .ZN(U3229) );
  INV_X1 U35500 ( .A(n4549), .ZN(n4524) );
  OR2_X1 U35510 ( .A1(n2754), .A2(n3598), .ZN(n2755) );
  NAND2_X1 U35520 ( .A1(n2756), .A2(n2755), .ZN(n2966) );
  NAND3_X1 U35530 ( .A1(n3019), .A2(n3598), .A3(n2534), .ZN(n2757) );
  NAND2_X1 U35540 ( .A1(n2758), .A2(n2757), .ZN(n2759) );
  NAND2_X1 U35550 ( .A1(n2759), .A2(n4040), .ZN(n2766) );
  INV_X1 U35560 ( .A(n4270), .ZN(n2760) );
  NAND2_X1 U35570 ( .A1(n2966), .A2(n2760), .ZN(n2765) );
  NAND2_X1 U35580 ( .A1(n4273), .A2(n4024), .ZN(n2762) );
  NAND2_X1 U35590 ( .A1(n3718), .A2(n4272), .ZN(n2761) );
  OAI211_X1 U35600 ( .C1(n4029), .C2(n2774), .A(n2762), .B(n2761), .ZN(n2763)
         );
  INV_X1 U35610 ( .A(n2763), .ZN(n2764) );
  NAND3_X1 U35620 ( .A1(n2766), .A2(n2765), .A3(n2764), .ZN(n2964) );
  AOI21_X1 U35630 ( .B1(n4524), .B2(n2966), .A(n2964), .ZN(n2868) );
  AND2_X1 U35640 ( .A1(n3017), .A2(n2793), .ZN(n2767) );
  OR2_X1 U35650 ( .A1(n2767), .A2(n2943), .ZN(n2969) );
  OAI22_X1 U35660 ( .A1(n4268), .A2(n2969), .B1(n4567), .B2(n2661), .ZN(n2768)
         );
  INV_X1 U35670 ( .A(n2768), .ZN(n2769) );
  OAI21_X1 U35680 ( .B1(n2868), .B2(n4564), .A(n2769), .ZN(U3520) );
  NAND2_X1 U35690 ( .A1(n2273), .A2(n2779), .ZN(n2771) );
  NAND2_X1 U35700 ( .A1(n3357), .A2(n2793), .ZN(n2770) );
  NAND2_X1 U35710 ( .A1(n2771), .A2(n2770), .ZN(n2773) );
  AND2_X2 U35720 ( .A1(n2772), .A2(n2725), .ZN(n3324) );
  XNOR2_X1 U35730 ( .A(n2773), .B(n3358), .ZN(n2798) );
  OAI22_X1 U35740 ( .A1(n2938), .A2(n3338), .B1(n2774), .B2(n3352), .ZN(n2797)
         );
  XNOR2_X1 U35750 ( .A(n2798), .B(n2797), .ZN(n2791) );
  INV_X1 U35760 ( .A(n2775), .ZN(n2776) );
  OR2_X1 U35770 ( .A1(n2776), .A2(n3358), .ZN(n2777) );
  NAND2_X1 U35780 ( .A1(n2778), .A2(n2777), .ZN(n3422) );
  NAND2_X1 U35790 ( .A1(n4273), .A2(n2779), .ZN(n2781) );
  NAND2_X1 U35800 ( .A1(n3357), .A2(n3419), .ZN(n2780) );
  OAI22_X1 U35810 ( .A1(n2257), .A2(n3338), .B1(n2005), .B2(n3023), .ZN(n2784)
         );
  XNOR2_X1 U3582 ( .A(n2783), .B(n2784), .ZN(n3423) );
  NAND2_X1 U3583 ( .A1(n3422), .A2(n3423), .ZN(n3421) );
  INV_X1 U3584 ( .A(n2783), .ZN(n2785) );
  NAND2_X1 U3585 ( .A1(n2785), .A2(n2784), .ZN(n2786) );
  NAND2_X1 U3586 ( .A1(n3421), .A2(n2786), .ZN(n2790) );
  INV_X1 U3587 ( .A(n2790), .ZN(n2788) );
  NAND2_X1 U3588 ( .A1(n2788), .A2(n2787), .ZN(n2800) );
  INV_X1 U3589 ( .A(n2800), .ZN(n2789) );
  AOI21_X1 U3590 ( .B1(n2791), .B2(n2790), .A(n2789), .ZN(n2796) );
  OR2_X2 U3591 ( .A1(n2792), .A2(n4335), .ZN(n3530) );
  INV_X1 U3592 ( .A(n3530), .ZN(n3497) );
  AOI22_X1 U3593 ( .A1(n2793), .A2(n3532), .B1(n3497), .B2(n4273), .ZN(n2795)
         );
  AOI22_X1 U3594 ( .A1(n3420), .A2(REG3_REG_2__SCAN_IN), .B1(n3498), .B2(n3718), .ZN(n2794) );
  OAI211_X1 U3595 ( .C1(n2796), .C2(n3536), .A(n2795), .B(n2794), .ZN(U3234)
         );
  OR2_X1 U3596 ( .A1(n2798), .A2(n2797), .ZN(n2799) );
  NAND2_X1 U3597 ( .A1(n2800), .A2(n2799), .ZN(n2836) );
  NAND2_X1 U3598 ( .A1(n3718), .A2(n2779), .ZN(n2802) );
  NAND2_X1 U3599 ( .A1(n3357), .A2(n2936), .ZN(n2801) );
  NAND2_X1 U3600 ( .A1(n2802), .A2(n2801), .ZN(n2803) );
  XNOR2_X1 U3601 ( .A(n2803), .B(n3324), .ZN(n2837) );
  OAI22_X1 U3602 ( .A1(n2848), .A2(n3353), .B1(n3352), .B2(n2942), .ZN(n2838)
         );
  XNOR2_X1 U3603 ( .A(n2837), .B(n2838), .ZN(n2835) );
  XOR2_X1 U3604 ( .A(n2836), .B(n2835), .Z(n2815) );
  OAI22_X1 U3605 ( .A1(n3517), .A2(n2942), .B1(n3530), .B2(n2938), .ZN(n2813)
         );
  INV_X1 U3606 ( .A(n2804), .ZN(n2807) );
  AND3_X1 U3607 ( .A1(n2807), .A2(n2806), .A3(n2805), .ZN(n2808) );
  AOI21_X1 U3608 ( .B1(n2809), .B2(n2808), .A(U3149), .ZN(n2811) );
  MUX2_X1 U3609 ( .A(n3533), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2812) );
  AOI211_X1 U3610 ( .C1(n3498), .C2(n3717), .A(n2813), .B(n2812), .ZN(n2814)
         );
  OAI21_X1 U3611 ( .B1(n3536), .B2(n2815), .A(n2814), .ZN(U3215) );
  NOR2_X1 U3612 ( .A1(n4335), .A2(n4327), .ZN(n2819) );
  INV_X1 U3613 ( .A(n3698), .ZN(n2817) );
  NAND2_X1 U3614 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3724) );
  OAI22_X1 U3615 ( .A1(n2817), .A2(n3724), .B1(n2816), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2818) );
  AOI211_X1 U3616 ( .C1(n2820), .C2(n2819), .A(n3719), .B(n2818), .ZN(n2861)
         );
  OAI211_X1 U3617 ( .C1(n2823), .C2(n2822), .A(n4437), .B(n2821), .ZN(n2832)
         );
  MUX2_X1 U3618 ( .A(REG1_REG_2__SCAN_IN), .B(n2661), .S(n2824), .Z(n2825) );
  NAND3_X1 U3619 ( .A1(n3721), .A2(n2826), .A3(n2825), .ZN(n2827) );
  NAND3_X1 U3620 ( .A1(n4435), .A2(n2828), .A3(n2827), .ZN(n2831) );
  NAND2_X1 U3621 ( .A1(n4450), .A2(n4332), .ZN(n2830) );
  AOI22_X1 U3622 ( .A1(n4427), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2829) );
  NAND4_X1 U3623 ( .A1(n2832), .A2(n2831), .A3(n2830), .A4(n2829), .ZN(n2833)
         );
  OR2_X1 U3624 ( .A1(n2861), .A2(n2833), .ZN(U3242) );
  INV_X1 U3625 ( .A(n2834), .ZN(n2960) );
  INV_X1 U3626 ( .A(n2837), .ZN(n2839) );
  OR2_X1 U3627 ( .A1(n2839), .A2(n2838), .ZN(n2840) );
  NAND2_X1 U3628 ( .A1(n3717), .A2(n2779), .ZN(n2842) );
  NAND2_X1 U3629 ( .A1(n3357), .A2(n2850), .ZN(n2841) );
  NAND2_X1 U3630 ( .A1(n2842), .A2(n2841), .ZN(n2843) );
  XNOR2_X1 U3631 ( .A(n2843), .B(n3358), .ZN(n2871) );
  INV_X1 U3632 ( .A(n3717), .ZN(n2973) );
  OAI22_X1 U3633 ( .A1(n2973), .A2(n3353), .B1(n3352), .B2(n2958), .ZN(n2870)
         );
  XNOR2_X1 U3634 ( .A(n2871), .B(n2870), .ZN(n2845) );
  AOI21_X1 U3635 ( .B1(n2844), .B2(n2845), .A(n3536), .ZN(n2847) );
  NAND2_X1 U3636 ( .A1(n2847), .A2(n2873), .ZN(n2852) );
  AND2_X1 U3637 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n2857) );
  OAI22_X1 U3638 ( .A1(n3048), .A2(n3529), .B1(n3530), .B2(n2848), .ZN(n2849)
         );
  AOI211_X1 U3639 ( .C1(n2850), .C2(n3532), .A(n2857), .B(n2849), .ZN(n2851)
         );
  OAI211_X1 U3640 ( .C1(n3114), .C2(n2960), .A(n2852), .B(n2851), .ZN(U3227)
         );
  XNOR2_X1 U3641 ( .A(n2853), .B(REG2_REG_4__SCAN_IN), .ZN(n2863) );
  XNOR2_X1 U3642 ( .A(n2854), .B(REG1_REG_4__SCAN_IN), .ZN(n2855) );
  NAND2_X1 U3643 ( .A1(n4435), .A2(n2855), .ZN(n2860) );
  NAND2_X1 U3644 ( .A1(n4450), .A2(n2856), .ZN(n2859) );
  AOI21_X1 U3645 ( .B1(n4427), .B2(ADDR_REG_4__SCAN_IN), .A(n2857), .ZN(n2858)
         );
  NAND3_X1 U3646 ( .A1(n2860), .A2(n2859), .A3(n2858), .ZN(n2862) );
  AOI211_X1 U3647 ( .C1(n4437), .C2(n2863), .A(n2862), .B(n2861), .ZN(n2864)
         );
  INV_X1 U3648 ( .A(n2864), .ZN(U3244) );
  INV_X1 U3649 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2865) );
  OAI22_X1 U3650 ( .A1(n4325), .A2(n2969), .B1(n4555), .B2(n2865), .ZN(n2866)
         );
  INV_X1 U3651 ( .A(n2866), .ZN(n2867) );
  OAI21_X1 U3652 ( .B1(n2868), .B2(n4553), .A(n2867), .ZN(U3471) );
  INV_X1 U3653 ( .A(n2869), .ZN(n2979) );
  NAND2_X1 U3654 ( .A1(n2871), .A2(n2870), .ZN(n2872) );
  NAND2_X1 U3655 ( .A1(n2873), .A2(n2872), .ZN(n2877) );
  OAI22_X1 U3656 ( .A1(n3048), .A2(n3352), .B1(n3348), .B2(n2875), .ZN(n2874)
         );
  XNOR2_X1 U3657 ( .A(n2874), .B(n3324), .ZN(n2898) );
  OAI22_X1 U3658 ( .A1(n3048), .A2(n3353), .B1(n3352), .B2(n2875), .ZN(n2899)
         );
  XNOR2_X1 U3659 ( .A(n2898), .B(n2899), .ZN(n2876) );
  INV_X1 U3660 ( .A(n3536), .ZN(n3495) );
  OAI211_X1 U3661 ( .C1(n2877), .C2(n2876), .A(n2902), .B(n3495), .ZN(n2881)
         );
  OAI22_X1 U3662 ( .A1(n2973), .A2(n3530), .B1(n3529), .B2(n2922), .ZN(n2878)
         );
  AOI211_X1 U3663 ( .C1(n2976), .C2(n3532), .A(n2879), .B(n2878), .ZN(n2880)
         );
  OAI211_X1 U3664 ( .C1(n3114), .C2(n2979), .A(n2881), .B(n2880), .ZN(U3224)
         );
  INV_X1 U3665 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4188) );
  INV_X1 U3666 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4354) );
  NOR2_X1 U3667 ( .A1(n4362), .A2(n2883), .ZN(n2884) );
  INV_X1 U3668 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U3669 ( .A1(REG1_REG_9__SCAN_IN), .A2(n4501), .B1(n2886), .B2(n4562), .ZN(n4364) );
  AOI211_X1 U3670 ( .C1(n4188), .C2(n2885), .A(n3751), .B(n4441), .ZN(n2897)
         );
  INV_X1 U3671 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2891) );
  AOI22_X1 U3672 ( .A1(REG2_REG_9__SCAN_IN), .A2(n2886), .B1(n4501), .B2(n2891), .ZN(n4369) );
  NAND2_X1 U3673 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4359), .ZN(n4358) );
  NAND2_X1 U3674 ( .A1(n4502), .A2(n2889), .ZN(n2890) );
  NAND2_X1 U3675 ( .A1(n4358), .A2(n2890), .ZN(n4368) );
  NAND2_X1 U3676 ( .A1(n4369), .A2(n4368), .ZN(n4367) );
  NAND2_X1 U3677 ( .A1(REG2_REG_10__SCAN_IN), .A2(n2893), .ZN(n3733) );
  OAI211_X1 U3678 ( .C1(n2893), .C2(REG2_REG_10__SCAN_IN), .A(n4437), .B(n3733), .ZN(n2895) );
  AND2_X1 U3679 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n3110) );
  AOI21_X1 U3680 ( .B1(n4427), .B2(ADDR_REG_10__SCAN_IN), .A(n3110), .ZN(n2894) );
  OAI211_X1 U3681 ( .C1(n4440), .C2(n2077), .A(n2895), .B(n2894), .ZN(n2896)
         );
  OR2_X1 U3682 ( .A1(n2897), .A2(n2896), .ZN(U3250) );
  INV_X1 U3683 ( .A(n2898), .ZN(n2900) );
  NAND2_X1 U3684 ( .A1(n2900), .A2(n2899), .ZN(n2901) );
  NAND2_X1 U3685 ( .A1(n3714), .A2(n2779), .ZN(n2904) );
  NAND2_X1 U3686 ( .A1(n3357), .A2(n2909), .ZN(n2903) );
  NAND2_X1 U3687 ( .A1(n2904), .A2(n2903), .ZN(n2905) );
  XNOR2_X1 U3688 ( .A(n2905), .B(n3358), .ZN(n2913) );
  OAI22_X1 U3689 ( .A1(n2922), .A2(n3353), .B1(n3352), .B2(n3055), .ZN(n2914)
         );
  XNOR2_X1 U3690 ( .A(n2913), .B(n2914), .ZN(n2906) );
  XNOR2_X1 U3691 ( .A(n2915), .B(n2906), .ZN(n2907) );
  NAND2_X1 U3692 ( .A1(n2907), .A2(n3495), .ZN(n2911) );
  AND2_X1 U3693 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n4347) );
  INV_X1 U3694 ( .A(n3713), .ZN(n3012) );
  OAI22_X1 U3695 ( .A1(n3048), .A2(n3530), .B1(n3529), .B2(n3012), .ZN(n2908)
         );
  AOI211_X1 U3696 ( .C1(n2909), .C2(n3532), .A(n4347), .B(n2908), .ZN(n2910)
         );
  OAI211_X1 U3697 ( .C1(n3114), .C2(n2912), .A(n2911), .B(n2910), .ZN(U3236)
         );
  NAND2_X1 U3698 ( .A1(n3713), .A2(n2779), .ZN(n2918) );
  NAND2_X1 U3699 ( .A1(n3357), .A2(n2916), .ZN(n2917) );
  NAND2_X1 U3700 ( .A1(n2918), .A2(n2917), .ZN(n2919) );
  XNOR2_X1 U3701 ( .A(n2919), .B(n3324), .ZN(n3000) );
  OAI22_X1 U3702 ( .A1(n3012), .A2(n3353), .B1(n3352), .B2(n2991), .ZN(n3001)
         );
  XNOR2_X1 U3703 ( .A(n3000), .B(n3001), .ZN(n2998) );
  XNOR2_X1 U3704 ( .A(n2999), .B(n2998), .ZN(n2926) );
  INV_X1 U3705 ( .A(n2920), .ZN(n2921) );
  OAI21_X1 U3706 ( .B1(n3517), .B2(n2991), .A(n2921), .ZN(n2924) );
  OAI22_X1 U3707 ( .A1(n3081), .A2(n3529), .B1(n3530), .B2(n2922), .ZN(n2923)
         );
  AOI211_X1 U3708 ( .C1(n2994), .C2(n3533), .A(n2924), .B(n2923), .ZN(n2925)
         );
  OAI21_X1 U3709 ( .B1(n2926), .B2(n3536), .A(n2925), .ZN(U3210) );
  XNOR2_X1 U3710 ( .A(n2927), .B(n2935), .ZN(n4516) );
  INV_X2 U3711 ( .A(n4470), .ZN(n4463) );
  NAND2_X1 U3712 ( .A1(n2932), .A2(n3769), .ZN(n2981) );
  INV_X1 U3713 ( .A(n4466), .ZN(n3028) );
  OAI21_X1 U3714 ( .B1(n2935), .B2(n2934), .A(n2933), .ZN(n2940) );
  INV_X1 U3715 ( .A(n4029), .ZN(n4064) );
  AOI22_X1 U3716 ( .A1(n3717), .A2(n4272), .B1(n4064), .B2(n2936), .ZN(n2937)
         );
  OAI21_X1 U3717 ( .B1(n2938), .B2(n4044), .A(n2937), .ZN(n2939) );
  AOI21_X1 U3718 ( .B1(n2940), .B2(n4040), .A(n2939), .ZN(n2941) );
  OAI21_X1 U3719 ( .B1(n4516), .B2(n4270), .A(n2941), .ZN(n4518) );
  NAND2_X1 U3720 ( .A1(n4518), .A2(n4470), .ZN(n2947) );
  NAND2_X1 U3721 ( .A1(n4470), .A2(n3780), .ZN(n3993) );
  NOR2_X1 U3722 ( .A1(n3993), .A2(n4548), .ZN(n4458) );
  OAI21_X1 U3723 ( .B1(n2943), .B2(n2942), .A(n2957), .ZN(n4515) );
  INV_X1 U3724 ( .A(n4515), .ZN(n2945) );
  OAI22_X1 U3725 ( .A1(n4470), .A2(n4122), .B1(REG3_REG_3__SCAN_IN), .B2(n4476), .ZN(n2944) );
  AOI21_X1 U3726 ( .B1(n4458), .B2(n2945), .A(n2944), .ZN(n2946) );
  OAI211_X1 U3727 ( .C1(n4516), .C2(n3028), .A(n2947), .B(n2946), .ZN(U3287)
         );
  INV_X1 U3728 ( .A(n2949), .ZN(n3589) );
  NAND2_X1 U3729 ( .A1(n2948), .A2(n3589), .ZN(n2950) );
  NAND2_X1 U3730 ( .A1(n2951), .A2(n2950), .ZN(n4520) );
  INV_X1 U3731 ( .A(n4040), .ZN(n4269) );
  XNOR2_X1 U3732 ( .A(n2952), .B(n2949), .ZN(n2956) );
  OAI22_X1 U3733 ( .A1(n3048), .A2(n3946), .B1(n2958), .B2(n4029), .ZN(n2954)
         );
  NOR2_X1 U3734 ( .A1(n4520), .A2(n4270), .ZN(n2953) );
  AOI211_X1 U3735 ( .C1(n4024), .C2(n3718), .A(n2954), .B(n2953), .ZN(n2955)
         );
  OAI21_X1 U3736 ( .B1(n4269), .B2(n2956), .A(n2955), .ZN(n4522) );
  INV_X1 U3737 ( .A(n2957), .ZN(n2959) );
  OAI211_X1 U3738 ( .C1(n2959), .C2(n2958), .A(n4545), .B(n2977), .ZN(n4521)
         );
  OAI22_X1 U3739 ( .A1(n4521), .A2(n3769), .B1(n4476), .B2(n2960), .ZN(n2961)
         );
  OAI21_X1 U3740 ( .B1(n4522), .B2(n2961), .A(n4470), .ZN(n2963) );
  NAND2_X1 U3741 ( .A1(n4463), .A2(REG2_REG_4__SCAN_IN), .ZN(n2962) );
  OAI211_X1 U3742 ( .C1(n4520), .C2(n3028), .A(n2963), .B(n2962), .ZN(U3286)
         );
  MUX2_X1 U3743 ( .A(n2964), .B(REG2_REG_2__SCAN_IN), .S(n4463), .Z(n2965) );
  INV_X1 U3744 ( .A(n2965), .ZN(n2968) );
  AOI22_X1 U3745 ( .A1(n4466), .A2(n2966), .B1(REG3_REG_2__SCAN_IN), .B2(n4453), .ZN(n2967) );
  OAI211_X1 U3746 ( .C1(n4050), .C2(n2969), .A(n2968), .B(n2967), .ZN(U3288)
         );
  INV_X1 U3747 ( .A(n2970), .ZN(n3635) );
  NAND2_X1 U3748 ( .A1(n3635), .A2(n3649), .ZN(n3575) );
  XNOR2_X1 U3749 ( .A(n2971), .B(n3575), .ZN(n2975) );
  AOI22_X1 U3750 ( .A1(n3714), .A2(n4272), .B1(n4064), .B2(n2976), .ZN(n2972)
         );
  OAI21_X1 U3751 ( .B1(n2973), .B2(n4044), .A(n2972), .ZN(n2974) );
  AOI21_X1 U3752 ( .B1(n2975), .B2(n4040), .A(n2974), .ZN(n4528) );
  AND2_X1 U3753 ( .A1(n2977), .A2(n2976), .ZN(n2978) );
  NOR2_X1 U3754 ( .A1(n3056), .A2(n2978), .ZN(n4531) );
  OAI22_X1 U3755 ( .A1(n4470), .A2(n4232), .B1(n2979), .B2(n4476), .ZN(n2984)
         );
  XNOR2_X1 U3756 ( .A(n2980), .B(n3575), .ZN(n4527) );
  NAND2_X1 U3757 ( .A1(n4270), .A2(n2981), .ZN(n2982) );
  NOR2_X1 U3758 ( .A1(n4527), .A2(n4054), .ZN(n2983) );
  AOI211_X1 U3759 ( .C1(n4531), .C2(n4458), .A(n2984), .B(n2983), .ZN(n2985)
         );
  OAI21_X1 U3760 ( .B1(n4463), .B2(n4528), .A(n2985), .ZN(U3285) );
  OAI22_X1 U3761 ( .A1(n3081), .A2(n3946), .B1(n2991), .B2(n4029), .ZN(n2989)
         );
  XNOR2_X1 U3762 ( .A(n2986), .B(n3638), .ZN(n2987) );
  NOR2_X1 U3763 ( .A1(n2987), .A2(n4269), .ZN(n2988) );
  AOI211_X1 U3764 ( .C1(n4024), .C2(n3714), .A(n2989), .B(n2988), .ZN(n4538)
         );
  NOR2_X1 U3765 ( .A1(n4470), .A2(n2990), .ZN(n2993) );
  OAI211_X1 U3766 ( .C1(n3058), .C2(n2991), .A(n4545), .B(n3039), .ZN(n4537)
         );
  NOR2_X1 U3767 ( .A1(n4537), .A2(n3993), .ZN(n2992) );
  AOI211_X1 U3768 ( .C1(n4453), .C2(n2994), .A(n2993), .B(n2992), .ZN(n2997)
         );
  OR2_X1 U3769 ( .A1(n2995), .A2(n3638), .ZN(n4535) );
  NAND2_X1 U3770 ( .A1(n2995), .A2(n3638), .ZN(n4534) );
  NAND3_X1 U3771 ( .A1(n4535), .A2(n3999), .A3(n4534), .ZN(n2996) );
  OAI211_X1 U3772 ( .C1(n4538), .C2(n4463), .A(n2997), .B(n2996), .ZN(U3283)
         );
  NAND2_X1 U3773 ( .A1(n2999), .A2(n2998), .ZN(n3004) );
  INV_X1 U3774 ( .A(n3000), .ZN(n3002) );
  NAND2_X1 U3775 ( .A1(n3002), .A2(n3001), .ZN(n3003) );
  NAND2_X1 U3776 ( .A1(n3004), .A2(n3003), .ZN(n3076) );
  OAI22_X1 U3777 ( .A1(n3081), .A2(n3352), .B1(n3348), .B2(n3032), .ZN(n3005)
         );
  XNOR2_X1 U3778 ( .A(n3005), .B(n3358), .ZN(n3009) );
  INV_X1 U3779 ( .A(n3009), .ZN(n3007) );
  OAI22_X1 U3780 ( .A1(n3081), .A2(n3353), .B1(n3352), .B2(n3032), .ZN(n3008)
         );
  INV_X1 U3781 ( .A(n3008), .ZN(n3006) );
  NAND2_X1 U3782 ( .A1(n3007), .A2(n3006), .ZN(n3074) );
  INV_X1 U3783 ( .A(n3074), .ZN(n3010) );
  AND2_X1 U3784 ( .A1(n3009), .A2(n3008), .ZN(n3075) );
  NOR2_X1 U3785 ( .A1(n3010), .A2(n3075), .ZN(n3011) );
  XNOR2_X1 U3786 ( .A(n3076), .B(n3011), .ZN(n3016) );
  NAND2_X1 U3787 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4355) );
  OAI21_X1 U3788 ( .B1(n3517), .B2(n3032), .A(n4355), .ZN(n3014) );
  INV_X1 U3789 ( .A(n3711), .ZN(n3119) );
  OAI22_X1 U3790 ( .A1(n3012), .A2(n3530), .B1(n3529), .B2(n3119), .ZN(n3013)
         );
  AOI211_X1 U3791 ( .C1(n3041), .C2(n3533), .A(n3014), .B(n3013), .ZN(n3015)
         );
  OAI21_X1 U3792 ( .B1(n3016), .B2(n3536), .A(n3015), .ZN(U3218) );
  OAI21_X1 U3793 ( .B1(n3601), .B2(n3023), .A(n3017), .ZN(n4510) );
  XNOR2_X1 U3794 ( .A(n2533), .B(n3018), .ZN(n4511) );
  OAI21_X1 U3795 ( .B1(n3020), .B2(n3626), .A(n3019), .ZN(n3025) );
  NAND2_X1 U3796 ( .A1(n3720), .A2(n4024), .ZN(n3022) );
  NAND2_X1 U3797 ( .A1(n2273), .A2(n4272), .ZN(n3021) );
  OAI211_X1 U3798 ( .C1(n4029), .C2(n3023), .A(n3022), .B(n3021), .ZN(n3024)
         );
  AOI21_X1 U3799 ( .B1(n3025), .B2(n4040), .A(n3024), .ZN(n3026) );
  OAI21_X1 U3800 ( .B1(n4511), .B2(n4270), .A(n3026), .ZN(n4513) );
  AOI22_X1 U3801 ( .A1(n4463), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4453), .ZN(n3027) );
  OAI21_X1 U3802 ( .B1(n3028), .B2(n4511), .A(n3027), .ZN(n3029) );
  AOI21_X1 U3803 ( .B1(n4470), .B2(n4513), .A(n3029), .ZN(n3030) );
  OAI21_X1 U3804 ( .B1(n4050), .B2(n4510), .A(n3030), .ZN(U3289) );
  NAND2_X1 U3805 ( .A1(n3643), .A2(n3652), .ZN(n3597) );
  XOR2_X1 U3806 ( .A(n3597), .B(n3031), .Z(n3035) );
  OAI22_X1 U3807 ( .A1(n3119), .A2(n3946), .B1(n4029), .B2(n3032), .ZN(n3033)
         );
  AOI21_X1 U3808 ( .B1(n4024), .B2(n3713), .A(n3033), .ZN(n3034) );
  OAI21_X1 U3809 ( .B1(n3035), .B2(n4269), .A(n3034), .ZN(n3066) );
  INV_X1 U3810 ( .A(n3066), .ZN(n3046) );
  NAND2_X1 U3811 ( .A1(n4534), .A2(n3036), .ZN(n3037) );
  XOR2_X1 U3812 ( .A(n3597), .B(n3037), .Z(n3067) );
  INV_X1 U3813 ( .A(n3090), .ZN(n3038) );
  AOI21_X1 U3814 ( .B1(n3040), .B2(n3039), .A(n3038), .ZN(n3071) );
  INV_X1 U3815 ( .A(n3071), .ZN(n3043) );
  AOI22_X1 U3816 ( .A1(n4463), .A2(REG2_REG_8__SCAN_IN), .B1(n3041), .B2(n4453), .ZN(n3042) );
  OAI21_X1 U3817 ( .B1(n3043), .B2(n4050), .A(n3042), .ZN(n3044) );
  AOI21_X1 U3818 ( .B1(n3067), .B2(n3999), .A(n3044), .ZN(n3045) );
  OAI21_X1 U3819 ( .B1(n3046), .B2(n4463), .A(n3045), .ZN(U3282) );
  NAND2_X1 U3820 ( .A1(n3639), .A2(n3651), .ZN(n3600) );
  XNOR2_X1 U3821 ( .A(n3047), .B(n3600), .ZN(n4455) );
  OAI22_X1 U3822 ( .A1(n3048), .A2(n4044), .B1(n3055), .B2(n4029), .ZN(n3052)
         );
  XNOR2_X1 U3823 ( .A(n3049), .B(n3600), .ZN(n3050) );
  NOR2_X1 U3824 ( .A1(n3050), .A2(n4269), .ZN(n3051) );
  AOI211_X1 U3825 ( .C1(n4272), .C2(n3713), .A(n3052), .B(n3051), .ZN(n3053)
         );
  OAI21_X1 U3826 ( .B1(n4270), .B2(n4455), .A(n3053), .ZN(n3054) );
  INV_X1 U3827 ( .A(n3054), .ZN(n4462) );
  OAI21_X1 U3828 ( .B1(n4549), .B2(n4455), .A(n4462), .ZN(n3064) );
  NOR2_X1 U3829 ( .A1(n3056), .A2(n3055), .ZN(n3057) );
  OR2_X1 U3830 ( .A1(n3058), .A2(n3057), .ZN(n4456) );
  INV_X1 U3831 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3059) );
  OAI22_X1 U3832 ( .A1(n4456), .A2(n4268), .B1(n4567), .B2(n3059), .ZN(n3060)
         );
  AOI21_X1 U3833 ( .B1(n3064), .B2(n4567), .A(n3060), .ZN(n3061) );
  INV_X1 U3834 ( .A(n3061), .ZN(U3524) );
  INV_X1 U3835 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3062) );
  OAI22_X1 U3836 ( .A1(n4456), .A2(n4325), .B1(n4555), .B2(n3062), .ZN(n3063)
         );
  AOI21_X1 U3837 ( .B1(n3064), .B2(n4555), .A(n3063), .ZN(n3065) );
  INV_X1 U3838 ( .A(n3065), .ZN(U3479) );
  AOI21_X1 U3839 ( .B1(n3067), .B2(n4533), .A(n3066), .ZN(n3073) );
  INV_X1 U3840 ( .A(n4325), .ZN(n3259) );
  INV_X1 U3841 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3068) );
  NOR2_X1 U3842 ( .A1(n4555), .A2(n3068), .ZN(n3069) );
  AOI21_X1 U3843 ( .B1(n3071), .B2(n3259), .A(n3069), .ZN(n3070) );
  OAI21_X1 U3844 ( .B1(n3073), .B2(n4553), .A(n3070), .ZN(U3483) );
  INV_X1 U3845 ( .A(n4268), .ZN(n3255) );
  AOI22_X1 U3846 ( .A1(n3071), .A2(n3255), .B1(n4564), .B2(REG1_REG_8__SCAN_IN), .ZN(n3072) );
  OAI21_X1 U3847 ( .B1(n3073), .B2(n4564), .A(n3072), .ZN(U3526) );
  OAI21_X2 U3848 ( .B1(n3076), .B2(n3075), .A(n3074), .ZN(n3097) );
  NAND2_X1 U3849 ( .A1(n3711), .A2(n2779), .ZN(n3078) );
  NAND2_X1 U3850 ( .A1(n3357), .A2(n3091), .ZN(n3077) );
  NAND2_X1 U3851 ( .A1(n3078), .A2(n3077), .ZN(n3079) );
  XNOR2_X1 U3852 ( .A(n3079), .B(n3324), .ZN(n3098) );
  OAI22_X1 U3853 ( .A1(n3119), .A2(n3353), .B1(n3352), .B2(n2081), .ZN(n3099)
         );
  XNOR2_X1 U3854 ( .A(n3098), .B(n3099), .ZN(n3096) );
  XNOR2_X1 U3855 ( .A(n3097), .B(n3096), .ZN(n3080) );
  NAND2_X1 U3856 ( .A1(n3080), .A2(n3495), .ZN(n3084) );
  NOR2_X1 U3857 ( .A1(STATE_REG_SCAN_IN), .A2(n4231), .ZN(n4365) );
  OAI22_X1 U3858 ( .A1(n3081), .A2(n3530), .B1(n3529), .B2(n3154), .ZN(n3082)
         );
  AOI211_X1 U3859 ( .C1(n3091), .C2(n3532), .A(n4365), .B(n3082), .ZN(n3083)
         );
  OAI211_X1 U3860 ( .C1(n3114), .C2(n3092), .A(n3084), .B(n3083), .ZN(U3228)
         );
  INV_X1 U3861 ( .A(n3646), .ZN(n3653) );
  NAND2_X1 U3862 ( .A1(n3653), .A2(n3644), .ZN(n3599) );
  XNOR2_X1 U3863 ( .A(n3085), .B(n3599), .ZN(n4541) );
  XOR2_X1 U3864 ( .A(n3599), .B(n3086), .Z(n3089) );
  OAI22_X1 U3865 ( .A1(n3154), .A2(n3946), .B1(n4029), .B2(n2081), .ZN(n3087)
         );
  AOI21_X1 U3866 ( .B1(n4024), .B2(n3712), .A(n3087), .ZN(n3088) );
  OAI21_X1 U3867 ( .B1(n3089), .B2(n4269), .A(n3088), .ZN(n4542) );
  NAND2_X1 U3868 ( .A1(n4542), .A2(n4470), .ZN(n3095) );
  AOI21_X1 U3869 ( .B1(n3091), .B2(n3090), .A(n3126), .ZN(n4544) );
  OAI22_X1 U3870 ( .A1(n4470), .A2(n2891), .B1(n3092), .B2(n4476), .ZN(n3093)
         );
  AOI21_X1 U3871 ( .B1(n4544), .B2(n4458), .A(n3093), .ZN(n3094) );
  OAI211_X1 U3872 ( .C1(n4541), .C2(n4054), .A(n3095), .B(n3094), .ZN(U3281)
         );
  INV_X1 U3873 ( .A(n3127), .ZN(n3113) );
  INV_X1 U3874 ( .A(n3098), .ZN(n3100) );
  OR2_X1 U3875 ( .A1(n3100), .A2(n3099), .ZN(n3101) );
  NAND2_X1 U3876 ( .A1(n3191), .A2(n2779), .ZN(n3103) );
  NAND2_X1 U3877 ( .A1(n3357), .A2(n3117), .ZN(n3102) );
  NAND2_X1 U3878 ( .A1(n3103), .A2(n3102), .ZN(n3104) );
  XNOR2_X1 U3879 ( .A(n3104), .B(n3358), .ZN(n3146) );
  OAI22_X1 U3880 ( .A1(n3154), .A2(n3353), .B1(n3352), .B2(n3125), .ZN(n3145)
         );
  XNOR2_X1 U3881 ( .A(n3146), .B(n3145), .ZN(n3106) );
  AOI21_X1 U3882 ( .B1(n3105), .B2(n3106), .A(n3536), .ZN(n3108) );
  NAND2_X1 U3883 ( .A1(n3108), .A2(n3148), .ZN(n3112) );
  OAI22_X1 U3884 ( .A1(n3119), .A2(n3530), .B1(n3529), .B2(n3173), .ZN(n3109)
         );
  AOI211_X1 U3885 ( .C1(n3117), .C2(n3532), .A(n3110), .B(n3109), .ZN(n3111)
         );
  OAI211_X1 U3886 ( .C1(n3114), .C2(n3113), .A(n3112), .B(n3111), .ZN(U3214)
         );
  NAND2_X1 U3887 ( .A1(n3655), .A2(n3661), .ZN(n3574) );
  XOR2_X1 U3888 ( .A(n3574), .B(n3115), .Z(n3123) );
  XOR2_X1 U3889 ( .A(n3574), .B(n3116), .Z(n3121) );
  AOI22_X1 U3890 ( .A1(n3710), .A2(n4272), .B1(n4064), .B2(n3117), .ZN(n3118)
         );
  OAI21_X1 U3891 ( .B1(n3119), .B2(n4044), .A(n3118), .ZN(n3120) );
  AOI21_X1 U3892 ( .B1(n3121), .B2(n4040), .A(n3120), .ZN(n3122) );
  OAI21_X1 U3893 ( .B1(n3123), .B2(n4270), .A(n3122), .ZN(n3179) );
  INV_X1 U3894 ( .A(n3179), .ZN(n3131) );
  INV_X1 U3895 ( .A(n3123), .ZN(n3180) );
  INV_X1 U3896 ( .A(n3196), .ZN(n3124) );
  OAI21_X1 U3897 ( .B1(n3126), .B2(n3125), .A(n3124), .ZN(n3185) );
  AOI22_X1 U3898 ( .A1(n4463), .A2(REG2_REG_10__SCAN_IN), .B1(n3127), .B2(
        n4453), .ZN(n3128) );
  OAI21_X1 U3899 ( .B1(n3185), .B2(n4050), .A(n3128), .ZN(n3129) );
  AOI21_X1 U3900 ( .B1(n3180), .B2(n4466), .A(n3129), .ZN(n3130) );
  OAI21_X1 U3901 ( .B1(n3131), .B2(n4463), .A(n3130), .ZN(U3280) );
  INV_X1 U3902 ( .A(n3220), .ZN(n3132) );
  OR2_X1 U3903 ( .A1(n3221), .A2(n3132), .ZN(n3576) );
  INV_X1 U3904 ( .A(n3576), .ZN(n3133) );
  XNOR2_X1 U3905 ( .A(n3222), .B(n3133), .ZN(n3137) );
  NAND2_X1 U3906 ( .A1(n3710), .A2(n4024), .ZN(n3135) );
  NAND2_X1 U3907 ( .A1(n3708), .A2(n4272), .ZN(n3134) );
  OAI211_X1 U3908 ( .C1(n4029), .C2(n3172), .A(n3135), .B(n3134), .ZN(n3136)
         );
  AOI21_X1 U3909 ( .B1(n3137), .B2(n4040), .A(n3136), .ZN(n3253) );
  XNOR2_X1 U3910 ( .A(n3138), .B(n3576), .ZN(n3251) );
  INV_X1 U3911 ( .A(n3139), .ZN(n3230) );
  AOI21_X1 U3912 ( .B1(n3140), .B2(n3194), .A(n3230), .ZN(n3260) );
  INV_X1 U3913 ( .A(n3260), .ZN(n3142) );
  AOI22_X1 U3914 ( .A1(n4463), .A2(REG2_REG_12__SCAN_IN), .B1(n3176), .B2(
        n4453), .ZN(n3141) );
  OAI21_X1 U3915 ( .B1(n3142), .B2(n4050), .A(n3141), .ZN(n3143) );
  AOI21_X1 U3916 ( .B1(n3251), .B2(n3999), .A(n3143), .ZN(n3144) );
  OAI21_X1 U3917 ( .B1(n3253), .B2(n4463), .A(n3144), .ZN(U3278) );
  NAND2_X1 U3918 ( .A1(n3146), .A2(n3145), .ZN(n3147) );
  NAND2_X2 U3919 ( .A1(n3148), .A2(n3147), .ZN(n3162) );
  OAI22_X1 U3920 ( .A1(n3173), .A2(n3353), .B1(n3352), .B2(n3195), .ZN(n3161)
         );
  NAND2_X1 U3921 ( .A1(n3710), .A2(n2779), .ZN(n3150) );
  INV_X1 U3922 ( .A(n3195), .ZN(n3156) );
  NAND2_X1 U3923 ( .A1(n3357), .A2(n3156), .ZN(n3149) );
  NAND2_X1 U3924 ( .A1(n3150), .A2(n3149), .ZN(n3151) );
  XNOR2_X1 U3925 ( .A(n3151), .B(n3358), .ZN(n3160) );
  XOR2_X1 U3926 ( .A(n3161), .B(n3160), .Z(n3152) );
  XNOR2_X1 U3927 ( .A(n3162), .B(n3152), .ZN(n3159) );
  INV_X1 U3928 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3153) );
  NOR2_X1 U3929 ( .A1(STATE_REG_SCAN_IN), .A2(n3153), .ZN(n4376) );
  OAI22_X1 U3930 ( .A1(n3244), .A2(n3529), .B1(n3530), .B2(n3154), .ZN(n3155)
         );
  AOI211_X1 U3931 ( .C1(n3156), .C2(n3532), .A(n4376), .B(n3155), .ZN(n3158)
         );
  NAND2_X1 U3932 ( .A1(n3533), .A2(n3197), .ZN(n3157) );
  OAI211_X1 U3933 ( .C1(n3159), .C2(n3536), .A(n3158), .B(n3157), .ZN(U3233)
         );
  OAI21_X1 U3934 ( .B1(n3162), .B2(n3161), .A(n3160), .ZN(n3164) );
  NAND2_X1 U3935 ( .A1(n3162), .A2(n3161), .ZN(n3163) );
  NAND2_X1 U3936 ( .A1(n3164), .A2(n3163), .ZN(n3237) );
  OAI22_X1 U3937 ( .A1(n3244), .A2(n3352), .B1(n3348), .B2(n3172), .ZN(n3165)
         );
  XNOR2_X1 U3938 ( .A(n3165), .B(n3358), .ZN(n3169) );
  INV_X1 U3939 ( .A(n3169), .ZN(n3167) );
  OAI22_X1 U3940 ( .A1(n3244), .A2(n3353), .B1(n3352), .B2(n3172), .ZN(n3168)
         );
  INV_X1 U3941 ( .A(n3168), .ZN(n3166) );
  NAND2_X1 U3942 ( .A1(n3167), .A2(n3166), .ZN(n3235) );
  INV_X1 U3943 ( .A(n3235), .ZN(n3170) );
  AND2_X1 U3944 ( .A1(n3169), .A2(n3168), .ZN(n3236) );
  NOR2_X1 U3945 ( .A1(n3170), .A2(n3236), .ZN(n3171) );
  XNOR2_X1 U3946 ( .A(n3237), .B(n3171), .ZN(n3178) );
  NAND2_X1 U3947 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4386) );
  OAI21_X1 U3948 ( .B1(n3517), .B2(n3172), .A(n4386), .ZN(n3175) );
  INV_X1 U3949 ( .A(n3708), .ZN(n3389) );
  OAI22_X1 U3950 ( .A1(n3173), .A2(n3530), .B1(n3529), .B2(n3389), .ZN(n3174)
         );
  AOI211_X1 U3951 ( .C1(n3176), .C2(n3533), .A(n3175), .B(n3174), .ZN(n3177)
         );
  OAI21_X1 U3952 ( .B1(n3178), .B2(n3536), .A(n3177), .ZN(U3221) );
  AOI21_X1 U3953 ( .B1(n4524), .B2(n3180), .A(n3179), .ZN(n3182) );
  MUX2_X1 U3954 ( .A(n4188), .B(n3182), .S(n4567), .Z(n3181) );
  OAI21_X1 U3955 ( .B1(n3185), .B2(n4268), .A(n3181), .ZN(U3528) );
  INV_X1 U3956 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3183) );
  MUX2_X1 U3957 ( .A(n3183), .B(n3182), .S(n4555), .Z(n3184) );
  OAI21_X1 U3958 ( .B1(n3185), .B2(n4325), .A(n3184), .ZN(U3487) );
  XNOR2_X1 U3959 ( .A(n3187), .B(n3186), .ZN(n3193) );
  OAI22_X1 U3960 ( .A1(n3244), .A2(n3946), .B1(n3195), .B2(n4029), .ZN(n3190)
         );
  AOI21_X1 U3961 ( .B1(n3590), .B2(n3188), .A(n2036), .ZN(n4550) );
  NOR2_X1 U3962 ( .A1(n4550), .A2(n4270), .ZN(n3189) );
  AOI211_X1 U3963 ( .C1(n4024), .C2(n3191), .A(n3190), .B(n3189), .ZN(n3192)
         );
  OAI21_X1 U3964 ( .B1(n4269), .B2(n3193), .A(n3192), .ZN(n4552) );
  INV_X1 U3965 ( .A(n4552), .ZN(n3202) );
  INV_X1 U3966 ( .A(n4550), .ZN(n3200) );
  OAI21_X1 U3967 ( .B1(n3196), .B2(n3195), .A(n3194), .ZN(n4547) );
  AOI22_X1 U3968 ( .A1(n4463), .A2(REG2_REG_11__SCAN_IN), .B1(n3197), .B2(
        n4453), .ZN(n3198) );
  OAI21_X1 U3969 ( .B1(n4547), .B2(n4050), .A(n3198), .ZN(n3199) );
  AOI21_X1 U3970 ( .B1(n3200), .B2(n4466), .A(n3199), .ZN(n3201) );
  OAI21_X1 U3971 ( .B1(n3202), .B2(n4463), .A(n3201), .ZN(U3279) );
  XNOR2_X1 U3972 ( .A(n3550), .B(n3591), .ZN(n3203) );
  NAND2_X1 U3973 ( .A1(n3203), .A2(n4040), .ZN(n3206) );
  OAI22_X1 U3974 ( .A1(n3455), .A2(n3946), .B1(n3388), .B2(n4029), .ZN(n3204)
         );
  INV_X1 U3975 ( .A(n3204), .ZN(n3205) );
  OAI211_X1 U3976 ( .C1(n3389), .C2(n4044), .A(n3206), .B(n3205), .ZN(n4261)
         );
  INV_X1 U3977 ( .A(n4261), .ZN(n3215) );
  OAI21_X1 U3978 ( .B1(n3207), .B2(n3209), .A(n3208), .ZN(n4262) );
  INV_X1 U3979 ( .A(n3229), .ZN(n3211) );
  INV_X1 U3980 ( .A(n4047), .ZN(n3210) );
  OAI21_X1 U3981 ( .B1(n3211), .B2(n3388), .A(n3210), .ZN(n4321) );
  AOI22_X1 U3982 ( .A1(n4463), .A2(REG2_REG_14__SCAN_IN), .B1(n3392), .B2(
        n4453), .ZN(n3212) );
  OAI21_X1 U3983 ( .B1(n4321), .B2(n4050), .A(n3212), .ZN(n3213) );
  AOI21_X1 U3984 ( .B1(n4262), .B2(n3999), .A(n3213), .ZN(n3214) );
  OAI21_X1 U3985 ( .B1(n4463), .B2(n3215), .A(n3214), .ZN(U3276) );
  INV_X1 U3986 ( .A(n3216), .ZN(n3218) );
  NAND2_X1 U3987 ( .A1(n3218), .A2(n3217), .ZN(n3588) );
  XOR2_X1 U3988 ( .A(n3588), .B(n3219), .Z(n3228) );
  OAI21_X1 U3989 ( .B1(n3222), .B2(n3221), .A(n3220), .ZN(n3223) );
  XOR2_X1 U3990 ( .A(n3588), .B(n3223), .Z(n3226) );
  AOI22_X1 U3991 ( .A1(n3707), .A2(n4272), .B1(n4064), .B2(n3246), .ZN(n3224)
         );
  OAI21_X1 U3992 ( .B1(n3244), .B2(n4044), .A(n3224), .ZN(n3225) );
  AOI21_X1 U3993 ( .B1(n3226), .B2(n4040), .A(n3225), .ZN(n3227) );
  OAI21_X1 U3994 ( .B1(n3228), .B2(n4270), .A(n3227), .ZN(n4264) );
  INV_X1 U3995 ( .A(n4264), .ZN(n3234) );
  INV_X1 U3996 ( .A(n3228), .ZN(n4265) );
  OAI21_X1 U3997 ( .B1(n3230), .B2(n3238), .A(n3229), .ZN(n4326) );
  AOI22_X1 U3998 ( .A1(n4463), .A2(REG2_REG_13__SCAN_IN), .B1(n3247), .B2(
        n4453), .ZN(n3231) );
  OAI21_X1 U3999 ( .B1(n4326), .B2(n4050), .A(n3231), .ZN(n3232) );
  AOI21_X1 U4000 ( .B1(n4265), .B2(n4466), .A(n3232), .ZN(n3233) );
  OAI21_X1 U4001 ( .B1(n3234), .B2(n4463), .A(n3233), .ZN(U3277) );
  OAI21_X2 U4002 ( .B1(n3237), .B2(n3236), .A(n3235), .ZN(n3263) );
  OAI22_X1 U4003 ( .A1(n3389), .A2(n3353), .B1(n3352), .B2(n3238), .ZN(n3262)
         );
  NAND2_X1 U4004 ( .A1(n3708), .A2(n2779), .ZN(n3240) );
  NAND2_X1 U4005 ( .A1(n3357), .A2(n3246), .ZN(n3239) );
  NAND2_X1 U4006 ( .A1(n3240), .A2(n3239), .ZN(n3241) );
  XNOR2_X1 U4007 ( .A(n3241), .B(n3324), .ZN(n3264) );
  XOR2_X1 U4008 ( .A(n3262), .B(n3264), .Z(n3242) );
  XNOR2_X1 U4009 ( .A(n3263), .B(n3242), .ZN(n3250) );
  NOR2_X1 U4010 ( .A1(STATE_REG_SCAN_IN), .A2(n3243), .ZN(n4396) );
  INV_X1 U4011 ( .A(n3707), .ZN(n4045) );
  OAI22_X1 U4012 ( .A1(n3244), .A2(n3530), .B1(n3529), .B2(n4045), .ZN(n3245)
         );
  AOI211_X1 U4013 ( .C1(n3246), .C2(n3532), .A(n4396), .B(n3245), .ZN(n3249)
         );
  NAND2_X1 U4014 ( .A1(n3533), .A2(n3247), .ZN(n3248) );
  OAI211_X1 U4015 ( .C1(n3250), .C2(n3536), .A(n3249), .B(n3248), .ZN(U3231)
         );
  NAND2_X1 U4016 ( .A1(n3251), .A2(n4533), .ZN(n3252) );
  NAND2_X1 U4017 ( .A1(n3253), .A2(n3252), .ZN(n3257) );
  MUX2_X1 U4018 ( .A(REG1_REG_12__SCAN_IN), .B(n3257), .S(n4567), .Z(n3254) );
  AOI21_X1 U4019 ( .B1(n3255), .B2(n3260), .A(n3254), .ZN(n3256) );
  INV_X1 U4020 ( .A(n3256), .ZN(U3530) );
  MUX2_X1 U4021 ( .A(REG0_REG_12__SCAN_IN), .B(n3257), .S(n4555), .Z(n3258) );
  AOI21_X1 U4022 ( .B1(n3260), .B2(n3259), .A(n3258), .ZN(n3261) );
  INV_X1 U4023 ( .A(n3261), .ZN(U3491) );
  INV_X1 U4024 ( .A(n3264), .ZN(n3265) );
  NAND2_X1 U4025 ( .A1(n3707), .A2(n2779), .ZN(n3268) );
  NAND2_X1 U4026 ( .A1(n3357), .A2(n3266), .ZN(n3267) );
  NAND2_X1 U4027 ( .A1(n3268), .A2(n3267), .ZN(n3269) );
  XNOR2_X1 U4028 ( .A(n3269), .B(n3324), .ZN(n3274) );
  INV_X1 U4029 ( .A(n3274), .ZN(n3272) );
  NOR2_X1 U4030 ( .A1(n3352), .A2(n3388), .ZN(n3270) );
  AOI21_X1 U4031 ( .B1(n3356), .B2(n3707), .A(n3270), .ZN(n3273) );
  INV_X1 U4032 ( .A(n3273), .ZN(n3271) );
  NAND2_X1 U4033 ( .A1(n3272), .A2(n3271), .ZN(n3385) );
  OAI22_X1 U4034 ( .A1(n3455), .A2(n3352), .B1(n3348), .B2(n3275), .ZN(n3276)
         );
  XNOR2_X1 U4035 ( .A(n3276), .B(n3358), .ZN(n3279) );
  OR2_X1 U4036 ( .A1(n3353), .A2(n3455), .ZN(n3278) );
  NAND2_X1 U4037 ( .A1(n2779), .A2(n4046), .ZN(n3277) );
  NAND2_X1 U4038 ( .A1(n3278), .A2(n3277), .ZN(n3526) );
  INV_X1 U4039 ( .A(n3526), .ZN(n3452) );
  NOR2_X1 U4040 ( .A1(n3451), .A2(n3452), .ZN(n3287) );
  NAND2_X1 U4041 ( .A1(n3280), .A2(n3279), .ZN(n3450) );
  OAI22_X1 U4042 ( .A1(n4014), .A2(n3352), .B1(n4028), .B2(n3348), .ZN(n3281)
         );
  XNOR2_X1 U40430 ( .A(n3281), .B(n3358), .ZN(n3283) );
  OAI22_X1 U4044 ( .A1(n4014), .A2(n3353), .B1(n4028), .B2(n3352), .ZN(n3282)
         );
  NOR2_X1 U4045 ( .A1(n3283), .A2(n3282), .ZN(n3284) );
  AOI21_X1 U4046 ( .B1(n3283), .B2(n3282), .A(n3284), .ZN(n3453) );
  NAND2_X1 U4047 ( .A1(n3450), .A2(n3453), .ZN(n3286) );
  INV_X1 U4048 ( .A(n3284), .ZN(n3285) );
  OAI21_X1 U4049 ( .B1(n3287), .B2(n3286), .A(n3285), .ZN(n3460) );
  OAI22_X1 U4050 ( .A1(n3985), .A2(n3352), .B1(n3348), .B2(n3467), .ZN(n3288)
         );
  XNOR2_X1 U4051 ( .A(n3288), .B(n3358), .ZN(n3290) );
  OAI22_X1 U4052 ( .A1(n3985), .A2(n3353), .B1(n3352), .B2(n3467), .ZN(n3289)
         );
  NAND2_X1 U4053 ( .A1(n3290), .A2(n3289), .ZN(n3462) );
  NOR2_X1 U4054 ( .A1(n3290), .A2(n3289), .ZN(n3461) );
  AOI21_X1 U4055 ( .B1(n3460), .B2(n3462), .A(n3461), .ZN(n3405) );
  NAND2_X1 U4056 ( .A1(n3983), .A2(n2779), .ZN(n3292) );
  NAND2_X1 U4057 ( .A1(n3357), .A2(n3415), .ZN(n3291) );
  NAND2_X1 U4058 ( .A1(n3292), .A2(n3291), .ZN(n3293) );
  XNOR2_X1 U4059 ( .A(n3293), .B(n3324), .ZN(n3303) );
  NOR2_X1 U4060 ( .A1(n3352), .A2(n3973), .ZN(n3294) );
  AOI21_X1 U4061 ( .B1(n3356), .B2(n3983), .A(n3294), .ZN(n3304) );
  NOR2_X1 U4062 ( .A1(n3303), .A2(n3304), .ZN(n3410) );
  NAND2_X1 U4063 ( .A1(n4011), .A2(n2779), .ZN(n3296) );
  NAND2_X1 U4064 ( .A1(n3357), .A2(n3991), .ZN(n3295) );
  NAND2_X1 U4065 ( .A1(n3296), .A2(n3295), .ZN(n3297) );
  XNOR2_X1 U4066 ( .A(n3297), .B(n3358), .ZN(n3503) );
  NAND2_X1 U4067 ( .A1(n3356), .A2(n4011), .ZN(n3299) );
  NAND2_X1 U4068 ( .A1(n2779), .A2(n3991), .ZN(n3298) );
  NAND2_X1 U4069 ( .A1(n3299), .A2(n3298), .ZN(n3406) );
  NOR2_X1 U4070 ( .A1(n3405), .A2(n3302), .ZN(n3308) );
  NOR3_X1 U4071 ( .A1(n3410), .A2(n3406), .A3(n3503), .ZN(n3307) );
  INV_X1 U4072 ( .A(n3303), .ZN(n3306) );
  INV_X1 U4073 ( .A(n3304), .ZN(n3305) );
  NOR2_X1 U4074 ( .A1(n3306), .A2(n3305), .ZN(n3409) );
  NAND2_X1 U4075 ( .A1(n3969), .A2(n2779), .ZN(n3310) );
  OR2_X1 U4076 ( .A1(n3348), .A2(n3953), .ZN(n3309) );
  NAND2_X1 U4077 ( .A1(n3310), .A2(n3309), .ZN(n3311) );
  XNOR2_X1 U4078 ( .A(n3311), .B(n3324), .ZN(n3314) );
  NOR2_X1 U4079 ( .A1(n3352), .A2(n3953), .ZN(n3312) );
  AOI21_X1 U4080 ( .B1(n3356), .B2(n3969), .A(n3312), .ZN(n3313) );
  NOR2_X1 U4081 ( .A1(n3314), .A2(n3313), .ZN(n3483) );
  AND2_X1 U4082 ( .A1(n3314), .A2(n3313), .ZN(n3430) );
  NAND2_X1 U4083 ( .A1(n3706), .A2(n2779), .ZN(n3316) );
  OR2_X1 U4084 ( .A1(n3348), .A2(n3932), .ZN(n3315) );
  NAND2_X1 U4085 ( .A1(n3316), .A2(n3315), .ZN(n3317) );
  XNOR2_X1 U4086 ( .A(n3317), .B(n3324), .ZN(n3320) );
  NOR2_X1 U4087 ( .A1(n3352), .A2(n3932), .ZN(n3318) );
  AOI21_X1 U4088 ( .B1(n3706), .B2(n3356), .A(n3318), .ZN(n3319) );
  AND2_X1 U4089 ( .A1(n3320), .A2(n3319), .ZN(n3427) );
  NOR2_X1 U4090 ( .A1(n3320), .A2(n3319), .ZN(n3428) );
  OAI22_X1 U4091 ( .A1(n3898), .A2(n3353), .B1(n3910), .B2(n3352), .ZN(n3327)
         );
  OAI22_X1 U4092 ( .A1(n3898), .A2(n3352), .B1(n3910), .B2(n3348), .ZN(n3321)
         );
  XNOR2_X1 U4093 ( .A(n3321), .B(n3358), .ZN(n3326) );
  XOR2_X1 U4094 ( .A(n3327), .B(n3326), .Z(n3494) );
  NAND2_X1 U4095 ( .A1(n3493), .A2(n3494), .ZN(n3396) );
  NAND2_X1 U4096 ( .A1(n3869), .A2(n2779), .ZN(n3323) );
  OR2_X1 U4097 ( .A1(n3348), .A2(n3901), .ZN(n3322) );
  NAND2_X1 U4098 ( .A1(n3323), .A2(n3322), .ZN(n3325) );
  XNOR2_X1 U4099 ( .A(n3325), .B(n3324), .ZN(n3331) );
  OAI22_X1 U4100 ( .A1(n3911), .A2(n3338), .B1(n3352), .B2(n3901), .ZN(n3332)
         );
  XNOR2_X1 U4101 ( .A(n3331), .B(n3332), .ZN(n3397) );
  INV_X1 U4102 ( .A(n3326), .ZN(n3329) );
  INV_X1 U4103 ( .A(n3327), .ZN(n3328) );
  NAND2_X1 U4104 ( .A1(n3329), .A2(n3328), .ZN(n3398) );
  NAND3_X2 U4105 ( .A1(n3396), .A2(n3397), .A3(n3398), .ZN(n3395) );
  NOR2_X1 U4106 ( .A1(n3352), .A2(n3876), .ZN(n3330) );
  AOI21_X1 U4107 ( .B1(n3356), .B2(n3895), .A(n3330), .ZN(n3335) );
  INV_X1 U4108 ( .A(n3331), .ZN(n3333) );
  NAND2_X1 U4109 ( .A1(n3333), .A2(n3332), .ZN(n3336) );
  NAND3_X1 U4110 ( .A1(n3395), .A2(n3335), .A3(n3336), .ZN(n3473) );
  OAI22_X1 U4111 ( .A1(n3855), .A2(n3352), .B1(n3348), .B2(n3876), .ZN(n3334)
         );
  XNOR2_X1 U4112 ( .A(n3334), .B(n3358), .ZN(n3476) );
  AOI21_X2 U4113 ( .B1(n3395), .B2(n3336), .A(n3335), .ZN(n3475) );
  AOI21_X2 U4114 ( .B1(n3473), .B2(n3476), .A(n3475), .ZN(n3443) );
  OAI22_X1 U4115 ( .A1(n3839), .A2(n3352), .B1(n3348), .B2(n3857), .ZN(n3337)
         );
  XNOR2_X1 U4116 ( .A(n3337), .B(n3358), .ZN(n3340) );
  OAI22_X1 U4117 ( .A1(n3839), .A2(n3338), .B1(n3352), .B2(n3857), .ZN(n3339)
         );
  NOR2_X1 U4118 ( .A1(n3340), .A2(n3339), .ZN(n3440) );
  NAND2_X1 U4119 ( .A1(n3340), .A2(n3339), .ZN(n3441) );
  NAND2_X1 U4120 ( .A1(n3852), .A2(n2779), .ZN(n3342) );
  OR2_X1 U4121 ( .A1(n3348), .A2(n3841), .ZN(n3341) );
  NAND2_X1 U4122 ( .A1(n3342), .A2(n3341), .ZN(n3343) );
  XNOR2_X1 U4123 ( .A(n3343), .B(n3358), .ZN(n3344) );
  INV_X1 U4124 ( .A(n3852), .ZN(n3445) );
  OAI22_X1 U4125 ( .A1(n3445), .A2(n3353), .B1(n3841), .B2(n3352), .ZN(n3345)
         );
  AND2_X1 U4126 ( .A1(n3344), .A2(n3345), .ZN(n3513) );
  INV_X1 U4127 ( .A(n3344), .ZN(n3347) );
  INV_X1 U4128 ( .A(n3345), .ZN(n3346) );
  NAND2_X1 U4129 ( .A1(n3347), .A2(n3346), .ZN(n3512) );
  NAND2_X1 U4130 ( .A1(n3836), .A2(n2779), .ZN(n3350) );
  OR2_X1 U4131 ( .A1(n3348), .A2(n3823), .ZN(n3349) );
  NAND2_X1 U4132 ( .A1(n3350), .A2(n3349), .ZN(n3351) );
  XNOR2_X1 U4133 ( .A(n3351), .B(n3358), .ZN(n3355) );
  OAI22_X1 U4134 ( .A1(n3518), .A2(n3353), .B1(n3352), .B2(n3823), .ZN(n3354)
         );
  XNOR2_X1 U4135 ( .A(n3355), .B(n3354), .ZN(n3378) );
  INV_X1 U4136 ( .A(n3364), .ZN(n3796) );
  AOI22_X1 U4137 ( .A1(n3356), .A2(n3820), .B1(n3796), .B2(n2779), .ZN(n3361)
         );
  AOI22_X1 U4138 ( .A1(n2779), .A2(n3820), .B1(n3357), .B2(n3796), .ZN(n3359)
         );
  XNOR2_X1 U4139 ( .A(n3359), .B(n3358), .ZN(n3360) );
  XOR2_X1 U4140 ( .A(n3361), .B(n3360), .Z(n3362) );
  INV_X1 U4141 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3363) );
  OAI22_X1 U4142 ( .A1(n3517), .A2(n3364), .B1(STATE_REG_SCAN_IN), .B2(n3363), 
        .ZN(n3367) );
  INV_X1 U4143 ( .A(n3705), .ZN(n3365) );
  OAI22_X1 U4144 ( .A1(n3518), .A2(n3530), .B1(n3529), .B2(n3365), .ZN(n3366)
         );
  AOI211_X1 U4145 ( .C1(n3371), .C2(n3533), .A(n3367), .B(n3366), .ZN(n3368)
         );
  OAI21_X1 U4146 ( .B1(n3369), .B2(n3536), .A(n3368), .ZN(U3217) );
  INV_X1 U4147 ( .A(n3370), .ZN(n3375) );
  AOI22_X1 U4148 ( .A1(n4463), .A2(REG2_REG_28__SCAN_IN), .B1(n3371), .B2(
        n4453), .ZN(n3372) );
  OAI21_X1 U4149 ( .B1(n3373), .B2(n4050), .A(n3372), .ZN(n3374) );
  AOI21_X1 U4150 ( .B1(n3375), .B2(n4470), .A(n3374), .ZN(n3376) );
  OAI21_X1 U4151 ( .B1(n3377), .B2(n4054), .A(n3376), .ZN(U3262) );
  XNOR2_X1 U4152 ( .A(n3379), .B(n3378), .ZN(n3384) );
  OAI22_X1 U4153 ( .A1(n3517), .A2(n3823), .B1(STATE_REG_SCAN_IN), .B2(n4179), 
        .ZN(n3382) );
  INV_X1 U4154 ( .A(n3820), .ZN(n3380) );
  OAI22_X1 U4155 ( .A1(n3445), .A2(n3530), .B1(n3529), .B2(n3380), .ZN(n3381)
         );
  AOI211_X1 U4156 ( .C1(n3814), .C2(n3533), .A(n3382), .B(n3381), .ZN(n3383)
         );
  OAI21_X1 U4157 ( .B1(n3384), .B2(n3536), .A(n3383), .ZN(U3211) );
  NAND2_X1 U4158 ( .A1(n2046), .A2(n3385), .ZN(n3386) );
  XNOR2_X1 U4159 ( .A(n3387), .B(n3386), .ZN(n3394) );
  NAND2_X1 U4160 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4412) );
  OAI21_X1 U4161 ( .B1(n3517), .B2(n3388), .A(n4412), .ZN(n3391) );
  OAI22_X1 U4162 ( .A1(n3455), .A2(n3529), .B1(n3530), .B2(n3389), .ZN(n3390)
         );
  AOI211_X1 U4163 ( .C1(n3392), .C2(n3533), .A(n3391), .B(n3390), .ZN(n3393)
         );
  OAI21_X1 U4164 ( .B1(n3394), .B2(n3536), .A(n3393), .ZN(U3212) );
  NAND2_X1 U4165 ( .A1(n3395), .A2(n3495), .ZN(n3404) );
  AOI21_X1 U4166 ( .B1(n3396), .B2(n3398), .A(n3397), .ZN(n3403) );
  INV_X1 U4167 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3399) );
  OAI22_X1 U4168 ( .A1(n3517), .A2(n3901), .B1(STATE_REG_SCAN_IN), .B2(n3399), 
        .ZN(n3401) );
  OAI22_X1 U4169 ( .A1(n3898), .A2(n3530), .B1(n3529), .B2(n3855), .ZN(n3400)
         );
  AOI211_X1 U4170 ( .C1(n3902), .C2(n3533), .A(n3401), .B(n3400), .ZN(n3402)
         );
  OAI21_X1 U4171 ( .B1(n3404), .B2(n3403), .A(n3402), .ZN(U3213) );
  INV_X1 U4172 ( .A(n3506), .ZN(n3408) );
  INV_X1 U4173 ( .A(n3406), .ZN(n3504) );
  OAI21_X1 U4174 ( .B1(n3506), .B2(n3406), .A(n3503), .ZN(n3407) );
  OAI21_X1 U4175 ( .B1(n3408), .B2(n3504), .A(n3407), .ZN(n3412) );
  NOR2_X1 U4176 ( .A1(n3410), .A2(n3409), .ZN(n3411) );
  XNOR2_X1 U4177 ( .A(n3412), .B(n3411), .ZN(n3418) );
  NOR2_X1 U4178 ( .A1(n3413), .A2(STATE_REG_SCAN_IN), .ZN(n3778) );
  INV_X1 U4179 ( .A(n3969), .ZN(n3435) );
  OAI22_X1 U4180 ( .A1(n3972), .A2(n3530), .B1(n3529), .B2(n3435), .ZN(n3414)
         );
  AOI211_X1 U4181 ( .C1(n3415), .C2(n3532), .A(n3778), .B(n3414), .ZN(n3417)
         );
  NAND2_X1 U4182 ( .A1(n3533), .A2(n3977), .ZN(n3416) );
  OAI211_X1 U4183 ( .C1(n3418), .C2(n3536), .A(n3417), .B(n3416), .ZN(U3216)
         );
  AOI22_X1 U4184 ( .A1(n3419), .A2(n3532), .B1(n3497), .B2(n3720), .ZN(n3426)
         );
  AOI22_X1 U4185 ( .A1(n3420), .A2(REG3_REG_1__SCAN_IN), .B1(n3498), .B2(n2273), .ZN(n3425) );
  OAI211_X1 U4186 ( .C1(n3423), .C2(n3422), .A(n3421), .B(n3495), .ZN(n3424)
         );
  NAND3_X1 U4187 ( .A1(n3426), .A2(n3425), .A3(n3424), .ZN(U3219) );
  NOR2_X1 U4188 ( .A1(n3428), .A2(n3427), .ZN(n3432) );
  INV_X1 U4189 ( .A(n3430), .ZN(n3486) );
  AOI21_X1 U4190 ( .B1(n3429), .B2(n3486), .A(n3483), .ZN(n3431) );
  XOR2_X1 U4191 ( .A(n3432), .B(n3431), .Z(n3439) );
  INV_X1 U4192 ( .A(n3433), .ZN(n3934) );
  OAI22_X1 U4193 ( .A1(n3517), .A2(n3932), .B1(STATE_REG_SCAN_IN), .B2(n3434), 
        .ZN(n3437) );
  OAI22_X1 U4194 ( .A1(n3435), .A2(n3530), .B1(n3529), .B2(n3898), .ZN(n3436)
         );
  AOI211_X1 U4195 ( .C1(n3934), .C2(n3533), .A(n3437), .B(n3436), .ZN(n3438)
         );
  OAI21_X1 U4196 ( .B1(n3439), .B2(n3536), .A(n3438), .ZN(U3220) );
  NAND2_X1 U4197 ( .A1(n2199), .A2(n3441), .ZN(n3442) );
  XNOR2_X1 U4198 ( .A(n3443), .B(n3442), .ZN(n3449) );
  INV_X1 U4199 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3444) );
  OAI22_X1 U4200 ( .A1(n3517), .A2(n3857), .B1(STATE_REG_SCAN_IN), .B2(n3444), 
        .ZN(n3447) );
  OAI22_X1 U4201 ( .A1(n3855), .A2(n3530), .B1(n3529), .B2(n3445), .ZN(n3446)
         );
  AOI211_X1 U4202 ( .C1(n3859), .C2(n3533), .A(n3447), .B(n3446), .ZN(n3448)
         );
  OAI21_X1 U4203 ( .B1(n3449), .B2(n3536), .A(n3448), .ZN(U3222) );
  AOI21_X1 U4204 ( .B1(n3452), .B2(n3523), .A(n3525), .ZN(n3454) );
  XNOR2_X1 U4205 ( .A(n3454), .B(n3453), .ZN(n3459) );
  NAND2_X1 U4206 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4425) );
  OAI21_X1 U4207 ( .B1(n3517), .B2(n4028), .A(n4425), .ZN(n3457) );
  OAI22_X1 U4208 ( .A1(n3985), .A2(n3529), .B1(n3530), .B2(n3455), .ZN(n3456)
         );
  AOI211_X1 U4209 ( .C1(n4033), .C2(n3533), .A(n3457), .B(n3456), .ZN(n3458)
         );
  OAI21_X1 U4210 ( .B1(n3459), .B2(n3536), .A(n3458), .ZN(U3223) );
  INV_X1 U4211 ( .A(n3461), .ZN(n3463) );
  NAND2_X1 U4212 ( .A1(n3463), .A2(n3462), .ZN(n3464) );
  XNOR2_X1 U4213 ( .A(n3465), .B(n3464), .ZN(n3472) );
  INV_X1 U4214 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4230) );
  NOR2_X1 U4215 ( .A1(STATE_REG_SCAN_IN), .A2(n4230), .ZN(n3748) );
  INV_X1 U4216 ( .A(n3748), .ZN(n3466) );
  OAI21_X1 U4217 ( .B1(n3517), .B2(n3467), .A(n3466), .ZN(n3469) );
  OAI22_X1 U4218 ( .A1(n4014), .A2(n3530), .B1(n3529), .B2(n3972), .ZN(n3468)
         );
  AOI211_X1 U4219 ( .C1(n3470), .C2(n3533), .A(n3469), .B(n3468), .ZN(n3471)
         );
  OAI21_X1 U4220 ( .B1(n3472), .B2(n3536), .A(n3471), .ZN(U3225) );
  INV_X1 U4221 ( .A(n3473), .ZN(n3474) );
  NOR2_X1 U4222 ( .A1(n3475), .A2(n3474), .ZN(n3477) );
  XNOR2_X1 U4223 ( .A(n3477), .B(n3476), .ZN(n3482) );
  INV_X1 U4224 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3478) );
  OAI22_X1 U4225 ( .A1(n3517), .A2(n3876), .B1(STATE_REG_SCAN_IN), .B2(n3478), 
        .ZN(n3480) );
  OAI22_X1 U4226 ( .A1(n3911), .A2(n3530), .B1(n3529), .B2(n3839), .ZN(n3479)
         );
  AOI211_X1 U4227 ( .C1(n3877), .C2(n3533), .A(n3480), .B(n3479), .ZN(n3481)
         );
  OAI21_X1 U4228 ( .B1(n3482), .B2(n3536), .A(n3481), .ZN(U3226) );
  INV_X1 U4229 ( .A(n3483), .ZN(n3484) );
  NAND2_X1 U4230 ( .A1(n3484), .A2(n3486), .ZN(n3485) );
  AOI22_X1 U4231 ( .A1(n2017), .A2(n3486), .B1(n3429), .B2(n3485), .ZN(n3492)
         );
  INV_X1 U4232 ( .A(n3487), .ZN(n3954) );
  OAI22_X1 U4233 ( .A1(n3517), .A2(n3953), .B1(STATE_REG_SCAN_IN), .B2(n3488), 
        .ZN(n3490) );
  INV_X1 U4234 ( .A(n3983), .ZN(n3507) );
  OAI22_X1 U4235 ( .A1(n3947), .A2(n3529), .B1(n3530), .B2(n3507), .ZN(n3489)
         );
  AOI211_X1 U4236 ( .C1(n3954), .C2(n3533), .A(n3490), .B(n3489), .ZN(n3491)
         );
  OAI21_X1 U4237 ( .B1(n3492), .B2(n3536), .A(n3491), .ZN(U3230) );
  OAI21_X1 U4238 ( .B1(n3494), .B2(n3493), .A(n3396), .ZN(n3496) );
  NAND2_X1 U4239 ( .A1(n3496), .A2(n3495), .ZN(n3502) );
  AOI22_X1 U4240 ( .A1(n3532), .A2(n3917), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3501) );
  AOI22_X1 U4241 ( .A1(n3498), .A2(n3869), .B1(n3497), .B2(n3706), .ZN(n3500)
         );
  NAND2_X1 U4242 ( .A1(n3533), .A2(n3915), .ZN(n3499) );
  NAND4_X1 U4243 ( .A1(n3502), .A2(n3501), .A3(n3500), .A4(n3499), .ZN(U3232)
         );
  XNOR2_X1 U4244 ( .A(n3504), .B(n3503), .ZN(n3505) );
  XNOR2_X1 U4245 ( .A(n3506), .B(n3505), .ZN(n3511) );
  OAI22_X1 U4246 ( .A1(n3985), .A2(n3530), .B1(n3529), .B2(n3507), .ZN(n3508)
         );
  AOI211_X1 U4247 ( .C1(n3991), .C2(n3532), .A(n2049), .B(n3508), .ZN(n3510)
         );
  NAND2_X1 U4248 ( .A1(n3533), .A2(n3994), .ZN(n3509) );
  OAI211_X1 U4249 ( .C1(n3511), .C2(n3536), .A(n3510), .B(n3509), .ZN(U3235)
         );
  NOR2_X1 U4250 ( .A1(n2195), .A2(n3513), .ZN(n3514) );
  XNOR2_X1 U4251 ( .A(n3515), .B(n3514), .ZN(n3522) );
  INV_X1 U4252 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3516) );
  OAI22_X1 U4253 ( .A1(n3517), .A2(n3841), .B1(STATE_REG_SCAN_IN), .B2(n3516), 
        .ZN(n3520) );
  OAI22_X1 U4254 ( .A1(n3839), .A2(n3530), .B1(n3529), .B2(n3518), .ZN(n3519)
         );
  AOI211_X1 U4255 ( .C1(n3842), .C2(n3533), .A(n3520), .B(n3519), .ZN(n3521)
         );
  OAI21_X1 U4256 ( .B1(n3522), .B2(n3536), .A(n3521), .ZN(U3237) );
  INV_X1 U4257 ( .A(n3523), .ZN(n3524) );
  NOR2_X1 U4258 ( .A1(n3525), .A2(n3524), .ZN(n3527) );
  XNOR2_X1 U4259 ( .A(n3527), .B(n3526), .ZN(n3537) );
  NOR2_X1 U4260 ( .A1(STATE_REG_SCAN_IN), .A2(n3528), .ZN(n4418) );
  OAI22_X1 U4261 ( .A1(n4045), .A2(n3530), .B1(n3529), .B2(n4014), .ZN(n3531)
         );
  AOI211_X1 U4262 ( .C1(n4046), .C2(n3532), .A(n4418), .B(n3531), .ZN(n3535)
         );
  NAND2_X1 U4263 ( .A1(n3533), .A2(n4048), .ZN(n3534) );
  OAI211_X1 U4264 ( .C1(n3537), .C2(n3536), .A(n3535), .B(n3534), .ZN(U3238)
         );
  NAND2_X1 U4265 ( .A1(n3538), .A2(REG1_REG_30__SCAN_IN), .ZN(n3541) );
  NAND2_X1 U4266 ( .A1(n2497), .A2(REG2_REG_30__SCAN_IN), .ZN(n3540) );
  NAND2_X1 U4267 ( .A1(n2258), .A2(REG0_REG_30__SCAN_IN), .ZN(n3539) );
  NAND3_X1 U4268 ( .A1(n3541), .A2(n3540), .A3(n3539), .ZN(n3790) );
  INV_X1 U4269 ( .A(n3790), .ZN(n3557) );
  NAND2_X1 U4270 ( .A1(n2295), .A2(DATAI_30_), .ZN(n3607) );
  NOR2_X1 U4271 ( .A1(n3557), .A2(n4065), .ZN(n3690) );
  NAND2_X1 U4272 ( .A1(n3538), .A2(REG1_REG_31__SCAN_IN), .ZN(n3544) );
  NAND2_X1 U4273 ( .A1(n2497), .A2(REG2_REG_31__SCAN_IN), .ZN(n3543) );
  NAND2_X1 U4274 ( .A1(n2258), .A2(REG0_REG_31__SCAN_IN), .ZN(n3542) );
  NAND3_X1 U4275 ( .A1(n3544), .A2(n3543), .A3(n3542), .ZN(n4057) );
  INV_X1 U4276 ( .A(n4057), .ZN(n3545) );
  NOR2_X1 U4277 ( .A1(n3690), .A2(n3545), .ZN(n3573) );
  NAND2_X1 U4278 ( .A1(n2006), .A2(DATAI_31_), .ZN(n4055) );
  NAND2_X1 U4279 ( .A1(n3604), .A2(n3583), .ZN(n3678) );
  NAND2_X1 U4280 ( .A1(n3546), .A2(n3549), .ZN(n3618) );
  NAND2_X1 U4281 ( .A1(n3548), .A2(n3547), .ZN(n3647) );
  NAND2_X1 U4282 ( .A1(n3647), .A2(n3549), .ZN(n3668) );
  OAI21_X1 U4283 ( .B1(n3550), .B2(n3618), .A(n3668), .ZN(n3552) );
  INV_X1 U4284 ( .A(n3551), .ZN(n3670) );
  AOI21_X1 U4285 ( .B1(n3552), .B2(n3669), .A(n3670), .ZN(n3555) );
  OAI21_X1 U4286 ( .B1(n3555), .B2(n3554), .A(n3553), .ZN(n3558) );
  NAND2_X1 U4287 ( .A1(n4057), .A2(n4055), .ZN(n3688) );
  INV_X1 U4288 ( .A(n3688), .ZN(n3556) );
  AOI21_X1 U4289 ( .B1(n3557), .B2(n4065), .A(n3556), .ZN(n3567) );
  OAI221_X1 U4290 ( .B1(n3678), .B2(n3681), .C1(n3678), .C2(n3558), .A(n3567), 
        .ZN(n3563) );
  NAND2_X1 U4291 ( .A1(n2006), .A2(DATAI_29_), .ZN(n3803) );
  OR2_X1 U4292 ( .A1(n3705), .A2(n3803), .ZN(n3603) );
  INV_X1 U4293 ( .A(n3603), .ZN(n3562) );
  INV_X1 U4294 ( .A(n3785), .ZN(n3560) );
  NOR2_X1 U4295 ( .A1(n3560), .A2(n3559), .ZN(n3569) );
  INV_X1 U4296 ( .A(n3569), .ZN(n3561) );
  NOR4_X1 U4297 ( .A1(n3563), .A2(n3562), .A3(n3685), .A4(n3561), .ZN(n3571)
         );
  NAND2_X1 U4298 ( .A1(n3705), .A2(n3803), .ZN(n3602) );
  INV_X1 U4299 ( .A(n3602), .ZN(n3565) );
  INV_X1 U4300 ( .A(n3566), .ZN(n3786) );
  NOR3_X1 U4301 ( .A1(n3565), .A2(n3786), .A3(n3564), .ZN(n3682) );
  NAND2_X1 U4302 ( .A1(n3602), .A2(n3566), .ZN(n3568) );
  OAI211_X1 U4303 ( .C1(n3569), .C2(n3568), .A(n3567), .B(n3603), .ZN(n3692)
         );
  AOI21_X1 U4304 ( .B1(n3818), .B2(n3682), .A(n3692), .ZN(n3570) );
  OAI22_X1 U4305 ( .A1(n3571), .A2(n3570), .B1(n4057), .B2(n3607), .ZN(n3572)
         );
  OAI21_X1 U4306 ( .B1(n3573), .B2(n4055), .A(n3572), .ZN(n3616) );
  NAND2_X1 U4307 ( .A1(n3960), .A2(n3883), .ZN(n4007) );
  OR4_X1 U4308 ( .A1(n4007), .A2(n3576), .A3(n3575), .A4(n3574), .ZN(n3595) );
  INV_X1 U4309 ( .A(n3577), .ZN(n3889) );
  NOR2_X1 U4310 ( .A1(n3889), .A2(n3676), .ZN(n3923) );
  INV_X1 U4311 ( .A(n3578), .ZN(n3579) );
  OR2_X1 U4312 ( .A1(n3580), .A2(n3579), .ZN(n3942) );
  INV_X1 U4313 ( .A(n3942), .ZN(n3585) );
  AND2_X1 U4314 ( .A1(n2126), .A2(n3582), .ZN(n3965) );
  XNOR2_X1 U4315 ( .A(n3869), .B(n3901), .ZN(n3892) );
  NAND2_X1 U4316 ( .A1(n3584), .A2(n3583), .ZN(n3866) );
  NOR4_X1 U4317 ( .A1(n3585), .A2(n3965), .A3(n3892), .A4(n3866), .ZN(n3586)
         );
  OR2_X1 U4318 ( .A1(n4057), .A2(n4055), .ZN(n3687) );
  NAND4_X1 U4319 ( .A1(n3923), .A2(n3586), .A3(n3687), .A4(n3688), .ZN(n3594)
         );
  NOR2_X1 U4320 ( .A1(n3587), .A2(n2016), .ZN(n3828) );
  INV_X1 U4321 ( .A(n3828), .ZN(n3832) );
  NAND3_X1 U4322 ( .A1(n4021), .A2(n3832), .A3(n3588), .ZN(n3593) );
  NAND4_X1 U4323 ( .A1(n3990), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3592)
         );
  NOR4_X1 U4324 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3613)
         );
  NOR4_X1 U4325 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3612)
         );
  NOR4_X1 U4326 ( .A1(n3908), .A2(n3638), .A3(n3600), .A4(n2533), .ZN(n3611)
         );
  AND2_X1 U4327 ( .A1(n3720), .A2(n3601), .ZN(n3622) );
  NOR2_X1 U4328 ( .A1(n3626), .A2(n3622), .ZN(n4464) );
  NAND2_X1 U4329 ( .A1(n3603), .A2(n3602), .ZN(n3799) );
  INV_X1 U4330 ( .A(n3799), .ZN(n3606) );
  NAND2_X1 U4331 ( .A1(n3830), .A2(n3604), .ZN(n3848) );
  INV_X1 U4332 ( .A(n3848), .ZN(n3605) );
  NAND4_X1 U4333 ( .A1(n4464), .A2(n3606), .A3(n2043), .A4(n3605), .ZN(n3609)
         );
  XNOR2_X1 U4334 ( .A(n3790), .B(n3607), .ZN(n3608) );
  NOR4_X1 U4335 ( .A1(n3609), .A2(n3797), .A3(n3810), .A4(n3608), .ZN(n3610)
         );
  NAND4_X1 U4336 ( .A1(n3613), .A2(n3612), .A3(n3611), .A4(n3610), .ZN(n3615)
         );
  MUX2_X1 U4337 ( .A(n3616), .B(n3615), .S(n3614), .Z(n3696) );
  INV_X1 U4338 ( .A(n3617), .ZN(n3662) );
  INV_X1 U4339 ( .A(n3618), .ZN(n3619) );
  OAI211_X1 U4340 ( .C1(n3621), .C2(n3662), .A(n3620), .B(n3619), .ZN(n3667)
         );
  INV_X1 U4341 ( .A(n3622), .ZN(n3624) );
  OAI211_X1 U4342 ( .C1(n3626), .C2(n3625), .A(n3624), .B(n3623), .ZN(n3628)
         );
  NAND3_X1 U4343 ( .A1(n3628), .A2(n3627), .A3(n2534), .ZN(n3631) );
  NAND3_X1 U4344 ( .A1(n3631), .A2(n3630), .A3(n3629), .ZN(n3634) );
  NAND3_X1 U4345 ( .A1(n3634), .A2(n3633), .A3(n3632), .ZN(n3637) );
  NAND4_X1 U4346 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3651), .ZN(n3641)
         );
  INV_X1 U4347 ( .A(n3638), .ZN(n3640) );
  NAND3_X1 U4348 ( .A1(n3641), .A2(n3640), .A3(n3639), .ZN(n3642) );
  NAND3_X1 U4349 ( .A1(n3642), .A2(n3648), .A3(n3652), .ZN(n3645) );
  NAND3_X1 U4350 ( .A1(n3645), .A2(n3644), .A3(n3643), .ZN(n3659) );
  NOR2_X1 U4351 ( .A1(n3647), .A2(n3646), .ZN(n3658) );
  INV_X1 U4352 ( .A(n3648), .ZN(n3650) );
  NOR2_X1 U4353 ( .A1(n3650), .A2(n3649), .ZN(n3654) );
  NAND4_X1 U4354 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3656)
         );
  NAND2_X1 U4355 ( .A1(n3656), .A2(n3655), .ZN(n3657) );
  AOI22_X1 U4356 ( .A1(n3659), .A2(n3658), .B1(n3668), .B2(n3657), .ZN(n3665)
         );
  INV_X1 U4357 ( .A(n3660), .ZN(n3664) );
  INV_X1 U4358 ( .A(n3661), .ZN(n3663) );
  NOR4_X1 U4359 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3666)
         );
  AOI21_X1 U4360 ( .B1(n3668), .B2(n3667), .A(n3666), .ZN(n3671) );
  OAI21_X1 U4361 ( .B1(n3671), .B2(n3670), .A(n3669), .ZN(n3673) );
  NAND2_X1 U4362 ( .A1(n3673), .A2(n3672), .ZN(n3675) );
  OAI221_X1 U4363 ( .B1(n3676), .B2(n3887), .C1(n3676), .C2(n3675), .A(n3674), 
        .ZN(n3677) );
  INV_X1 U4364 ( .A(n3677), .ZN(n3679) );
  AOI221_X1 U4365 ( .B1(n3681), .B2(n3680), .C1(n3681), .C2(n3679), .A(n3678), 
        .ZN(n3684) );
  OAI211_X1 U4366 ( .C1(n3685), .C2(n3684), .A(n3683), .B(n3682), .ZN(n3686)
         );
  INV_X1 U4367 ( .A(n3686), .ZN(n3693) );
  INV_X1 U4368 ( .A(n3687), .ZN(n3689) );
  OAI21_X1 U4369 ( .B1(n3690), .B2(n3689), .A(n3688), .ZN(n3691) );
  OAI21_X1 U4370 ( .B1(n3693), .B2(n3692), .A(n3691), .ZN(n3695) );
  MUX2_X1 U4371 ( .A(n3696), .B(n3695), .S(n3694), .Z(n3697) );
  XNOR2_X1 U4372 ( .A(n3697), .B(n3780), .ZN(n3704) );
  NAND2_X1 U4373 ( .A1(n3699), .A2(n3698), .ZN(n3700) );
  OAI211_X1 U4374 ( .C1(n3701), .C2(n3703), .A(n3700), .B(B_REG_SCAN_IN), .ZN(
        n3702) );
  OAI21_X1 U4375 ( .B1(n3704), .B2(n3703), .A(n3702), .ZN(U3239) );
  MUX2_X1 U4376 ( .A(n4057), .B(DATAO_REG_31__SCAN_IN), .S(n3719), .Z(U3581)
         );
  MUX2_X1 U4377 ( .A(n3790), .B(DATAO_REG_30__SCAN_IN), .S(n3719), .Z(U3580)
         );
  MUX2_X1 U4378 ( .A(n3705), .B(DATAO_REG_29__SCAN_IN), .S(n3719), .Z(U3579)
         );
  MUX2_X1 U4379 ( .A(n3820), .B(DATAO_REG_28__SCAN_IN), .S(n3719), .Z(U3578)
         );
  MUX2_X1 U4380 ( .A(n3836), .B(DATAO_REG_27__SCAN_IN), .S(n3716), .Z(U3577)
         );
  MUX2_X1 U4381 ( .A(n3852), .B(DATAO_REG_26__SCAN_IN), .S(n3719), .Z(U3576)
         );
  MUX2_X1 U4382 ( .A(n3895), .B(DATAO_REG_24__SCAN_IN), .S(n3719), .Z(U3574)
         );
  MUX2_X1 U4383 ( .A(n3869), .B(DATAO_REG_23__SCAN_IN), .S(n3716), .Z(U3573)
         );
  MUX2_X1 U4384 ( .A(n3706), .B(DATAO_REG_21__SCAN_IN), .S(n3719), .Z(U3571)
         );
  MUX2_X1 U4385 ( .A(n3969), .B(DATAO_REG_20__SCAN_IN), .S(n3719), .Z(U3570)
         );
  MUX2_X1 U4386 ( .A(n4011), .B(DATAO_REG_18__SCAN_IN), .S(n3716), .Z(U3568)
         );
  MUX2_X1 U4387 ( .A(n4023), .B(DATAO_REG_17__SCAN_IN), .S(n3719), .Z(U3567)
         );
  MUX2_X1 U4388 ( .A(n4041), .B(DATAO_REG_16__SCAN_IN), .S(n3719), .Z(U3566)
         );
  MUX2_X1 U4389 ( .A(DATAO_REG_15__SCAN_IN), .B(n4025), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4390 ( .A(n3707), .B(DATAO_REG_14__SCAN_IN), .S(n3716), .Z(U3564)
         );
  MUX2_X1 U4391 ( .A(n3708), .B(DATAO_REG_13__SCAN_IN), .S(n3719), .Z(U3563)
         );
  MUX2_X1 U4392 ( .A(DATAO_REG_12__SCAN_IN), .B(n3709), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4393 ( .A(n3710), .B(DATAO_REG_11__SCAN_IN), .S(n3719), .Z(U3561)
         );
  MUX2_X1 U4394 ( .A(n3711), .B(DATAO_REG_9__SCAN_IN), .S(n3716), .Z(U3559) );
  MUX2_X1 U4395 ( .A(DATAO_REG_8__SCAN_IN), .B(n3712), .S(U4043), .Z(U3558) );
  MUX2_X1 U4396 ( .A(n3713), .B(DATAO_REG_7__SCAN_IN), .S(n3719), .Z(U3557) );
  MUX2_X1 U4397 ( .A(n3714), .B(DATAO_REG_6__SCAN_IN), .S(n3716), .Z(U3556) );
  MUX2_X1 U4398 ( .A(DATAO_REG_5__SCAN_IN), .B(n3715), .S(U4043), .Z(U3555) );
  MUX2_X1 U4399 ( .A(n3717), .B(DATAO_REG_4__SCAN_IN), .S(n3716), .Z(U3554) );
  MUX2_X1 U4400 ( .A(n3718), .B(DATAO_REG_3__SCAN_IN), .S(n3719), .Z(U3553) );
  MUX2_X1 U4401 ( .A(n2273), .B(DATAO_REG_2__SCAN_IN), .S(n3719), .Z(U3552) );
  MUX2_X1 U4402 ( .A(n3720), .B(DATAO_REG_0__SCAN_IN), .S(n3719), .Z(U3550) );
  OAI211_X1 U4403 ( .C1(n3723), .C2(n3722), .A(n4435), .B(n3721), .ZN(n3730)
         );
  OAI211_X1 U4404 ( .C1(n3726), .C2(n2669), .A(n4437), .B(n3725), .ZN(n3729)
         );
  AOI22_X1 U4405 ( .A1(n4427), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3728) );
  NAND2_X1 U4406 ( .A1(n4450), .A2(n4333), .ZN(n3727) );
  NAND4_X1 U4407 ( .A1(n3730), .A2(n3729), .A3(n3728), .A4(n3727), .ZN(U3241)
         );
  XNOR2_X1 U4408 ( .A(n3749), .B(REG2_REG_17__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U4409 ( .A1(n4498), .A2(REG2_REG_11__SCAN_IN), .ZN(n3735) );
  INV_X1 U4410 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4411 ( .A1(n4498), .A2(REG2_REG_11__SCAN_IN), .B1(n3731), .B2(
        n4382), .ZN(n4379) );
  NAND2_X1 U4412 ( .A1(n3732), .A2(n4331), .ZN(n3734) );
  NAND2_X1 U4413 ( .A1(n3734), .A2(n3733), .ZN(n4378) );
  NAND2_X1 U4414 ( .A1(n4379), .A2(n4378), .ZN(n4377) );
  NAND2_X1 U4415 ( .A1(n3753), .A2(n3736), .ZN(n3737) );
  AND2_X1 U4416 ( .A1(n4398), .A2(REG2_REG_13__SCAN_IN), .ZN(n3739) );
  NOR2_X1 U4417 ( .A1(n3757), .A2(n3740), .ZN(n3741) );
  INV_X1 U4418 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4409) );
  INV_X1 U4419 ( .A(n3759), .ZN(n4492) );
  INV_X1 U4420 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4421 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4492), .B1(n3759), .B2(
        n3742), .ZN(n4416) );
  NAND2_X1 U4422 ( .A1(n3743), .A2(n4490), .ZN(n3744) );
  XOR2_X1 U4423 ( .A(n3743), .B(n4490), .Z(n4430) );
  INV_X1 U4424 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4429) );
  NAND2_X1 U4425 ( .A1(n4430), .A2(n4429), .ZN(n4428) );
  NAND2_X1 U4426 ( .A1(n3744), .A2(n4428), .ZN(n3745) );
  OAI21_X1 U4427 ( .B1(n3746), .B2(n3745), .A(n3773), .ZN(n3747) );
  AOI22_X1 U4428 ( .A1(n3774), .A2(n4450), .B1(n4437), .B2(n3747), .ZN(n3767)
         );
  AOI21_X1 U4429 ( .B1(n4427), .B2(ADDR_REG_17__SCAN_IN), .A(n3748), .ZN(n3766) );
  XNOR2_X1 U4430 ( .A(n3749), .B(REG1_REG_17__SCAN_IN), .ZN(n3763) );
  INV_X1 U4431 ( .A(n3750), .ZN(n3752) );
  INV_X1 U4432 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U4433 ( .A1(n4498), .A2(n4565), .B1(REG1_REG_11__SCAN_IN), .B2(
        n4382), .ZN(n4373) );
  NOR2_X1 U4434 ( .A1(n4374), .A2(n4373), .ZN(n4372) );
  NOR2_X1 U4435 ( .A1(n3754), .A2(n2093), .ZN(n3755) );
  INV_X1 U4436 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4385) );
  INV_X1 U4437 ( .A(n4398), .ZN(n4496) );
  INV_X1 U4438 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4266) );
  AOI22_X1 U4439 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4496), .B1(n4398), .B2(
        n4266), .ZN(n4394) );
  NOR2_X1 U4440 ( .A1(n3756), .A2(n3757), .ZN(n3758) );
  INV_X1 U4441 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4406) );
  XNOR2_X1 U4442 ( .A(n3757), .B(n3756), .ZN(n4405) );
  NOR2_X1 U4443 ( .A1(n4406), .A2(n4405), .ZN(n4404) );
  INV_X1 U4444 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U4445 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4492), .B1(n3759), .B2(
        n4221), .ZN(n4421) );
  NAND2_X1 U4446 ( .A1(n3760), .A2(n4490), .ZN(n3761) );
  INV_X1 U4447 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4432) );
  NAND2_X1 U4448 ( .A1(n4433), .A2(n4432), .ZN(n4431) );
  NAND2_X1 U4449 ( .A1(n3761), .A2(n4431), .ZN(n3762) );
  OAI21_X1 U4450 ( .B1(n3763), .B2(n3762), .A(n3768), .ZN(n3764) );
  NAND2_X1 U4451 ( .A1(n4435), .A2(n3764), .ZN(n3765) );
  NAND3_X1 U4452 ( .A1(n3767), .A2(n3766), .A3(n3765), .ZN(U3257) );
  INV_X1 U4453 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4244) );
  AOI22_X1 U4454 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4488), .B1(n4449), .B2(
        n4244), .ZN(n4444) );
  XNOR2_X1 U4455 ( .A(n3769), .B(REG1_REG_19__SCAN_IN), .ZN(n3770) );
  XNOR2_X1 U4456 ( .A(n3771), .B(n3770), .ZN(n3784) );
  NAND2_X1 U4457 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4449), .ZN(n3772) );
  OAI21_X1 U4458 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4449), .A(n3772), .ZN(n4447) );
  INV_X1 U4459 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3775) );
  MUX2_X1 U4460 ( .A(n3775), .B(REG2_REG_19__SCAN_IN), .S(n3780), .Z(n3776) );
  XNOR2_X1 U4461 ( .A(n3777), .B(n3776), .ZN(n3782) );
  AOI21_X1 U4462 ( .B1(n4427), .B2(ADDR_REG_19__SCAN_IN), .A(n3778), .ZN(n3779) );
  OAI21_X1 U4463 ( .B1(n4440), .B2(n3780), .A(n3779), .ZN(n3781) );
  OAI21_X1 U4464 ( .B1(n3784), .B2(n4441), .A(n3783), .ZN(U3259) );
  OAI21_X1 U4465 ( .B1(n3787), .B2(n3786), .A(n3785), .ZN(n3788) );
  NAND2_X1 U4466 ( .A1(n3820), .A2(n4024), .ZN(n3792) );
  AND2_X1 U4467 ( .A1(n4327), .A2(B_REG_SCAN_IN), .ZN(n3789) );
  NOR2_X1 U4468 ( .A1(n3946), .A2(n3789), .ZN(n4056) );
  NAND2_X1 U4469 ( .A1(n3790), .A2(n4056), .ZN(n3791) );
  OAI211_X1 U4470 ( .C1(n3803), .C2(n4029), .A(n3792), .B(n3791), .ZN(n3793)
         );
  INV_X1 U4471 ( .A(n4070), .ZN(n3794) );
  AOI21_X1 U4472 ( .B1(n3795), .B2(n4453), .A(n3794), .ZN(n3808) );
  AOI22_X1 U4473 ( .A1(n3798), .A2(n3797), .B1(n3796), .B2(n3820), .ZN(n3800)
         );
  XNOR2_X1 U4474 ( .A(n3800), .B(n3799), .ZN(n4068) );
  NAND2_X1 U4475 ( .A1(n4068), .A2(n3999), .ZN(n3807) );
  INV_X1 U4476 ( .A(n3802), .ZN(n3804) );
  INV_X1 U4477 ( .A(n3803), .ZN(n3801) );
  INV_X1 U4478 ( .A(n4069), .ZN(n3805) );
  AOI22_X1 U4479 ( .A1(n3805), .A2(n4458), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4463), .ZN(n3806) );
  OAI211_X1 U4480 ( .C1(n4463), .C2(n3808), .A(n3807), .B(n3806), .ZN(U3354)
         );
  XNOR2_X1 U4481 ( .A(n3809), .B(n3810), .ZN(n4075) );
  AND2_X1 U4482 ( .A1(n3840), .A2(n3811), .ZN(n3812) );
  NOR2_X1 U4483 ( .A1(n3813), .A2(n3812), .ZN(n4072) );
  INV_X1 U4484 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3816) );
  INV_X1 U4485 ( .A(n3814), .ZN(n3815) );
  OAI22_X1 U4486 ( .A1(n4470), .A2(n3816), .B1(n3815), .B2(n4476), .ZN(n3817)
         );
  AOI21_X1 U4487 ( .B1(n4072), .B2(n4458), .A(n3817), .ZN(n3827) );
  XNOR2_X1 U4488 ( .A(n3819), .B(n3818), .ZN(n3825) );
  NAND2_X1 U4489 ( .A1(n3852), .A2(n4024), .ZN(n3822) );
  NAND2_X1 U4490 ( .A1(n3820), .A2(n4272), .ZN(n3821) );
  OAI211_X1 U4491 ( .C1(n4029), .C2(n3823), .A(n3822), .B(n3821), .ZN(n3824)
         );
  AOI21_X1 U4492 ( .B1(n3825), .B2(n4040), .A(n3824), .ZN(n4074) );
  OR2_X1 U4493 ( .A1(n4074), .A2(n4463), .ZN(n3826) );
  OAI211_X1 U4494 ( .C1(n4075), .C2(n4054), .A(n3827), .B(n3826), .ZN(U3263)
         );
  XNOR2_X1 U4495 ( .A(n3829), .B(n3828), .ZN(n4077) );
  INV_X1 U4496 ( .A(n4077), .ZN(n3846) );
  NAND2_X1 U4497 ( .A1(n3831), .A2(n3830), .ZN(n3833) );
  XNOR2_X1 U4498 ( .A(n3833), .B(n3832), .ZN(n3834) );
  NAND2_X1 U4499 ( .A1(n3834), .A2(n4040), .ZN(n3838) );
  NOR2_X1 U4500 ( .A1(n4029), .A2(n3841), .ZN(n3835) );
  AOI21_X1 U4501 ( .B1(n3836), .B2(n4272), .A(n3835), .ZN(n3837) );
  OAI211_X1 U4502 ( .C1(n3839), .C2(n4044), .A(n3838), .B(n3837), .ZN(n4076)
         );
  OAI21_X1 U4503 ( .B1(n2085), .B2(n3841), .A(n3840), .ZN(n4290) );
  AOI22_X1 U4504 ( .A1(n4463), .A2(REG2_REG_26__SCAN_IN), .B1(n3842), .B2(
        n4453), .ZN(n3843) );
  OAI21_X1 U4505 ( .B1(n4290), .B2(n4050), .A(n3843), .ZN(n3844) );
  AOI21_X1 U4506 ( .B1(n4076), .B2(n4470), .A(n3844), .ZN(n3845) );
  OAI21_X1 U4507 ( .B1(n3846), .B2(n4054), .A(n3845), .ZN(U3264) );
  XOR2_X1 U4508 ( .A(n3848), .B(n3847), .Z(n4080) );
  INV_X1 U4509 ( .A(n4080), .ZN(n3863) );
  XNOR2_X1 U4510 ( .A(n3849), .B(n3848), .ZN(n3850) );
  NAND2_X1 U4511 ( .A1(n3850), .A2(n4040), .ZN(n3854) );
  NOR2_X1 U4512 ( .A1(n4029), .A2(n3857), .ZN(n3851) );
  AOI21_X1 U4513 ( .B1(n3852), .B2(n4272), .A(n3851), .ZN(n3853) );
  OAI211_X1 U4514 ( .C1(n3855), .C2(n4044), .A(n3854), .B(n3853), .ZN(n4079)
         );
  INV_X1 U4515 ( .A(n3875), .ZN(n3858) );
  OAI21_X1 U4516 ( .B1(n3858), .B2(n3857), .A(n3856), .ZN(n4294) );
  AOI22_X1 U4517 ( .A1(n4463), .A2(REG2_REG_25__SCAN_IN), .B1(n3859), .B2(
        n4453), .ZN(n3860) );
  OAI21_X1 U4518 ( .B1(n4294), .B2(n4050), .A(n3860), .ZN(n3861) );
  AOI21_X1 U4519 ( .B1(n4079), .B2(n4470), .A(n3861), .ZN(n3862) );
  OAI21_X1 U4520 ( .B1(n3863), .B2(n4054), .A(n3862), .ZN(U3265) );
  XOR2_X1 U4521 ( .A(n3866), .B(n2026), .Z(n4084) );
  NAND2_X1 U4522 ( .A1(n3865), .A2(n3864), .ZN(n3868) );
  INV_X1 U4523 ( .A(n3866), .ZN(n3867) );
  XNOR2_X1 U4524 ( .A(n3868), .B(n3867), .ZN(n3874) );
  NAND2_X1 U4525 ( .A1(n3869), .A2(n4024), .ZN(n3872) );
  NAND2_X1 U4526 ( .A1(n3870), .A2(n4272), .ZN(n3871) );
  OAI211_X1 U4527 ( .C1(n4029), .C2(n3876), .A(n3872), .B(n3871), .ZN(n3873)
         );
  AOI21_X1 U4528 ( .B1(n3874), .B2(n4040), .A(n3873), .ZN(n4083) );
  INV_X1 U4529 ( .A(n4083), .ZN(n3880) );
  OAI21_X1 U4530 ( .B1(n3899), .B2(n3876), .A(n3875), .ZN(n4299) );
  AOI22_X1 U4531 ( .A1(n4463), .A2(REG2_REG_24__SCAN_IN), .B1(n3877), .B2(
        n4453), .ZN(n3878) );
  OAI21_X1 U4532 ( .B1(n4299), .B2(n4050), .A(n3878), .ZN(n3879) );
  AOI21_X1 U4533 ( .B1(n3880), .B2(n4470), .A(n3879), .ZN(n3881) );
  OAI21_X1 U4534 ( .B1(n4084), .B2(n4054), .A(n3881), .ZN(U3266) );
  INV_X1 U4535 ( .A(n3884), .ZN(n3885) );
  INV_X1 U4536 ( .A(n3886), .ZN(n3888) );
  OAI21_X1 U4537 ( .B1(n3909), .B2(n3908), .A(n3890), .ZN(n3891) );
  XOR2_X1 U4538 ( .A(n3892), .B(n3891), .Z(n3893) );
  NAND2_X1 U4539 ( .A1(n3893), .A2(n4040), .ZN(n3897) );
  NOR2_X1 U4540 ( .A1(n4029), .A2(n3901), .ZN(n3894) );
  AOI21_X1 U4541 ( .B1(n3895), .B2(n4272), .A(n3894), .ZN(n3896) );
  INV_X1 U4542 ( .A(n3899), .ZN(n3900) );
  OAI21_X1 U4543 ( .B1(n3916), .B2(n3901), .A(n3900), .ZN(n4303) );
  AOI22_X1 U4544 ( .A1(n4463), .A2(REG2_REG_23__SCAN_IN), .B1(n3902), .B2(
        n4453), .ZN(n3903) );
  OAI21_X1 U4545 ( .B1(n4303), .B2(n4050), .A(n3903), .ZN(n3904) );
  AOI21_X1 U4546 ( .B1(n4087), .B2(n4470), .A(n3904), .ZN(n3905) );
  OAI21_X1 U4547 ( .B1(n2008), .B2(n4054), .A(n3905), .ZN(U3267) );
  OAI21_X1 U4548 ( .B1(n3906), .B2(n3908), .A(n3907), .ZN(n4092) );
  XNOR2_X1 U4549 ( .A(n3909), .B(n3908), .ZN(n3914) );
  NOR2_X1 U4550 ( .A1(n3947), .A2(n4044), .ZN(n3913) );
  OAI22_X1 U4551 ( .A1(n3911), .A2(n3946), .B1(n3910), .B2(n4029), .ZN(n3912)
         );
  AOI211_X1 U4552 ( .C1(n3914), .C2(n4040), .A(n3913), .B(n3912), .ZN(n4091)
         );
  AOI22_X1 U4553 ( .A1(n4463), .A2(REG2_REG_22__SCAN_IN), .B1(n3915), .B2(
        n4453), .ZN(n3919) );
  INV_X1 U4554 ( .A(n3916), .ZN(n4089) );
  NAND2_X1 U4555 ( .A1(n3931), .A2(n3917), .ZN(n4088) );
  NAND3_X1 U4556 ( .A1(n4089), .A2(n4458), .A3(n4088), .ZN(n3918) );
  OAI211_X1 U4557 ( .C1(n4091), .C2(n4463), .A(n3919), .B(n3918), .ZN(n3920)
         );
  INV_X1 U4558 ( .A(n3920), .ZN(n3921) );
  OAI21_X1 U4559 ( .B1(n4092), .B2(n4054), .A(n3921), .ZN(U3268) );
  XNOR2_X1 U4560 ( .A(n3922), .B(n3923), .ZN(n4093) );
  XNOR2_X1 U4561 ( .A(n3924), .B(n3923), .ZN(n3930) );
  NAND2_X1 U4562 ( .A1(n3969), .A2(n4024), .ZN(n3928) );
  NOR2_X1 U4563 ( .A1(n4029), .A2(n3932), .ZN(n3925) );
  AOI21_X1 U4564 ( .B1(n3926), .B2(n4272), .A(n3925), .ZN(n3927) );
  NAND2_X1 U4565 ( .A1(n3928), .A2(n3927), .ZN(n3929) );
  AOI21_X1 U4566 ( .B1(n3930), .B2(n4040), .A(n3929), .ZN(n4094) );
  NOR2_X1 U4567 ( .A1(n4094), .A2(n4463), .ZN(n3937) );
  INV_X1 U4568 ( .A(n3952), .ZN(n3933) );
  OAI21_X1 U4569 ( .B1(n3933), .B2(n3932), .A(n3931), .ZN(n4096) );
  AOI22_X1 U4570 ( .A1(n4463), .A2(REG2_REG_21__SCAN_IN), .B1(n3934), .B2(
        n4453), .ZN(n3935) );
  OAI21_X1 U4571 ( .B1(n4096), .B2(n4050), .A(n3935), .ZN(n3936) );
  AOI211_X1 U4572 ( .C1(n4093), .C2(n3999), .A(n3937), .B(n3936), .ZN(n3938)
         );
  INV_X1 U4573 ( .A(n3938), .ZN(U3269) );
  XNOR2_X1 U4574 ( .A(n3939), .B(n3942), .ZN(n3951) );
  NAND2_X1 U4575 ( .A1(n3941), .A2(n3940), .ZN(n3943) );
  XNOR2_X1 U4576 ( .A(n3943), .B(n3942), .ZN(n3949) );
  AOI22_X1 U4577 ( .A1(n3983), .A2(n4024), .B1(n3944), .B2(n4064), .ZN(n3945)
         );
  OAI21_X1 U4578 ( .B1(n3947), .B2(n3946), .A(n3945), .ZN(n3948) );
  AOI21_X1 U4579 ( .B1(n3949), .B2(n4040), .A(n3948), .ZN(n3950) );
  OAI21_X1 U4580 ( .B1(n3951), .B2(n4270), .A(n3950), .ZN(n4097) );
  INV_X1 U4581 ( .A(n4097), .ZN(n3958) );
  INV_X1 U4582 ( .A(n3951), .ZN(n4098) );
  OAI21_X1 U4583 ( .B1(n3976), .B2(n3953), .A(n3952), .ZN(n4309) );
  AOI22_X1 U4584 ( .A1(n4463), .A2(REG2_REG_20__SCAN_IN), .B1(n3954), .B2(
        n4453), .ZN(n3955) );
  OAI21_X1 U4585 ( .B1(n4309), .B2(n4050), .A(n3955), .ZN(n3956) );
  AOI21_X1 U4586 ( .B1(n4098), .B2(n4466), .A(n3956), .ZN(n3957) );
  OAI21_X1 U4587 ( .B1(n3958), .B2(n4463), .A(n3957), .ZN(U3270) );
  XOR2_X1 U4588 ( .A(n3965), .B(n3959), .Z(n4101) );
  INV_X1 U4589 ( .A(n4101), .ZN(n3981) );
  NAND2_X1 U4590 ( .A1(n3961), .A2(n3960), .ZN(n3982) );
  INV_X1 U4591 ( .A(n3962), .ZN(n3964) );
  OAI21_X1 U4592 ( .B1(n3982), .B2(n3964), .A(n3963), .ZN(n3966) );
  XNOR2_X1 U4593 ( .A(n3966), .B(n3965), .ZN(n3967) );
  NAND2_X1 U4594 ( .A1(n3967), .A2(n4040), .ZN(n3971) );
  NOR2_X1 U4595 ( .A1(n3973), .A2(n4029), .ZN(n3968) );
  AOI21_X1 U4596 ( .B1(n3969), .B2(n4272), .A(n3968), .ZN(n3970) );
  OAI211_X1 U4597 ( .C1(n3972), .C2(n4044), .A(n3971), .B(n3970), .ZN(n4100)
         );
  AOI21_X1 U4598 ( .B1(n4003), .B2(n3974), .A(n3973), .ZN(n3975) );
  OR2_X1 U4599 ( .A1(n3976), .A2(n3975), .ZN(n4313) );
  AOI22_X1 U4600 ( .A1(n4463), .A2(REG2_REG_19__SCAN_IN), .B1(n3977), .B2(
        n4453), .ZN(n3978) );
  OAI21_X1 U4601 ( .B1(n4313), .B2(n4050), .A(n3978), .ZN(n3979) );
  AOI21_X1 U4602 ( .B1(n4100), .B2(n4470), .A(n3979), .ZN(n3980) );
  OAI21_X1 U4603 ( .B1(n3981), .B2(n4054), .A(n3980), .ZN(U3271) );
  XNOR2_X1 U4604 ( .A(n3982), .B(n3990), .ZN(n3987) );
  AOI22_X1 U4605 ( .A1(n3983), .A2(n4272), .B1(n4064), .B2(n3991), .ZN(n3984)
         );
  OAI21_X1 U4606 ( .B1(n3985), .B2(n4044), .A(n3984), .ZN(n3986) );
  AOI21_X1 U4607 ( .B1(n3987), .B2(n4040), .A(n3986), .ZN(n4105) );
  AOI21_X1 U4608 ( .B1(n3990), .B2(n3989), .A(n3988), .ZN(n4106) );
  INV_X1 U4609 ( .A(n4106), .ZN(n4000) );
  XNOR2_X1 U4610 ( .A(n4003), .B(n3991), .ZN(n3992) );
  NAND2_X1 U4611 ( .A1(n3992), .A2(n4545), .ZN(n4104) );
  NOR2_X1 U4612 ( .A1(n4104), .A2(n3993), .ZN(n3998) );
  INV_X1 U4613 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3996) );
  INV_X1 U4614 ( .A(n3994), .ZN(n3995) );
  OAI22_X1 U4615 ( .A1(n4470), .A2(n3996), .B1(n3995), .B2(n4476), .ZN(n3997)
         );
  AOI211_X1 U4616 ( .C1(n4000), .C2(n3999), .A(n3998), .B(n3997), .ZN(n4001)
         );
  OAI21_X1 U4617 ( .B1(n4463), .B2(n4105), .A(n4001), .ZN(U3272) );
  XNOR2_X1 U4618 ( .A(n4002), .B(n4007), .ZN(n4110) );
  AOI21_X1 U4619 ( .B1(n4010), .B2(n4030), .A(n4003), .ZN(n4108) );
  INV_X1 U4620 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4005) );
  OAI22_X1 U4621 ( .A1(n4470), .A2(n4005), .B1(n4004), .B2(n4476), .ZN(n4006)
         );
  AOI21_X1 U4622 ( .B1(n4108), .B2(n4458), .A(n4006), .ZN(n4016) );
  XNOR2_X1 U4623 ( .A(n4008), .B(n4007), .ZN(n4009) );
  NAND2_X1 U4624 ( .A1(n4009), .A2(n4040), .ZN(n4013) );
  AOI22_X1 U4625 ( .A1(n4011), .A2(n4272), .B1(n4064), .B2(n4010), .ZN(n4012)
         );
  OAI211_X1 U4626 ( .C1(n4014), .C2(n4044), .A(n4013), .B(n4012), .ZN(n4107)
         );
  NAND2_X1 U4627 ( .A1(n4107), .A2(n4470), .ZN(n4015) );
  OAI211_X1 U4628 ( .C1(n4110), .C2(n4054), .A(n4016), .B(n4015), .ZN(U3273)
         );
  OAI21_X1 U4629 ( .B1(n4019), .B2(n4018), .A(n4017), .ZN(n4256) );
  OAI211_X1 U4630 ( .C1(n4022), .C2(n4021), .A(n4020), .B(n4040), .ZN(n4027)
         );
  AOI22_X1 U4631 ( .A1(n4025), .A2(n4024), .B1(n4272), .B2(n4023), .ZN(n4026)
         );
  OAI211_X1 U4632 ( .C1(n4029), .C2(n4028), .A(n4027), .B(n4026), .ZN(n4253)
         );
  INV_X1 U4633 ( .A(n4030), .ZN(n4031) );
  AOI21_X1 U4634 ( .B1(n2433), .B2(n4032), .A(n4031), .ZN(n4254) );
  INV_X1 U4635 ( .A(n4254), .ZN(n4035) );
  AOI22_X1 U4636 ( .A1(n4463), .A2(REG2_REG_16__SCAN_IN), .B1(n4033), .B2(
        n4453), .ZN(n4034) );
  OAI21_X1 U4637 ( .B1(n4035), .B2(n4050), .A(n4034), .ZN(n4036) );
  AOI21_X1 U4638 ( .B1(n4253), .B2(n4470), .A(n4036), .ZN(n4037) );
  OAI21_X1 U4639 ( .B1(n4256), .B2(n4054), .A(n4037), .ZN(U3274) );
  XNOR2_X1 U4640 ( .A(n4038), .B(n2043), .ZN(n4260) );
  OAI211_X1 U4641 ( .C1(n2037), .C2(n2043), .A(n4040), .B(n4039), .ZN(n4043)
         );
  AOI22_X1 U4642 ( .A1(n4041), .A2(n4272), .B1(n4064), .B2(n4046), .ZN(n4042)
         );
  OAI211_X1 U4643 ( .C1(n4045), .C2(n4044), .A(n4043), .B(n4042), .ZN(n4257)
         );
  XNOR2_X1 U4644 ( .A(n4047), .B(n4046), .ZN(n4258) );
  INV_X1 U4645 ( .A(n4258), .ZN(n4051) );
  AOI22_X1 U4646 ( .A1(n4463), .A2(REG2_REG_15__SCAN_IN), .B1(n4048), .B2(
        n4453), .ZN(n4049) );
  OAI21_X1 U4647 ( .B1(n4051), .B2(n4050), .A(n4049), .ZN(n4052) );
  AOI21_X1 U4648 ( .B1(n4257), .B2(n4470), .A(n4052), .ZN(n4053) );
  OAI21_X1 U4649 ( .B1(n4260), .B2(n4054), .A(n4053), .ZN(U3275) );
  XOR2_X1 U4650 ( .A(n4055), .B(n4061), .Z(n4336) );
  INV_X1 U4651 ( .A(n4336), .ZN(n4281) );
  INV_X1 U4652 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4059) );
  INV_X1 U4653 ( .A(n4055), .ZN(n4058) );
  AND2_X1 U4654 ( .A1(n4057), .A2(n4056), .ZN(n4063) );
  AOI21_X1 U4655 ( .B1(n4058), .B2(n4064), .A(n4063), .ZN(n4338) );
  MUX2_X1 U4656 ( .A(n4059), .B(n4338), .S(n4567), .Z(n4060) );
  OAI21_X1 U4657 ( .B1(n4281), .B2(n4268), .A(n4060), .ZN(U3549) );
  AOI21_X1 U4658 ( .B1(n4065), .B2(n4062), .A(n4061), .ZN(n4339) );
  INV_X1 U4659 ( .A(n4339), .ZN(n4284) );
  INV_X1 U4660 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4066) );
  AOI21_X1 U4661 ( .B1(n4065), .B2(n4064), .A(n4063), .ZN(n4341) );
  MUX2_X1 U4662 ( .A(n4066), .B(n4341), .S(n4567), .Z(n4067) );
  OAI21_X1 U4663 ( .B1(n4284), .B2(n4268), .A(n4067), .ZN(U3548) );
  NAND2_X1 U4664 ( .A1(n4068), .A2(n4533), .ZN(n4071) );
  MUX2_X1 U4665 ( .A(REG1_REG_29__SCAN_IN), .B(n4285), .S(n4567), .Z(U3547) );
  NAND2_X1 U4666 ( .A1(n4072), .A2(n4545), .ZN(n4073) );
  OAI211_X1 U4667 ( .C1(n4075), .C2(n4540), .A(n4074), .B(n4073), .ZN(n4286)
         );
  MUX2_X1 U4668 ( .A(REG1_REG_27__SCAN_IN), .B(n4286), .S(n4567), .Z(U3545) );
  INV_X1 U4669 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4124) );
  AOI21_X1 U4670 ( .B1(n4077), .B2(n4533), .A(n4076), .ZN(n4287) );
  MUX2_X1 U4671 ( .A(n4124), .B(n4287), .S(n4567), .Z(n4078) );
  OAI21_X1 U4672 ( .B1(n4268), .B2(n4290), .A(n4078), .ZN(U3544) );
  INV_X1 U4673 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4081) );
  AOI21_X1 U4674 ( .B1(n4080), .B2(n4533), .A(n4079), .ZN(n4291) );
  MUX2_X1 U4675 ( .A(n4081), .B(n4291), .S(n4567), .Z(n4082) );
  OAI21_X1 U4676 ( .B1(n4268), .B2(n4294), .A(n4082), .ZN(U3543) );
  OAI21_X1 U4677 ( .B1(n4084), .B2(n4540), .A(n4083), .ZN(n4295) );
  MUX2_X1 U4678 ( .A(REG1_REG_24__SCAN_IN), .B(n4295), .S(n4567), .Z(n4085) );
  INV_X1 U4679 ( .A(n4085), .ZN(n4086) );
  OAI21_X1 U4680 ( .B1(n4268), .B2(n4299), .A(n4086), .ZN(U3542) );
  INV_X1 U4681 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4191) );
  NAND3_X1 U4682 ( .A1(n4089), .A2(n4545), .A3(n4088), .ZN(n4090) );
  OAI211_X1 U4683 ( .C1(n4092), .C2(n4540), .A(n4091), .B(n4090), .ZN(n4304)
         );
  MUX2_X1 U4684 ( .A(REG1_REG_22__SCAN_IN), .B(n4304), .S(n4567), .Z(U3540) );
  NAND2_X1 U4685 ( .A1(n4093), .A2(n4533), .ZN(n4095) );
  OAI211_X1 U4686 ( .C1(n4548), .C2(n4096), .A(n4095), .B(n4094), .ZN(n4305)
         );
  MUX2_X1 U4687 ( .A(REG1_REG_21__SCAN_IN), .B(n4305), .S(n4567), .Z(U3539) );
  INV_X1 U4688 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4192) );
  AOI21_X1 U4689 ( .B1(n4524), .B2(n4098), .A(n4097), .ZN(n4306) );
  MUX2_X1 U4690 ( .A(n4192), .B(n4306), .S(n4567), .Z(n4099) );
  OAI21_X1 U4691 ( .B1(n4268), .B2(n4309), .A(n4099), .ZN(U3538) );
  INV_X1 U4692 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4102) );
  AOI21_X1 U4693 ( .B1(n4101), .B2(n4533), .A(n4100), .ZN(n4310) );
  MUX2_X1 U4694 ( .A(n4102), .B(n4310), .S(n4567), .Z(n4103) );
  OAI21_X1 U4695 ( .B1(n4268), .B2(n4313), .A(n4103), .ZN(U3537) );
  OAI211_X1 U4696 ( .C1(n4106), .C2(n4540), .A(n4105), .B(n4104), .ZN(n4314)
         );
  MUX2_X1 U4697 ( .A(REG1_REG_18__SCAN_IN), .B(n4314), .S(n4567), .Z(U3536) );
  AOI21_X1 U4698 ( .B1(n4545), .B2(n4108), .A(n4107), .ZN(n4109) );
  OAI21_X1 U4699 ( .B1(n4110), .B2(n4540), .A(n4109), .ZN(n4315) );
  MUX2_X1 U4700 ( .A(REG1_REG_17__SCAN_IN), .B(n4315), .S(n4567), .Z(n4252) );
  INV_X1 U4701 ( .A(D_REG_21__SCAN_IN), .ZN(n4477) );
  INV_X1 U4702 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4514) );
  AOI22_X1 U4703 ( .A1(n4477), .A2(keyinput17), .B1(keyinput26), .B2(n4514), 
        .ZN(n4111) );
  OAI221_X1 U4704 ( .B1(n4477), .B2(keyinput17), .C1(n4514), .C2(keyinput26), 
        .A(n4111), .ZN(n4120) );
  INV_X1 U4705 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4532) );
  INV_X1 U4706 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4707 ( .A1(n4532), .A2(keyinput49), .B1(n4113), .B2(keyinput46), 
        .ZN(n4112) );
  OAI221_X1 U4708 ( .B1(n4532), .B2(keyinput49), .C1(n4113), .C2(keyinput46), 
        .A(n4112), .ZN(n4119) );
  INV_X1 U4709 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4319) );
  INV_X1 U4710 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U4711 ( .A1(n4319), .A2(keyinput13), .B1(n4115), .B2(keyinput10), 
        .ZN(n4114) );
  OAI221_X1 U4712 ( .B1(n4319), .B2(keyinput13), .C1(n4115), .C2(keyinput10), 
        .A(n4114), .ZN(n4118) );
  INV_X1 U4713 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4307) );
  INV_X1 U4714 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U4715 ( .A1(n4307), .A2(keyinput29), .B1(keyinput36), .B2(n4297), 
        .ZN(n4116) );
  OAI221_X1 U4716 ( .B1(n4307), .B2(keyinput29), .C1(n4297), .C2(keyinput36), 
        .A(n4116), .ZN(n4117) );
  NOR4_X1 U4717 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4171)
         );
  INV_X1 U4718 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U4719 ( .A1(n4122), .A2(keyinput11), .B1(n2667), .B2(keyinput35), 
        .ZN(n4121) );
  OAI221_X1 U4720 ( .B1(n4122), .B2(keyinput11), .C1(n2667), .C2(keyinput35), 
        .A(n4121), .ZN(n4130) );
  INV_X1 U4721 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U4722 ( .A1(n4213), .A2(keyinput31), .B1(n4124), .B2(keyinput50), 
        .ZN(n4123) );
  OAI221_X1 U4723 ( .B1(n4213), .B2(keyinput31), .C1(n4124), .C2(keyinput50), 
        .A(n4123), .ZN(n4129) );
  XNOR2_X1 U4724 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput57), .ZN(n4127) );
  XNOR2_X1 U4725 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput16), .ZN(n4126) );
  XNOR2_X1 U4726 ( .A(keyinput40), .B(IR_REG_24__SCAN_IN), .ZN(n4125) );
  NAND3_X1 U4727 ( .A1(n4127), .A2(n4126), .A3(n4125), .ZN(n4128) );
  NOR3_X1 U4728 ( .A1(n4130), .A2(n4129), .A3(n4128), .ZN(n4170) );
  INV_X1 U4729 ( .A(D_REG_4__SCAN_IN), .ZN(n4482) );
  AOI22_X1 U4730 ( .A1(n4132), .A2(keyinput28), .B1(n4482), .B2(keyinput37), 
        .ZN(n4131) );
  OAI221_X1 U4731 ( .B1(n4132), .B2(keyinput28), .C1(n4482), .C2(keyinput37), 
        .A(n4131), .ZN(n4139) );
  INV_X1 U4732 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n4212) );
  XNOR2_X1 U4733 ( .A(n4212), .B(keyinput23), .ZN(n4138) );
  XNOR2_X1 U4734 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput2), .ZN(n4136) );
  XNOR2_X1 U4735 ( .A(IR_REG_2__SCAN_IN), .B(keyinput30), .ZN(n4135) );
  XNOR2_X1 U4736 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput12), .ZN(n4134) );
  XNOR2_X1 U4737 ( .A(keyinput44), .B(IR_REG_16__SCAN_IN), .ZN(n4133) );
  NAND4_X1 U4738 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4137)
         );
  NOR3_X1 U4739 ( .A1(n4139), .A2(n4138), .A3(n4137), .ZN(n4154) );
  AOI22_X1 U4740 ( .A1(n4142), .A2(keyinput52), .B1(keyinput61), .B2(n4141), 
        .ZN(n4140) );
  OAI221_X1 U4741 ( .B1(n4142), .B2(keyinput52), .C1(n4141), .C2(keyinput61), 
        .A(n4140), .ZN(n4147) );
  AOI22_X1 U4742 ( .A1(n4145), .A2(keyinput27), .B1(keyinput39), .B2(n4144), 
        .ZN(n4143) );
  OAI221_X1 U4743 ( .B1(n4145), .B2(keyinput27), .C1(n4144), .C2(keyinput39), 
        .A(n4143), .ZN(n4146) );
  NOR2_X1 U4744 ( .A1(n4147), .A2(n4146), .ZN(n4153) );
  INV_X1 U4745 ( .A(D_REG_16__SCAN_IN), .ZN(n4479) );
  INV_X1 U4746 ( .A(D_REG_18__SCAN_IN), .ZN(n4478) );
  AOI22_X1 U4747 ( .A1(n4479), .A2(keyinput47), .B1(keyinput1), .B2(n4478), 
        .ZN(n4148) );
  OAI221_X1 U4748 ( .B1(n4479), .B2(keyinput47), .C1(n4478), .C2(keyinput1), 
        .A(n4148), .ZN(n4151) );
  INV_X1 U4749 ( .A(D_REG_6__SCAN_IN), .ZN(n4481) );
  INV_X1 U4750 ( .A(D_REG_12__SCAN_IN), .ZN(n4480) );
  AOI22_X1 U4751 ( .A1(n4481), .A2(keyinput6), .B1(keyinput42), .B2(n4480), 
        .ZN(n4149) );
  OAI221_X1 U4752 ( .B1(n4481), .B2(keyinput6), .C1(n4480), .C2(keyinput42), 
        .A(n4149), .ZN(n4150) );
  NOR2_X1 U4753 ( .A1(n4151), .A2(n4150), .ZN(n4152) );
  AND3_X1 U4754 ( .A1(n4154), .A2(n4153), .A3(n4152), .ZN(n4169) );
  INV_X1 U4755 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U4756 ( .A1(n4156), .A2(keyinput56), .B1(keyinput5), .B2(n4232), 
        .ZN(n4155) );
  OAI221_X1 U4757 ( .B1(n4156), .B2(keyinput56), .C1(n4232), .C2(keyinput5), 
        .A(n4155), .ZN(n4167) );
  XNOR2_X1 U4758 ( .A(IR_REG_1__SCAN_IN), .B(keyinput15), .ZN(n4160) );
  XNOR2_X1 U4759 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput55), .ZN(n4159) );
  XNOR2_X1 U4760 ( .A(IR_REG_14__SCAN_IN), .B(keyinput14), .ZN(n4158) );
  XNOR2_X1 U4761 ( .A(IR_REG_8__SCAN_IN), .B(keyinput45), .ZN(n4157) );
  NAND4_X1 U4762 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), .ZN(n4166)
         );
  XNOR2_X1 U4763 ( .A(IR_REG_22__SCAN_IN), .B(keyinput51), .ZN(n4164) );
  XNOR2_X1 U4764 ( .A(REG1_REG_28__SCAN_IN), .B(keyinput21), .ZN(n4163) );
  XNOR2_X1 U4765 ( .A(IR_REG_27__SCAN_IN), .B(keyinput19), .ZN(n4162) );
  XNOR2_X1 U4766 ( .A(B_REG_SCAN_IN), .B(keyinput54), .ZN(n4161) );
  NAND4_X1 U4767 ( .A1(n4164), .A2(n4163), .A3(n4162), .A4(n4161), .ZN(n4165)
         );
  NOR3_X1 U4768 ( .A1(n4167), .A2(n4166), .A3(n4165), .ZN(n4168) );
  AND4_X1 U4769 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4211)
         );
  INV_X1 U4770 ( .A(DATAI_28_), .ZN(n4334) );
  AOI22_X1 U4771 ( .A1(n4334), .A2(keyinput41), .B1(keyinput9), .B2(n4173), 
        .ZN(n4172) );
  OAI221_X1 U4772 ( .B1(n4334), .B2(keyinput41), .C1(n4173), .C2(keyinput9), 
        .A(n4172), .ZN(n4184) );
  INV_X1 U4773 ( .A(DATAI_20_), .ZN(n4175) );
  AOI22_X1 U4774 ( .A1(n4175), .A2(keyinput59), .B1(keyinput63), .B2(n2439), 
        .ZN(n4174) );
  OAI221_X1 U4775 ( .B1(n4175), .B2(keyinput59), .C1(n2439), .C2(keyinput63), 
        .A(n4174), .ZN(n4183) );
  AOI22_X1 U4776 ( .A1(n4177), .A2(keyinput25), .B1(keyinput20), .B2(n2307), 
        .ZN(n4176) );
  OAI221_X1 U4777 ( .B1(n4177), .B2(keyinput25), .C1(n2307), .C2(keyinput20), 
        .A(n4176), .ZN(n4182) );
  AOI22_X1 U4778 ( .A1(n4180), .A2(keyinput38), .B1(n4179), .B2(keyinput8), 
        .ZN(n4178) );
  OAI221_X1 U4779 ( .B1(n4180), .B2(keyinput38), .C1(n4179), .C2(keyinput8), 
        .A(n4178), .ZN(n4181) );
  NOR4_X1 U4780 ( .A1(n4184), .A2(n4183), .A3(n4182), .A4(n4181), .ZN(n4210)
         );
  INV_X1 U4781 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4288) );
  INV_X1 U4782 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U4783 ( .A1(n4288), .A2(keyinput34), .B1(n4186), .B2(keyinput48), 
        .ZN(n4185) );
  OAI221_X1 U4784 ( .B1(n4288), .B2(keyinput34), .C1(n4186), .C2(keyinput48), 
        .A(n4185), .ZN(n4196) );
  AOI22_X1 U4785 ( .A1(n4266), .A2(keyinput53), .B1(keyinput60), .B2(n4188), 
        .ZN(n4187) );
  OAI221_X1 U4786 ( .B1(n4266), .B2(keyinput53), .C1(n4188), .C2(keyinput60), 
        .A(n4187), .ZN(n4195) );
  AOI22_X1 U4787 ( .A1(n4244), .A2(keyinput3), .B1(n4221), .B2(keyinput62), 
        .ZN(n4189) );
  OAI221_X1 U4788 ( .B1(n4244), .B2(keyinput3), .C1(n4221), .C2(keyinput62), 
        .A(n4189), .ZN(n4194) );
  AOI22_X1 U4789 ( .A1(n4192), .A2(keyinput22), .B1(n4191), .B2(keyinput7), 
        .ZN(n4190) );
  OAI221_X1 U4790 ( .B1(n4192), .B2(keyinput22), .C1(n4191), .C2(keyinput7), 
        .A(n4190), .ZN(n4193) );
  NOR4_X1 U4791 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(n4209)
         );
  INV_X1 U4792 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4215) );
  INV_X1 U4793 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4397) );
  AOI22_X1 U4794 ( .A1(n4215), .A2(keyinput0), .B1(keyinput43), .B2(n4397), 
        .ZN(n4197) );
  OAI221_X1 U4795 ( .B1(n4215), .B2(keyinput0), .C1(n4397), .C2(keyinput43), 
        .A(n4197), .ZN(n4207) );
  INV_X1 U4796 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4452) );
  INV_X1 U4797 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U4798 ( .A1(n4452), .A2(keyinput33), .B1(keyinput58), .B2(n4199), 
        .ZN(n4198) );
  OAI221_X1 U4799 ( .B1(n4452), .B2(keyinput33), .C1(n4199), .C2(keyinput58), 
        .A(n4198), .ZN(n4206) );
  INV_X1 U4800 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4345) );
  INV_X1 U4801 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U4802 ( .A1(n4345), .A2(keyinput4), .B1(keyinput18), .B2(n4201), 
        .ZN(n4200) );
  OAI221_X1 U4803 ( .B1(n4345), .B2(keyinput4), .C1(n4201), .C2(keyinput18), 
        .A(n4200), .ZN(n4205) );
  AOI22_X1 U4804 ( .A1(n2660), .A2(keyinput32), .B1(n4203), .B2(keyinput24), 
        .ZN(n4202) );
  OAI221_X1 U4805 ( .B1(n2660), .B2(keyinput32), .C1(n4203), .C2(keyinput24), 
        .A(n4202), .ZN(n4204) );
  NOR4_X1 U4806 ( .A1(n4207), .A2(n4206), .A3(n4205), .A4(n4204), .ZN(n4208)
         );
  NAND4_X1 U4807 ( .A1(n4211), .A2(n4210), .A3(n4209), .A4(n4208), .ZN(n4250)
         );
  INV_X1 U4808 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4214) );
  NAND4_X1 U4809 ( .A1(n4214), .A2(n4307), .A3(n4213), .A4(n4212), .ZN(n4219)
         );
  NAND4_X1 U4810 ( .A1(DATAI_28_), .A2(ADDR_REG_0__SCAN_IN), .A3(
        ADDR_REG_13__SCAN_IN), .A4(n4215), .ZN(n4218) );
  NAND4_X1 U4811 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG0_REG_28__SCAN_IN), .A3(
        REG0_REG_26__SCAN_IN), .A4(REG1_REG_26__SCAN_IN), .ZN(n4217) );
  NAND4_X1 U4812 ( .A1(REG1_REG_23__SCAN_IN), .A2(REG1_REG_20__SCAN_IN), .A3(
        DATAI_20_), .A4(REG0_REG_24__SCAN_IN), .ZN(n4216) );
  NOR4_X1 U4813 ( .A1(n4219), .A2(n4218), .A3(n4217), .A4(n4216), .ZN(n4248)
         );
  NOR4_X1 U4814 ( .A1(DATAO_REG_25__SCAN_IN), .A2(DATAO_REG_10__SCAN_IN), .A3(
        DATAO_REG_19__SCAN_IN), .A4(ADDR_REG_18__SCAN_IN), .ZN(n4243) );
  NAND4_X1 U4815 ( .A1(n4478), .A2(n4481), .A3(REG0_REG_5__SCAN_IN), .A4(
        D_REG_0__SCAN_IN), .ZN(n4223) );
  NAND4_X1 U4816 ( .A1(n4221), .A2(n4220), .A3(REG0_REG_16__SCAN_IN), .A4(
        REG0_REG_14__SCAN_IN), .ZN(n4222) );
  NOR2_X1 U4817 ( .A1(n4223), .A2(n4222), .ZN(n4242) );
  INV_X1 U4818 ( .A(IR_REG_24__SCAN_IN), .ZN(n4226) );
  INV_X1 U4819 ( .A(B_REG_SCAN_IN), .ZN(n4224) );
  NAND4_X1 U4820 ( .A1(n4226), .A2(n4225), .A3(n4224), .A4(IR_REG_8__SCAN_IN), 
        .ZN(n4240) );
  NAND3_X1 U4821 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .ZN(n4239) );
  NOR4_X1 U4822 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .A3(
        IR_REG_2__SCAN_IN), .A4(IR_REG_1__SCAN_IN), .ZN(n4229) );
  NOR3_X1 U4823 ( .A1(REG1_REG_10__SCAN_IN), .A2(DATAI_7_), .A3(DATAI_5_), 
        .ZN(n4228) );
  NOR4_X1 U4824 ( .A1(REG0_REG_12__SCAN_IN), .A2(REG2_REG_13__SCAN_IN), .A3(
        REG2_REG_12__SCAN_IN), .A4(n4266), .ZN(n4227) );
  NAND3_X1 U4825 ( .A1(n4229), .A2(n4228), .A3(n4227), .ZN(n4236) );
  NOR4_X1 U4826 ( .A1(REG3_REG_7__SCAN_IN), .A2(DATAI_17_), .A3(n4231), .A4(
        n4230), .ZN(n4234) );
  NOR4_X1 U4827 ( .A1(REG3_REG_2__SCAN_IN), .A2(REG0_REG_1__SCAN_IN), .A3(
        n4232), .A4(n2667), .ZN(n4233) );
  NAND2_X1 U4828 ( .A1(n4234), .A2(n4233), .ZN(n4235) );
  NOR2_X1 U4829 ( .A1(n4236), .A2(n4235), .ZN(n4237) );
  NAND3_X1 U4830 ( .A1(n2248), .A2(D_REG_12__SCAN_IN), .A3(n4237), .ZN(n4238)
         );
  NOR3_X1 U4831 ( .A1(n4240), .A2(n4239), .A3(n4238), .ZN(n4241) );
  AND3_X1 U4832 ( .A1(n4243), .A2(n4242), .A3(n4241), .ZN(n4247) );
  NOR4_X1 U4833 ( .A1(REG2_REG_1__SCAN_IN), .A2(REG2_REG_3__SCAN_IN), .A3(
        DATAO_REG_22__SCAN_IN), .A4(n4244), .ZN(n4246) );
  NOR4_X1 U4834 ( .A1(DATAI_26_), .A2(DATAO_REG_1__SCAN_IN), .A3(
        ADDR_REG_6__SCAN_IN), .A4(ADDR_REG_2__SCAN_IN), .ZN(n4245) );
  NAND4_X1 U4835 ( .A1(n4248), .A2(n4247), .A3(n4246), .A4(n4245), .ZN(n4249)
         );
  XNOR2_X1 U4836 ( .A(n4250), .B(n4249), .ZN(n4251) );
  XNOR2_X1 U4837 ( .A(n4252), .B(n4251), .ZN(U3535) );
  AOI21_X1 U4838 ( .B1(n4545), .B2(n4254), .A(n4253), .ZN(n4255) );
  OAI21_X1 U4839 ( .B1(n4256), .B2(n4540), .A(n4255), .ZN(n4316) );
  MUX2_X1 U4840 ( .A(REG1_REG_16__SCAN_IN), .B(n4316), .S(n4567), .Z(U3534) );
  AOI21_X1 U4841 ( .B1(n4545), .B2(n4258), .A(n4257), .ZN(n4259) );
  OAI21_X1 U4842 ( .B1(n4260), .B2(n4540), .A(n4259), .ZN(n4317) );
  MUX2_X1 U4843 ( .A(REG1_REG_15__SCAN_IN), .B(n4317), .S(n4567), .Z(U3533) );
  AOI21_X1 U4844 ( .B1(n4262), .B2(n4533), .A(n4261), .ZN(n4318) );
  MUX2_X1 U4845 ( .A(n4406), .B(n4318), .S(n4567), .Z(n4263) );
  OAI21_X1 U4846 ( .B1(n4268), .B2(n4321), .A(n4263), .ZN(U3532) );
  AOI21_X1 U4847 ( .B1(n4524), .B2(n4265), .A(n4264), .ZN(n4322) );
  MUX2_X1 U4848 ( .A(n4266), .B(n4322), .S(n4567), .Z(n4267) );
  OAI21_X1 U4849 ( .B1(n4268), .B2(n4326), .A(n4267), .ZN(U3531) );
  AND2_X1 U4850 ( .A1(n4270), .A2(n4269), .ZN(n4271) );
  OR2_X1 U4851 ( .A1(n4464), .A2(n4271), .ZN(n4275) );
  NAND2_X1 U4852 ( .A1(n4273), .A2(n4272), .ZN(n4274) );
  NAND2_X1 U4853 ( .A1(n4275), .A2(n4274), .ZN(n4471) );
  NAND2_X1 U4854 ( .A1(n4277), .A2(n4276), .ZN(n4469) );
  OAI21_X1 U4855 ( .B1(n4464), .B2(n4549), .A(n4469), .ZN(n4278) );
  OR2_X1 U4856 ( .A1(n4471), .A2(n4278), .ZN(n4507) );
  MUX2_X1 U4857 ( .A(REG1_REG_0__SCAN_IN), .B(n4507), .S(n4567), .Z(U3518) );
  INV_X1 U4858 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4279) );
  MUX2_X1 U4859 ( .A(n4279), .B(n4338), .S(n4555), .Z(n4280) );
  OAI21_X1 U4860 ( .B1(n4281), .B2(n4325), .A(n4280), .ZN(U3517) );
  INV_X1 U4861 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4282) );
  MUX2_X1 U4862 ( .A(n4282), .B(n4341), .S(n4555), .Z(n4283) );
  OAI21_X1 U4863 ( .B1(n4284), .B2(n4325), .A(n4283), .ZN(U3516) );
  MUX2_X1 U4864 ( .A(REG0_REG_29__SCAN_IN), .B(n4285), .S(n4555), .Z(U3515) );
  MUX2_X1 U4865 ( .A(REG0_REG_27__SCAN_IN), .B(n4286), .S(n4555), .Z(U3513) );
  MUX2_X1 U4866 ( .A(n4288), .B(n4287), .S(n4555), .Z(n4289) );
  OAI21_X1 U4867 ( .B1(n4290), .B2(n4325), .A(n4289), .ZN(U3512) );
  INV_X1 U4868 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4292) );
  MUX2_X1 U4869 ( .A(n4292), .B(n4291), .S(n4555), .Z(n4293) );
  OAI21_X1 U4870 ( .B1(n4294), .B2(n4325), .A(n4293), .ZN(U3511) );
  INV_X1 U4871 ( .A(n4295), .ZN(n4296) );
  MUX2_X1 U4872 ( .A(n4297), .B(n4296), .S(n4555), .Z(n4298) );
  OAI21_X1 U4873 ( .B1(n4299), .B2(n4325), .A(n4298), .ZN(U3510) );
  INV_X1 U4874 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4301) );
  MUX2_X1 U4875 ( .A(n4301), .B(n4300), .S(n4555), .Z(n4302) );
  OAI21_X1 U4876 ( .B1(n4303), .B2(n4325), .A(n4302), .ZN(U3509) );
  MUX2_X1 U4877 ( .A(REG0_REG_22__SCAN_IN), .B(n4304), .S(n4555), .Z(U3508) );
  MUX2_X1 U4878 ( .A(REG0_REG_21__SCAN_IN), .B(n4305), .S(n4555), .Z(U3507) );
  MUX2_X1 U4879 ( .A(n4307), .B(n4306), .S(n4555), .Z(n4308) );
  OAI21_X1 U4880 ( .B1(n4309), .B2(n4325), .A(n4308), .ZN(U3506) );
  INV_X1 U4881 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4311) );
  MUX2_X1 U4882 ( .A(n4311), .B(n4310), .S(n4555), .Z(n4312) );
  OAI21_X1 U4883 ( .B1(n4313), .B2(n4325), .A(n4312), .ZN(U3505) );
  MUX2_X1 U4884 ( .A(REG0_REG_18__SCAN_IN), .B(n4314), .S(n4555), .Z(U3503) );
  MUX2_X1 U4885 ( .A(REG0_REG_17__SCAN_IN), .B(n4315), .S(n4555), .Z(U3501) );
  MUX2_X1 U4886 ( .A(REG0_REG_16__SCAN_IN), .B(n4316), .S(n4555), .Z(U3499) );
  MUX2_X1 U4887 ( .A(REG0_REG_15__SCAN_IN), .B(n4317), .S(n4555), .Z(U3497) );
  MUX2_X1 U4888 ( .A(n4319), .B(n4318), .S(n4555), .Z(n4320) );
  OAI21_X1 U4889 ( .B1(n4321), .B2(n4325), .A(n4320), .ZN(U3495) );
  INV_X1 U4890 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4323) );
  MUX2_X1 U4891 ( .A(n4323), .B(n4322), .S(n4555), .Z(n4324) );
  OAI21_X1 U4892 ( .B1(n4326), .B2(n4325), .A(n4324), .ZN(U3493) );
  MUX2_X1 U4893 ( .A(n2240), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4894 ( .A(n4327), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4895 ( .A(DATAI_25_), .B(n4328), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4896 ( .A(n4329), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4897 ( .A(DATAI_20_), .B(n4330), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4898 ( .A(n4331), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U4899 ( .A(n2702), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4900 ( .A(n4332), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4901 ( .A(n4333), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4902 ( .A1(STATE_REG_SCAN_IN), .A2(n4335), .B1(n4334), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U4903 ( .A1(n4336), .A2(n4458), .B1(n4463), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4337) );
  OAI21_X1 U4904 ( .B1(n4463), .B2(n4338), .A(n4337), .ZN(U3260) );
  AOI22_X1 U4905 ( .A1(n4339), .A2(n4458), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4463), .ZN(n4340) );
  OAI21_X1 U4906 ( .B1(n4463), .B2(n4341), .A(n4340), .ZN(U3261) );
  OAI211_X1 U4907 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4343), .A(n4437), .B(n4342), 
        .ZN(n4344) );
  OAI21_X1 U4908 ( .B1(n4451), .B2(n4345), .A(n4344), .ZN(n4346) );
  NOR2_X1 U4909 ( .A1(n4347), .A2(n4346), .ZN(n4351) );
  OAI211_X1 U4910 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4349), .A(n4435), .B(n4348), 
        .ZN(n4350) );
  OAI211_X1 U4911 ( .C1(n4440), .C2(n4505), .A(n4351), .B(n4350), .ZN(U3246)
         );
  AOI211_X1 U4912 ( .C1(n4354), .C2(n4353), .A(n4352), .B(n4441), .ZN(n4357)
         );
  INV_X1 U4913 ( .A(n4355), .ZN(n4356) );
  AOI211_X1 U4914 ( .C1(n4427), .C2(ADDR_REG_8__SCAN_IN), .A(n4357), .B(n4356), 
        .ZN(n4361) );
  OAI211_X1 U4915 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4359), .A(n4437), .B(n4358), 
        .ZN(n4360) );
  OAI211_X1 U4916 ( .C1(n4440), .C2(n4362), .A(n4361), .B(n4360), .ZN(U3248)
         );
  AOI211_X1 U4917 ( .C1(n2045), .C2(n4364), .A(n4363), .B(n4441), .ZN(n4366)
         );
  AOI211_X1 U4918 ( .C1(n4427), .C2(ADDR_REG_9__SCAN_IN), .A(n4366), .B(n4365), 
        .ZN(n4371) );
  OAI211_X1 U4919 ( .C1(n4369), .C2(n4368), .A(n4437), .B(n4367), .ZN(n4370)
         );
  OAI211_X1 U4920 ( .C1(n4440), .C2(n4501), .A(n4371), .B(n4370), .ZN(U3249)
         );
  AOI211_X1 U4921 ( .C1(n4374), .C2(n4373), .A(n4372), .B(n4441), .ZN(n4375)
         );
  AOI211_X1 U4922 ( .C1(n4427), .C2(ADDR_REG_11__SCAN_IN), .A(n4376), .B(n4375), .ZN(n4381) );
  OAI211_X1 U4923 ( .C1(n4379), .C2(n4378), .A(n4437), .B(n4377), .ZN(n4380)
         );
  OAI211_X1 U4924 ( .C1(n4440), .C2(n4382), .A(n4381), .B(n4380), .ZN(U3251)
         );
  AOI211_X1 U4925 ( .C1(n4385), .C2(n4384), .A(n4383), .B(n4441), .ZN(n4388)
         );
  INV_X1 U4926 ( .A(n4386), .ZN(n4387) );
  AOI211_X1 U4927 ( .C1(n4427), .C2(ADDR_REG_12__SCAN_IN), .A(n4388), .B(n4387), .ZN(n4392) );
  OAI211_X1 U4928 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4390), .A(n4437), .B(n4389), .ZN(n4391) );
  OAI211_X1 U4929 ( .C1(n4440), .C2(n2093), .A(n4392), .B(n4391), .ZN(U3252)
         );
  AOI211_X1 U4930 ( .C1(n2038), .C2(n4394), .A(n4393), .B(n4441), .ZN(n4395)
         );
  AOI211_X1 U4931 ( .C1(ADDR_REG_13__SCAN_IN), .C2(n4427), .A(n4396), .B(n4395), .ZN(n4403) );
  AOI22_X1 U4932 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4398), .B1(n4496), .B2(
        n4397), .ZN(n4401) );
  AOI21_X1 U4933 ( .B1(n4401), .B2(n4400), .A(n4445), .ZN(n4399) );
  OAI21_X1 U4934 ( .B1(n4401), .B2(n4400), .A(n4399), .ZN(n4402) );
  OAI211_X1 U4935 ( .C1(n4440), .C2(n4496), .A(n4403), .B(n4402), .ZN(U3253)
         );
  NAND2_X1 U4936 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4427), .ZN(n4414) );
  AOI211_X1 U4937 ( .C1(n4406), .C2(n4405), .A(n4404), .B(n4441), .ZN(n4411)
         );
  AOI211_X1 U4938 ( .C1(n4409), .C2(n4408), .A(n4407), .B(n4445), .ZN(n4410)
         );
  AOI211_X1 U4939 ( .C1(n4450), .C2(n4493), .A(n4411), .B(n4410), .ZN(n4413)
         );
  NAND3_X1 U4940 ( .A1(n4414), .A2(n4413), .A3(n4412), .ZN(U3254) );
  AOI211_X1 U4941 ( .C1(n2034), .C2(n4416), .A(n4415), .B(n4445), .ZN(n4417)
         );
  AOI211_X1 U4942 ( .C1(n4427), .C2(ADDR_REG_15__SCAN_IN), .A(n4418), .B(n4417), .ZN(n4424) );
  AOI21_X1 U4943 ( .B1(n4421), .B2(n4420), .A(n4419), .ZN(n4422) );
  NAND2_X1 U4944 ( .A1(n4435), .A2(n4422), .ZN(n4423) );
  OAI211_X1 U4945 ( .C1(n4440), .C2(n4492), .A(n4424), .B(n4423), .ZN(U3255)
         );
  INV_X1 U4946 ( .A(n4425), .ZN(n4426) );
  AOI21_X1 U4947 ( .B1(n4427), .B2(ADDR_REG_16__SCAN_IN), .A(n4426), .ZN(n4439) );
  OAI21_X1 U4948 ( .B1(n4430), .B2(n4429), .A(n4428), .ZN(n4436) );
  OAI21_X1 U4949 ( .B1(n4433), .B2(n4432), .A(n4431), .ZN(n4434) );
  AOI22_X1 U4950 ( .A1(n4437), .A2(n4436), .B1(n4435), .B2(n4434), .ZN(n4438)
         );
  OAI211_X1 U4951 ( .C1(n4490), .C2(n4440), .A(n4439), .B(n4438), .ZN(U3256)
         );
  AOI211_X1 U4952 ( .C1(n4447), .C2(n4446), .A(n2028), .B(n4445), .ZN(n4448)
         );
  AOI22_X1 U4953 ( .A1(n4454), .A2(n4453), .B1(REG2_REG_6__SCAN_IN), .B2(n4463), .ZN(n4461) );
  INV_X1 U4954 ( .A(n4455), .ZN(n4459) );
  INV_X1 U4955 ( .A(n4456), .ZN(n4457) );
  AOI22_X1 U4956 ( .A1(n4459), .A2(n4466), .B1(n4458), .B2(n4457), .ZN(n4460)
         );
  OAI211_X1 U4957 ( .C1(n4463), .C2(n4462), .A(n4461), .B(n4460), .ZN(U3284)
         );
  INV_X1 U4958 ( .A(n4464), .ZN(n4465) );
  AOI22_X1 U4959 ( .A1(n4466), .A2(n4465), .B1(REG2_REG_0__SCAN_IN), .B2(n4463), .ZN(n4474) );
  INV_X1 U4960 ( .A(n4467), .ZN(n4468) );
  NOR2_X1 U4961 ( .A1(n4469), .A2(n4468), .ZN(n4472) );
  OAI21_X1 U4962 ( .B1(n4472), .B2(n4471), .A(n4470), .ZN(n4473) );
  OAI211_X1 U4963 ( .C1(n4476), .C2(n4475), .A(n4474), .B(n4473), .ZN(U3290)
         );
  AND2_X1 U4964 ( .A1(D_REG_31__SCAN_IN), .A2(n4484), .ZN(U3291) );
  AND2_X1 U4965 ( .A1(D_REG_30__SCAN_IN), .A2(n4484), .ZN(U3292) );
  AND2_X1 U4966 ( .A1(D_REG_29__SCAN_IN), .A2(n4484), .ZN(U3293) );
  AND2_X1 U4967 ( .A1(D_REG_28__SCAN_IN), .A2(n4484), .ZN(U3294) );
  AND2_X1 U4968 ( .A1(D_REG_27__SCAN_IN), .A2(n4484), .ZN(U3295) );
  AND2_X1 U4969 ( .A1(D_REG_26__SCAN_IN), .A2(n4484), .ZN(U3296) );
  AND2_X1 U4970 ( .A1(D_REG_25__SCAN_IN), .A2(n4484), .ZN(U3297) );
  AND2_X1 U4971 ( .A1(D_REG_24__SCAN_IN), .A2(n4484), .ZN(U3298) );
  AND2_X1 U4972 ( .A1(D_REG_23__SCAN_IN), .A2(n4484), .ZN(U3299) );
  AND2_X1 U4973 ( .A1(D_REG_22__SCAN_IN), .A2(n4484), .ZN(U3300) );
  NOR2_X1 U4974 ( .A1(n4483), .A2(n4477), .ZN(U3301) );
  AND2_X1 U4975 ( .A1(D_REG_20__SCAN_IN), .A2(n4484), .ZN(U3302) );
  AND2_X1 U4976 ( .A1(D_REG_19__SCAN_IN), .A2(n4484), .ZN(U3303) );
  NOR2_X1 U4977 ( .A1(n4483), .A2(n4478), .ZN(U3304) );
  AND2_X1 U4978 ( .A1(D_REG_17__SCAN_IN), .A2(n4484), .ZN(U3305) );
  NOR2_X1 U4979 ( .A1(n4483), .A2(n4479), .ZN(U3306) );
  AND2_X1 U4980 ( .A1(D_REG_15__SCAN_IN), .A2(n4484), .ZN(U3307) );
  AND2_X1 U4981 ( .A1(D_REG_14__SCAN_IN), .A2(n4484), .ZN(U3308) );
  AND2_X1 U4982 ( .A1(D_REG_13__SCAN_IN), .A2(n4484), .ZN(U3309) );
  NOR2_X1 U4983 ( .A1(n4483), .A2(n4480), .ZN(U3310) );
  AND2_X1 U4984 ( .A1(D_REG_11__SCAN_IN), .A2(n4484), .ZN(U3311) );
  AND2_X1 U4985 ( .A1(D_REG_10__SCAN_IN), .A2(n4484), .ZN(U3312) );
  AND2_X1 U4986 ( .A1(D_REG_9__SCAN_IN), .A2(n4484), .ZN(U3313) );
  AND2_X1 U4987 ( .A1(D_REG_8__SCAN_IN), .A2(n4484), .ZN(U3314) );
  AND2_X1 U4988 ( .A1(D_REG_7__SCAN_IN), .A2(n4484), .ZN(U3315) );
  NOR2_X1 U4989 ( .A1(n4483), .A2(n4481), .ZN(U3316) );
  AND2_X1 U4990 ( .A1(D_REG_5__SCAN_IN), .A2(n4484), .ZN(U3317) );
  NOR2_X1 U4991 ( .A1(n4483), .A2(n4482), .ZN(U3318) );
  AND2_X1 U4992 ( .A1(D_REG_3__SCAN_IN), .A2(n4484), .ZN(U3319) );
  AND2_X1 U4993 ( .A1(D_REG_2__SCAN_IN), .A2(n4484), .ZN(U3320) );
  INV_X1 U4994 ( .A(DATAI_23_), .ZN(n4486) );
  AOI21_X1 U4995 ( .B1(U3149), .B2(n4486), .A(n4485), .ZN(U3329) );
  AOI22_X1 U4996 ( .A1(STATE_REG_SCAN_IN), .A2(n4488), .B1(n4487), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U4997 ( .A1(STATE_REG_SCAN_IN), .A2(n4490), .B1(n4489), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U4998 ( .A(DATAI_15_), .ZN(n4491) );
  AOI22_X1 U4999 ( .A1(STATE_REG_SCAN_IN), .A2(n4492), .B1(n4491), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5000 ( .A1(U3149), .A2(n4493), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4494) );
  INV_X1 U5001 ( .A(n4494), .ZN(U3338) );
  INV_X1 U5002 ( .A(DATAI_13_), .ZN(n4495) );
  AOI22_X1 U5003 ( .A1(STATE_REG_SCAN_IN), .A2(n4496), .B1(n4495), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5004 ( .A(DATAI_12_), .ZN(n4497) );
  AOI22_X1 U5005 ( .A1(STATE_REG_SCAN_IN), .A2(n2093), .B1(n4497), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5006 ( .A1(U3149), .A2(n4498), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4499) );
  INV_X1 U5007 ( .A(n4499), .ZN(U3341) );
  INV_X1 U5008 ( .A(DATAI_9_), .ZN(n4500) );
  AOI22_X1 U5009 ( .A1(STATE_REG_SCAN_IN), .A2(n4501), .B1(n4500), .B2(U3149), 
        .ZN(U3343) );
  OAI22_X1 U5010 ( .A1(U3149), .A2(n4502), .B1(DATAI_8_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4503) );
  INV_X1 U5011 ( .A(n4503), .ZN(U3344) );
  INV_X1 U5012 ( .A(DATAI_6_), .ZN(n4504) );
  AOI22_X1 U5013 ( .A1(STATE_REG_SCAN_IN), .A2(n4505), .B1(n4504), .B2(U3149), 
        .ZN(U3346) );
  OAI22_X1 U5014 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4506) );
  INV_X1 U5015 ( .A(n4506), .ZN(U3352) );
  INV_X1 U5016 ( .A(n4507), .ZN(n4509) );
  INV_X1 U5017 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4508) );
  AOI22_X1 U5018 ( .A1(n4555), .A2(n4509), .B1(n4508), .B2(n4553), .ZN(U3467)
         );
  OAI22_X1 U5019 ( .A1(n4511), .A2(n4549), .B1(n4548), .B2(n4510), .ZN(n4512)
         );
  NOR2_X1 U5020 ( .A1(n4513), .A2(n4512), .ZN(n4556) );
  AOI22_X1 U5021 ( .A1(n4555), .A2(n4556), .B1(n4514), .B2(n4553), .ZN(U3469)
         );
  OAI22_X1 U5022 ( .A1(n4516), .A2(n4549), .B1(n4548), .B2(n4515), .ZN(n4517)
         );
  NOR2_X1 U5023 ( .A1(n4518), .A2(n4517), .ZN(n4558) );
  INV_X1 U5024 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4519) );
  AOI22_X1 U5025 ( .A1(n4555), .A2(n4558), .B1(n4519), .B2(n4553), .ZN(U3473)
         );
  INV_X1 U5026 ( .A(n4520), .ZN(n4525) );
  INV_X1 U5027 ( .A(n4521), .ZN(n4523) );
  AOI211_X1 U5028 ( .C1(n4525), .C2(n4524), .A(n4523), .B(n4522), .ZN(n4559)
         );
  INV_X1 U5029 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U5030 ( .A1(n4555), .A2(n4559), .B1(n4526), .B2(n4553), .ZN(U3475)
         );
  NOR2_X1 U5031 ( .A1(n4527), .A2(n4540), .ZN(n4530) );
  INV_X1 U5032 ( .A(n4528), .ZN(n4529) );
  AOI211_X1 U5033 ( .C1(n4545), .C2(n4531), .A(n4530), .B(n4529), .ZN(n4560)
         );
  AOI22_X1 U5034 ( .A1(n4555), .A2(n4560), .B1(n4532), .B2(n4553), .ZN(U3477)
         );
  NAND3_X1 U5035 ( .A1(n4535), .A2(n4534), .A3(n4533), .ZN(n4536) );
  AND3_X1 U5036 ( .A1(n4538), .A2(n4537), .A3(n4536), .ZN(n4561) );
  INV_X1 U5037 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5038 ( .A1(n4555), .A2(n4561), .B1(n4539), .B2(n4553), .ZN(U3481)
         );
  NOR2_X1 U5039 ( .A1(n4541), .A2(n4540), .ZN(n4543) );
  AOI211_X1 U5040 ( .C1(n4545), .C2(n4544), .A(n4543), .B(n4542), .ZN(n4563)
         );
  INV_X1 U5041 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4546) );
  AOI22_X1 U5042 ( .A1(n4555), .A2(n4563), .B1(n4546), .B2(n4553), .ZN(U3485)
         );
  OAI22_X1 U5043 ( .A1(n4550), .A2(n4549), .B1(n4548), .B2(n4547), .ZN(n4551)
         );
  NOR2_X1 U5044 ( .A1(n4552), .A2(n4551), .ZN(n4566) );
  INV_X1 U5045 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U5046 ( .A1(n4555), .A2(n4566), .B1(n4554), .B2(n4553), .ZN(U3489)
         );
  AOI22_X1 U5047 ( .A1(n4567), .A2(n4556), .B1(n2253), .B2(n4564), .ZN(U3519)
         );
  INV_X1 U5048 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4557) );
  AOI22_X1 U5049 ( .A1(n4567), .A2(n4558), .B1(n4557), .B2(n4564), .ZN(U3521)
         );
  AOI22_X1 U5050 ( .A1(n4567), .A2(n4559), .B1(n2073), .B2(n4564), .ZN(U3522)
         );
  AOI22_X1 U5051 ( .A1(n4567), .A2(n4560), .B1(n2701), .B2(n4564), .ZN(U3523)
         );
  AOI22_X1 U5052 ( .A1(n4567), .A2(n4561), .B1(n2700), .B2(n4564), .ZN(U3525)
         );
  AOI22_X1 U5053 ( .A1(n4567), .A2(n4563), .B1(n4562), .B2(n4564), .ZN(U3527)
         );
  AOI22_X1 U5054 ( .A1(n4567), .A2(n4566), .B1(n4565), .B2(n4564), .ZN(U3529)
         );
  OR2_X1 U33090 ( .A1(n3849), .A2(n2559), .ZN(n3831) );
endmodule

