

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972;

  OAI21_X1 U2295 ( .B1(n2971), .B2(n2970), .A(n4928), .ZN(n4954) );
  BUF_X2 U2296 ( .A(n2711), .Z(n2262) );
  AND2_X1 U2298 ( .A1(n2676), .A2(n2675), .ZN(n2712) );
  INV_X1 U2300 ( .A(n2734), .ZN(n3066) );
  MUX2_X1 U2301 ( .A(IR_REG_31__SCAN_IN), .B(n2670), .S(IR_REG_29__SCAN_IN), 
        .Z(n2672) );
  NAND2_X1 U2302 ( .A1(n3167), .A2(n3166), .ZN(n3533) );
  NAND2_X1 U2303 ( .A1(n2533), .A2(IR_REG_31__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U2304 ( .A1(n4094), .A2(n4096), .ZN(n4095) );
  XNOR2_X1 U2305 ( .A(n2535), .B(n2534), .ZN(n3257) );
  NAND4_X1 U2306 ( .A1(n2745), .A2(n2744), .A3(n2743), .A4(n2742), .ZN(n4064)
         );
  OAI21_X1 U2307 ( .B1(n3252), .B2(n4912), .A(n2356), .ZN(n3253) );
  NOR2_X2 U2308 ( .A1(n2277), .A2(n2934), .ZN(n4865) );
  OAI21_X2 U2309 ( .B1(n3385), .B2(n2314), .A(n2312), .ZN(n2647) );
  AOI21_X2 U2310 ( .B1(n4159), .B2(n3191), .A(n4168), .ZN(n3193) );
  XNOR2_X2 U2311 ( .A(n2576), .B(IR_REG_2__SCAN_IN), .ZN(n4386) );
  INV_X4 U2312 ( .A(n2726), .ZN(n2810) );
  AND2_X4 U2313 ( .A1(n2688), .A2(n4874), .ZN(n2737) );
  NOR2_X2 U2314 ( .A1(n2804), .A2(n2452), .ZN(n2451) );
  CLKBUF_X1 U2315 ( .A(n3078), .Z(n2260) );
  OR2_X1 U2316 ( .A1(n3976), .A2(n3977), .ZN(n2344) );
  NAND2_X1 U2317 ( .A1(n3147), .A2(n4827), .ZN(n4960) );
  NAND4_X1 U2318 ( .A1(n2761), .A2(n2760), .A3(n2759), .A4(n2758), .ZN(n4063)
         );
  INV_X2 U2319 ( .A(n2762), .ZN(n3738) );
  NOR2_X1 U2320 ( .A1(n2334), .A2(n2333), .ZN(n2332) );
  NAND2_X1 U2321 ( .A1(n2344), .A2(n2296), .ZN(n3985) );
  AND2_X1 U2322 ( .A1(n2464), .A2(n2463), .ZN(n3194) );
  NAND2_X1 U2323 ( .A1(n2469), .A2(n2468), .ZN(n4185) );
  OAI21_X1 U2324 ( .B1(n3897), .B2(n3220), .A(n3728), .ZN(n4246) );
  NAND2_X1 U2325 ( .A1(n2422), .A2(n2420), .ZN(n3650) );
  NAND2_X1 U2326 ( .A1(n3579), .A2(n2423), .ZN(n2422) );
  NOR2_X1 U2327 ( .A1(n2467), .A2(n2466), .ZN(n2463) );
  AND2_X1 U2328 ( .A1(n4127), .A2(n4145), .ZN(n2467) );
  AND2_X1 U2329 ( .A1(n2421), .A2(n4583), .ZN(n2420) );
  AND2_X1 U2330 ( .A1(n2299), .A2(n2268), .ZN(n2426) );
  NAND2_X1 U2331 ( .A1(n2336), .A2(n2335), .ZN(n2773) );
  NOR2_X1 U2332 ( .A1(n2481), .A2(n3165), .ZN(n2480) );
  NAND2_X1 U2333 ( .A1(n3998), .A2(n2957), .ZN(n2427) );
  NAND2_X1 U2334 ( .A1(n3433), .A2(n4827), .ZN(n4825) );
  NAND3_X1 U2335 ( .A1(n2731), .A2(n2730), .A3(n2496), .ZN(n4065) );
  NAND2_X2 U2336 ( .A1(n3142), .A2(n3140), .ZN(n2734) );
  AND2_X1 U2337 ( .A1(n2675), .A2(n3263), .ZN(n2727) );
  OAI21_X1 U2338 ( .B1(n2746), .B2(n2399), .A(n2398), .ZN(n4732) );
  INV_X1 U2339 ( .A(n3434), .ZN(n3142) );
  AND2_X1 U2340 ( .A1(n2687), .A2(n3800), .ZN(n3434) );
  XNOR2_X1 U2341 ( .A(n2532), .B(IR_REG_26__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U2342 ( .A1(n2681), .A2(IR_REG_31__SCAN_IN), .ZN(n2683) );
  INV_X1 U2343 ( .A(n2543), .ZN(n2667) );
  AND2_X1 U2344 ( .A1(n2514), .A2(n2294), .ZN(n2375) );
  AND2_X1 U2345 ( .A1(n2513), .A2(n2512), .ZN(n2515) );
  NAND2_X1 U2346 ( .A1(n2575), .A2(n2499), .ZN(n2579) );
  AND2_X1 U2347 ( .A1(n2557), .A2(n2504), .ZN(n2513) );
  AND4_X1 U2348 ( .A1(n2503), .A2(n2502), .A3(n2501), .A4(n2592), .ZN(n2557)
         );
  INV_X1 U2349 ( .A(IR_REG_20__SCAN_IN), .ZN(n2682) );
  INV_X1 U2350 ( .A(IR_REG_13__SCAN_IN), .ZN(n2558) );
  NOR2_X1 U2351 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2502)
         );
  NOR2_X1 U2352 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2501)
         );
  NAND2_X1 U2353 ( .A1(n2439), .A2(n2437), .ZN(n2681) );
  INV_X1 U2354 ( .A(n2438), .ZN(n2437) );
  OR2_X1 U2355 ( .A1(n2553), .A2(n2440), .ZN(n2439) );
  OAI21_X1 U2356 ( .B1(n2264), .B2(n2440), .A(n2508), .ZN(n2438) );
  NOR2_X1 U2357 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2493)
         );
  NOR2_X1 U2358 ( .A1(n2773), .A2(n2418), .ZN(n2417) );
  INV_X1 U2359 ( .A(n3055), .ZN(n2462) );
  INV_X1 U2360 ( .A(n4635), .ZN(n2314) );
  NAND2_X1 U2361 ( .A1(n2474), .A2(n2473), .ZN(n2472) );
  INV_X1 U2362 ( .A(n4205), .ZN(n2473) );
  NAND2_X1 U2363 ( .A1(n2476), .A2(n2282), .ZN(n2474) );
  INV_X1 U2364 ( .A(n2483), .ZN(n2478) );
  AOI21_X1 U2365 ( .B1(n4124), .B2(n3746), .A(n3229), .ZN(n3230) );
  INV_X1 U2366 ( .A(IR_REG_28__SCAN_IN), .ZN(n2544) );
  INV_X1 U2367 ( .A(IR_REG_2__SCAN_IN), .ZN(n2499) );
  INV_X1 U2368 ( .A(n2323), .ZN(n2575) );
  AND2_X1 U2369 ( .A1(n2458), .A2(n2297), .ZN(n2457) );
  INV_X1 U2370 ( .A(n3964), .ZN(n2452) );
  XNOR2_X1 U2371 ( .A(n2750), .B(n2734), .ZN(n2751) );
  AND2_X1 U2372 ( .A1(n2676), .A2(n2674), .ZN(n2756) );
  OR2_X1 U2373 ( .A1(n4616), .A2(n4617), .ZN(n2380) );
  AND2_X1 U2374 ( .A1(n2405), .A2(n2404), .ZN(n4630) );
  OAI21_X1 U2375 ( .B1(n4648), .B2(n2409), .A(n2407), .ZN(n2610) );
  AND2_X1 U2376 ( .A1(n4646), .A2(REG1_REG_11__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U2377 ( .A1(n4822), .A2(n2408), .ZN(n2407) );
  OR2_X1 U2378 ( .A1(n4093), .A2(n4092), .ZN(n2324) );
  NAND2_X1 U2379 ( .A1(n4694), .A2(n2656), .ZN(n4094) );
  INV_X1 U2380 ( .A(n2316), .ZN(n2655) );
  NAND2_X1 U2381 ( .A1(n2324), .A2(n2310), .ZN(n2622) );
  OR2_X1 U2382 ( .A1(n3193), .A2(n2291), .ZN(n2464) );
  OAI22_X1 U2383 ( .A1(n3267), .A2(D_REG_0__SCAN_IN), .B1(n3270), .B2(n3269), 
        .ZN(n3429) );
  AND2_X1 U2384 ( .A1(n2545), .A2(n2544), .ZN(n2664) );
  NAND2_X1 U2385 ( .A1(n2681), .A2(n2509), .ZN(n4787) );
  NAND2_X1 U2386 ( .A1(n2553), .A2(n2264), .ZN(n2436) );
  INV_X1 U2387 ( .A(n4731), .ZN(n3155) );
  INV_X1 U2388 ( .A(n2766), .ZN(n2717) );
  AND2_X1 U2389 ( .A1(n2338), .A2(n3693), .ZN(n2337) );
  NAND2_X1 U2390 ( .A1(n3650), .A2(n2340), .ZN(n2339) );
  NAND2_X1 U2391 ( .A1(n2340), .A2(n2343), .ZN(n2338) );
  INV_X1 U2392 ( .A(n4084), .ZN(n2378) );
  INV_X1 U2393 ( .A(n2653), .ZN(n2377) );
  NOR2_X1 U2394 ( .A1(n2366), .A2(n4142), .ZN(n2365) );
  INV_X1 U2395 ( .A(n2368), .ZN(n2366) );
  OR2_X1 U2396 ( .A1(n3744), .A2(n3766), .ZN(n2370) );
  INV_X1 U2397 ( .A(n2471), .ZN(n2470) );
  OAI21_X1 U2398 ( .B1(n2472), .B2(n2283), .A(n2265), .ZN(n2471) );
  AOI21_X1 U2399 ( .B1(n4893), .B2(n3184), .A(n2286), .ZN(n2490) );
  NAND2_X1 U2400 ( .A1(n3169), .A2(n2495), .ZN(n2486) );
  INV_X1 U2401 ( .A(n3164), .ZN(n2481) );
  NOR2_X1 U2402 ( .A1(n3993), .A2(n4160), .ZN(n2354) );
  INV_X1 U2403 ( .A(n4235), .ZN(n4239) );
  NAND2_X1 U2404 ( .A1(n3908), .A2(n3926), .ZN(n2353) );
  AND2_X1 U2405 ( .A1(n2524), .A2(n2520), .ZN(n2492) );
  AND2_X1 U2406 ( .A1(n2541), .A2(n2540), .ZN(n2545) );
  NOR2_X1 U2407 ( .A1(IR_REG_25__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2541)
         );
  INV_X1 U2408 ( .A(IR_REG_21__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U2409 ( .A1(n2493), .A2(n2327), .ZN(n2328) );
  AND2_X1 U2410 ( .A1(n2558), .A2(n2500), .ZN(n2327) );
  INV_X1 U2411 ( .A(IR_REG_14__SCAN_IN), .ZN(n2500) );
  INV_X1 U2412 ( .A(IR_REG_5__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U2413 ( .A1(n2414), .A2(n2493), .ZN(n2556) );
  INV_X1 U2414 ( .A(n2579), .ZN(n2414) );
  NOR2_X1 U2415 ( .A1(n2451), .A2(n3496), .ZN(n2447) );
  AOI21_X1 U2416 ( .B1(n2451), .B2(n2449), .A(n2279), .ZN(n2448) );
  INV_X1 U2417 ( .A(n2497), .ZN(n2449) );
  NAND2_X1 U2418 ( .A1(n2626), .A2(n2517), .ZN(n2518) );
  INV_X1 U2419 ( .A(n2425), .ZN(n2424) );
  OAI21_X1 U2420 ( .B1(n2870), .B2(n2263), .A(n2885), .ZN(n2425) );
  INV_X1 U2421 ( .A(n2945), .ZN(n2435) );
  NAND2_X1 U2422 ( .A1(n4863), .A2(n2429), .ZN(n2432) );
  NOR2_X1 U2423 ( .A1(n4882), .A2(n2430), .ZN(n2429) );
  INV_X1 U2424 ( .A(n4866), .ZN(n2430) );
  AOI21_X1 U2425 ( .B1(n2419), .B2(n3401), .A(n2417), .ZN(n2416) );
  NAND2_X1 U2426 ( .A1(n2418), .A2(n2773), .ZN(n2419) );
  NOR2_X1 U2427 ( .A1(n3429), .A2(n3112), .ZN(n3144) );
  NAND2_X1 U2428 ( .A1(n3934), .A2(n2634), .ZN(n2635) );
  NAND2_X1 U2429 ( .A1(n4610), .A2(n2589), .ZN(n2590) );
  NOR2_X1 U2430 ( .A1(n4605), .A2(n2281), .ZN(n2639) );
  AOI22_X1 U2431 ( .A1(n2642), .A2(REG2_REG_7__SCAN_IN), .B1(n2641), .B2(n4383), .ZN(n2644) );
  NAND2_X1 U2432 ( .A1(n2321), .A2(n4382), .ZN(n2404) );
  INV_X1 U2433 ( .A(n2597), .ZN(n2321) );
  NAND2_X1 U2434 ( .A1(n2406), .A2(REG1_REG_8__SCAN_IN), .ZN(n2405) );
  INV_X1 U2435 ( .A(n2313), .ZN(n2312) );
  OAI21_X1 U2436 ( .B1(n2645), .B2(n2314), .A(n2646), .ZN(n2313) );
  AND2_X1 U2437 ( .A1(n2320), .A2(n2319), .ZN(n2614) );
  NAND2_X1 U2438 ( .A1(n4839), .A2(n4845), .ZN(n2319) );
  NAND2_X1 U2439 ( .A1(n4669), .A2(n4667), .ZN(n2320) );
  NAND2_X1 U2440 ( .A1(n4080), .A2(n2403), .ZN(n2618) );
  NAND2_X1 U2441 ( .A1(n4381), .A2(REG1_REG_15__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U2442 ( .A1(n2762), .A2(DATAI_22_), .ZN(n4235) );
  NAND2_X1 U2443 ( .A1(n2491), .A2(n4905), .ZN(n4904) );
  NOR2_X1 U2444 ( .A1(n3163), .A2(n2484), .ZN(n2483) );
  NAND2_X1 U2445 ( .A1(n4725), .A2(n4719), .ZN(n4718) );
  AOI21_X1 U2446 ( .B1(n3240), .B2(n4891), .A(n2360), .ZN(n3961) );
  NAND2_X1 U2447 ( .A1(n2361), .A2(n2307), .ZN(n2360) );
  NOR2_X1 U2448 ( .A1(n4144), .A2(n3249), .ZN(n4120) );
  NAND2_X1 U2449 ( .A1(n4120), .A2(n3740), .ZN(n4288) );
  XNOR2_X1 U2450 ( .A(n2668), .B(n3956), .ZN(n2676) );
  NAND2_X1 U2451 ( .A1(n2671), .A2(IR_REG_31__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U2452 ( .A1(n2672), .A2(n2671), .ZN(n2674) );
  NOR2_X1 U2453 ( .A1(n2556), .A2(IR_REG_5__SCAN_IN), .ZN(n2571) );
  INV_X1 U2454 ( .A(IR_REG_3__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U2455 ( .A1(n4704), .A2(n2322), .ZN(n2323) );
  NAND2_X1 U2456 ( .A1(n2456), .A2(n2454), .ZN(n3949) );
  AND2_X1 U2457 ( .A1(n2455), .A2(n4042), .ZN(n2454) );
  NAND2_X1 U2458 ( .A1(n2854), .A2(n2853), .ZN(n3581) );
  NOR2_X1 U2459 ( .A1(n3991), .A2(n3990), .ZN(n2334) );
  INV_X1 U2460 ( .A(n4008), .ZN(n2333) );
  NOR2_X1 U2461 ( .A1(n4044), .A2(n3991), .ZN(n2331) );
  AND2_X1 U2462 ( .A1(n3131), .A2(n3130), .ZN(n4966) );
  NAND4_X1 U2463 ( .A1(n3062), .A2(n3061), .A3(n3060), .A4(n3059), .ZN(n4175)
         );
  NOR2_X1 U2464 ( .A1(n4603), .A2(n4704), .ZN(n2402) );
  NOR2_X1 U2465 ( .A1(n4607), .A2(n4606), .ZN(n4605) );
  XNOR2_X1 U2466 ( .A(n2639), .B(n4624), .ZN(n4616) );
  NAND2_X1 U2467 ( .A1(n3386), .A2(REG2_REG_8__SCAN_IN), .ZN(n3385) );
  NAND2_X1 U2468 ( .A1(n3385), .A2(n2645), .ZN(n4634) );
  XNOR2_X1 U2469 ( .A(n2647), .B(n4813), .ZN(n4639) );
  NAND2_X1 U2470 ( .A1(n4639), .A2(REG2_REG_10__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U2471 ( .A1(n4640), .A2(n2606), .ZN(n4648) );
  XNOR2_X1 U2472 ( .A(n2610), .B(n2609), .ZN(n4658) );
  NOR2_X1 U2473 ( .A1(n4658), .A2(n4659), .ZN(n4657) );
  XNOR2_X1 U2474 ( .A(n2614), .B(n4690), .ZN(n4687) );
  NAND2_X1 U2475 ( .A1(n4687), .A2(REG1_REG_14__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U2476 ( .A1(n4081), .A2(n2617), .ZN(n4080) );
  XNOR2_X1 U2477 ( .A(n2618), .B(n2940), .ZN(n4699) );
  INV_X1 U2478 ( .A(n2388), .ZN(n2384) );
  AOI21_X1 U2479 ( .B1(n4697), .B2(ADDR_REG_18__SCAN_IN), .A(n4105), .ZN(n2388) );
  NAND2_X1 U2480 ( .A1(n4601), .A2(n3325), .ZN(n4703) );
  XNOR2_X1 U2481 ( .A(n2625), .B(n2624), .ZN(n2393) );
  AND2_X1 U2482 ( .A1(n4601), .A2(n3886), .ZN(n4698) );
  AOI21_X1 U2483 ( .B1(n4095), .B2(n2386), .A(n2309), .ZN(n2661) );
  INV_X1 U2484 ( .A(n2630), .ZN(n2396) );
  OR2_X1 U2485 ( .A1(n3962), .A2(n4280), .ZN(n2347) );
  NAND2_X1 U2486 ( .A1(n4972), .A2(REG2_REG_29__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U2487 ( .A1(n3961), .A2(n2350), .ZN(n2349) );
  NAND2_X1 U2488 ( .A1(n3959), .A2(n4917), .ZN(n2350) );
  AND2_X1 U2489 ( .A1(n2341), .A2(n2303), .ZN(n2340) );
  NOR2_X1 U2490 ( .A1(n4203), .A2(n4202), .ZN(n2476) );
  XNOR2_X1 U2491 ( .A(n2397), .B(IR_REG_0__SCAN_IN), .ZN(n4473) );
  INV_X1 U2492 ( .A(keyinput_119), .ZN(n2397) );
  INV_X1 U2493 ( .A(IR_REG_6__SCAN_IN), .ZN(n4572) );
  INV_X1 U2494 ( .A(IR_REG_19__SCAN_IN), .ZN(n2508) );
  INV_X1 U2495 ( .A(n2442), .ZN(n2440) );
  AND2_X1 U2496 ( .A1(n2506), .A2(n2547), .ZN(n2507) );
  AND2_X1 U2497 ( .A1(n2369), .A2(n3867), .ZN(n2368) );
  OR2_X1 U2498 ( .A1(n3744), .A2(n3863), .ZN(n2369) );
  OR2_X1 U2499 ( .A1(n4187), .A2(n3766), .ZN(n2371) );
  INV_X1 U2500 ( .A(n2746), .ZN(n2762) );
  INV_X1 U2501 ( .A(n3461), .ZN(n3767) );
  INV_X1 U2502 ( .A(n3239), .ZN(n2361) );
  AOI21_X1 U2503 ( .B1(n3483), .B2(n3832), .A(n3836), .ZN(n4778) );
  NAND2_X1 U2504 ( .A1(n2522), .A2(n2492), .ZN(n2526) );
  INV_X1 U2505 ( .A(IR_REG_22__SCAN_IN), .ZN(n2520) );
  OR2_X1 U2506 ( .A1(n3648), .A2(n2342), .ZN(n2341) );
  INV_X1 U2507 ( .A(n3647), .ZN(n2342) );
  NOR2_X1 U2508 ( .A1(n2913), .A2(n3647), .ZN(n2343) );
  NOR2_X1 U2509 ( .A1(n3738), .A2(n3092), .ZN(n3249) );
  INV_X1 U2510 ( .A(n2772), .ZN(n2336) );
  INV_X1 U2511 ( .A(n2771), .ZN(n2335) );
  INV_X1 U2512 ( .A(n3985), .ZN(n3988) );
  NOR2_X1 U2513 ( .A1(n3738), .A2(n3036), .ZN(n4012) );
  AOI21_X1 U2514 ( .B1(n4063), .B2(n2737), .A(n2768), .ZN(n2772) );
  NOR2_X1 U2515 ( .A1(n3421), .A2(n2767), .ZN(n2768) );
  INV_X1 U2516 ( .A(n2741), .ZN(n2412) );
  AOI21_X1 U2517 ( .B1(n4064), .B2(n2737), .A(n2747), .ZN(n2752) );
  NAND2_X1 U2518 ( .A1(n2770), .A2(n2769), .ZN(n3389) );
  AND2_X1 U2519 ( .A1(REG3_REG_19__SCAN_IN), .A2(n2972), .ZN(n2973) );
  AND2_X1 U2520 ( .A1(n2304), .A2(n2424), .ZN(n2423) );
  INV_X1 U2521 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2871) );
  NOR2_X1 U2522 ( .A1(n2872), .A2(n2871), .ZN(n2886) );
  AOI21_X1 U2523 ( .B1(n4066), .B2(n2737), .A(n2718), .ZN(n2723) );
  XNOR2_X1 U2524 ( .A(n2735), .B(n3066), .ZN(n2740) );
  AOI21_X1 U2525 ( .B1(n4065), .B2(n2737), .A(n2736), .ZN(n2739) );
  AND2_X1 U2526 ( .A1(n3477), .A2(n2766), .ZN(n2736) );
  NAND2_X1 U2527 ( .A1(n2413), .A2(n2738), .ZN(n3297) );
  INV_X1 U2528 ( .A(n3299), .ZN(n2413) );
  NAND2_X1 U2529 ( .A1(n2462), .A2(n2461), .ZN(n2458) );
  NAND2_X1 U2530 ( .A1(n3056), .A2(n2296), .ZN(n2461) );
  NAND2_X1 U2531 ( .A1(n2462), .A2(n2460), .ZN(n2459) );
  INV_X1 U2532 ( .A(n3977), .ZN(n2460) );
  OR2_X1 U2533 ( .A1(n3042), .A2(n4483), .ZN(n3057) );
  AND2_X1 U2534 ( .A1(n3889), .A2(n3800), .ZN(n3237) );
  NAND2_X1 U2535 ( .A1(n2507), .A2(n2443), .ZN(n2442) );
  AOI21_X1 U2536 ( .B1(n4069), .B2(n3938), .A(n3939), .ZN(n3937) );
  NAND2_X1 U2537 ( .A1(n4072), .A2(n2633), .ZN(n3935) );
  NAND2_X1 U2538 ( .A1(n3936), .A2(n3935), .ZN(n3934) );
  XNOR2_X1 U2539 ( .A(n2637), .B(n3316), .ZN(n3309) );
  NAND2_X1 U2540 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U2541 ( .A1(n3309), .A2(REG2_REG_4__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U2542 ( .A1(n4620), .A2(n2591), .ZN(n3291) );
  OAI21_X1 U2543 ( .B1(n4630), .B2(n4625), .A(n4627), .ZN(n2605) );
  NAND2_X1 U2544 ( .A1(n2391), .A2(REG1_REG_10__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U2545 ( .A1(n4652), .A2(n2649), .ZN(n2650) );
  NAND2_X1 U2546 ( .A1(n2318), .A2(n2317), .ZN(n4082) );
  OAI21_X1 U2547 ( .B1(n2653), .B2(REG2_REG_14__SCAN_IN), .A(n2378), .ZN(n2376) );
  NAND2_X1 U2548 ( .A1(n4082), .A2(n2654), .ZN(n2316) );
  OR2_X1 U2549 ( .A1(n4380), .A2(REG2_REG_17__SCAN_IN), .ZN(n2390) );
  NOR2_X1 U2550 ( .A1(n4104), .A2(n2387), .ZN(n2386) );
  INV_X1 U2551 ( .A(n2390), .ZN(n2387) );
  AND2_X1 U2552 ( .A1(n2629), .A2(n2627), .ZN(n4601) );
  NAND2_X1 U2553 ( .A1(n2364), .A2(n2362), .ZN(n4124) );
  AOI21_X1 U2554 ( .B1(n2365), .B2(n2370), .A(n2363), .ZN(n2362) );
  INV_X1 U2555 ( .A(n3741), .ZN(n2363) );
  AND2_X1 U2556 ( .A1(n3742), .A2(n3746), .ZN(n4123) );
  NAND2_X1 U2557 ( .A1(n2367), .A2(n2368), .ZN(n4134) );
  OR2_X1 U2558 ( .A1(n4187), .A2(n2370), .ZN(n2367) );
  OR2_X1 U2559 ( .A1(n3057), .A2(n4045), .ZN(n3085) );
  NOR2_X1 U2560 ( .A1(n4159), .A2(n3191), .ZN(n3192) );
  AOI21_X1 U2561 ( .B1(n2470), .B2(n2472), .A(n2285), .ZN(n2468) );
  INV_X1 U2562 ( .A(n4232), .ZN(n4188) );
  NAND2_X1 U2563 ( .A1(n2986), .A2(REG3_REG_21__SCAN_IN), .ZN(n3016) );
  NAND2_X1 U2564 ( .A1(n4244), .A2(n3189), .ZN(n2475) );
  INV_X1 U2565 ( .A(n2374), .ZN(n4210) );
  OAI21_X1 U2566 ( .B1(n4246), .B2(n3784), .A(n3851), .ZN(n2374) );
  AOI21_X1 U2567 ( .B1(n2490), .B2(n2488), .A(n2298), .ZN(n2487) );
  INV_X1 U2568 ( .A(n2490), .ZN(n2489) );
  INV_X1 U2569 ( .A(n3184), .ZN(n2488) );
  NAND2_X1 U2570 ( .A1(n2946), .A2(REG3_REG_17__SCAN_IN), .ZN(n2958) );
  NAND2_X1 U2571 ( .A1(n4892), .A2(n3218), .ZN(n3897) );
  INV_X1 U2572 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4691) );
  NOR2_X1 U2573 ( .A1(n2935), .A2(n4691), .ZN(n2946) );
  INV_X1 U2574 ( .A(n4054), .ZN(n4902) );
  NAND2_X1 U2575 ( .A1(n3616), .A2(n2355), .ZN(n4890) );
  AND2_X1 U2576 ( .A1(n2267), .A2(n4857), .ZN(n2355) );
  OR2_X1 U2577 ( .A1(n2917), .A2(n2690), .ZN(n2935) );
  OR2_X1 U2578 ( .A1(n3660), .A2(n3788), .ZN(n3658) );
  OAI21_X1 U2579 ( .B1(n3509), .B2(n3841), .A(n3843), .ZN(n3627) );
  OR2_X1 U2580 ( .A1(n2855), .A2(n4486), .ZN(n2872) );
  INV_X1 U2581 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U2582 ( .A1(n2486), .A2(n3170), .ZN(n3626) );
  OR2_X1 U2583 ( .A1(n2838), .A2(n2837), .ZN(n2855) );
  NAND2_X1 U2584 ( .A1(n2373), .A2(n3802), .ZN(n3509) );
  NAND2_X1 U2585 ( .A1(n3534), .A2(n3842), .ZN(n2373) );
  AOI21_X1 U2586 ( .B1(n2480), .B2(n2478), .A(n2273), .ZN(n2477) );
  INV_X1 U2587 ( .A(n2480), .ZN(n2479) );
  OAI21_X1 U2588 ( .B1(n3370), .B2(n3369), .A(n3805), .ZN(n3483) );
  NAND2_X1 U2589 ( .A1(n2372), .A2(n3833), .ZN(n3370) );
  NAND2_X1 U2590 ( .A1(n3417), .A2(n3828), .ZN(n2372) );
  INV_X1 U2591 ( .A(n3409), .ZN(n3421) );
  NAND2_X1 U2592 ( .A1(n3878), .A2(n4705), .ZN(n4780) );
  INV_X1 U2593 ( .A(n4065), .ZN(n4723) );
  OR2_X1 U2594 ( .A1(n4725), .A2(n4724), .ZN(n4727) );
  NOR2_X1 U2595 ( .A1(n4288), .A2(n4289), .ZN(n4287) );
  INV_X1 U2596 ( .A(n4780), .ZN(n4896) );
  NAND2_X1 U2597 ( .A1(n4195), .A2(n2269), .ZN(n4144) );
  NOR2_X1 U2598 ( .A1(n3738), .A2(n3063), .ZN(n4160) );
  NAND2_X1 U2599 ( .A1(n4195), .A2(n2354), .ZN(n4162) );
  NAND2_X1 U2600 ( .A1(n4195), .A2(n3191), .ZN(n4178) );
  AND2_X1 U2601 ( .A1(n4219), .A2(n4193), .ZN(n4195) );
  INV_X1 U2602 ( .A(n4012), .ZN(n4193) );
  OR2_X1 U2603 ( .A1(n4942), .A2(n4239), .ZN(n2352) );
  NOR2_X1 U2604 ( .A1(n4319), .A2(n3971), .ZN(n4219) );
  INV_X1 U2605 ( .A(n4959), .ZN(n3926) );
  NOR3_X1 U2606 ( .A1(n4265), .A2(n4942), .A3(n4926), .ZN(n4256) );
  OR2_X1 U2607 ( .A1(n4264), .A2(n4036), .ZN(n4265) );
  NOR2_X1 U2608 ( .A1(n4265), .A2(n4926), .ZN(n4254) );
  NOR2_X1 U2609 ( .A1(n4890), .A2(n4895), .ZN(n4889) );
  INV_X1 U2610 ( .A(n4001), .ZN(n3706) );
  NAND2_X1 U2611 ( .A1(n3616), .A2(n2267), .ZN(n3676) );
  NAND2_X1 U2612 ( .A1(n3616), .A2(n3615), .ZN(n3675) );
  AND2_X1 U2613 ( .A1(n3588), .A2(n4587), .ZN(n3616) );
  INV_X1 U2614 ( .A(n3209), .ZN(n4587) );
  NOR2_X1 U2615 ( .A1(n3623), .A2(n3594), .ZN(n3588) );
  OR2_X1 U2616 ( .A1(n3622), .A2(n3628), .ZN(n3623) );
  INV_X1 U2617 ( .A(n3523), .ZN(n3514) );
  OR2_X1 U2618 ( .A1(n4775), .A2(n4774), .ZN(n4776) );
  NOR2_X1 U2619 ( .A1(n4776), .A2(n3501), .ZN(n3530) );
  OR2_X1 U2620 ( .A1(n3375), .A2(n3454), .ZN(n4775) );
  NOR2_X1 U2621 ( .A1(n3410), .A2(n3409), .ZN(n3413) );
  AND2_X1 U2622 ( .A1(n4730), .A2(n3469), .ZN(n3475) );
  AND3_X1 U2623 ( .A1(n3430), .A2(n3244), .A3(n3428), .ZN(n3251) );
  INV_X1 U2624 ( .A(n3145), .ZN(n3268) );
  NAND2_X1 U2625 ( .A1(n3099), .A2(n3269), .ZN(n3267) );
  NAND2_X1 U2626 ( .A1(n2345), .A2(IR_REG_31__SCAN_IN), .ZN(n2626) );
  INV_X1 U2627 ( .A(IR_REG_25__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U2628 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U2629 ( .A1(n2441), .A2(IR_REG_31__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U2630 ( .A1(n2553), .A2(n2271), .ZN(n2441) );
  NAND2_X1 U2631 ( .A1(n2553), .A2(n2552), .ZN(n2554) );
  AND2_X1 U2632 ( .A1(n2573), .A2(n2572), .ZN(n2783) );
  AND2_X1 U2633 ( .A1(n2453), .A2(n3451), .ZN(n3965) );
  NAND2_X1 U2634 ( .A1(n2805), .A2(n2497), .ZN(n2453) );
  NAND2_X1 U2635 ( .A1(n3012), .A2(n3011), .ZN(n3013) );
  INV_X1 U2636 ( .A(n3009), .ZN(n3012) );
  INV_X1 U2637 ( .A(n2344), .ZN(n3974) );
  OAI21_X1 U2638 ( .B1(n2805), .B2(n2450), .A(n2448), .ZN(n3499) );
  XNOR2_X1 U2639 ( .A(n2722), .B(n2723), .ZN(n2410) );
  NOR2_X1 U2640 ( .A1(n3738), .A2(n2993), .ZN(n4959) );
  OAI21_X1 U2641 ( .B1(n3579), .B2(n2263), .A(n2424), .ZN(n4585) );
  AND2_X1 U2642 ( .A1(n4863), .A2(n4866), .ZN(n2434) );
  NAND2_X1 U2643 ( .A1(n2300), .A2(n2432), .ZN(n4000) );
  NAND2_X1 U2644 ( .A1(n2445), .A2(n2325), .ZN(n3522) );
  AOI21_X1 U2645 ( .B1(n2447), .B2(n2448), .A(n2446), .ZN(n2445) );
  INV_X1 U2646 ( .A(n3497), .ZN(n2446) );
  NAND2_X1 U2647 ( .A1(n2746), .A2(IR_REG_0__SCAN_IN), .ZN(n2398) );
  AND2_X1 U2648 ( .A1(n3144), .A2(n3138), .ZN(n4948) );
  NAND2_X1 U2649 ( .A1(n3579), .A2(n2870), .ZN(n3573) );
  INV_X1 U2650 ( .A(n3477), .ZN(n3469) );
  AND2_X1 U2651 ( .A1(n3144), .A2(n3143), .ZN(n4957) );
  NAND4_X1 U2652 ( .A1(n2980), .A2(n2979), .A3(n2978), .A4(n2977), .ZN(n4958)
         );
  NAND4_X1 U2653 ( .A1(n2680), .A2(n2679), .A3(n2678), .A4(n2677), .ZN(n4944)
         );
  NAND4_X1 U2654 ( .A1(n2701), .A2(n2700), .A3(n2699), .A4(n2698), .ZN(n4721)
         );
  NAND2_X1 U2655 ( .A1(n4070), .A2(n4071), .ZN(n4069) );
  XNOR2_X1 U2656 ( .A(n2635), .B(n3279), .ZN(n3282) );
  AND2_X1 U2657 ( .A1(n3313), .A2(n2379), .ZN(n4607) );
  NAND2_X1 U2658 ( .A1(n2637), .A2(n4384), .ZN(n2379) );
  XNOR2_X1 U2659 ( .A(n2590), .B(n4624), .ZN(n4621) );
  NAND2_X1 U2660 ( .A1(n4621), .A2(REG1_REG_6__SCAN_IN), .ZN(n4620) );
  INV_X1 U2661 ( .A(n2380), .ZN(n4615) );
  AND2_X1 U2662 ( .A1(n2380), .A2(n2292), .ZN(n3288) );
  NAND2_X1 U2663 ( .A1(n2404), .A2(n2406), .ZN(n3382) );
  NOR2_X1 U2664 ( .A1(n2405), .A2(n2599), .ZN(n3381) );
  INV_X1 U2665 ( .A(n2404), .ZN(n2599) );
  NAND2_X1 U2666 ( .A1(n4638), .A2(n2648), .ZN(n4653) );
  NAND2_X1 U2667 ( .A1(n4653), .A2(n4654), .ZN(n4652) );
  NOR2_X1 U2668 ( .A1(n4657), .A2(n2611), .ZN(n4669) );
  NOR2_X1 U2669 ( .A1(n4682), .A2(n4683), .ZN(n4681) );
  NAND2_X1 U2670 ( .A1(n4686), .A2(n2615), .ZN(n4081) );
  XNOR2_X1 U2671 ( .A(n2316), .B(n2315), .ZN(n4695) );
  NAND2_X1 U2672 ( .A1(n4695), .A2(n4693), .ZN(n4694) );
  NOR2_X1 U2673 ( .A1(n4700), .A2(n2619), .ZN(n4093) );
  INV_X1 U2674 ( .A(n2324), .ZN(n4091) );
  INV_X1 U2675 ( .A(n2622), .ZN(n4106) );
  NOR2_X1 U2676 ( .A1(n2384), .A2(n2383), .ZN(n2382) );
  INV_X1 U2677 ( .A(n2386), .ZN(n2383) );
  AND2_X1 U2678 ( .A1(n4663), .A2(n2308), .ZN(n2385) );
  NOR2_X1 U2679 ( .A1(n4703), .A2(n4787), .ZN(n2395) );
  NAND2_X1 U2680 ( .A1(n2464), .A2(n2465), .ZN(n4143) );
  NAND2_X1 U2681 ( .A1(n4904), .A2(n3184), .ZN(n3702) );
  INV_X1 U2682 ( .A(n4968), .ZN(n4259) );
  NAND2_X1 U2683 ( .A1(n2482), .A2(n3164), .ZN(n3482) );
  NAND2_X1 U2684 ( .A1(n3162), .A2(n2483), .ZN(n2482) );
  AND2_X1 U2685 ( .A1(n4825), .A2(n3435), .ZN(n4832) );
  AND2_X2 U2686 ( .A1(n3251), .A2(n3245), .ZN(n4911) );
  INV_X1 U2687 ( .A(n4911), .ZN(n4909) );
  INV_X1 U2688 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2357) );
  NAND2_X1 U2689 ( .A1(n3961), .A2(n2358), .ZN(n3252) );
  NAND2_X1 U2690 ( .A1(n2359), .A2(n4877), .ZN(n2358) );
  INV_X1 U2691 ( .A(n3962), .ZN(n2359) );
  INV_X1 U2692 ( .A(n3257), .ZN(n3270) );
  NAND2_X1 U2693 ( .A1(n3268), .A2(n3267), .ZN(n4389) );
  INV_X1 U2694 ( .A(IR_REG_30__SCAN_IN), .ZN(n3956) );
  AND2_X1 U2695 ( .A1(n2665), .A2(n2664), .ZN(n2666) );
  INV_X1 U2696 ( .A(IR_REG_29__SCAN_IN), .ZN(n2665) );
  AND2_X1 U2697 ( .A1(n2585), .A2(n2582), .ZN(n4385) );
  NAND2_X1 U2698 ( .A1(n2323), .A2(IR_REG_31__SCAN_IN), .ZN(n2576) );
  XNOR2_X1 U2699 ( .A(n2311), .B(IR_REG_1__SCAN_IN), .ZN(n4387) );
  NAND2_X1 U2700 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2311)
         );
  OAI21_X1 U2701 ( .B1(n2330), .B2(n3975), .A(n2329), .ZN(U3222) );
  INV_X1 U2702 ( .A(n3996), .ZN(n2329) );
  AOI21_X1 U2703 ( .B1(n3989), .B2(n2332), .A(n2331), .ZN(n2330) );
  NAND2_X1 U2704 ( .A1(n4602), .A2(n2400), .ZN(U3240) );
  NOR2_X1 U2705 ( .A1(n2402), .A2(n2401), .ZN(n2400) );
  NOR2_X1 U2706 ( .A1(n4604), .A2(IR_REG_0__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U2707 ( .A1(n4634), .A2(n4635), .ZN(n4633) );
  NOR2_X1 U2708 ( .A1(n2396), .A2(n2395), .ZN(n2394) );
  NAND2_X1 U2709 ( .A1(n2393), .A2(n4698), .ZN(n2392) );
  OAI21_X1 U2710 ( .B1(n2348), .B2(n4972), .A(n2289), .ZN(U3354) );
  AOI21_X1 U2711 ( .B1(n3960), .B2(n4968), .A(n2349), .ZN(n2348) );
  INV_X1 U2712 ( .A(n2767), .ZN(n3078) );
  AND2_X1 U2713 ( .A1(n2475), .A2(n2275), .ZN(n3921) );
  AND2_X1 U2714 ( .A1(n3571), .A2(n3570), .ZN(n2263) );
  AND2_X1 U2715 ( .A1(n2271), .A2(n2507), .ZN(n2264) );
  OR2_X1 U2716 ( .A1(n4232), .A2(n3971), .ZN(n2265) );
  OR3_X1 U2717 ( .A1(n4265), .A2(n2353), .A3(n4942), .ZN(n2266) );
  AND2_X1 U2718 ( .A1(n3615), .A2(n3683), .ZN(n2267) );
  INV_X1 U2719 ( .A(n4903), .ZN(n2491) );
  NAND2_X1 U2720 ( .A1(n2435), .A2(n2944), .ZN(n2268) );
  AND2_X1 U2721 ( .A1(n2354), .A2(n4145), .ZN(n2269) );
  OR2_X1 U2722 ( .A1(n2384), .A2(n2385), .ZN(n2270) );
  INV_X1 U2723 ( .A(n2940), .ZN(n2315) );
  INV_X1 U2724 ( .A(n4663), .ZN(n4692) );
  AND2_X1 U2725 ( .A1(n4601), .A2(n2662), .ZN(n4663) );
  NAND3_X1 U2726 ( .A1(n3269), .A2(n3270), .A3(n4378), .ZN(n2704) );
  AND2_X1 U2727 ( .A1(n3263), .A2(n2674), .ZN(n2711) );
  XNOR2_X1 U2728 ( .A(n2683), .B(n2682), .ZN(n2687) );
  AND2_X1 U2729 ( .A1(n2552), .A2(n2444), .ZN(n2271) );
  NOR2_X1 U2730 ( .A1(n3193), .A2(n3192), .ZN(n2272) );
  INV_X1 U2731 ( .A(n3400), .ZN(n2418) );
  AND2_X1 U2732 ( .A1(n4783), .A2(n3454), .ZN(n2273) );
  NAND2_X1 U2733 ( .A1(n2519), .A2(n2518), .ZN(n2746) );
  OR2_X1 U2734 ( .A1(n3401), .A2(n3400), .ZN(n2274) );
  XNOR2_X1 U2735 ( .A(n2721), .B(n2734), .ZN(n2722) );
  NAND2_X1 U2736 ( .A1(n4958), .A2(n4942), .ZN(n2275) );
  NOR2_X1 U2737 ( .A1(n4140), .A2(n3227), .ZN(n2276) );
  AND2_X1 U2738 ( .A1(n2339), .A2(n2337), .ZN(n2277) );
  INV_X1 U2739 ( .A(n2451), .ZN(n2450) );
  NAND2_X1 U2740 ( .A1(n4058), .A2(n3628), .ZN(n2278) );
  AND2_X1 U2741 ( .A1(n2821), .A2(n2820), .ZN(n2279) );
  OR2_X1 U2742 ( .A1(n3321), .A2(n2734), .ZN(n2280) );
  AND2_X1 U2743 ( .A1(n2783), .A2(REG2_REG_5__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2744 ( .A1(n4201), .A2(n2275), .ZN(n2282) );
  AND2_X1 U2745 ( .A1(n2476), .A2(n3189), .ZN(n2283) );
  NOR2_X1 U2746 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2284)
         );
  NOR2_X1 U2747 ( .A1(n4188), .A2(n4221), .ZN(n2285) );
  INV_X1 U2748 ( .A(n2466), .ZN(n2465) );
  NOR2_X1 U2749 ( .A1(n4175), .A2(n4160), .ZN(n2466) );
  AND2_X1 U2750 ( .A1(n4902), .A2(n3706), .ZN(n2286) );
  AND2_X1 U2751 ( .A1(n2515), .A2(n2514), .ZN(n2522) );
  NAND2_X1 U2752 ( .A1(n2522), .A2(n2524), .ZN(n2287) );
  AND2_X1 U2753 ( .A1(n2436), .A2(n2442), .ZN(n2288) );
  AND2_X1 U2754 ( .A1(n2347), .A2(n2346), .ZN(n2289) );
  NAND2_X1 U2755 ( .A1(n2663), .A2(n4663), .ZN(n2290) );
  OR2_X1 U2756 ( .A1(n2276), .A2(n3192), .ZN(n2291) );
  OR2_X1 U2757 ( .A1(n2639), .A2(n4624), .ZN(n2292) );
  AND2_X1 U2758 ( .A1(n2769), .A2(n2274), .ZN(n2293) );
  AND4_X1 U2759 ( .A1(n2716), .A2(n2715), .A3(n2713), .A4(n2714), .ZN(n3156)
         );
  INV_X1 U2760 ( .A(IR_REG_16__SCAN_IN), .ZN(n2444) );
  AND2_X1 U2761 ( .A1(n2492), .A2(n2284), .ZN(n2294) );
  AND2_X1 U2762 ( .A1(n2371), .A2(n3863), .ZN(n2295) );
  INV_X1 U2763 ( .A(IR_REG_27__SCAN_IN), .ZN(n2540) );
  OR2_X1 U2764 ( .A1(n3028), .A2(n3027), .ZN(n2296) );
  OAI21_X1 U2765 ( .B1(n3650), .B2(n2343), .A(n2341), .ZN(n3692) );
  OR2_X1 U2766 ( .A1(n3070), .A2(n3069), .ZN(n2297) );
  AND2_X1 U2767 ( .A1(n4054), .A2(n4001), .ZN(n2298) );
  NOR3_X1 U2768 ( .A1(n4265), .A2(n2352), .A3(n2353), .ZN(n2351) );
  INV_X1 U2769 ( .A(n4882), .ZN(n2433) );
  OR2_X1 U2770 ( .A1(n3998), .A2(n2957), .ZN(n2299) );
  INV_X1 U2771 ( .A(IR_REG_31__SCAN_IN), .ZN(n2443) );
  AND2_X1 U2772 ( .A1(n2431), .A2(n2268), .ZN(n2300) );
  NOR2_X1 U2773 ( .A1(n2434), .A2(n4865), .ZN(n2301) );
  NOR2_X1 U2774 ( .A1(n4681), .A2(n2653), .ZN(n2302) );
  INV_X1 U2775 ( .A(n4942), .ZN(n4253) );
  INV_X1 U2776 ( .A(n2737), .ZN(n2689) );
  NAND2_X1 U2777 ( .A1(n3389), .A2(n2773), .ZN(n3399) );
  NAND2_X1 U2778 ( .A1(n2453), .A2(n2451), .ZN(n3963) );
  OR2_X1 U2779 ( .A1(n3581), .A2(n3582), .ZN(n3579) );
  INV_X1 U2780 ( .A(n4905), .ZN(n4893) );
  OR2_X1 U2781 ( .A1(n3848), .A2(n3854), .ZN(n4905) );
  NAND2_X1 U2782 ( .A1(n2927), .A2(n2928), .ZN(n2303) );
  NAND2_X1 U2783 ( .A1(n2898), .A2(n2899), .ZN(n2304) );
  NAND2_X1 U2784 ( .A1(n2667), .A2(n2545), .ZN(n2305) );
  OR2_X1 U2785 ( .A1(n2384), .A2(n2389), .ZN(n2306) );
  INV_X1 U2786 ( .A(n2805), .ZN(n3450) );
  INV_X1 U2787 ( .A(DATAI_0_), .ZN(n2399) );
  AND2_X2 U2788 ( .A1(n3251), .A2(n3429), .ZN(n4915) );
  NOR2_X1 U2789 ( .A1(n3738), .A2(n3076), .ZN(n4136) );
  NAND2_X1 U2790 ( .A1(n3297), .A2(n2741), .ZN(n3342) );
  INV_X1 U2791 ( .A(n4104), .ZN(n2389) );
  AND2_X1 U2792 ( .A1(n3358), .A2(n4251), .ZN(n4906) );
  INV_X1 U2793 ( .A(n4906), .ZN(n4877) );
  INV_X1 U2794 ( .A(n3496), .ZN(n2326) );
  OR2_X1 U2795 ( .A1(n3753), .A2(n4113), .ZN(n2307) );
  OR2_X1 U2796 ( .A1(n2389), .A2(n2390), .ZN(n2308) );
  AND2_X1 U2797 ( .A1(n3259), .A2(REG2_REG_18__SCAN_IN), .ZN(n2309) );
  OR2_X1 U2798 ( .A1(n4380), .A2(REG1_REG_17__SCAN_IN), .ZN(n2310) );
  INV_X1 U2799 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2408) );
  XNOR2_X1 U2800 ( .A(n4387), .B(n2632), .ZN(n4074) );
  NAND2_X1 U2801 ( .A1(n2377), .A2(n4682), .ZN(n2317) );
  INV_X1 U2802 ( .A(n2376), .ZN(n2318) );
  INV_X1 U2803 ( .A(IR_REG_1__SCAN_IN), .ZN(n2322) );
  NAND3_X1 U2804 ( .A1(n2448), .A2(n2805), .A3(n2326), .ZN(n2325) );
  AND2_X2 U2805 ( .A1(n2415), .A2(n2416), .ZN(n2805) );
  NOR2_X2 U2806 ( .A1(n2579), .A2(n2328), .ZN(n2514) );
  MUX2_X1 U2807 ( .A(n4384), .B(DATAI_4_), .S(n2762), .Z(n3409) );
  NAND3_X1 U2808 ( .A1(n2375), .A2(n2515), .A3(n2541), .ZN(n2345) );
  NAND2_X1 U2809 ( .A1(n2375), .A2(n2515), .ZN(n2543) );
  INV_X1 U2810 ( .A(n2351), .ZN(n4319) );
  NAND2_X1 U2811 ( .A1(n4912), .A2(n2357), .ZN(n2356) );
  NAND2_X1 U2812 ( .A1(n4187), .A2(n2365), .ZN(n2364) );
  INV_X1 U2813 ( .A(n2371), .ZN(n4170) );
  NAND2_X2 U2814 ( .A1(n3824), .A2(n3821), .ZN(n4725) );
  NAND3_X1 U2815 ( .A1(n2375), .A2(n2515), .A3(n2666), .ZN(n2671) );
  NAND2_X1 U2816 ( .A1(n4095), .A2(n2382), .ZN(n2381) );
  OAI211_X1 U2817 ( .C1(n4095), .C2(n2306), .A(n2270), .B(n2381), .ZN(n4110)
         );
  NAND2_X1 U2818 ( .A1(n3215), .A2(n3813), .ZN(n3725) );
  MUX2_X1 U2819 ( .A(DATAI_1_), .B(n4387), .S(n2746), .Z(n4731) );
  OAI211_X1 U2820 ( .C1(n2391), .C2(REG1_REG_10__SCAN_IN), .A(n4640), .B(n4698), .ZN(n4641) );
  XNOR2_X1 U2821 ( .A(n2605), .B(n4813), .ZN(n2391) );
  NAND3_X1 U2822 ( .A1(n2290), .A2(n2394), .A3(n2392), .ZN(U3259) );
  INV_X2 U2823 ( .A(IR_REG_0__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U2824 ( .A1(n2597), .A2(n2598), .ZN(n2406) );
  OAI211_X1 U2825 ( .C1(n3332), .C2(n2410), .A(n3331), .B(n4961), .ZN(n3335)
         );
  NAND2_X1 U2826 ( .A1(n3332), .A2(n2410), .ZN(n3331) );
  NAND2_X1 U2827 ( .A1(n4066), .A2(n2766), .ZN(n2720) );
  AND2_X2 U2828 ( .A1(n3434), .A2(n2704), .ZN(n2766) );
  OAI211_X1 U2829 ( .C1(n2738), .C2(n2412), .A(n2411), .B(n3343), .ZN(n2755)
         );
  NAND2_X1 U2830 ( .A1(n3299), .A2(n2741), .ZN(n2411) );
  NAND2_X1 U2831 ( .A1(n2514), .A2(n2513), .ZN(n2505) );
  NAND2_X1 U2832 ( .A1(n2770), .A2(n2293), .ZN(n2415) );
  NAND3_X1 U2833 ( .A1(n2304), .A2(n2424), .A3(n2263), .ZN(n2421) );
  NAND3_X1 U2834 ( .A1(n2431), .A2(n2432), .A3(n2426), .ZN(n2428) );
  NAND2_X1 U2835 ( .A1(n4865), .A2(n2433), .ZN(n2431) );
  AOI21_X2 U2836 ( .B1(n4033), .B2(n4030), .A(n4029), .ZN(n4929) );
  NAND2_X1 U2837 ( .A1(n2428), .A2(n2427), .ZN(n4033) );
  OAI21_X1 U2838 ( .B1(n3976), .B2(n2459), .A(n2458), .ZN(n4044) );
  NAND3_X1 U2839 ( .A1(n2458), .A2(n2459), .A3(n2297), .ZN(n2455) );
  NAND2_X1 U2840 ( .A1(n3976), .A2(n2457), .ZN(n2456) );
  NAND2_X1 U2841 ( .A1(n4244), .A2(n2470), .ZN(n2469) );
  OAI21_X2 U2842 ( .B1(n3162), .B2(n2479), .A(n2477), .ZN(n4788) );
  NAND2_X1 U2843 ( .A1(n3162), .A2(n3161), .ZN(n3368) );
  INV_X1 U2844 ( .A(n3161), .ZN(n2484) );
  NAND2_X1 U2845 ( .A1(n2486), .A2(n2485), .ZN(n3172) );
  AND2_X1 U2846 ( .A1(n2278), .A2(n3170), .ZN(n2485) );
  OAI21_X1 U2847 ( .B1(n4903), .B2(n2489), .A(n2487), .ZN(n4278) );
  AOI21_X1 U2848 ( .B1(n4386), .B2(REG1_REG_2__SCAN_IN), .A(n3937), .ZN(n2583)
         );
  NAND2_X1 U2849 ( .A1(n2711), .A2(REG2_REG_1__SCAN_IN), .ZN(n2715) );
  AND2_X1 U2850 ( .A1(n2729), .A2(n2728), .ZN(n2496) );
  AND2_X2 U2851 ( .A1(n3820), .A2(n3827), .ZN(n3461) );
  CLKBUF_X1 U2852 ( .A(n4788), .Z(n4790) );
  NAND2_X1 U2853 ( .A1(n4065), .A2(n2766), .ZN(n2733) );
  NOR2_X1 U2854 ( .A1(n3002), .A2(n4951), .ZN(n4020) );
  OR2_X1 U2855 ( .A1(n3958), .A2(n4334), .ZN(n2494) );
  OAI21_X1 U2856 ( .B1(n4381), .B2(REG1_REG_15__SCAN_IN), .A(n2616), .ZN(n4079) );
  NOR2_X1 U2857 ( .A1(n3738), .A2(n4408), .ZN(n3993) );
  OR2_X1 U2858 ( .A1(n4059), .A2(n3523), .ZN(n2495) );
  NAND2_X1 U2859 ( .A1(n2800), .A2(n2801), .ZN(n2497) );
  INV_X1 U2860 ( .A(n2712), .ZN(n2726) );
  OR2_X1 U2861 ( .A1(n3958), .A2(n4374), .ZN(n2498) );
  AND4_X1 U2862 ( .A1(n2511), .A2(n2510), .A3(n2444), .A4(n2552), .ZN(n2512)
         );
  AND2_X1 U2863 ( .A1(n3180), .A2(n3667), .ZN(n3177) );
  AND2_X1 U2864 ( .A1(n3679), .A2(n3177), .ZN(n3178) );
  INV_X1 U2865 ( .A(n3010), .ZN(n3011) );
  AND2_X1 U2866 ( .A1(n2544), .A2(n2540), .ZN(n2517) );
  INV_X1 U2867 ( .A(n3993), .ZN(n3191) );
  INV_X1 U2868 ( .A(n4927), .ZN(n3903) );
  INV_X1 U2869 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2837) );
  AND2_X1 U2870 ( .A1(n4055), .A2(n3183), .ZN(n3848) );
  AND2_X1 U2871 ( .A1(n2886), .A2(REG3_REG_12__SCAN_IN), .ZN(n2902) );
  INV_X1 U2872 ( .A(n2892), .ZN(n2609) );
  AND2_X1 U2873 ( .A1(n3228), .A2(n3741), .ZN(n3761) );
  AND2_X1 U2874 ( .A1(n2902), .A2(REG3_REG_13__SCAN_IN), .ZN(n2914) );
  AND3_X1 U2875 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2774) );
  INV_X1 U2876 ( .A(n4156), .ZN(n4127) );
  INV_X1 U2877 ( .A(n3651), .ZN(n3615) );
  INV_X1 U2878 ( .A(n3354), .ZN(n3360) );
  INV_X1 U2879 ( .A(IR_REG_23__SCAN_IN), .ZN(n2527) );
  OR3_X1 U2880 ( .A1(n2567), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2600) );
  INV_X1 U2881 ( .A(n3451), .ZN(n2804) );
  AND2_X1 U2882 ( .A1(n2973), .A2(REG3_REG_20__SCAN_IN), .ZN(n2986) );
  INV_X1 U2883 ( .A(n4948), .ZN(n4931) );
  INV_X1 U2884 ( .A(n4811), .ZN(n2845) );
  INV_X1 U2885 ( .A(n4079), .ZN(n2617) );
  INV_X1 U2886 ( .A(n3761), .ZN(n4142) );
  INV_X1 U2887 ( .A(n4175), .ZN(n4140) );
  AND2_X1 U2888 ( .A1(n3225), .A2(n4211), .ZN(n4203) );
  NAND2_X1 U2889 ( .A1(n2914), .A2(REG3_REG_14__SCAN_IN), .ZN(n2917) );
  INV_X1 U2890 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2806) );
  NOR2_X1 U2891 ( .A1(n3738), .A2(n4419), .ZN(n3971) );
  AND2_X1 U2892 ( .A1(n3325), .A2(n3237), .ZN(n4274) );
  INV_X1 U2893 ( .A(n4891), .ZN(n4785) );
  INV_X1 U2894 ( .A(n4274), .ZN(n4901) );
  INV_X1 U2895 ( .A(n3124), .ZN(n4705) );
  INV_X1 U2896 ( .A(IR_REG_24__SCAN_IN), .ZN(n2534) );
  INV_X1 U2897 ( .A(IR_REG_15__SCAN_IN), .ZN(n2552) );
  NOR2_X1 U2898 ( .A1(n2600), .A2(IR_REG_9__SCAN_IN), .ZN(n2602) );
  AND2_X1 U2899 ( .A1(n2539), .A2(STATE_REG_SCAN_IN), .ZN(n3254) );
  NOR2_X1 U2900 ( .A1(n2958), .A2(n4035), .ZN(n2972) );
  NOR2_X1 U2901 ( .A1(n3738), .A2(n2981), .ZN(n4942) );
  AND4_X1 U2902 ( .A1(n3136), .A2(n3135), .A3(n3134), .A4(n3133), .ZN(n4125)
         );
  AND4_X1 U2903 ( .A1(n3006), .A2(n3005), .A3(n3004), .A4(n3003), .ZN(n4214)
         );
  INV_X1 U2904 ( .A(n3933), .ZN(n4697) );
  AND2_X1 U2905 ( .A1(n3132), .A2(n3086), .ZN(n4119) );
  INV_X1 U2906 ( .A(n4203), .ZN(n4230) );
  INV_X1 U2907 ( .A(n4268), .ZN(n4897) );
  NAND2_X1 U2908 ( .A1(n3756), .A2(n3232), .ZN(n4891) );
  NOR2_X1 U2909 ( .A1(n2807), .A2(n2806), .ZN(n2822) );
  AND2_X1 U2910 ( .A1(n4825), .A2(n3441), .ZN(n4968) );
  INV_X1 U2911 ( .A(n4827), .ZN(n4917) );
  NAND2_X1 U2912 ( .A1(n4889), .A2(n3706), .ZN(n4264) );
  INV_X1 U2913 ( .A(n4874), .ZN(n4908) );
  AND2_X1 U2914 ( .A1(n4710), .A2(n3231), .ZN(n4844) );
  INV_X1 U2915 ( .A(n3818), .ZN(n3800) );
  AND2_X1 U2916 ( .A1(n2607), .A2(n2565), .ZN(n4646) );
  AND2_X1 U2917 ( .A1(n3151), .A2(n3150), .ZN(n3152) );
  NAND4_X1 U2918 ( .A1(n3075), .A2(n3074), .A3(n3073), .A4(n3072), .ZN(n4156)
         );
  NAND4_X1 U2919 ( .A1(n3035), .A2(n3034), .A3(n3033), .A4(n3032), .ZN(n4216)
         );
  INV_X1 U2920 ( .A(n4698), .ZN(n4680) );
  NAND2_X1 U2921 ( .A1(n4825), .A2(n4791), .ZN(n4280) );
  NAND2_X1 U2922 ( .A1(n3146), .A2(n4844), .ZN(n4827) );
  NAND2_X1 U2923 ( .A1(n4911), .A2(n4908), .ZN(n4334) );
  NAND2_X1 U2924 ( .A1(n4915), .A2(n4908), .ZN(n4374) );
  INV_X1 U2925 ( .A(n4915), .ZN(n4912) );
  INV_X1 U2926 ( .A(n4787), .ZN(n4379) );
  AND2_X1 U2927 ( .A1(n2595), .A2(n2594), .ZN(n4383) );
  INV_X2 U2928 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U2929 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2503)
         );
  INV_X1 U2930 ( .A(IR_REG_7__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U2931 ( .A1(n2505), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U2932 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U2933 ( .A1(n2288), .A2(IR_REG_19__SCAN_IN), .ZN(n2509) );
  NOR2_X1 U2934 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2511)
         );
  NOR2_X1 U2935 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2510)
         );
  NOR2_X1 U2936 ( .A1(n2626), .A2(n2544), .ZN(n2516) );
  NAND2_X1 U2937 ( .A1(n2516), .A2(IR_REG_27__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U2938 ( .A1(n2287), .A2(IR_REG_31__SCAN_IN), .ZN(n2521) );
  XNOR2_X1 U2939 ( .A(n2521), .B(n2520), .ZN(n3231) );
  INV_X1 U2940 ( .A(n3231), .ZN(n3889) );
  INV_X1 U2941 ( .A(n2522), .ZN(n2523) );
  NAND2_X1 U2942 ( .A1(n2523), .A2(IR_REG_31__SCAN_IN), .ZN(n2525) );
  XNOR2_X1 U2943 ( .A(n2525), .B(n2524), .ZN(n3818) );
  NAND2_X1 U2944 ( .A1(n2526), .A2(IR_REG_31__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U2945 ( .A1(n2528), .A2(n2527), .ZN(n2533) );
  OR2_X1 U2946 ( .A1(n2528), .A2(n2527), .ZN(n2529) );
  NAND2_X1 U2947 ( .A1(n2533), .A2(n2529), .ZN(n2539) );
  AND2_X1 U2948 ( .A1(n3237), .A2(n2539), .ZN(n2530) );
  NOR2_X1 U2949 ( .A1(n3738), .A2(n2530), .ZN(n2629) );
  NAND2_X1 U2950 ( .A1(n2667), .A2(n2531), .ZN(n2537) );
  NAND2_X1 U2951 ( .A1(n2537), .A2(IR_REG_31__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U2952 ( .A1(n2543), .A2(IR_REG_31__SCAN_IN), .ZN(n2536) );
  MUX2_X1 U2953 ( .A(IR_REG_31__SCAN_IN), .B(n2536), .S(IR_REG_25__SCAN_IN), 
        .Z(n2538) );
  NAND2_X1 U2954 ( .A1(n2538), .A2(n2537), .ZN(n3110) );
  INV_X1 U2955 ( .A(n3110), .ZN(n4378) );
  NAND2_X1 U2956 ( .A1(n2704), .A2(n3254), .ZN(n3145) );
  OR2_X1 U2957 ( .A1(n2539), .A2(U3149), .ZN(n4388) );
  NAND2_X1 U2958 ( .A1(n3145), .A2(n4388), .ZN(n2627) );
  NAND2_X1 U2959 ( .A1(n2305), .A2(IR_REG_31__SCAN_IN), .ZN(n2542) );
  MUX2_X1 U2960 ( .A(IR_REG_31__SCAN_IN), .B(n2542), .S(IR_REG_28__SCAN_IN), 
        .Z(n2546) );
  NAND2_X1 U2961 ( .A1(n2667), .A2(n2664), .ZN(n2669) );
  NAND2_X1 U2962 ( .A1(n2546), .A2(n2669), .ZN(n3325) );
  NAND2_X1 U2963 ( .A1(n2550), .A2(n2547), .ZN(n2549) );
  INV_X1 U2964 ( .A(IR_REG_18__SCAN_IN), .ZN(n2548) );
  XNOR2_X1 U2965 ( .A(n2549), .B(n2548), .ZN(n3259) );
  XNOR2_X1 U2966 ( .A(n3259), .B(REG1_REG_18__SCAN_IN), .ZN(n4107) );
  XNOR2_X1 U2967 ( .A(n2550), .B(IR_REG_17__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U2968 ( .A1(n2554), .A2(IR_REG_31__SCAN_IN), .ZN(n2551) );
  XNOR2_X1 U2969 ( .A(n2551), .B(IR_REG_16__SCAN_IN), .ZN(n2940) );
  INV_X1 U2970 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4878) );
  OR2_X1 U2971 ( .A1(n2553), .A2(n2552), .ZN(n2555) );
  AND2_X1 U2972 ( .A1(n2555), .A2(n2554), .ZN(n4381) );
  INV_X1 U2973 ( .A(n4381), .ZN(n4086) );
  AND2_X1 U2974 ( .A1(n2557), .A2(n2571), .ZN(n2612) );
  NAND2_X1 U2975 ( .A1(n2612), .A2(n2558), .ZN(n2559) );
  NAND2_X1 U2976 ( .A1(n2559), .A2(IR_REG_31__SCAN_IN), .ZN(n2560) );
  XNOR2_X1 U2977 ( .A(n2560), .B(IR_REG_14__SCAN_IN), .ZN(n4848) );
  INV_X1 U2978 ( .A(n4848), .ZN(n4690) );
  NAND2_X1 U2979 ( .A1(n2571), .A2(n4572), .ZN(n2567) );
  INV_X1 U2980 ( .A(IR_REG_10__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U2981 ( .A1(n2602), .A2(n2561), .ZN(n2562) );
  NAND2_X1 U2982 ( .A1(n2562), .A2(IR_REG_31__SCAN_IN), .ZN(n2564) );
  INV_X1 U2983 ( .A(IR_REG_11__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U2984 ( .A1(n2564), .A2(n2563), .ZN(n2607) );
  OR2_X1 U2985 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  OR2_X1 U2986 ( .A1(n2602), .A2(n2443), .ZN(n2566) );
  XNOR2_X1 U2987 ( .A(n2566), .B(IR_REG_10__SCAN_IN), .ZN(n2861) );
  INV_X1 U2988 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3542) );
  NAND2_X1 U2989 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U2990 ( .A1(n2593), .A2(n2592), .ZN(n2595) );
  NAND2_X1 U2991 ( .A1(n2595), .A2(IR_REG_31__SCAN_IN), .ZN(n2568) );
  XNOR2_X1 U2992 ( .A(n2568), .B(IR_REG_8__SCAN_IN), .ZN(n4382) );
  INV_X1 U2993 ( .A(n4382), .ZN(n2598) );
  OR2_X1 U2994 ( .A1(n2571), .A2(n2443), .ZN(n2569) );
  XNOR2_X1 U2995 ( .A(n2569), .B(IR_REG_6__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U2996 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2570) );
  MUX2_X1 U2997 ( .A(IR_REG_31__SCAN_IN), .B(n2570), .S(IR_REG_5__SCAN_IN), 
        .Z(n2573) );
  INV_X1 U2998 ( .A(n2571), .ZN(n2572) );
  NAND2_X1 U2999 ( .A1(n2783), .A2(REG1_REG_5__SCAN_IN), .ZN(n2589) );
  INV_X1 U3000 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2574) );
  INV_X1 U3001 ( .A(n2783), .ZN(n4764) );
  AOI22_X1 U3002 ( .A1(n2783), .A2(REG1_REG_5__SCAN_IN), .B1(n2574), .B2(n4764), .ZN(n4612) );
  INV_X1 U3003 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2577) );
  MUX2_X1 U3004 ( .A(REG1_REG_1__SCAN_IN), .B(n2577), .S(n4387), .Z(n4070) );
  INV_X1 U3005 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4707) );
  NOR2_X1 U3006 ( .A1(n4704), .A2(n4707), .ZN(n4071) );
  NAND2_X1 U3007 ( .A1(n4387), .A2(REG1_REG_1__SCAN_IN), .ZN(n3938) );
  INV_X1 U3008 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2578) );
  MUX2_X1 U3009 ( .A(n2578), .B(REG1_REG_2__SCAN_IN), .S(n4386), .Z(n3939) );
  NAND2_X1 U3010 ( .A1(n2579), .A2(IR_REG_31__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U3011 ( .A1(n2581), .A2(n2580), .ZN(n2585) );
  OR2_X1 U3012 ( .A1(n2581), .A2(n2580), .ZN(n2582) );
  XNOR2_X1 U3013 ( .A(n2583), .B(n4385), .ZN(n3278) );
  INV_X1 U3014 ( .A(n2583), .ZN(n2584) );
  AOI22_X1 U3015 ( .A1(n3278), .A2(REG1_REG_3__SCAN_IN), .B1(n4385), .B2(n2584), .ZN(n2588) );
  NAND2_X1 U3016 ( .A1(n2585), .A2(IR_REG_31__SCAN_IN), .ZN(n2586) );
  XNOR2_X1 U3017 ( .A(n2586), .B(IR_REG_4__SCAN_IN), .ZN(n4384) );
  INV_X1 U3018 ( .A(n4384), .ZN(n3316) );
  XNOR2_X1 U3019 ( .A(n2588), .B(n4384), .ZN(n3308) );
  NAND2_X1 U3020 ( .A1(n3308), .A2(REG1_REG_4__SCAN_IN), .ZN(n2587) );
  OAI21_X1 U3021 ( .B1(n2588), .B2(n3316), .A(n2587), .ZN(n4611) );
  NAND2_X1 U3022 ( .A1(n4612), .A2(n4611), .ZN(n4610) );
  NAND2_X1 U3023 ( .A1(n4765), .A2(n2590), .ZN(n2591) );
  INV_X1 U3024 ( .A(n4765), .ZN(n4624) );
  AND2_X1 U3025 ( .A1(n3291), .A2(REG1_REG_7__SCAN_IN), .ZN(n2596) );
  OR2_X1 U3026 ( .A1(n2593), .A2(n2592), .ZN(n2594) );
  OAI22_X1 U3027 ( .A1(n2596), .A2(n4383), .B1(REG1_REG_7__SCAN_IN), .B2(n3291), .ZN(n2597) );
  NAND2_X1 U3028 ( .A1(n2600), .A2(IR_REG_31__SCAN_IN), .ZN(n2601) );
  MUX2_X1 U3029 ( .A(IR_REG_31__SCAN_IN), .B(n2601), .S(IR_REG_9__SCAN_IN), 
        .Z(n2604) );
  INV_X1 U3030 ( .A(n2602), .ZN(n2603) );
  NAND2_X1 U3031 ( .A1(n2604), .A2(n2603), .ZN(n4811) );
  NOR2_X1 U3032 ( .A1(n2845), .A2(REG1_REG_9__SCAN_IN), .ZN(n4625) );
  NAND2_X1 U3033 ( .A1(n2845), .A2(REG1_REG_9__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U3034 ( .A1(n2861), .A2(n2605), .ZN(n2606) );
  INV_X1 U3035 ( .A(n2861), .ZN(n4813) );
  NAND2_X1 U3036 ( .A1(n2607), .A2(IR_REG_31__SCAN_IN), .ZN(n2608) );
  XNOR2_X1 U3037 ( .A(n2608), .B(IR_REG_12__SCAN_IN), .ZN(n2892) );
  NOR2_X1 U3038 ( .A1(n2610), .A2(n2609), .ZN(n2611) );
  INV_X1 U3039 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4659) );
  OR2_X1 U3040 ( .A1(n2612), .A2(n2443), .ZN(n2613) );
  XNOR2_X1 U3041 ( .A(n2613), .B(IR_REG_13__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U3042 ( .A1(n4668), .A2(REG1_REG_13__SCAN_IN), .ZN(n4667) );
  INV_X1 U3043 ( .A(n4668), .ZN(n4839) );
  INV_X1 U3044 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4845) );
  NAND2_X1 U3045 ( .A1(n4848), .A2(n2614), .ZN(n2615) );
  NAND2_X1 U3046 ( .A1(n4381), .A2(REG1_REG_15__SCAN_IN), .ZN(n2616) );
  NOR2_X1 U3047 ( .A1(n2940), .A2(n2618), .ZN(n2619) );
  NOR2_X1 U3048 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4699), .ZN(n4700) );
  INV_X1 U3049 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2620) );
  INV_X1 U3050 ( .A(n4380), .ZN(n4100) );
  OAI21_X1 U3051 ( .B1(n2620), .B2(n4100), .A(n2310), .ZN(n4092) );
  INV_X1 U3052 ( .A(n3259), .ZN(n4111) );
  INV_X1 U3053 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2621) );
  OAI22_X1 U3054 ( .A1(n4107), .A2(n2622), .B1(n4111), .B2(n2621), .ZN(n2625)
         );
  INV_X1 U3055 ( .A(REG1_REG_19__SCAN_IN), .ZN(n2623) );
  MUX2_X1 U3056 ( .A(REG1_REG_19__SCAN_IN), .B(n2623), .S(n4787), .Z(n2624) );
  XNOR2_X1 U3057 ( .A(n2626), .B(IR_REG_27__SCAN_IN), .ZN(n4599) );
  INV_X1 U3058 ( .A(n4599), .ZN(n3886) );
  INV_X1 U3059 ( .A(n2627), .ZN(n2628) );
  OR2_X1 U3060 ( .A1(n2629), .A2(n2628), .ZN(n3933) );
  AND2_X1 U3061 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4933) );
  AOI21_X1 U3062 ( .B1(n4697), .B2(ADDR_REG_19__SCAN_IN), .A(n4933), .ZN(n2630) );
  INV_X1 U3063 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4672) );
  NOR2_X1 U3064 ( .A1(n4839), .A2(n4672), .ZN(n4671) );
  NAND2_X1 U3065 ( .A1(n4646), .A2(REG2_REG_11__SCAN_IN), .ZN(n2649) );
  INV_X1 U3066 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4826) );
  INV_X1 U3067 ( .A(n4646), .ZN(n4822) );
  AOI22_X1 U3068 ( .A1(n4646), .A2(REG2_REG_11__SCAN_IN), .B1(n4826), .B2(
        n4822), .ZN(n4654) );
  NAND2_X1 U3069 ( .A1(n2845), .A2(REG2_REG_9__SCAN_IN), .ZN(n2646) );
  INV_X1 U3070 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U3071 ( .A1(n2845), .A2(REG2_REG_9__SCAN_IN), .B1(n3515), .B2(n4811), .ZN(n4635) );
  INV_X1 U3072 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2631) );
  MUX2_X1 U3073 ( .A(REG2_REG_2__SCAN_IN), .B(n2631), .S(n4386), .Z(n3936) );
  INV_X1 U3074 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2632) );
  INV_X1 U3075 ( .A(n3326), .ZN(n4073) );
  NAND2_X1 U3076 ( .A1(n4074), .A2(n4073), .ZN(n4072) );
  NAND2_X1 U3077 ( .A1(n4387), .A2(REG2_REG_1__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3078 ( .A1(n4386), .A2(REG2_REG_2__SCAN_IN), .ZN(n2634) );
  INV_X1 U3079 ( .A(n4385), .ZN(n3279) );
  NAND2_X1 U3080 ( .A1(n3282), .A2(REG2_REG_3__SCAN_IN), .ZN(n3281) );
  NAND2_X1 U3081 ( .A1(n2635), .A2(n4385), .ZN(n2636) );
  NAND2_X1 U3082 ( .A1(n3281), .A2(n2636), .ZN(n2637) );
  NAND2_X1 U3083 ( .A1(n2783), .A2(REG2_REG_5__SCAN_IN), .ZN(n2638) );
  OAI21_X1 U3084 ( .B1(n2783), .B2(REG2_REG_5__SCAN_IN), .A(n2638), .ZN(n4606)
         );
  INV_X1 U3085 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4617) );
  INV_X1 U3086 ( .A(n3288), .ZN(n2642) );
  INV_X1 U3087 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U3088 ( .A1(n3288), .A2(n2640), .ZN(n2641) );
  INV_X1 U3089 ( .A(n2644), .ZN(n2643) );
  NAND2_X1 U3090 ( .A1(n2643), .A2(n4382), .ZN(n2645) );
  XNOR2_X1 U3091 ( .A(n2644), .B(n4382), .ZN(n3386) );
  NAND2_X1 U3092 ( .A1(n2861), .A2(n2647), .ZN(n2648) );
  NAND2_X1 U3093 ( .A1(n2892), .A2(n2650), .ZN(n2651) );
  XNOR2_X1 U3094 ( .A(n2650), .B(n2609), .ZN(n4664) );
  NAND2_X1 U3095 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4664), .ZN(n4662) );
  NAND2_X1 U3096 ( .A1(n2651), .A2(n4662), .ZN(n4673) );
  OAI22_X1 U3097 ( .A1(n4671), .A2(n4673), .B1(n4668), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n2652) );
  NOR2_X1 U3098 ( .A1(n4690), .A2(n2652), .ZN(n2653) );
  INV_X1 U3099 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4683) );
  XOR2_X1 U3100 ( .A(n4848), .B(n2652), .Z(n4682) );
  NAND2_X1 U3101 ( .A1(n4381), .A2(REG2_REG_15__SCAN_IN), .ZN(n2654) );
  OAI21_X1 U3102 ( .B1(n4381), .B2(REG2_REG_15__SCAN_IN), .A(n2654), .ZN(n4084) );
  NAND2_X1 U3103 ( .A1(n2655), .A2(n2315), .ZN(n2656) );
  INV_X1 U3104 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4693) );
  XOR2_X1 U3105 ( .A(REG2_REG_17__SCAN_IN), .B(n4380), .Z(n4096) );
  INV_X1 U3106 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2658) );
  NOR2_X1 U3107 ( .A1(n3259), .A2(n2658), .ZN(n2657) );
  AOI21_X1 U3108 ( .B1(n2658), .B2(n3259), .A(n2657), .ZN(n4104) );
  INV_X1 U3109 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2659) );
  MUX2_X1 U3110 ( .A(n2659), .B(REG2_REG_19__SCAN_IN), .S(n4787), .Z(n2660) );
  XNOR2_X1 U3111 ( .A(n2661), .B(n2660), .ZN(n2663) );
  NOR2_X1 U3112 ( .A1(n3325), .A2(n3886), .ZN(n2662) );
  NAND2_X1 U3113 ( .A1(n2669), .A2(IR_REG_31__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U3114 ( .A1(n3081), .A2(REG0_REG_19__SCAN_IN), .ZN(n2680) );
  INV_X1 U3115 ( .A(n2676), .ZN(n3263) );
  CLKBUF_X3 U3116 ( .A(n2727), .Z(n3071) );
  NAND2_X1 U3117 ( .A1(n2774), .A2(REG3_REG_6__SCAN_IN), .ZN(n2807) );
  NAND2_X1 U3118 ( .A1(n2822), .A2(REG3_REG_8__SCAN_IN), .ZN(n2838) );
  INV_X1 U3119 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2690) );
  INV_X1 U3120 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4035) );
  XNOR2_X1 U3121 ( .A(REG3_REG_19__SCAN_IN), .B(n2972), .ZN(n4938) );
  INV_X1 U3122 ( .A(n4938), .ZN(n2673) );
  NAND2_X1 U3123 ( .A1(n3071), .A2(n2673), .ZN(n2679) );
  NAND2_X1 U3124 ( .A1(n2262), .A2(REG2_REG_19__SCAN_IN), .ZN(n2678) );
  INV_X1 U3125 ( .A(n2674), .ZN(n2675) );
  NAND2_X1 U3126 ( .A1(n2810), .A2(REG1_REG_19__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U3127 ( .A1(n4944), .A2(n2261), .ZN(n2685) );
  MUX2_X1 U3128 ( .A(DATAI_19_), .B(n4379), .S(n3738), .Z(n4926) );
  AND2_X1 U3129 ( .A1(n3142), .A2(n2704), .ZN(n2688) );
  INV_X2 U3130 ( .A(n3007), .ZN(n3077) );
  NAND2_X1 U3131 ( .A1(n4926), .A2(n3077), .ZN(n2684) );
  NAND2_X1 U3132 ( .A1(n2685), .A2(n2684), .ZN(n2686) );
  NAND2_X1 U3133 ( .A1(n4787), .A2(n3889), .ZN(n3140) );
  XNOR2_X1 U3134 ( .A(n2686), .B(n2734), .ZN(n2971) );
  NAND2_X1 U3135 ( .A1(n3231), .A2(n3818), .ZN(n3124) );
  NAND2_X1 U3136 ( .A1(n2687), .A2(n4705), .ZN(n4874) );
  AOI22_X1 U3137 ( .A1(n4944), .A2(n2737), .B1(n2261), .B2(n4926), .ZN(n2969)
         );
  INV_X1 U3138 ( .A(n2969), .ZN(n2970) );
  NAND2_X1 U3139 ( .A1(n3081), .A2(REG0_REG_15__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3140 ( .A1(n2917), .A2(n2690), .ZN(n2691) );
  NAND2_X1 U3141 ( .A1(n2935), .A2(n2691), .ZN(n4871) );
  INV_X1 U3142 ( .A(n4871), .ZN(n2692) );
  NAND2_X1 U3143 ( .A1(n3071), .A2(n2692), .ZN(n2695) );
  NAND2_X1 U3144 ( .A1(n2262), .A2(REG2_REG_15__SCAN_IN), .ZN(n2694) );
  NAND2_X1 U3145 ( .A1(n2810), .A2(REG1_REG_15__SCAN_IN), .ZN(n2693) );
  NAND4_X1 U3146 ( .A1(n2696), .A2(n2695), .A3(n2694), .A4(n2693), .ZN(n4898)
         );
  MUX2_X1 U3147 ( .A(DATAI_15_), .B(n4381), .S(n3738), .Z(n3248) );
  INV_X1 U31480 ( .A(n3248), .ZN(n4857) );
  NOR2_X1 U31490 ( .A1(n4857), .A2(n2717), .ZN(n2697) );
  AOI21_X1 U3150 ( .B1(n4898), .B2(n2737), .A(n2697), .ZN(n4866) );
  NAND2_X1 U3151 ( .A1(n2756), .A2(REG0_REG_0__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U3152 ( .A1(n2727), .A2(REG3_REG_0__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U3153 ( .A1(n2711), .A2(REG2_REG_0__SCAN_IN), .ZN(n2699) );
  NAND2_X1 U3154 ( .A1(n2712), .A2(REG1_REG_0__SCAN_IN), .ZN(n2698) );
  NAND2_X1 U3155 ( .A1(n4721), .A2(n2737), .ZN(n2703) );
  NAND2_X1 U3156 ( .A1(n4732), .A2(n2766), .ZN(n2702) );
  NAND2_X1 U3157 ( .A1(n2703), .A2(n2702), .ZN(n3320) );
  NAND2_X1 U3158 ( .A1(n4721), .A2(n2766), .ZN(n2706) );
  NAND2_X1 U3159 ( .A1(n3142), .A2(n2704), .ZN(n3007) );
  NAND2_X1 U3160 ( .A1(n4732), .A2(n3077), .ZN(n2705) );
  NAND2_X1 U3161 ( .A1(n2706), .A2(n2705), .ZN(n3321) );
  NAND2_X1 U3162 ( .A1(n3320), .A2(n3321), .ZN(n2709) );
  INV_X1 U3163 ( .A(n2704), .ZN(n2707) );
  NAND2_X1 U3164 ( .A1(n2707), .A2(n4071), .ZN(n2708) );
  NAND2_X1 U3165 ( .A1(n2709), .A2(n2708), .ZN(n3322) );
  INV_X1 U3166 ( .A(n3322), .ZN(n2710) );
  NAND2_X1 U3167 ( .A1(n2710), .A2(n2280), .ZN(n3332) );
  NAND2_X1 U3168 ( .A1(n2727), .A2(REG3_REG_1__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U3169 ( .A1(n2756), .A2(REG0_REG_1__SCAN_IN), .ZN(n2714) );
  NAND2_X1 U3170 ( .A1(n2712), .A2(REG1_REG_1__SCAN_IN), .ZN(n2713) );
  INV_X2 U3171 ( .A(n3156), .ZN(n4066) );
  NOR2_X1 U3172 ( .A1(n3155), .A2(n2717), .ZN(n2718) );
  NAND2_X1 U3173 ( .A1(n4731), .A2(n2688), .ZN(n2719) );
  NAND2_X1 U3174 ( .A1(n2720), .A2(n2719), .ZN(n2721) );
  INV_X1 U3175 ( .A(n2723), .ZN(n2724) );
  NAND2_X1 U3176 ( .A1(n2722), .A2(n2724), .ZN(n2725) );
  NAND2_X1 U3177 ( .A1(n3331), .A2(n2725), .ZN(n3299) );
  NAND2_X1 U3178 ( .A1(n2712), .A2(REG1_REG_2__SCAN_IN), .ZN(n2731) );
  NAND2_X1 U3179 ( .A1(n2711), .A2(REG2_REG_2__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U3180 ( .A1(n2727), .A2(REG3_REG_2__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U3181 ( .A1(n2756), .A2(REG0_REG_2__SCAN_IN), .ZN(n2728) );
  MUX2_X1 U3182 ( .A(DATAI_2_), .B(n4386), .S(n2746), .Z(n3477) );
  NAND2_X1 U3183 ( .A1(n3477), .A2(n3077), .ZN(n2732) );
  NAND2_X1 U3184 ( .A1(n2733), .A2(n2732), .ZN(n2735) );
  XNOR2_X1 U3185 ( .A(n2740), .B(n2739), .ZN(n3300) );
  INV_X1 U3186 ( .A(n3300), .ZN(n2738) );
  NAND2_X1 U3187 ( .A1(n2740), .A2(n2739), .ZN(n2741) );
  INV_X1 U3188 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U3189 ( .A1(n3071), .A2(n2757), .ZN(n2745) );
  NAND2_X1 U3190 ( .A1(n2262), .A2(REG2_REG_3__SCAN_IN), .ZN(n2744) );
  NAND2_X1 U3191 ( .A1(n2810), .A2(REG1_REG_3__SCAN_IN), .ZN(n2743) );
  NAND2_X1 U3192 ( .A1(n3081), .A2(REG0_REG_3__SCAN_IN), .ZN(n2742) );
  MUX2_X1 U3193 ( .A(DATAI_3_), .B(n4385), .S(n2746), .Z(n3354) );
  NOR2_X1 U3194 ( .A1(n3360), .A2(n2717), .ZN(n2747) );
  NAND2_X1 U3195 ( .A1(n4064), .A2(n3091), .ZN(n2749) );
  NAND2_X1 U3196 ( .A1(n3354), .A2(n3077), .ZN(n2748) );
  NAND2_X1 U3197 ( .A1(n2749), .A2(n2748), .ZN(n2750) );
  XNOR2_X1 U3198 ( .A(n2752), .B(n2751), .ZN(n3343) );
  INV_X1 U3199 ( .A(n2751), .ZN(n2753) );
  NAND2_X1 U3200 ( .A1(n2753), .A2(n2752), .ZN(n2754) );
  NAND2_X1 U3201 ( .A1(n2755), .A2(n2754), .ZN(n3391) );
  INV_X1 U3202 ( .A(n3391), .ZN(n2770) );
  NAND2_X1 U3203 ( .A1(n3081), .A2(REG0_REG_4__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U3204 ( .A1(n2262), .A2(REG2_REG_4__SCAN_IN), .ZN(n2760) );
  XNOR2_X1 U3205 ( .A(n2757), .B(REG3_REG_4__SCAN_IN), .ZN(n3427) );
  NAND2_X1 U3206 ( .A1(n3071), .A2(n3427), .ZN(n2759) );
  NAND2_X1 U3207 ( .A1(n2810), .A2(REG1_REG_4__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U3208 ( .A1(n4063), .A2(n2260), .ZN(n2764) );
  NAND2_X1 U3209 ( .A1(n3409), .A2(n3077), .ZN(n2763) );
  NAND2_X1 U32100 ( .A1(n2764), .A2(n2763), .ZN(n2765) );
  XNOR2_X1 U32110 ( .A(n2765), .B(n3066), .ZN(n2771) );
  INV_X2 U32120 ( .A(n2766), .ZN(n2767) );
  XNOR2_X1 U32130 ( .A(n2771), .B(n2772), .ZN(n3392) );
  INV_X1 U32140 ( .A(n3392), .ZN(n2769) );
  NAND2_X1 U32150 ( .A1(n3081), .A2(REG0_REG_5__SCAN_IN), .ZN(n2782) );
  INV_X1 U32160 ( .A(n2774), .ZN(n2789) );
  INV_X1 U32170 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U32180 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2775) );
  NAND2_X1 U32190 ( .A1(n2776), .A2(n2775), .ZN(n2777) );
  NAND2_X1 U32200 ( .A1(n2789), .A2(n2777), .ZN(n3442) );
  INV_X1 U32210 ( .A(n3442), .ZN(n2778) );
  NAND2_X1 U32220 ( .A1(n3071), .A2(n2778), .ZN(n2781) );
  NAND2_X1 U32230 ( .A1(n2262), .A2(REG2_REG_5__SCAN_IN), .ZN(n2780) );
  NAND2_X1 U32240 ( .A1(n2810), .A2(REG1_REG_5__SCAN_IN), .ZN(n2779) );
  NAND4_X1 U32250 ( .A1(n2782), .A2(n2781), .A3(n2780), .A4(n2779), .ZN(n4062)
         );
  NAND2_X1 U32260 ( .A1(n4062), .A2(n2737), .ZN(n2785) );
  MUX2_X1 U32270 ( .A(DATAI_5_), .B(n2783), .S(n3738), .Z(n3403) );
  INV_X2 U32280 ( .A(n2767), .ZN(n3091) );
  NAND2_X1 U32290 ( .A1(n3403), .A2(n3091), .ZN(n2784) );
  NAND2_X1 U32300 ( .A1(n2785), .A2(n2784), .ZN(n3400) );
  NAND2_X1 U32310 ( .A1(n4062), .A2(n2261), .ZN(n2787) );
  NAND2_X1 U32320 ( .A1(n3403), .A2(n3077), .ZN(n2786) );
  NAND2_X1 U32330 ( .A1(n2787), .A2(n2786), .ZN(n2788) );
  XNOR2_X1 U32340 ( .A(n2788), .B(n2734), .ZN(n3401) );
  INV_X1 U32350 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3453) );
  NAND2_X1 U32360 ( .A1(n2789), .A2(n3453), .ZN(n2790) );
  AND2_X1 U32370 ( .A1(n2790), .A2(n2807), .ZN(n4767) );
  NAND2_X1 U32380 ( .A1(n3071), .A2(n4767), .ZN(n2794) );
  NAND2_X1 U32390 ( .A1(n2262), .A2(REG2_REG_6__SCAN_IN), .ZN(n2793) );
  NAND2_X1 U32400 ( .A1(n2810), .A2(REG1_REG_6__SCAN_IN), .ZN(n2792) );
  NAND2_X1 U32410 ( .A1(n3081), .A2(REG0_REG_6__SCAN_IN), .ZN(n2791) );
  NAND4_X1 U32420 ( .A1(n2794), .A2(n2793), .A3(n2792), .A4(n2791), .ZN(n4783)
         );
  NAND2_X1 U32430 ( .A1(n4783), .A2(n3091), .ZN(n2796) );
  MUX2_X1 U32440 ( .A(DATAI_6_), .B(n4765), .S(n3738), .Z(n3454) );
  NAND2_X1 U32450 ( .A1(n3454), .A2(n3077), .ZN(n2795) );
  NAND2_X1 U32460 ( .A1(n2796), .A2(n2795), .ZN(n2797) );
  XNOR2_X1 U32470 ( .A(n2797), .B(n2734), .ZN(n2800) );
  NAND2_X1 U32480 ( .A1(n4783), .A2(n2737), .ZN(n2799) );
  NAND2_X1 U32490 ( .A1(n3454), .A2(n3091), .ZN(n2798) );
  NAND2_X1 U32500 ( .A1(n2799), .A2(n2798), .ZN(n2801) );
  INV_X1 U32510 ( .A(n2800), .ZN(n2803) );
  INV_X1 U32520 ( .A(n2801), .ZN(n2802) );
  NAND2_X1 U32530 ( .A1(n2803), .A2(n2802), .ZN(n3451) );
  AND2_X1 U32540 ( .A1(n2807), .A2(n2806), .ZN(n2808) );
  OR2_X1 U32550 ( .A1(n2808), .A2(n2822), .ZN(n4796) );
  INV_X1 U32560 ( .A(n4796), .ZN(n2809) );
  NAND2_X1 U32570 ( .A1(n3071), .A2(n2809), .ZN(n2814) );
  NAND2_X1 U32580 ( .A1(n2262), .A2(REG2_REG_7__SCAN_IN), .ZN(n2813) );
  NAND2_X1 U32590 ( .A1(n2810), .A2(REG1_REG_7__SCAN_IN), .ZN(n2812) );
  NAND2_X1 U32600 ( .A1(n3081), .A2(REG0_REG_7__SCAN_IN), .ZN(n2811) );
  NAND4_X1 U32610 ( .A1(n2814), .A2(n2813), .A3(n2812), .A4(n2811), .ZN(n4061)
         );
  NAND2_X1 U32620 ( .A1(n4061), .A2(n3091), .ZN(n2816) );
  MUX2_X1 U32630 ( .A(DATAI_7_), .B(n4383), .S(n3738), .Z(n4774) );
  NAND2_X1 U32640 ( .A1(n4774), .A2(n3077), .ZN(n2815) );
  NAND2_X1 U32650 ( .A1(n2816), .A2(n2815), .ZN(n2817) );
  XNOR2_X1 U32660 ( .A(n2817), .B(n2734), .ZN(n2821) );
  INV_X1 U32670 ( .A(n4774), .ZN(n4779) );
  NOR2_X1 U32680 ( .A1(n4779), .A2(n2767), .ZN(n2818) );
  AOI21_X1 U32690 ( .B1(n4061), .B2(n2737), .A(n2818), .ZN(n2819) );
  XNOR2_X1 U32700 ( .A(n2821), .B(n2819), .ZN(n3964) );
  INV_X1 U32710 ( .A(n2819), .ZN(n2820) );
  NAND2_X1 U32720 ( .A1(n3081), .A2(REG0_REG_8__SCAN_IN), .ZN(n2827) );
  OR2_X1 U32730 ( .A1(n2822), .A2(REG3_REG_8__SCAN_IN), .ZN(n2823) );
  AND2_X1 U32740 ( .A1(n2838), .A2(n2823), .ZN(n4803) );
  NAND2_X1 U32750 ( .A1(n3071), .A2(n4803), .ZN(n2826) );
  NAND2_X1 U32760 ( .A1(n2262), .A2(REG2_REG_8__SCAN_IN), .ZN(n2825) );
  NAND2_X1 U32770 ( .A1(n2810), .A2(REG1_REG_8__SCAN_IN), .ZN(n2824) );
  NAND4_X1 U32780 ( .A1(n2827), .A2(n2826), .A3(n2825), .A4(n2824), .ZN(n4060)
         );
  NAND2_X1 U32790 ( .A1(n4060), .A2(n3091), .ZN(n2829) );
  MUX2_X1 U32800 ( .A(DATAI_8_), .B(n4382), .S(n3738), .Z(n3501) );
  NAND2_X1 U32810 ( .A1(n3501), .A2(n3077), .ZN(n2828) );
  NAND2_X1 U32820 ( .A1(n2829), .A2(n2828), .ZN(n2830) );
  XNOR2_X1 U32830 ( .A(n2830), .B(n2734), .ZN(n2833) );
  NAND2_X1 U32840 ( .A1(n4060), .A2(n2737), .ZN(n2832) );
  NAND2_X1 U32850 ( .A1(n3501), .A2(n2261), .ZN(n2831) );
  NAND2_X1 U32860 ( .A1(n2832), .A2(n2831), .ZN(n2834) );
  AND2_X1 U32870 ( .A1(n2833), .A2(n2834), .ZN(n3496) );
  INV_X1 U32880 ( .A(n2833), .ZN(n2836) );
  INV_X1 U32890 ( .A(n2834), .ZN(n2835) );
  NAND2_X1 U32900 ( .A1(n2836), .A2(n2835), .ZN(n3497) );
  NAND2_X1 U32910 ( .A1(n2838), .A2(n2837), .ZN(n2839) );
  NAND2_X1 U32920 ( .A1(n2855), .A2(n2839), .ZN(n3526) );
  INV_X1 U32930 ( .A(n3526), .ZN(n2840) );
  NAND2_X1 U32940 ( .A1(n3071), .A2(n2840), .ZN(n2844) );
  NAND2_X1 U32950 ( .A1(n2262), .A2(REG2_REG_9__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U32960 ( .A1(n2810), .A2(REG1_REG_9__SCAN_IN), .ZN(n2842) );
  NAND2_X1 U32970 ( .A1(n3081), .A2(REG0_REG_9__SCAN_IN), .ZN(n2841) );
  NAND4_X1 U32980 ( .A1(n2844), .A2(n2843), .A3(n2842), .A4(n2841), .ZN(n4059)
         );
  NAND2_X1 U32990 ( .A1(n4059), .A2(n3091), .ZN(n2847) );
  MUX2_X1 U33000 ( .A(DATAI_9_), .B(n2845), .S(n3738), .Z(n3523) );
  NAND2_X1 U33010 ( .A1(n3523), .A2(n3077), .ZN(n2846) );
  NAND2_X1 U33020 ( .A1(n2847), .A2(n2846), .ZN(n2848) );
  XNOR2_X1 U33030 ( .A(n2848), .B(n2734), .ZN(n2850) );
  NOR2_X1 U33040 ( .A1(n3514), .A2(n2717), .ZN(n2849) );
  AOI21_X1 U33050 ( .B1(n4059), .B2(n2737), .A(n2849), .ZN(n2851) );
  XNOR2_X1 U33060 ( .A(n2850), .B(n2851), .ZN(n3521) );
  NAND2_X1 U33070 ( .A1(n3522), .A2(n3521), .ZN(n2854) );
  INV_X1 U33080 ( .A(n2850), .ZN(n2852) );
  NAND2_X1 U33090 ( .A1(n2852), .A2(n2851), .ZN(n2853) );
  NAND2_X1 U33100 ( .A1(n3081), .A2(REG0_REG_10__SCAN_IN), .ZN(n2860) );
  NAND2_X1 U33110 ( .A1(n2855), .A2(n4486), .ZN(n2856) );
  AND2_X1 U33120 ( .A1(n2872), .A2(n2856), .ZN(n4814) );
  NAND2_X1 U33130 ( .A1(n3071), .A2(n4814), .ZN(n2859) );
  NAND2_X1 U33140 ( .A1(n2262), .A2(REG2_REG_10__SCAN_IN), .ZN(n2858) );
  NAND2_X1 U33150 ( .A1(n2810), .A2(REG1_REG_10__SCAN_IN), .ZN(n2857) );
  NAND4_X1 U33160 ( .A1(n2860), .A2(n2859), .A3(n2858), .A4(n2857), .ZN(n4058)
         );
  NAND2_X1 U33170 ( .A1(n4058), .A2(n3091), .ZN(n2863) );
  MUX2_X1 U33180 ( .A(DATAI_10_), .B(n2861), .S(n3738), .Z(n3628) );
  NAND2_X1 U33190 ( .A1(n3628), .A2(n3077), .ZN(n2862) );
  NAND2_X1 U33200 ( .A1(n2863), .A2(n2862), .ZN(n2864) );
  XNOR2_X1 U33210 ( .A(n2864), .B(n3066), .ZN(n2866) );
  INV_X1 U33220 ( .A(n3628), .ZN(n3624) );
  NOR2_X1 U33230 ( .A1(n3624), .A2(n2717), .ZN(n2865) );
  AOI21_X1 U33240 ( .B1(n4058), .B2(n2737), .A(n2865), .ZN(n2867) );
  XNOR2_X1 U33250 ( .A(n2866), .B(n2867), .ZN(n3582) );
  INV_X1 U33260 ( .A(n2866), .ZN(n2869) );
  INV_X1 U33270 ( .A(n2867), .ZN(n2868) );
  NAND2_X1 U33280 ( .A1(n2869), .A2(n2868), .ZN(n2870) );
  NAND2_X1 U33290 ( .A1(n3081), .A2(REG0_REG_11__SCAN_IN), .ZN(n2878) );
  AND2_X1 U33300 ( .A1(n2872), .A2(n2871), .ZN(n2873) );
  OR2_X1 U33310 ( .A1(n2873), .A2(n2886), .ZN(n4828) );
  INV_X1 U33320 ( .A(n4828), .ZN(n2874) );
  NAND2_X1 U33330 ( .A1(n3071), .A2(n2874), .ZN(n2877) );
  NAND2_X1 U33340 ( .A1(n2262), .A2(REG2_REG_11__SCAN_IN), .ZN(n2876) );
  NAND2_X1 U33350 ( .A1(n2810), .A2(REG1_REG_11__SCAN_IN), .ZN(n2875) );
  NAND4_X1 U33360 ( .A1(n2878), .A2(n2877), .A3(n2876), .A4(n2875), .ZN(n4057)
         );
  NAND2_X1 U33370 ( .A1(n4057), .A2(n3091), .ZN(n2880) );
  MUX2_X1 U33380 ( .A(DATAI_11_), .B(n4646), .S(n3738), .Z(n3594) );
  NAND2_X1 U33390 ( .A1(n3594), .A2(n3077), .ZN(n2879) );
  NAND2_X1 U33400 ( .A1(n2880), .A2(n2879), .ZN(n2881) );
  XNOR2_X1 U33410 ( .A(n2881), .B(n3066), .ZN(n3571) );
  INV_X1 U33420 ( .A(n3594), .ZN(n3590) );
  NOR2_X1 U33430 ( .A1(n3590), .A2(n2717), .ZN(n2882) );
  AOI21_X1 U33440 ( .B1(n4057), .B2(n2737), .A(n2882), .ZN(n3570) );
  INV_X1 U33450 ( .A(n3571), .ZN(n2884) );
  INV_X1 U33460 ( .A(n3570), .ZN(n2883) );
  NAND2_X1 U33470 ( .A1(n2884), .A2(n2883), .ZN(n2885) );
  NAND2_X1 U33480 ( .A1(n3081), .A2(REG0_REG_12__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U33490 ( .A1(n2262), .A2(REG2_REG_12__SCAN_IN), .ZN(n2890) );
  NOR2_X1 U33500 ( .A1(n2886), .A2(REG3_REG_12__SCAN_IN), .ZN(n2887) );
  OR2_X1 U33510 ( .A1(n2902), .A2(n2887), .ZN(n4593) );
  INV_X1 U33520 ( .A(n4593), .ZN(n3565) );
  NAND2_X1 U3353 ( .A1(n3071), .A2(n3565), .ZN(n2889) );
  NAND2_X1 U33540 ( .A1(n2810), .A2(REG1_REG_12__SCAN_IN), .ZN(n2888) );
  NAND4_X1 U3355 ( .A1(n2891), .A2(n2890), .A3(n2889), .A4(n2888), .ZN(n4056)
         );
  NAND2_X1 U3356 ( .A1(n4056), .A2(n2261), .ZN(n2894) );
  MUX2_X1 U3357 ( .A(DATAI_12_), .B(n2892), .S(n3738), .Z(n3209) );
  NAND2_X1 U3358 ( .A1(n3209), .A2(n3077), .ZN(n2893) );
  NAND2_X1 U3359 ( .A1(n2894), .A2(n2893), .ZN(n2895) );
  XNOR2_X1 U3360 ( .A(n2895), .B(n2734), .ZN(n2898) );
  NAND2_X1 U3361 ( .A1(n4056), .A2(n2737), .ZN(n2897) );
  NAND2_X1 U3362 ( .A1(n3209), .A2(n2766), .ZN(n2896) );
  NAND2_X1 U3363 ( .A1(n2897), .A2(n2896), .ZN(n2899) );
  INV_X1 U3364 ( .A(n2898), .ZN(n2901) );
  INV_X1 U3365 ( .A(n2899), .ZN(n2900) );
  NAND2_X1 U3366 ( .A1(n2901), .A2(n2900), .ZN(n4583) );
  NAND2_X1 U3367 ( .A1(n3081), .A2(REG0_REG_13__SCAN_IN), .ZN(n2907) );
  NOR2_X1 U3368 ( .A1(n2902), .A2(REG3_REG_13__SCAN_IN), .ZN(n2903) );
  OR2_X1 U3369 ( .A1(n2914), .A2(n2903), .ZN(n3654) );
  INV_X1 U3370 ( .A(n3654), .ZN(n3617) );
  NAND2_X1 U3371 ( .A1(n3071), .A2(n3617), .ZN(n2906) );
  NAND2_X1 U3372 ( .A1(n2262), .A2(REG2_REG_13__SCAN_IN), .ZN(n2905) );
  NAND2_X1 U3373 ( .A1(n2810), .A2(REG1_REG_13__SCAN_IN), .ZN(n2904) );
  NAND4_X1 U3374 ( .A1(n2907), .A2(n2906), .A3(n2905), .A4(n2904), .ZN(n4591)
         );
  NAND2_X1 U3375 ( .A1(n4591), .A2(n2261), .ZN(n2909) );
  MUX2_X1 U3376 ( .A(DATAI_13_), .B(n4668), .S(n3738), .Z(n3651) );
  NAND2_X1 U3377 ( .A1(n3651), .A2(n3077), .ZN(n2908) );
  NAND2_X1 U3378 ( .A1(n2909), .A2(n2908), .ZN(n2910) );
  XNOR2_X1 U3379 ( .A(n2910), .B(n3066), .ZN(n3648) );
  NAND2_X1 U3380 ( .A1(n4591), .A2(n2737), .ZN(n2912) );
  NAND2_X1 U3381 ( .A1(n3651), .A2(n2261), .ZN(n2911) );
  NAND2_X1 U3382 ( .A1(n2912), .A2(n2911), .ZN(n3647) );
  INV_X1 U3383 ( .A(n3648), .ZN(n2913) );
  INV_X1 U3384 ( .A(n2914), .ZN(n2915) );
  INV_X1 U3385 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4536) );
  NAND2_X1 U3386 ( .A1(n2915), .A2(n4536), .ZN(n2916) );
  AND2_X1 U3387 ( .A1(n2917), .A2(n2916), .ZN(n4850) );
  NAND2_X1 U3388 ( .A1(n3071), .A2(n4850), .ZN(n2921) );
  NAND2_X1 U3389 ( .A1(n2262), .A2(REG2_REG_14__SCAN_IN), .ZN(n2920) );
  NAND2_X1 U3390 ( .A1(n2810), .A2(REG1_REG_14__SCAN_IN), .ZN(n2919) );
  NAND2_X1 U3391 ( .A1(n3081), .A2(REG0_REG_14__SCAN_IN), .ZN(n2918) );
  NAND4_X1 U3392 ( .A1(n2921), .A2(n2920), .A3(n2919), .A4(n2918), .ZN(n4862)
         );
  NAND2_X1 U3393 ( .A1(n4862), .A2(n3091), .ZN(n2923) );
  MUX2_X1 U3394 ( .A(DATAI_14_), .B(n4848), .S(n3738), .Z(n3695) );
  NAND2_X1 U3395 ( .A1(n3695), .A2(n3077), .ZN(n2922) );
  NAND2_X1 U3396 ( .A1(n2923), .A2(n2922), .ZN(n2924) );
  XNOR2_X1 U3397 ( .A(n2924), .B(n2734), .ZN(n2927) );
  NAND2_X1 U3398 ( .A1(n4862), .A2(n2737), .ZN(n2926) );
  NAND2_X1 U3399 ( .A1(n3695), .A2(n2766), .ZN(n2925) );
  NAND2_X1 U3400 ( .A1(n2926), .A2(n2925), .ZN(n2928) );
  INV_X1 U3401 ( .A(n2927), .ZN(n2930) );
  INV_X1 U3402 ( .A(n2928), .ZN(n2929) );
  NAND2_X1 U3403 ( .A1(n2930), .A2(n2929), .ZN(n3693) );
  NAND2_X1 U3404 ( .A1(n4898), .A2(n2261), .ZN(n2932) );
  NAND2_X1 U3405 ( .A1(n3248), .A2(n3077), .ZN(n2931) );
  NAND2_X1 U3406 ( .A1(n2932), .A2(n2931), .ZN(n2933) );
  XNOR2_X1 U3407 ( .A(n2933), .B(n2734), .ZN(n2934) );
  NAND2_X1 U3408 ( .A1(n2277), .A2(n2934), .ZN(n4863) );
  NAND2_X1 U3409 ( .A1(n3081), .A2(REG0_REG_16__SCAN_IN), .ZN(n2939) );
  AOI21_X1 U3410 ( .B1(n2935), .B2(n4691), .A(n2946), .ZN(n4918) );
  NAND2_X1 U3411 ( .A1(n3071), .A2(n4918), .ZN(n2938) );
  NAND2_X1 U3412 ( .A1(n2262), .A2(REG2_REG_16__SCAN_IN), .ZN(n2937) );
  NAND2_X1 U3413 ( .A1(n2810), .A2(REG1_REG_16__SCAN_IN), .ZN(n2936) );
  NAND4_X1 U3414 ( .A1(n2939), .A2(n2938), .A3(n2937), .A4(n2936), .ZN(n4055)
         );
  MUX2_X1 U3415 ( .A(DATAI_16_), .B(n2940), .S(n3738), .Z(n4895) );
  AOI22_X1 U3416 ( .A1(n4055), .A2(n2737), .B1(n3091), .B2(n4895), .ZN(n2944)
         );
  NAND2_X1 U3417 ( .A1(n4055), .A2(n2261), .ZN(n2942) );
  NAND2_X1 U3418 ( .A1(n4895), .A2(n3077), .ZN(n2941) );
  NAND2_X1 U3419 ( .A1(n2942), .A2(n2941), .ZN(n2943) );
  XNOR2_X1 U3420 ( .A(n2943), .B(n2734), .ZN(n2945) );
  XOR2_X1 U3421 ( .A(n2944), .B(n2945), .Z(n4882) );
  NAND2_X1 U3422 ( .A1(n3081), .A2(REG0_REG_17__SCAN_IN), .ZN(n2951) );
  NAND2_X1 U3423 ( .A1(n2262), .A2(REG2_REG_17__SCAN_IN), .ZN(n2950) );
  OAI21_X1 U3424 ( .B1(REG3_REG_17__SCAN_IN), .B2(n2946), .A(n2958), .ZN(n4004) );
  INV_X1 U3425 ( .A(n4004), .ZN(n2947) );
  NAND2_X1 U3426 ( .A1(n3071), .A2(n2947), .ZN(n2949) );
  NAND2_X1 U3427 ( .A1(n2810), .A2(REG1_REG_17__SCAN_IN), .ZN(n2948) );
  NAND4_X1 U3428 ( .A1(n2951), .A2(n2950), .A3(n2949), .A4(n2948), .ZN(n4054)
         );
  NAND2_X1 U3429 ( .A1(n4054), .A2(n3091), .ZN(n2953) );
  MUX2_X1 U3430 ( .A(DATAI_17_), .B(n4380), .S(n3738), .Z(n4001) );
  NAND2_X1 U3431 ( .A1(n4001), .A2(n3077), .ZN(n2952) );
  NAND2_X1 U3432 ( .A1(n2953), .A2(n2952), .ZN(n2954) );
  XNOR2_X1 U3433 ( .A(n2954), .B(n2734), .ZN(n3998) );
  NAND2_X1 U3434 ( .A1(n4054), .A2(n2737), .ZN(n2956) );
  NAND2_X1 U3435 ( .A1(n4001), .A2(n2766), .ZN(n2955) );
  NAND2_X1 U3436 ( .A1(n2956), .A2(n2955), .ZN(n2957) );
  INV_X1 U3437 ( .A(n2957), .ZN(n3997) );
  NAND2_X1 U3438 ( .A1(n3081), .A2(REG0_REG_18__SCAN_IN), .ZN(n2962) );
  NAND2_X1 U3439 ( .A1(n2262), .A2(REG2_REG_18__SCAN_IN), .ZN(n2961) );
  AOI21_X1 U3440 ( .B1(n4035), .B2(n2958), .A(n2972), .ZN(n4034) );
  NAND2_X1 U3441 ( .A1(n3071), .A2(n4034), .ZN(n2960) );
  NAND2_X1 U3442 ( .A1(n2810), .A2(REG1_REG_18__SCAN_IN), .ZN(n2959) );
  NAND4_X1 U3443 ( .A1(n2962), .A2(n2961), .A3(n2960), .A4(n2959), .ZN(n4927)
         );
  NAND2_X1 U3444 ( .A1(n4927), .A2(n2261), .ZN(n2964) );
  MUX2_X1 U3445 ( .A(DATAI_18_), .B(n3259), .S(n3738), .Z(n4036) );
  NAND2_X1 U3446 ( .A1(n4036), .A2(n3077), .ZN(n2963) );
  NAND2_X1 U3447 ( .A1(n2964), .A2(n2963), .ZN(n2965) );
  XNOR2_X1 U3448 ( .A(n2965), .B(n3066), .ZN(n2968) );
  INV_X1 U3449 ( .A(n4036), .ZN(n4267) );
  NOR2_X1 U3450 ( .A1(n4267), .A2(n2717), .ZN(n2966) );
  AOI21_X1 U3451 ( .B1(n4927), .B2(n2737), .A(n2966), .ZN(n2967) );
  NAND2_X1 U3452 ( .A1(n2968), .A2(n2967), .ZN(n4030) );
  NOR2_X1 U3453 ( .A1(n2968), .A2(n2967), .ZN(n4029) );
  XNOR2_X1 U3454 ( .A(n2971), .B(n2969), .ZN(n4930) );
  NAND2_X1 U3455 ( .A1(n4929), .A2(n4930), .ZN(n4928) );
  INV_X1 U3456 ( .A(n2986), .ZN(n2987) );
  INV_X1 U3457 ( .A(n2973), .ZN(n2975) );
  INV_X1 U34580 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2974) );
  NAND2_X1 U34590 ( .A1(n2975), .A2(n2974), .ZN(n2976) );
  NAND2_X1 U3460 ( .A1(n2987), .A2(n2976), .ZN(n4947) );
  INV_X1 U3461 ( .A(n4947), .ZN(n4257) );
  NAND2_X1 U3462 ( .A1(n3071), .A2(n4257), .ZN(n2980) );
  NAND2_X1 U3463 ( .A1(n2262), .A2(REG2_REG_20__SCAN_IN), .ZN(n2979) );
  NAND2_X1 U3464 ( .A1(n2810), .A2(REG1_REG_20__SCAN_IN), .ZN(n2978) );
  NAND2_X1 U3465 ( .A1(n3081), .A2(REG0_REG_20__SCAN_IN), .ZN(n2977) );
  NAND2_X1 U3466 ( .A1(n4958), .A2(n2261), .ZN(n2983) );
  INV_X1 U34670 ( .A(DATAI_20_), .ZN(n2981) );
  NAND2_X1 U3468 ( .A1(n4942), .A2(n3077), .ZN(n2982) );
  NAND2_X1 U34690 ( .A1(n2983), .A2(n2982), .ZN(n2984) );
  XNOR2_X1 U3470 ( .A(n2984), .B(n3066), .ZN(n2999) );
  NOR2_X1 U34710 ( .A1(n4253), .A2(n2767), .ZN(n2985) );
  AOI21_X1 U3472 ( .B1(n4958), .B2(n2737), .A(n2985), .ZN(n2998) );
  OR2_X1 U34730 ( .A1(n2999), .A2(n2998), .ZN(n4952) );
  NAND2_X1 U3474 ( .A1(n3081), .A2(REG0_REG_21__SCAN_IN), .ZN(n2992) );
  NAND2_X1 U34750 ( .A1(n2262), .A2(REG2_REG_21__SCAN_IN), .ZN(n2991) );
  INV_X1 U3476 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4548) );
  NAND2_X1 U34770 ( .A1(n2987), .A2(n4548), .ZN(n2988) );
  NAND2_X1 U3478 ( .A1(n3016), .A2(n2988), .ZN(n4965) );
  INV_X1 U34790 ( .A(n4965), .ZN(n3928) );
  NAND2_X1 U3480 ( .A1(n3071), .A2(n3928), .ZN(n2990) );
  NAND2_X1 U34810 ( .A1(n2810), .A2(REG1_REG_21__SCAN_IN), .ZN(n2989) );
  NAND4_X1 U3482 ( .A1(n2992), .A2(n2991), .A3(n2990), .A4(n2989), .ZN(n4939)
         );
  NAND2_X1 U34830 ( .A1(n4939), .A2(n3091), .ZN(n2995) );
  INV_X1 U3484 ( .A(DATAI_21_), .ZN(n2993) );
  NAND2_X1 U34850 ( .A1(n4959), .A2(n3077), .ZN(n2994) );
  NAND2_X1 U3486 ( .A1(n2995), .A2(n2994), .ZN(n2996) );
  XNOR2_X1 U34870 ( .A(n2996), .B(n3066), .ZN(n3001) );
  NOR2_X1 U3488 ( .A1(n3926), .A2(n2717), .ZN(n2997) );
  AOI21_X1 U34890 ( .B1(n4939), .B2(n2737), .A(n2997), .ZN(n3000) );
  AND2_X1 U3490 ( .A1(n3001), .A2(n3000), .ZN(n4950) );
  AND2_X1 U34910 ( .A1(n2999), .A2(n2998), .ZN(n4953) );
  AOI211_X1 U3492 ( .C1(n4954), .C2(n4952), .A(n4950), .B(n4953), .ZN(n3002)
         );
  NOR2_X1 U34930 ( .A1(n3001), .A2(n3000), .ZN(n4951) );
  NAND2_X1 U3494 ( .A1(n3081), .A2(REG0_REG_22__SCAN_IN), .ZN(n3006) );
  NAND2_X1 U34950 ( .A1(n2810), .A2(REG1_REG_22__SCAN_IN), .ZN(n3005) );
  XNOR2_X1 U3496 ( .A(n3016), .B(REG3_REG_22__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U34970 ( .A1(n3071), .A2(n4238), .ZN(n3004) );
  NAND2_X1 U3498 ( .A1(n2262), .A2(REG2_REG_22__SCAN_IN), .ZN(n3003) );
  OAI22_X1 U34990 ( .A1(n4214), .A2(n2689), .B1(n2717), .B2(n4235), .ZN(n3010)
         );
  OAI22_X1 U3500 ( .A1(n4214), .A2(n2767), .B1(n3007), .B2(n4235), .ZN(n3008)
         );
  XNOR2_X1 U35010 ( .A(n3008), .B(n2734), .ZN(n3009) );
  XOR2_X1 U3502 ( .A(n3010), .B(n3009), .Z(n4021) );
  NAND2_X1 U35030 ( .A1(n4020), .A2(n4021), .ZN(n4019) );
  NAND2_X1 U3504 ( .A1(n4019), .A2(n3013), .ZN(n3976) );
  NAND2_X1 U35050 ( .A1(n2810), .A2(REG1_REG_23__SCAN_IN), .ZN(n3021) );
  NAND2_X1 U35060 ( .A1(n3081), .A2(REG0_REG_23__SCAN_IN), .ZN(n3020) );
  INV_X1 U35070 ( .A(n3016), .ZN(n3015) );
  AND2_X1 U35080 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n3014) );
  NAND2_X1 U35090 ( .A1(n3015), .A2(n3014), .ZN(n3030) );
  INV_X1 U35100 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4023) );
  INV_X1 U35110 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4394) );
  OAI21_X1 U35120 ( .B1(n3016), .B2(n4023), .A(n4394), .ZN(n3017) );
  AND2_X1 U35130 ( .A1(n3030), .A2(n3017), .ZN(n4222) );
  NAND2_X1 U35140 ( .A1(n3071), .A2(n4222), .ZN(n3019) );
  NAND2_X1 U35150 ( .A1(n2262), .A2(REG2_REG_23__SCAN_IN), .ZN(n3018) );
  NAND4_X1 U35160 ( .A1(n3021), .A2(n3020), .A3(n3019), .A4(n3018), .ZN(n4232)
         );
  INV_X1 U35170 ( .A(DATAI_23_), .ZN(n4419) );
  INV_X1 U35180 ( .A(n3971), .ZN(n4221) );
  NOR2_X1 U35190 ( .A1(n4221), .A2(n2767), .ZN(n3022) );
  AOI21_X1 U35200 ( .B1(n4232), .B2(n2737), .A(n3022), .ZN(n3027) );
  NAND2_X1 U35210 ( .A1(n4232), .A2(n2766), .ZN(n3024) );
  NAND2_X1 U35220 ( .A1(n3971), .A2(n3077), .ZN(n3023) );
  NAND2_X1 U35230 ( .A1(n3024), .A2(n3023), .ZN(n3025) );
  XNOR2_X1 U35240 ( .A(n3025), .B(n2734), .ZN(n3026) );
  XOR2_X1 U35250 ( .A(n3027), .B(n3026), .Z(n3977) );
  INV_X1 U35260 ( .A(n3026), .ZN(n3028) );
  NAND2_X1 U35270 ( .A1(n2810), .A2(REG1_REG_24__SCAN_IN), .ZN(n3035) );
  NAND2_X1 U35280 ( .A1(n3081), .A2(REG0_REG_24__SCAN_IN), .ZN(n3034) );
  INV_X1 U35290 ( .A(n3030), .ZN(n3029) );
  NAND2_X1 U35300 ( .A1(n3029), .A2(REG3_REG_24__SCAN_IN), .ZN(n3042) );
  INV_X1 U35310 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4557) );
  NAND2_X1 U35320 ( .A1(n3030), .A2(n4557), .ZN(n3031) );
  AND2_X1 U35330 ( .A1(n3042), .A2(n3031), .ZN(n4196) );
  NAND2_X1 U35340 ( .A1(n3071), .A2(n4196), .ZN(n3033) );
  NAND2_X1 U35350 ( .A1(n2262), .A2(REG2_REG_24__SCAN_IN), .ZN(n3032) );
  NAND2_X1 U35360 ( .A1(n4216), .A2(n2737), .ZN(n3038) );
  INV_X1 U35370 ( .A(DATAI_24_), .ZN(n3036) );
  NAND2_X1 U35380 ( .A1(n4012), .A2(n3091), .ZN(n3037) );
  NAND2_X1 U35390 ( .A1(n3038), .A2(n3037), .ZN(n4010) );
  NAND2_X1 U35400 ( .A1(n4216), .A2(n3091), .ZN(n3040) );
  NAND2_X1 U35410 ( .A1(n4012), .A2(n3077), .ZN(n3039) );
  NAND2_X1 U35420 ( .A1(n3040), .A2(n3039), .ZN(n3041) );
  XNOR2_X1 U35430 ( .A(n3041), .B(n2734), .ZN(n3984) );
  NAND2_X1 U35440 ( .A1(n3081), .A2(REG0_REG_25__SCAN_IN), .ZN(n3047) );
  NAND2_X1 U35450 ( .A1(n2810), .A2(REG1_REG_25__SCAN_IN), .ZN(n3046) );
  INV_X1 U35460 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4483) );
  NAND2_X1 U35470 ( .A1(n3042), .A2(n4483), .ZN(n3043) );
  AND2_X1 U35480 ( .A1(n3057), .A2(n3043), .ZN(n3992) );
  NAND2_X1 U35490 ( .A1(n3071), .A2(n3992), .ZN(n3045) );
  NAND2_X1 U35500 ( .A1(n2262), .A2(REG2_REG_25__SCAN_IN), .ZN(n3044) );
  NAND4_X1 U35510 ( .A1(n3047), .A2(n3046), .A3(n3045), .A4(n3044), .ZN(n4190)
         );
  NAND2_X1 U35520 ( .A1(n4190), .A2(n2766), .ZN(n3049) );
  INV_X1 U35530 ( .A(DATAI_25_), .ZN(n4408) );
  NAND2_X1 U35540 ( .A1(n3993), .A2(n3077), .ZN(n3048) );
  NAND2_X1 U35550 ( .A1(n3049), .A2(n3048), .ZN(n3050) );
  XNOR2_X1 U35560 ( .A(n3050), .B(n3066), .ZN(n3052) );
  NOR2_X1 U35570 ( .A1(n3191), .A2(n2767), .ZN(n3051) );
  AOI21_X1 U35580 ( .B1(n4190), .B2(n2737), .A(n3051), .ZN(n3981) );
  NOR2_X1 U35590 ( .A1(n3052), .A2(n3981), .ZN(n3990) );
  AOI21_X1 U35600 ( .B1(n4010), .B2(n3984), .A(n3990), .ZN(n3056) );
  INV_X1 U35610 ( .A(n3984), .ZN(n3987) );
  INV_X1 U35620 ( .A(n4010), .ZN(n3986) );
  AOI21_X1 U35630 ( .B1(n3987), .B2(n3986), .A(n3981), .ZN(n3054) );
  INV_X1 U35640 ( .A(n3052), .ZN(n3983) );
  NAND2_X1 U35650 ( .A1(n3986), .A2(n3981), .ZN(n3053) );
  OAI22_X1 U35660 ( .A1(n3054), .A2(n3983), .B1(n3984), .B2(n3053), .ZN(n3055)
         );
  NAND2_X1 U35670 ( .A1(n2810), .A2(REG1_REG_26__SCAN_IN), .ZN(n3062) );
  NAND2_X1 U35680 ( .A1(n3081), .A2(REG0_REG_26__SCAN_IN), .ZN(n3061) );
  INV_X1 U35690 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U35700 ( .A1(n3057), .A2(n4045), .ZN(n3058) );
  NAND2_X1 U35710 ( .A1(n3085), .A2(n3058), .ZN(n4049) );
  INV_X1 U35720 ( .A(n4049), .ZN(n4163) );
  NAND2_X1 U35730 ( .A1(n3071), .A2(n4163), .ZN(n3060) );
  NAND2_X1 U35740 ( .A1(n2262), .A2(REG2_REG_26__SCAN_IN), .ZN(n3059) );
  NAND2_X1 U35750 ( .A1(n4175), .A2(n2261), .ZN(n3065) );
  INV_X1 U35760 ( .A(DATAI_26_), .ZN(n3063) );
  NAND2_X1 U35770 ( .A1(n4160), .A2(n3077), .ZN(n3064) );
  NAND2_X1 U35780 ( .A1(n3065), .A2(n3064), .ZN(n3067) );
  XNOR2_X1 U35790 ( .A(n3067), .B(n3066), .ZN(n3070) );
  INV_X1 U35800 ( .A(n4160), .ZN(n3227) );
  NOR2_X1 U35810 ( .A1(n3227), .A2(n2717), .ZN(n3068) );
  AOI21_X1 U3582 ( .B1(n4175), .B2(n2737), .A(n3068), .ZN(n3069) );
  NAND2_X1 U3583 ( .A1(n3070), .A2(n3069), .ZN(n4042) );
  INV_X1 U3584 ( .A(n3949), .ZN(n3080) );
  NAND2_X1 U3585 ( .A1(n3081), .A2(REG0_REG_27__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U3586 ( .A1(n2810), .A2(REG1_REG_27__SCAN_IN), .ZN(n3074) );
  XNOR2_X1 U3587 ( .A(n3085), .B(REG3_REG_27__SCAN_IN), .ZN(n4141) );
  NAND2_X1 U3588 ( .A1(n3071), .A2(n4141), .ZN(n3073) );
  NAND2_X1 U3589 ( .A1(n2262), .A2(REG2_REG_27__SCAN_IN), .ZN(n3072) );
  INV_X1 U3590 ( .A(DATAI_27_), .ZN(n3076) );
  AOI22_X1 U3591 ( .A1(n4156), .A2(n2737), .B1(n2766), .B2(n4136), .ZN(n3116)
         );
  AOI22_X1 U3592 ( .A1(n4156), .A2(n2261), .B1(n4136), .B2(n3077), .ZN(n3079)
         );
  XNOR2_X1 U3593 ( .A(n3079), .B(n2734), .ZN(n3117) );
  XOR2_X1 U3594 ( .A(n3116), .B(n3117), .Z(n3948) );
  NAND2_X1 U3595 ( .A1(n3080), .A2(n3948), .ZN(n3119) );
  INV_X1 U3596 ( .A(n3119), .ZN(n3115) );
  NAND2_X1 U3597 ( .A1(n2810), .A2(REG1_REG_28__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3598 ( .A1(n3081), .A2(REG0_REG_28__SCAN_IN), .ZN(n3089) );
  INV_X1 U3599 ( .A(n3085), .ZN(n3083) );
  AND2_X1 U3600 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n3082) );
  NAND2_X1 U3601 ( .A1(n3083), .A2(n3082), .ZN(n3132) );
  INV_X1 U3602 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3084) );
  INV_X1 U3603 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3139) );
  OAI21_X1 U3604 ( .B1(n3085), .B2(n3084), .A(n3139), .ZN(n3086) );
  NAND2_X1 U3605 ( .A1(n3071), .A2(n4119), .ZN(n3088) );
  NAND2_X1 U3606 ( .A1(n2262), .A2(REG2_REG_28__SCAN_IN), .ZN(n3087) );
  NAND4_X1 U3607 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .ZN(n4137)
         );
  NAND2_X1 U3608 ( .A1(n4137), .A2(n3091), .ZN(n3094) );
  INV_X1 U3609 ( .A(DATAI_28_), .ZN(n3092) );
  NAND2_X1 U3610 ( .A1(n3249), .A2(n3077), .ZN(n3093) );
  NAND2_X1 U3611 ( .A1(n3094), .A2(n3093), .ZN(n3095) );
  XNOR2_X1 U3612 ( .A(n3095), .B(n2734), .ZN(n3097) );
  AOI22_X1 U3613 ( .A1(n4137), .A2(n2737), .B1(n2766), .B2(n3249), .ZN(n3096)
         );
  XNOR2_X1 U3614 ( .A(n3097), .B(n3096), .ZN(n3118) );
  INV_X1 U3615 ( .A(n3118), .ZN(n3121) );
  NAND2_X1 U3616 ( .A1(n3110), .A2(n3257), .ZN(n3098) );
  MUX2_X1 U3617 ( .A(n3257), .B(n3098), .S(B_REG_SCAN_IN), .Z(n3099) );
  NOR4_X1 U3618 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n3108) );
  NOR4_X1 U3619 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n3107) );
  OR4_X1 U3620 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n3105) );
  NOR4_X1 U3621 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n3103) );
  NOR4_X1 U3622 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n3102) );
  NOR4_X1 U3623 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n3101) );
  NOR4_X1 U3624 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n3100) );
  NAND4_X1 U3625 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n3104)
         );
  NOR4_X1 U3626 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(n3105), 
        .A4(n3104), .ZN(n3106) );
  AND3_X1 U3627 ( .A1(n3108), .A2(n3107), .A3(n3106), .ZN(n3109) );
  NOR2_X1 U3628 ( .A1(n3267), .A2(n3109), .ZN(n3241) );
  INV_X1 U3629 ( .A(n3269), .ZN(n3111) );
  NAND2_X1 U3630 ( .A1(n3111), .A2(n3110), .ZN(n4377) );
  OAI21_X1 U3631 ( .B1(n3267), .B2(D_REG_1__SCAN_IN), .A(n4377), .ZN(n3428) );
  NOR2_X1 U3632 ( .A1(n3241), .A2(n3428), .ZN(n3123) );
  NAND2_X1 U3633 ( .A1(n3268), .A2(n3123), .ZN(n3112) );
  NAND2_X1 U3634 ( .A1(n2687), .A2(n4787), .ZN(n3126) );
  AOI21_X1 U3635 ( .B1(n3126), .B2(n4705), .A(n3237), .ZN(n3113) );
  AND2_X2 U3636 ( .A1(n3144), .A2(n3113), .ZN(n4961) );
  AND2_X1 U3637 ( .A1(n3121), .A2(n4961), .ZN(n3114) );
  NAND2_X1 U3638 ( .A1(n3115), .A2(n3114), .ZN(n3154) );
  OR2_X1 U3639 ( .A1(n3117), .A2(n3116), .ZN(n3120) );
  NAND4_X1 U3640 ( .A1(n3119), .A2(n4961), .A3(n3118), .A4(n3120), .ZN(n3153)
         );
  INV_X1 U3641 ( .A(n3120), .ZN(n3122) );
  NAND3_X1 U3642 ( .A1(n3122), .A2(n4961), .A3(n3121), .ZN(n3151) );
  INV_X1 U3643 ( .A(n3429), .ZN(n3245) );
  NAND2_X1 U3644 ( .A1(n3245), .A2(n3123), .ZN(n3129) );
  OR2_X1 U3645 ( .A1(n4787), .A2(n3124), .ZN(n3125) );
  NAND2_X1 U3646 ( .A1(n3129), .A2(n3125), .ZN(n3303) );
  NAND2_X1 U3647 ( .A1(n3126), .A2(n3237), .ZN(n3242) );
  NAND3_X1 U3648 ( .A1(n3303), .A2(n2704), .A3(n3242), .ZN(n3127) );
  NAND2_X1 U3649 ( .A1(n3127), .A2(STATE_REG_SCAN_IN), .ZN(n3131) );
  INV_X1 U3650 ( .A(n2687), .ZN(n3878) );
  NOR2_X1 U3651 ( .A1(n4780), .A2(U3149), .ZN(n3128) );
  NAND2_X1 U3652 ( .A1(n3129), .A2(n3128), .ZN(n3302) );
  AND2_X1 U3653 ( .A1(n3302), .A2(n4388), .ZN(n3130) );
  INV_X1 U3654 ( .A(n4966), .ZN(n4026) );
  NAND2_X1 U3655 ( .A1(n2810), .A2(REG1_REG_29__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U3656 ( .A1(n3081), .A2(REG0_REG_29__SCAN_IN), .ZN(n3135) );
  INV_X1 U3657 ( .A(n3132), .ZN(n3959) );
  NAND2_X1 U3658 ( .A1(n3071), .A2(n3959), .ZN(n3134) );
  NAND2_X1 U3659 ( .A1(n2262), .A2(REG2_REG_29__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U3660 ( .A1(n3325), .A2(n4787), .ZN(n3137) );
  OR2_X1 U3661 ( .A1(n3142), .A2(n3231), .ZN(n3197) );
  NOR2_X1 U3662 ( .A1(n3137), .A2(n3197), .ZN(n3138) );
  OAI22_X1 U3663 ( .A1(n4125), .A2(n4931), .B1(STATE_REG_SCAN_IN), .B2(n3139), 
        .ZN(n3149) );
  INV_X1 U3664 ( .A(n3325), .ZN(n3318) );
  INV_X1 U3665 ( .A(n3140), .ZN(n3141) );
  NAND2_X1 U3666 ( .A1(n3318), .A2(n3141), .ZN(n3888) );
  NOR2_X1 U3667 ( .A1(n3888), .A2(n3142), .ZN(n3143) );
  INV_X1 U3668 ( .A(n4957), .ZN(n4588) );
  NAND2_X1 U3669 ( .A1(n3144), .A2(n4896), .ZN(n3147) );
  NOR2_X1 U3670 ( .A1(n3145), .A2(n3800), .ZN(n3146) );
  AND2_X1 U3671 ( .A1(n2687), .A2(n4379), .ZN(n4710) );
  INV_X1 U3672 ( .A(n4960), .ZN(n4858) );
  INV_X1 U3673 ( .A(n3249), .ZN(n4126) );
  OAI22_X1 U3674 ( .A1(n4127), .A2(n4588), .B1(n4858), .B2(n4126), .ZN(n3148)
         );
  AOI211_X1 U3675 ( .C1(n4119), .C2(n4026), .A(n3149), .B(n3148), .ZN(n3150)
         );
  NAND3_X1 U3676 ( .A1(n3154), .A2(n3153), .A3(n3152), .ZN(U3217) );
  INV_X1 U3677 ( .A(n4136), .ZN(n4145) );
  INV_X1 U3678 ( .A(n4190), .ZN(n4159) );
  NAND2_X1 U3679 ( .A1(n4066), .A2(n3155), .ZN(n3824) );
  NAND2_X1 U3680 ( .A1(n3156), .A2(n4731), .ZN(n3821) );
  AND2_X1 U3681 ( .A1(n4721), .A2(n4732), .ZN(n4719) );
  NAND2_X1 U3682 ( .A1(n4066), .A2(n4731), .ZN(n3157) );
  NAND2_X1 U3683 ( .A1(n4718), .A2(n3157), .ZN(n3462) );
  INV_X1 U3684 ( .A(n3462), .ZN(n3158) );
  NAND2_X1 U3685 ( .A1(n4723), .A2(n3477), .ZN(n3820) );
  NAND2_X1 U3686 ( .A1(n4065), .A2(n3469), .ZN(n3827) );
  NAND2_X1 U3687 ( .A1(n3158), .A2(n3767), .ZN(n3464) );
  NAND2_X1 U3688 ( .A1(n4723), .A2(n3469), .ZN(n3159) );
  NAND2_X1 U3689 ( .A1(n3464), .A2(n3159), .ZN(n3350) );
  NOR2_X1 U3690 ( .A1(n4064), .A2(n3354), .ZN(n3160) );
  INV_X1 U3691 ( .A(n4064), .ZN(n3201) );
  OAI22_X2 U3692 ( .A1(n3350), .A2(n3160), .B1(n3201), .B2(n3360), .ZN(n3415)
         );
  INV_X1 U3693 ( .A(n4063), .ZN(n3374) );
  NAND2_X1 U3694 ( .A1(n3374), .A2(n3409), .ZN(n3202) );
  NAND2_X1 U3695 ( .A1(n4063), .A2(n3421), .ZN(n3833) );
  NAND2_X1 U3696 ( .A1(n3202), .A2(n3833), .ZN(n3414) );
  NAND2_X1 U3697 ( .A1(n3415), .A2(n3414), .ZN(n3162) );
  NAND2_X1 U3698 ( .A1(n4063), .A2(n3409), .ZN(n3161) );
  AND2_X1 U3699 ( .A1(n4062), .A2(n3403), .ZN(n3163) );
  INV_X1 U3700 ( .A(n4062), .ZN(n3485) );
  INV_X1 U3701 ( .A(n3403), .ZN(n3247) );
  NAND2_X1 U3702 ( .A1(n3485), .A2(n3247), .ZN(n3164) );
  NOR2_X1 U3703 ( .A1(n4783), .A2(n3454), .ZN(n3165) );
  INV_X1 U3704 ( .A(n4061), .ZN(n3536) );
  NAND2_X1 U3705 ( .A1(n3536), .A2(n4774), .ZN(n3835) );
  NAND2_X1 U3706 ( .A1(n4061), .A2(n4779), .ZN(n3803) );
  NAND2_X1 U3707 ( .A1(n3835), .A2(n3803), .ZN(n4789) );
  NAND2_X1 U3708 ( .A1(n4788), .A2(n4789), .ZN(n3167) );
  NAND2_X1 U3709 ( .A1(n4061), .A2(n4774), .ZN(n3166) );
  AND2_X1 U3710 ( .A1(n4060), .A2(n3501), .ZN(n3168) );
  OAI22_X1 U3711 ( .A1(n3533), .A2(n3168), .B1(n3501), .B2(n4060), .ZN(n3508)
         );
  INV_X1 U3712 ( .A(n3508), .ZN(n3169) );
  NAND2_X1 U3713 ( .A1(n4059), .A2(n3523), .ZN(n3170) );
  INV_X1 U3714 ( .A(n4058), .ZN(n3205) );
  NAND2_X1 U3715 ( .A1(n3205), .A2(n3624), .ZN(n3171) );
  NAND2_X1 U3716 ( .A1(n3172), .A2(n3171), .ZN(n3592) );
  INV_X1 U3717 ( .A(n4057), .ZN(n4589) );
  NAND2_X1 U3718 ( .A1(n4589), .A2(n3594), .ZN(n3557) );
  NAND2_X1 U3719 ( .A1(n4057), .A2(n3590), .ZN(n3559) );
  NAND2_X1 U3720 ( .A1(n3557), .A2(n3559), .ZN(n3777) );
  NOR2_X1 U3721 ( .A1(n4057), .A2(n3594), .ZN(n3173) );
  AOI21_X2 U3722 ( .B1(n3592), .B2(n3777), .A(n3173), .ZN(n3556) );
  INV_X1 U3723 ( .A(n4056), .ZN(n3210) );
  NAND2_X1 U3724 ( .A1(n3210), .A2(n4587), .ZN(n3174) );
  NAND2_X1 U3725 ( .A1(n3556), .A2(n3174), .ZN(n3176) );
  NAND2_X1 U3726 ( .A1(n4056), .A2(n3209), .ZN(n3175) );
  NAND2_X1 U3727 ( .A1(n3176), .A2(n3175), .ZN(n3602) );
  INV_X1 U3728 ( .A(n4591), .ZN(n3560) );
  NAND2_X1 U3729 ( .A1(n3560), .A2(n3615), .ZN(n3668) );
  NAND2_X1 U3730 ( .A1(n3602), .A2(n3668), .ZN(n3179) );
  INV_X1 U3731 ( .A(n4862), .ZN(n3610) );
  NAND2_X1 U3732 ( .A1(n3610), .A2(n3695), .ZN(n3720) );
  INV_X1 U3733 ( .A(n3695), .ZN(n3683) );
  NAND2_X1 U3734 ( .A1(n4862), .A2(n3683), .ZN(n3721) );
  NAND2_X1 U3735 ( .A1(n3720), .A2(n3721), .ZN(n3679) );
  NAND2_X1 U3736 ( .A1(n4898), .A2(n3248), .ZN(n3180) );
  NAND2_X1 U3737 ( .A1(n4591), .A2(n3651), .ZN(n3667) );
  NAND2_X1 U3738 ( .A1(n3179), .A2(n3178), .ZN(n3182) );
  NOR2_X1 U3739 ( .A1(n4862), .A2(n3695), .ZN(n3670) );
  INV_X1 U3740 ( .A(n4898), .ZN(n3217) );
  AOI22_X1 U3741 ( .A1(n3670), .A2(n3180), .B1(n3217), .B2(n4857), .ZN(n3181)
         );
  NAND2_X1 U3742 ( .A1(n3182), .A2(n3181), .ZN(n4903) );
  INV_X1 U3743 ( .A(n4895), .ZN(n3183) );
  NOR2_X1 U3744 ( .A1(n4055), .A2(n3183), .ZN(n3854) );
  NAND2_X1 U3745 ( .A1(n4055), .A2(n4895), .ZN(n3184) );
  INV_X1 U3746 ( .A(n4278), .ZN(n3185) );
  NAND2_X1 U3747 ( .A1(n3903), .A2(n4036), .ZN(n3898) );
  NAND2_X1 U3748 ( .A1(n4927), .A2(n4267), .ZN(n3899) );
  NAND2_X1 U3749 ( .A1(n3898), .A2(n3899), .ZN(n4269) );
  INV_X1 U3750 ( .A(n4269), .ZN(n4279) );
  NAND2_X1 U3751 ( .A1(n3185), .A2(n4269), .ZN(n4276) );
  NAND2_X1 U3752 ( .A1(n3903), .A2(n4267), .ZN(n3186) );
  NAND2_X1 U3753 ( .A1(n4276), .A2(n3186), .ZN(n3893) );
  NAND2_X1 U3754 ( .A1(n4944), .A2(n4926), .ZN(n3188) );
  NOR2_X1 U3755 ( .A1(n4944), .A2(n4926), .ZN(n3187) );
  AOI21_X2 U3756 ( .B1(n3893), .B2(n3188), .A(n3187), .ZN(n4244) );
  INV_X1 U3757 ( .A(n4958), .ZN(n4932) );
  NAND2_X1 U3758 ( .A1(n4932), .A2(n4253), .ZN(n3189) );
  NAND2_X1 U3759 ( .A1(n4939), .A2(n4959), .ZN(n4201) );
  OR2_X1 U3760 ( .A1(n4214), .A2(n4239), .ZN(n3225) );
  NAND2_X1 U3761 ( .A1(n4214), .A2(n4239), .ZN(n4211) );
  NOR2_X1 U3762 ( .A1(n4939), .A2(n4959), .ZN(n4202) );
  NOR2_X1 U3763 ( .A1(n4214), .A2(n4235), .ZN(n4205) );
  INV_X1 U3764 ( .A(n4216), .ZN(n4173) );
  NOR2_X1 U3765 ( .A1(n4173), .A2(n4193), .ZN(n3190) );
  OAI22_X1 U3766 ( .A1(n4185), .A2(n3190), .B1(n4012), .B2(n4216), .ZN(n4168)
         );
  AOI21_X1 U3767 ( .B1(n4136), .B2(n4156), .A(n3194), .ZN(n4118) );
  INV_X1 U3768 ( .A(n4137), .ZN(n3238) );
  NAND2_X1 U3769 ( .A1(n3238), .A2(n3249), .ZN(n3742) );
  NAND2_X1 U3770 ( .A1(n4137), .A2(n4126), .ZN(n3746) );
  OAI22_X1 U3771 ( .A1(n4118), .A2(n4123), .B1(n3238), .B2(n4126), .ZN(n3196)
         );
  INV_X1 U3772 ( .A(DATAI_29_), .ZN(n3195) );
  NOR2_X1 U3773 ( .A1(n3738), .A2(n3195), .ZN(n3745) );
  XNOR2_X1 U3774 ( .A(n4125), .B(n3745), .ZN(n3199) );
  XNOR2_X1 U3775 ( .A(n3196), .B(n3199), .ZN(n3962) );
  INV_X1 U3776 ( .A(n4844), .ZN(n3358) );
  OR2_X1 U3777 ( .A1(n3434), .A2(n3889), .ZN(n3198) );
  NAND3_X1 U3778 ( .A1(n3198), .A2(n3197), .A3(n4787), .ZN(n4251) );
  INV_X1 U3779 ( .A(n3199), .ZN(n3798) );
  INV_X1 U3780 ( .A(n4721), .ZN(n3786) );
  NAND2_X1 U3781 ( .A1(n3786), .A2(n4732), .ZN(n4724) );
  NAND2_X1 U3782 ( .A1(n4727), .A2(n3821), .ZN(n3200) );
  NAND2_X1 U3783 ( .A1(n3200), .A2(n3461), .ZN(n3466) );
  NAND2_X1 U3784 ( .A1(n3466), .A2(n3820), .ZN(n3351) );
  NAND2_X1 U3785 ( .A1(n3201), .A2(n3354), .ZN(n3416) );
  NAND2_X1 U3786 ( .A1(n4064), .A2(n3360), .ZN(n3826) );
  NAND2_X1 U3787 ( .A1(n3416), .A2(n3826), .ZN(n3795) );
  INV_X1 U3788 ( .A(n3795), .ZN(n3352) );
  NAND2_X1 U3789 ( .A1(n3351), .A2(n3352), .ZN(n3417) );
  AND2_X1 U3790 ( .A1(n3416), .A2(n3202), .ZN(n3828) );
  AND2_X1 U3791 ( .A1(n4062), .A2(n3247), .ZN(n3369) );
  NAND2_X1 U3792 ( .A1(n3485), .A2(n3403), .ZN(n3805) );
  INV_X1 U3793 ( .A(n3454), .ZN(n3484) );
  NAND2_X1 U3794 ( .A1(n4783), .A2(n3484), .ZN(n3832) );
  NOR2_X1 U3795 ( .A1(n4783), .A2(n3484), .ZN(n3836) );
  NAND2_X1 U3796 ( .A1(n4778), .A2(n3835), .ZN(n3203) );
  NAND2_X1 U3797 ( .A1(n3203), .A2(n3803), .ZN(n3534) );
  INV_X1 U3798 ( .A(n4060), .ZN(n4781) );
  NAND2_X1 U3799 ( .A1(n4781), .A2(n3501), .ZN(n3842) );
  INV_X1 U3800 ( .A(n3501), .ZN(n3535) );
  NAND2_X1 U3801 ( .A1(n4060), .A2(n3535), .ZN(n3802) );
  AND2_X1 U3802 ( .A1(n4059), .A2(n3514), .ZN(n3841) );
  INV_X1 U3803 ( .A(n4059), .ZN(n3204) );
  NAND2_X1 U3804 ( .A1(n3204), .A2(n3523), .ZN(n3843) );
  NAND2_X1 U3805 ( .A1(n4058), .A2(n3624), .ZN(n3808) );
  NAND2_X1 U3806 ( .A1(n3627), .A2(n3808), .ZN(n3206) );
  NAND2_X1 U3807 ( .A1(n3205), .A2(n3628), .ZN(n3807) );
  NAND2_X1 U3808 ( .A1(n3206), .A2(n3807), .ZN(n3593) );
  NAND2_X1 U3809 ( .A1(n4056), .A2(n4587), .ZN(n3603) );
  NAND2_X1 U3810 ( .A1(n4591), .A2(n3615), .ZN(n3207) );
  NAND2_X1 U3811 ( .A1(n3603), .A2(n3207), .ZN(n3211) );
  INV_X1 U3812 ( .A(n3559), .ZN(n3208) );
  NOR2_X1 U3813 ( .A1(n3211), .A2(n3208), .ZN(n3809) );
  NAND2_X1 U3814 ( .A1(n3593), .A2(n3809), .ZN(n3215) );
  NAND2_X1 U3815 ( .A1(n3210), .A2(n3209), .ZN(n3605) );
  NAND2_X1 U3816 ( .A1(n3557), .A2(n3605), .ZN(n3214) );
  INV_X1 U3817 ( .A(n3211), .ZN(n3213) );
  NOR2_X1 U3818 ( .A1(n4591), .A2(n3615), .ZN(n3212) );
  AOI21_X1 U3819 ( .B1(n3214), .B2(n3213), .A(n3212), .ZN(n3813) );
  INV_X1 U3820 ( .A(n3679), .ZN(n3780) );
  NAND2_X1 U3821 ( .A1(n3725), .A2(n3780), .ZN(n3216) );
  NAND2_X1 U3822 ( .A1(n3216), .A2(n3720), .ZN(n3660) );
  NAND2_X1 U3823 ( .A1(n3217), .A2(n3248), .ZN(n3723) );
  NAND2_X1 U3824 ( .A1(n4898), .A2(n4857), .ZN(n3722) );
  NAND2_X1 U3825 ( .A1(n3723), .A2(n3722), .ZN(n3788) );
  NAND2_X1 U3826 ( .A1(n3658), .A2(n3722), .ZN(n4894) );
  NAND2_X1 U3827 ( .A1(n4894), .A2(n4893), .ZN(n4892) );
  INV_X1 U3828 ( .A(n3848), .ZN(n3218) );
  INV_X1 U3829 ( .A(n4926), .ZN(n3908) );
  NAND2_X1 U3830 ( .A1(n4944), .A2(n3908), .ZN(n3219) );
  AND2_X1 U3831 ( .A1(n3899), .A2(n3219), .ZN(n3222) );
  NAND2_X1 U3832 ( .A1(n4054), .A2(n3706), .ZN(n3894) );
  AND2_X1 U3833 ( .A1(n3222), .A2(n3894), .ZN(n3852) );
  INV_X1 U3834 ( .A(n3852), .ZN(n3220) );
  NAND2_X1 U3835 ( .A1(n4902), .A2(n4001), .ZN(n3895) );
  NAND2_X1 U3836 ( .A1(n3898), .A2(n3895), .ZN(n3223) );
  NOR2_X1 U3837 ( .A1(n4944), .A2(n3908), .ZN(n3221) );
  AOI21_X1 U3838 ( .B1(n3223), .B2(n3222), .A(n3221), .ZN(n3728) );
  NOR2_X1 U3839 ( .A1(n4958), .A2(n4253), .ZN(n3784) );
  NAND2_X1 U3840 ( .A1(n4958), .A2(n4253), .ZN(n3851) );
  INV_X1 U3841 ( .A(n4939), .ZN(n4245) );
  NAND2_X1 U3842 ( .A1(n4245), .A2(n4959), .ZN(n4207) );
  NAND2_X1 U3843 ( .A1(n4211), .A2(n4207), .ZN(n3858) );
  AND2_X1 U3844 ( .A1(n4939), .A2(n3926), .ZN(n3855) );
  NAND2_X1 U3845 ( .A1(n4232), .A2(n4221), .ZN(n3224) );
  NAND2_X1 U3846 ( .A1(n3225), .A2(n3224), .ZN(n3861) );
  AOI21_X1 U3847 ( .B1(n3855), .B2(n4211), .A(n3861), .ZN(n3732) );
  OAI21_X1 U3848 ( .B1(n4210), .B2(n3858), .A(n3732), .ZN(n3226) );
  NAND2_X1 U3849 ( .A1(n4188), .A2(n3971), .ZN(n3733) );
  NAND2_X1 U3850 ( .A1(n3226), .A2(n3733), .ZN(n4187) );
  NOR2_X1 U3851 ( .A1(n4216), .A2(n4193), .ZN(n3766) );
  NAND2_X1 U3852 ( .A1(n4216), .A2(n4193), .ZN(n3765) );
  NAND2_X1 U3853 ( .A1(n4190), .A2(n3191), .ZN(n3764) );
  AND2_X1 U3854 ( .A1(n3765), .A2(n3764), .ZN(n3863) );
  NAND2_X1 U3855 ( .A1(n4159), .A2(n3993), .ZN(n4151) );
  NAND2_X1 U3856 ( .A1(n4140), .A2(n4160), .ZN(n3763) );
  NAND2_X1 U3857 ( .A1(n4151), .A2(n3763), .ZN(n3744) );
  NAND2_X1 U3858 ( .A1(n4175), .A2(n3227), .ZN(n3867) );
  AND2_X1 U3859 ( .A1(n4156), .A2(n4145), .ZN(n3871) );
  INV_X1 U3860 ( .A(n3871), .ZN(n3228) );
  NAND2_X1 U3861 ( .A1(n4127), .A2(n4136), .ZN(n3741) );
  INV_X1 U3862 ( .A(n3742), .ZN(n3229) );
  XOR2_X1 U3863 ( .A(n3798), .B(n3230), .Z(n3240) );
  OR2_X1 U3864 ( .A1(n2687), .A2(n3818), .ZN(n3756) );
  OR2_X1 U3865 ( .A1(n4787), .A2(n3231), .ZN(n3232) );
  NAND2_X1 U3866 ( .A1(n2810), .A2(REG1_REG_30__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U3867 ( .A1(n2262), .A2(REG2_REG_30__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U3868 ( .A1(n3081), .A2(REG0_REG_30__SCAN_IN), .ZN(n3233) );
  AND3_X1 U3869 ( .A1(n3235), .A2(n3234), .A3(n3233), .ZN(n3753) );
  NAND2_X1 U3870 ( .A1(n4599), .A2(B_REG_SCAN_IN), .ZN(n3236) );
  NAND2_X1 U3871 ( .A1(n4274), .A2(n3236), .ZN(n4113) );
  NAND2_X1 U3872 ( .A1(n3318), .A2(n3237), .ZN(n4268) );
  INV_X1 U3873 ( .A(n3745), .ZN(n3740) );
  OAI22_X1 U3874 ( .A1(n3238), .A2(n4268), .B1(n4780), .B2(n3740), .ZN(n3239)
         );
  INV_X1 U3875 ( .A(n3241), .ZN(n3430) );
  AND2_X1 U3876 ( .A1(n4844), .A2(n3818), .ZN(n3243) );
  NAND2_X1 U3877 ( .A1(n3268), .A2(n3242), .ZN(n3301) );
  NOR2_X1 U3878 ( .A1(n3243), .A2(n3301), .ZN(n3244) );
  MUX2_X1 U3879 ( .A(REG1_REG_29__SCAN_IN), .B(n3252), .S(n4911), .Z(n3246) );
  INV_X1 U3880 ( .A(n3246), .ZN(n3250) );
  NOR2_X1 U3881 ( .A1(n4731), .A2(n4732), .ZN(n4730) );
  NAND2_X1 U3882 ( .A1(n3475), .A2(n3360), .ZN(n3410) );
  NAND2_X1 U3883 ( .A1(n3413), .A2(n3247), .ZN(n3375) );
  NAND2_X1 U3884 ( .A1(n3530), .A2(n3514), .ZN(n3622) );
  OAI21_X1 U3885 ( .B1(n4120), .B2(n3740), .A(n4288), .ZN(n3958) );
  NAND2_X1 U3886 ( .A1(n3250), .A2(n2494), .ZN(U3547) );
  NAND2_X1 U3887 ( .A1(n3253), .A2(n2498), .ZN(U3515) );
  INV_X1 U3888 ( .A(n3254), .ZN(n3887) );
  NOR2_X1 U3889 ( .A1(n2704), .A2(n3887), .ZN(U4043) );
  NAND2_X1 U3890 ( .A1(n3800), .A2(STATE_REG_SCAN_IN), .ZN(n3255) );
  OAI21_X1 U3891 ( .B1(STATE_REG_SCAN_IN), .B2(n2993), .A(n3255), .ZN(U3331)
         );
  INV_X1 U3892 ( .A(DATAI_22_), .ZN(n4490) );
  NAND2_X1 U3893 ( .A1(n3889), .A2(STATE_REG_SCAN_IN), .ZN(n3256) );
  OAI21_X1 U3894 ( .B1(STATE_REG_SCAN_IN), .B2(n4490), .A(n3256), .ZN(U3330)
         );
  MUX2_X1 U3895 ( .A(n3036), .B(n3257), .S(STATE_REG_SCAN_IN), .Z(n3258) );
  INV_X1 U3896 ( .A(n3258), .ZN(U3328) );
  INV_X1 U3897 ( .A(DATAI_18_), .ZN(n4400) );
  NAND2_X1 U3898 ( .A1(n3259), .A2(STATE_REG_SCAN_IN), .ZN(n3260) );
  OAI21_X1 U3899 ( .B1(STATE_REG_SCAN_IN), .B2(n4400), .A(n3260), .ZN(U3334)
         );
  NAND2_X1 U3900 ( .A1(n3269), .A2(STATE_REG_SCAN_IN), .ZN(n3261) );
  OAI21_X1 U3901 ( .B1(STATE_REG_SCAN_IN), .B2(n3063), .A(n3261), .ZN(U3326)
         );
  NAND2_X1 U3902 ( .A1(n2675), .A2(STATE_REG_SCAN_IN), .ZN(n3262) );
  OAI21_X1 U3903 ( .B1(STATE_REG_SCAN_IN), .B2(n3195), .A(n3262), .ZN(U3323)
         );
  INV_X1 U3904 ( .A(DATAI_30_), .ZN(n3719) );
  NAND2_X1 U3905 ( .A1(n3263), .A2(STATE_REG_SCAN_IN), .ZN(n3264) );
  OAI21_X1 U3906 ( .B1(STATE_REG_SCAN_IN), .B2(n3719), .A(n3264), .ZN(U3322)
         );
  NAND2_X1 U3907 ( .A1(n3878), .A2(STATE_REG_SCAN_IN), .ZN(n3265) );
  OAI21_X1 U3908 ( .B1(STATE_REG_SCAN_IN), .B2(n2981), .A(n3265), .ZN(U3332)
         );
  NAND2_X1 U3909 ( .A1(n3318), .A2(STATE_REG_SCAN_IN), .ZN(n3266) );
  OAI21_X1 U3910 ( .B1(STATE_REG_SCAN_IN), .B2(n3092), .A(n3266), .ZN(U3324)
         );
  INV_X1 U3911 ( .A(D_REG_0__SCAN_IN), .ZN(n3272) );
  NOR3_X1 U3912 ( .A1(n3270), .A2(n3269), .A3(n3887), .ZN(n3271) );
  AOI21_X1 U3913 ( .B1(n4389), .B2(n3272), .A(n3271), .ZN(U3458) );
  INV_X2 U3914 ( .A(U4043), .ZN(n4067) );
  NAND2_X1 U3915 ( .A1(n4067), .A2(DATAO_REG_30__SCAN_IN), .ZN(n3273) );
  OAI21_X1 U3916 ( .B1(n3753), .B2(n4067), .A(n3273), .ZN(U3580) );
  NAND2_X1 U3917 ( .A1(n2810), .A2(REG1_REG_31__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U3918 ( .A1(n2262), .A2(REG2_REG_31__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U3919 ( .A1(n3081), .A2(REG0_REG_31__SCAN_IN), .ZN(n3274) );
  AND3_X1 U3920 ( .A1(n3276), .A2(n3275), .A3(n3274), .ZN(n4114) );
  NAND2_X1 U3921 ( .A1(n4067), .A2(DATAO_REG_31__SCAN_IN), .ZN(n3277) );
  OAI21_X1 U3922 ( .B1(n4114), .B2(n4067), .A(n3277), .ZN(U3581) );
  XNOR2_X1 U3923 ( .A(n3278), .B(REG1_REG_3__SCAN_IN), .ZN(n3285) );
  NOR2_X1 U3924 ( .A1(STATE_REG_SCAN_IN), .A2(n2757), .ZN(n3344) );
  NOR2_X1 U3925 ( .A1(n4703), .A2(n3279), .ZN(n3280) );
  AOI211_X1 U3926 ( .C1(n4697), .C2(ADDR_REG_3__SCAN_IN), .A(n3344), .B(n3280), 
        .ZN(n3284) );
  OAI211_X1 U3927 ( .C1(REG2_REG_3__SCAN_IN), .C2(n3282), .A(n4663), .B(n3281), 
        .ZN(n3283) );
  OAI211_X1 U3928 ( .C1(n3285), .C2(n4680), .A(n3284), .B(n3283), .ZN(U3243)
         );
  MUX2_X1 U3929 ( .A(n2640), .B(REG2_REG_7__SCAN_IN), .S(n4383), .Z(n3287) );
  OAI21_X1 U3930 ( .B1(n3288), .B2(n3287), .A(n4663), .ZN(n3286) );
  AOI21_X1 U3931 ( .B1(n3288), .B2(n3287), .A(n3286), .ZN(n3296) );
  INV_X1 U3932 ( .A(n4383), .ZN(n3294) );
  MUX2_X1 U3933 ( .A(REG1_REG_7__SCAN_IN), .B(n4800), .S(n4383), .Z(n3290) );
  AOI21_X1 U3934 ( .B1(n3290), .B2(n3291), .A(n4680), .ZN(n3289) );
  OAI21_X1 U3935 ( .B1(n3291), .B2(n3290), .A(n3289), .ZN(n3293) );
  AND2_X1 U3936 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3966) );
  AOI21_X1 U3937 ( .B1(n4697), .B2(ADDR_REG_7__SCAN_IN), .A(n3966), .ZN(n3292)
         );
  OAI211_X1 U3938 ( .C1(n4703), .C2(n3294), .A(n3293), .B(n3292), .ZN(n3295)
         );
  OR2_X1 U3939 ( .A1(n3296), .A2(n3295), .ZN(U3247) );
  INV_X1 U3940 ( .A(n3297), .ZN(n3298) );
  AOI21_X1 U3941 ( .B1(n3300), .B2(n3299), .A(n3298), .ZN(n3307) );
  INV_X1 U3942 ( .A(n4961), .ZN(n3975) );
  INV_X1 U3943 ( .A(n3301), .ZN(n3431) );
  NAND3_X1 U3944 ( .A1(n3303), .A2(n3302), .A3(n3431), .ZN(n3338) );
  AOI22_X1 U3945 ( .A1(n4948), .A2(n4064), .B1(n4066), .B2(n4957), .ZN(n3304)
         );
  OAI21_X1 U3946 ( .B1(n4858), .B2(n3469), .A(n3304), .ZN(n3305) );
  AOI21_X1 U3947 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3338), .A(n3305), .ZN(n3306)
         );
  OAI21_X1 U3948 ( .B1(n3307), .B2(n3975), .A(n3306), .ZN(U3234) );
  XOR2_X1 U3949 ( .A(REG1_REG_4__SCAN_IN), .B(n3308), .Z(n3329) );
  INV_X1 U3950 ( .A(n3309), .ZN(n3311) );
  INV_X1 U3951 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U3952 ( .A1(n3311), .A2(n3310), .ZN(n3312) );
  NAND3_X1 U3953 ( .A1(n4663), .A2(n3313), .A3(n3312), .ZN(n3315) );
  AND2_X1 U3954 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3393) );
  AOI21_X1 U3955 ( .B1(n4697), .B2(ADDR_REG_4__SCAN_IN), .A(n3393), .ZN(n3314)
         );
  OAI211_X1 U3956 ( .C1(n4703), .C2(n3316), .A(n3315), .B(n3314), .ZN(n3328)
         );
  INV_X1 U3957 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4716) );
  NAND2_X1 U3958 ( .A1(n4599), .A2(n4716), .ZN(n3317) );
  NAND2_X1 U3959 ( .A1(n3318), .A2(n3317), .ZN(n4600) );
  AOI21_X1 U3960 ( .B1(n4704), .B2(n4707), .A(n2704), .ZN(n3319) );
  NOR3_X1 U3961 ( .A1(n3321), .A2(n3320), .A3(n3319), .ZN(n3323) );
  OR2_X1 U3962 ( .A1(n3323), .A2(n3322), .ZN(n3341) );
  NOR2_X1 U3963 ( .A1(n3341), .A2(n4599), .ZN(n3324) );
  AOI211_X1 U3964 ( .C1(n4599), .C2(n3326), .A(n3325), .B(n3324), .ZN(n3327)
         );
  AOI211_X1 U3965 ( .C1(n4704), .C2(n4600), .A(n4067), .B(n3327), .ZN(n3947)
         );
  AOI211_X1 U3966 ( .C1(n4698), .C2(n3329), .A(n3328), .B(n3947), .ZN(n3330)
         );
  INV_X1 U3967 ( .A(n3330), .ZN(U3244) );
  INV_X1 U3968 ( .A(n3338), .ZN(n3337) );
  INV_X1 U3969 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3336) );
  OAI22_X1 U3970 ( .A1(n3786), .A2(n4588), .B1(n4723), .B2(n4931), .ZN(n3333)
         );
  AOI21_X1 U3971 ( .B1(n4731), .B2(n4960), .A(n3333), .ZN(n3334) );
  OAI211_X1 U3972 ( .C1(n3337), .C2(n3336), .A(n3335), .B(n3334), .ZN(U3219)
         );
  AOI22_X1 U3973 ( .A1(n4066), .A2(n4948), .B1(n4960), .B2(n4732), .ZN(n3340)
         );
  NAND2_X1 U3974 ( .A1(n3338), .A2(REG3_REG_0__SCAN_IN), .ZN(n3339) );
  OAI211_X1 U3975 ( .C1(n3341), .C2(n3975), .A(n3340), .B(n3339), .ZN(U3229)
         );
  XNOR2_X1 U3976 ( .A(n3342), .B(n3343), .ZN(n3348) );
  AOI21_X1 U3977 ( .B1(n4063), .B2(n4948), .A(n3344), .ZN(n3346) );
  AOI22_X1 U3978 ( .A1(n4065), .A2(n4957), .B1(n4960), .B2(n3354), .ZN(n3345)
         );
  OAI211_X1 U3979 ( .C1(n4966), .C2(REG3_REG_3__SCAN_IN), .A(n3346), .B(n3345), 
        .ZN(n3347) );
  AOI21_X1 U3980 ( .B1(n3348), .B2(n4961), .A(n3347), .ZN(n3349) );
  INV_X1 U3981 ( .A(n3349), .ZN(U3215) );
  XNOR2_X1 U3982 ( .A(n3350), .B(n3795), .ZN(n4751) );
  INV_X1 U3983 ( .A(n4751), .ZN(n3359) );
  INV_X1 U3984 ( .A(n4251), .ZN(n4824) );
  OAI21_X1 U3985 ( .B1(n3352), .B2(n3351), .A(n3417), .ZN(n3353) );
  NAND2_X1 U3986 ( .A1(n3353), .A2(n4891), .ZN(n3356) );
  AOI22_X1 U3987 ( .A1(n4063), .A2(n4274), .B1(n4896), .B2(n3354), .ZN(n3355)
         );
  OAI211_X1 U3988 ( .C1(n4723), .C2(n4268), .A(n3356), .B(n3355), .ZN(n3357)
         );
  AOI21_X1 U3989 ( .B1(n4824), .B2(n4751), .A(n3357), .ZN(n4754) );
  OAI21_X1 U3990 ( .B1(n3359), .B2(n3358), .A(n4754), .ZN(n3366) );
  OAI21_X1 U3991 ( .B1(n3475), .B2(n3360), .A(n3410), .ZN(n4749) );
  INV_X1 U3992 ( .A(REG0_REG_3__SCAN_IN), .ZN(n3361) );
  OAI22_X1 U3993 ( .A1(n4749), .A2(n4374), .B1(n4915), .B2(n3361), .ZN(n3362)
         );
  AOI21_X1 U3994 ( .B1(n3366), .B2(n4915), .A(n3362), .ZN(n3363) );
  INV_X1 U3995 ( .A(n3363), .ZN(U3473) );
  INV_X1 U3996 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3364) );
  OAI22_X1 U3997 ( .A1(n4749), .A2(n4334), .B1(n4911), .B2(n3364), .ZN(n3365)
         );
  AOI21_X1 U3998 ( .B1(n3366), .B2(n4911), .A(n3365), .ZN(n3367) );
  INV_X1 U3999 ( .A(n3367), .ZN(U3521) );
  INV_X1 U4000 ( .A(n3369), .ZN(n3831) );
  NAND2_X1 U4001 ( .A1(n3831), .A2(n3805), .ZN(n3775) );
  XOR2_X1 U4002 ( .A(n3368), .B(n3775), .Z(n3440) );
  XNOR2_X1 U4003 ( .A(n3370), .B(n3775), .ZN(n3371) );
  NAND2_X1 U4004 ( .A1(n3371), .A2(n4891), .ZN(n3373) );
  AOI22_X1 U4005 ( .A1(n4783), .A2(n4274), .B1(n4896), .B2(n3403), .ZN(n3372)
         );
  OAI211_X1 U4006 ( .C1(n3374), .C2(n4268), .A(n3373), .B(n3372), .ZN(n3438)
         );
  AOI21_X1 U4007 ( .B1(n3440), .B2(n4877), .A(n3438), .ZN(n3379) );
  INV_X1 U4008 ( .A(n3413), .ZN(n3376) );
  INV_X1 U4009 ( .A(n3375), .ZN(n3481) );
  AOI21_X1 U4010 ( .B1(n3403), .B2(n3376), .A(n3481), .ZN(n3446) );
  INV_X1 U4011 ( .A(n4334), .ZN(n4743) );
  AOI22_X1 U4012 ( .A1(n3446), .A2(n4743), .B1(REG1_REG_5__SCAN_IN), .B2(n4909), .ZN(n3377) );
  OAI21_X1 U4013 ( .B1(n3379), .B2(n4909), .A(n3377), .ZN(U3523) );
  INV_X1 U4014 ( .A(n4374), .ZN(n4745) );
  AOI22_X1 U4015 ( .A1(n3446), .A2(n4745), .B1(REG0_REG_5__SCAN_IN), .B2(n4912), .ZN(n3378) );
  OAI21_X1 U4016 ( .B1(n3379), .B2(n4912), .A(n3378), .ZN(U3477) );
  INV_X1 U4017 ( .A(n4703), .ZN(n4068) );
  INV_X1 U4018 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4451) );
  NOR2_X1 U4019 ( .A1(STATE_REG_SCAN_IN), .A2(n4451), .ZN(n3500) );
  AOI21_X1 U4020 ( .B1(n4697), .B2(ADDR_REG_8__SCAN_IN), .A(n3500), .ZN(n3380)
         );
  INV_X1 U4021 ( .A(n3380), .ZN(n3384) );
  AOI211_X1 U4022 ( .C1(n3542), .C2(n3382), .A(n3381), .B(n4680), .ZN(n3383)
         );
  AOI211_X1 U4023 ( .C1(n4068), .C2(n4382), .A(n3384), .B(n3383), .ZN(n3388)
         );
  OAI211_X1 U4024 ( .C1(n3386), .C2(REG2_REG_8__SCAN_IN), .A(n4663), .B(n3385), 
        .ZN(n3387) );
  NAND2_X1 U4025 ( .A1(n3388), .A2(n3387), .ZN(U3248) );
  INV_X1 U4026 ( .A(n3389), .ZN(n3390) );
  AOI211_X1 U4027 ( .C1(n3392), .C2(n3391), .A(n3975), .B(n3390), .ZN(n3398)
         );
  INV_X1 U4028 ( .A(n3427), .ZN(n3396) );
  AOI21_X1 U4029 ( .B1(n4064), .B2(n4957), .A(n3393), .ZN(n3395) );
  AOI22_X1 U4030 ( .A1(n4062), .A2(n4948), .B1(n4960), .B2(n3409), .ZN(n3394)
         );
  OAI211_X1 U4031 ( .C1(n4966), .C2(n3396), .A(n3395), .B(n3394), .ZN(n3397)
         );
  OR2_X1 U4032 ( .A1(n3398), .A2(n3397), .ZN(U3227) );
  XNOR2_X1 U4033 ( .A(n3401), .B(n3400), .ZN(n3402) );
  XNOR2_X1 U4034 ( .A(n3399), .B(n3402), .ZN(n3407) );
  AND2_X1 U4035 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4608) );
  AOI21_X1 U4036 ( .B1(n4783), .B2(n4948), .A(n4608), .ZN(n3405) );
  AOI22_X1 U4037 ( .A1(n4063), .A2(n4957), .B1(n4960), .B2(n3403), .ZN(n3404)
         );
  OAI211_X1 U4038 ( .C1(n4966), .C2(n3442), .A(n3405), .B(n3404), .ZN(n3406)
         );
  AOI21_X1 U4039 ( .B1(n3407), .B2(n4961), .A(n3406), .ZN(n3408) );
  INV_X1 U4040 ( .A(n3408), .ZN(U3224) );
  NAND2_X1 U4041 ( .A1(n3410), .A2(n3409), .ZN(n3411) );
  NAND2_X1 U4042 ( .A1(n3411), .A2(n4908), .ZN(n3412) );
  OR2_X1 U40430 ( .A1(n3413), .A2(n3412), .ZN(n4756) );
  NOR2_X1 U4044 ( .A1(n4756), .A2(n4379), .ZN(n3426) );
  INV_X1 U4045 ( .A(n3414), .ZN(n3781) );
  XNOR2_X1 U4046 ( .A(n3415), .B(n3781), .ZN(n4755) );
  NAND2_X1 U4047 ( .A1(n4755), .A2(n4824), .ZN(n3425) );
  NAND2_X1 U4048 ( .A1(n3417), .A2(n3416), .ZN(n3418) );
  XNOR2_X1 U4049 ( .A(n3418), .B(n3781), .ZN(n3423) );
  NAND2_X1 U4050 ( .A1(n4064), .A2(n4897), .ZN(n3420) );
  NAND2_X1 U4051 ( .A1(n4062), .A2(n4274), .ZN(n3419) );
  OAI211_X1 U4052 ( .C1(n4780), .C2(n3421), .A(n3420), .B(n3419), .ZN(n3422)
         );
  AOI21_X1 U4053 ( .B1(n3423), .B2(n4891), .A(n3422), .ZN(n3424) );
  NAND2_X1 U4054 ( .A1(n3425), .A2(n3424), .ZN(n4759) );
  AOI211_X1 U4055 ( .C1(n4917), .C2(n3427), .A(n3426), .B(n4759), .ZN(n3437)
         );
  INV_X1 U4056 ( .A(n3428), .ZN(n3432) );
  NAND4_X1 U4057 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3433)
         );
  INV_X2 U4058 ( .A(n4825), .ZN(n4972) );
  NAND2_X1 U4059 ( .A1(n3434), .A2(n4379), .ZN(n3439) );
  INV_X1 U4060 ( .A(n3439), .ZN(n3435) );
  AOI22_X1 U4061 ( .A1(n4755), .A2(n4832), .B1(REG2_REG_4__SCAN_IN), .B2(n4972), .ZN(n3436) );
  OAI21_X1 U4062 ( .B1(n3437), .B2(n4972), .A(n3436), .ZN(U3286) );
  INV_X1 U4063 ( .A(n3438), .ZN(n3449) );
  NAND2_X1 U4064 ( .A1(n4251), .A2(n3439), .ZN(n4791) );
  INV_X1 U4065 ( .A(n4280), .ZN(n4921) );
  NAND2_X1 U4066 ( .A1(n3440), .A2(n4921), .ZN(n3448) );
  NOR2_X1 U4067 ( .A1(n4874), .A2(n4379), .ZN(n3441) );
  NOR2_X1 U4068 ( .A1(n3442), .A2(n4827), .ZN(n3445) );
  INV_X1 U4069 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3443) );
  NOR2_X1 U4070 ( .A1(n4825), .A2(n3443), .ZN(n3444) );
  AOI211_X1 U4071 ( .C1(n3446), .C2(n4968), .A(n3445), .B(n3444), .ZN(n3447)
         );
  OAI211_X1 U4072 ( .C1(n4972), .C2(n3449), .A(n3448), .B(n3447), .ZN(U3285)
         );
  NAND2_X1 U4073 ( .A1(n2497), .A2(n3451), .ZN(n3452) );
  XNOR2_X1 U4074 ( .A(n3450), .B(n3452), .ZN(n3459) );
  INV_X1 U4075 ( .A(n4767), .ZN(n3457) );
  NOR2_X1 U4076 ( .A1(STATE_REG_SCAN_IN), .A2(n3453), .ZN(n4618) );
  AOI21_X1 U4077 ( .B1(n4061), .B2(n4948), .A(n4618), .ZN(n3456) );
  AOI22_X1 U4078 ( .A1(n4062), .A2(n4957), .B1(n4960), .B2(n3454), .ZN(n3455)
         );
  OAI211_X1 U4079 ( .C1(n4966), .C2(n3457), .A(n3456), .B(n3455), .ZN(n3458)
         );
  AOI21_X1 U4080 ( .B1(n3459), .B2(n4961), .A(n3458), .ZN(n3460) );
  INV_X1 U4081 ( .A(n3460), .ZN(U3236) );
  NAND2_X1 U4082 ( .A1(n3462), .A2(n3461), .ZN(n3463) );
  NAND2_X1 U4083 ( .A1(n3464), .A2(n3463), .ZN(n4742) );
  INV_X1 U4084 ( .A(n4742), .ZN(n3480) );
  INV_X1 U4085 ( .A(n4832), .ZN(n3520) );
  NAND3_X1 U4086 ( .A1(n3767), .A2(n3821), .A3(n4727), .ZN(n3465) );
  NAND2_X1 U4087 ( .A1(n3466), .A2(n3465), .ZN(n3471) );
  NAND2_X1 U4088 ( .A1(n4066), .A2(n4897), .ZN(n3468) );
  NAND2_X1 U4089 ( .A1(n4064), .A2(n4274), .ZN(n3467) );
  OAI211_X1 U4090 ( .C1(n4780), .C2(n3469), .A(n3468), .B(n3467), .ZN(n3470)
         );
  AOI21_X1 U4091 ( .B1(n3471), .B2(n4891), .A(n3470), .ZN(n3473) );
  NAND2_X1 U4092 ( .A1(n4742), .A2(n4824), .ZN(n3472) );
  NAND2_X1 U4093 ( .A1(n3473), .A2(n3472), .ZN(n4741) );
  MUX2_X1 U4094 ( .A(n4741), .B(REG2_REG_2__SCAN_IN), .S(n4972), .Z(n3474) );
  INV_X1 U4095 ( .A(n3474), .ZN(n3479) );
  INV_X1 U4096 ( .A(n4730), .ZN(n3476) );
  AOI21_X1 U4097 ( .B1(n3477), .B2(n3476), .A(n3475), .ZN(n4746) );
  AOI22_X1 U4098 ( .A1(n4746), .A2(n4968), .B1(REG3_REG_2__SCAN_IN), .B2(n4917), .ZN(n3478) );
  OAI211_X1 U4099 ( .C1(n3480), .C2(n3520), .A(n3479), .B(n3478), .ZN(U3288)
         );
  OAI21_X1 U4100 ( .B1(n3481), .B2(n3484), .A(n4775), .ZN(n4768) );
  INV_X1 U4101 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3491) );
  INV_X1 U4102 ( .A(n3832), .ZN(n3806) );
  OR2_X1 U4103 ( .A1(n3806), .A2(n3836), .ZN(n3779) );
  XNOR2_X1 U4104 ( .A(n3482), .B(n3779), .ZN(n4770) );
  XNOR2_X1 U4105 ( .A(n3483), .B(n3779), .ZN(n3488) );
  OAI22_X1 U4106 ( .A1(n3485), .A2(n4268), .B1(n3484), .B2(n4780), .ZN(n3486)
         );
  AOI21_X1 U4107 ( .B1(n4274), .B2(n4061), .A(n3486), .ZN(n3487) );
  OAI21_X1 U4108 ( .B1(n3488), .B2(n4785), .A(n3487), .ZN(n3489) );
  AOI21_X1 U4109 ( .B1(n4770), .B2(n4824), .A(n3489), .ZN(n4773) );
  INV_X1 U4110 ( .A(n4773), .ZN(n3490) );
  AOI21_X1 U4111 ( .B1(n4844), .B2(n4770), .A(n3490), .ZN(n3493) );
  MUX2_X1 U4112 ( .A(n3491), .B(n3493), .S(n4911), .Z(n3492) );
  OAI21_X1 U4113 ( .B1(n4768), .B2(n4334), .A(n3492), .ZN(U3524) );
  INV_X1 U4114 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3494) );
  MUX2_X1 U4115 ( .A(n3494), .B(n3493), .S(n4915), .Z(n3495) );
  OAI21_X1 U4116 ( .B1(n4768), .B2(n4374), .A(n3495), .ZN(U3479) );
  NAND2_X1 U4117 ( .A1(n2326), .A2(n3497), .ZN(n3498) );
  XNOR2_X1 U4118 ( .A(n3499), .B(n3498), .ZN(n3506) );
  INV_X1 U4119 ( .A(n4803), .ZN(n3504) );
  AOI21_X1 U4120 ( .B1(n4061), .B2(n4957), .A(n3500), .ZN(n3503) );
  AOI22_X1 U4121 ( .A1(n4059), .A2(n4948), .B1(n4960), .B2(n3501), .ZN(n3502)
         );
  OAI211_X1 U4122 ( .C1(n4966), .C2(n3504), .A(n3503), .B(n3502), .ZN(n3505)
         );
  AOI21_X1 U4123 ( .B1(n3506), .B2(n4961), .A(n3505), .ZN(n3507) );
  INV_X1 U4124 ( .A(n3507), .ZN(U3218) );
  INV_X1 U4125 ( .A(n3841), .ZN(n3804) );
  NAND2_X1 U4126 ( .A1(n3804), .A2(n3843), .ZN(n3778) );
  XOR2_X1 U4127 ( .A(n3778), .B(n3508), .Z(n3547) );
  XNOR2_X1 U4128 ( .A(n3509), .B(n3778), .ZN(n3512) );
  AOI22_X1 U4129 ( .A1(n4058), .A2(n4274), .B1(n4896), .B2(n3523), .ZN(n3510)
         );
  OAI21_X1 U4130 ( .B1(n4781), .B2(n4268), .A(n3510), .ZN(n3511) );
  AOI21_X1 U4131 ( .B1(n3512), .B2(n4891), .A(n3511), .ZN(n3513) );
  OAI21_X1 U4132 ( .B1(n3547), .B2(n4251), .A(n3513), .ZN(n3548) );
  NAND2_X1 U4133 ( .A1(n3548), .A2(n4825), .ZN(n3519) );
  OAI21_X1 U4134 ( .B1(n3530), .B2(n3514), .A(n3622), .ZN(n3555) );
  INV_X1 U4135 ( .A(n3555), .ZN(n3517) );
  OAI22_X1 U4136 ( .A1(n3526), .A2(n4827), .B1(n3515), .B2(n4825), .ZN(n3516)
         );
  AOI21_X1 U4137 ( .B1(n3517), .B2(n4968), .A(n3516), .ZN(n3518) );
  OAI211_X1 U4138 ( .C1(n3547), .C2(n3520), .A(n3519), .B(n3518), .ZN(U3281)
         );
  XNOR2_X1 U4139 ( .A(n3522), .B(n3521), .ZN(n3528) );
  NOR2_X1 U4140 ( .A1(STATE_REG_SCAN_IN), .A2(n2837), .ZN(n4631) );
  AOI21_X1 U4141 ( .B1(n4058), .B2(n4948), .A(n4631), .ZN(n3525) );
  AOI22_X1 U4142 ( .A1(n4060), .A2(n4957), .B1(n4960), .B2(n3523), .ZN(n3524)
         );
  OAI211_X1 U4143 ( .C1(n4966), .C2(n3526), .A(n3525), .B(n3524), .ZN(n3527)
         );
  AOI21_X1 U4144 ( .B1(n3528), .B2(n4961), .A(n3527), .ZN(n3529) );
  INV_X1 U4145 ( .A(n3529), .ZN(U3228) );
  INV_X1 U4146 ( .A(n4776), .ZN(n3532) );
  INV_X1 U4147 ( .A(n3530), .ZN(n3531) );
  OAI21_X1 U4148 ( .B1(n3532), .B2(n3535), .A(n3531), .ZN(n4804) );
  NAND2_X1 U4149 ( .A1(n3842), .A2(n3802), .ZN(n3776) );
  XOR2_X1 U4150 ( .A(n3776), .B(n3533), .Z(n4806) );
  XOR2_X1 U4151 ( .A(n3776), .B(n3534), .Z(n3539) );
  OAI22_X1 U4152 ( .A1(n3536), .A2(n4268), .B1(n3535), .B2(n4780), .ZN(n3537)
         );
  AOI21_X1 U4153 ( .B1(n4274), .B2(n4059), .A(n3537), .ZN(n3538) );
  OAI21_X1 U4154 ( .B1(n3539), .B2(n4785), .A(n3538), .ZN(n3540) );
  AOI21_X1 U4155 ( .B1(n4806), .B2(n4824), .A(n3540), .ZN(n4809) );
  INV_X1 U4156 ( .A(n4809), .ZN(n3541) );
  AOI21_X1 U4157 ( .B1(n4844), .B2(n4806), .A(n3541), .ZN(n3544) );
  MUX2_X1 U4158 ( .A(n3542), .B(n3544), .S(n4911), .Z(n3543) );
  OAI21_X1 U4159 ( .B1(n4804), .B2(n4334), .A(n3543), .ZN(U3526) );
  INV_X1 U4160 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3545) );
  MUX2_X1 U4161 ( .A(n3545), .B(n3544), .S(n4915), .Z(n3546) );
  OAI21_X1 U4162 ( .B1(n4804), .B2(n4374), .A(n3546), .ZN(U3483) );
  INV_X1 U4163 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3550) );
  INV_X1 U4164 ( .A(n3547), .ZN(n3549) );
  AOI21_X1 U4165 ( .B1(n4844), .B2(n3549), .A(n3548), .ZN(n3552) );
  MUX2_X1 U4166 ( .A(n3550), .B(n3552), .S(n4911), .Z(n3551) );
  OAI21_X1 U4167 ( .B1(n4334), .B2(n3555), .A(n3551), .ZN(U3527) );
  INV_X1 U4168 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3553) );
  MUX2_X1 U4169 ( .A(n3553), .B(n3552), .S(n4915), .Z(n3554) );
  OAI21_X1 U4170 ( .B1(n3555), .B2(n4374), .A(n3554), .ZN(U3485) );
  NAND2_X1 U4171 ( .A1(n3605), .A2(n3603), .ZN(n3773) );
  XOR2_X1 U4172 ( .A(n3773), .B(n3556), .Z(n3641) );
  INV_X1 U4173 ( .A(n3641), .ZN(n3569) );
  INV_X1 U4174 ( .A(n3557), .ZN(n3558) );
  AOI21_X1 U4175 ( .B1(n3593), .B2(n3559), .A(n3558), .ZN(n3606) );
  XOR2_X1 U4176 ( .A(n3773), .B(n3606), .Z(n3563) );
  OAI22_X1 U4177 ( .A1(n3560), .A2(n4901), .B1(n4780), .B2(n4587), .ZN(n3561)
         );
  AOI21_X1 U4178 ( .B1(n4897), .B2(n4057), .A(n3561), .ZN(n3562) );
  OAI21_X1 U4179 ( .B1(n3563), .B2(n4785), .A(n3562), .ZN(n3640) );
  NOR2_X1 U4180 ( .A1(n3588), .A2(n4587), .ZN(n3564) );
  OR2_X1 U4181 ( .A1(n3616), .A2(n3564), .ZN(n3646) );
  AOI22_X1 U4182 ( .A1(n4972), .A2(REG2_REG_12__SCAN_IN), .B1(n3565), .B2(
        n4917), .ZN(n3566) );
  OAI21_X1 U4183 ( .B1(n3646), .B2(n4259), .A(n3566), .ZN(n3567) );
  AOI21_X1 U4184 ( .B1(n3640), .B2(n4825), .A(n3567), .ZN(n3568) );
  OAI21_X1 U4185 ( .B1(n3569), .B2(n4280), .A(n3568), .ZN(U3278) );
  XNOR2_X1 U4186 ( .A(n3571), .B(n3570), .ZN(n3572) );
  XNOR2_X1 U4187 ( .A(n3573), .B(n3572), .ZN(n3577) );
  AND2_X1 U4188 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4650) );
  AOI21_X1 U4189 ( .B1(n4056), .B2(n4948), .A(n4650), .ZN(n3575) );
  AOI22_X1 U4190 ( .A1(n4058), .A2(n4957), .B1(n4960), .B2(n3594), .ZN(n3574)
         );
  OAI211_X1 U4191 ( .C1(n4966), .C2(n4828), .A(n3575), .B(n3574), .ZN(n3576)
         );
  AOI21_X1 U4192 ( .B1(n3577), .B2(n4961), .A(n3576), .ZN(n3578) );
  INV_X1 U4193 ( .A(n3578), .ZN(U3233) );
  INV_X1 U4194 ( .A(n3579), .ZN(n3580) );
  AOI211_X1 U4195 ( .C1(n3582), .C2(n3581), .A(n3975), .B(n3580), .ZN(n3587)
         );
  INV_X1 U4196 ( .A(n4814), .ZN(n3585) );
  NOR2_X1 U4197 ( .A1(STATE_REG_SCAN_IN), .A2(n4486), .ZN(n4644) );
  AOI21_X1 U4198 ( .B1(n4057), .B2(n4948), .A(n4644), .ZN(n3584) );
  AOI22_X1 U4199 ( .A1(n4059), .A2(n4957), .B1(n4960), .B2(n3628), .ZN(n3583)
         );
  OAI211_X1 U4200 ( .C1(n4966), .C2(n3585), .A(n3584), .B(n3583), .ZN(n3586)
         );
  OR2_X1 U4201 ( .A1(n3587), .A2(n3586), .ZN(U3214) );
  INV_X1 U4202 ( .A(n3623), .ZN(n3591) );
  INV_X1 U4203 ( .A(n3588), .ZN(n3589) );
  OAI21_X1 U4204 ( .B1(n3591), .B2(n3590), .A(n3589), .ZN(n4830) );
  XNOR2_X1 U4205 ( .A(n3592), .B(n3777), .ZN(n4833) );
  XNOR2_X1 U4206 ( .A(n3593), .B(n3777), .ZN(n3597) );
  AOI22_X1 U4207 ( .A1(n4056), .A2(n4274), .B1(n4896), .B2(n3594), .ZN(n3596)
         );
  NAND2_X1 U4208 ( .A1(n4058), .A2(n4897), .ZN(n3595) );
  OAI211_X1 U4209 ( .C1(n3597), .C2(n4785), .A(n3596), .B(n3595), .ZN(n4823)
         );
  AOI21_X1 U4210 ( .B1(n4877), .B2(n4833), .A(n4823), .ZN(n3600) );
  INV_X1 U4211 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3598) );
  MUX2_X1 U4212 ( .A(n3600), .B(n3598), .S(n4912), .Z(n3599) );
  OAI21_X1 U4213 ( .B1(n4830), .B2(n4374), .A(n3599), .ZN(U3489) );
  MUX2_X1 U4214 ( .A(n3600), .B(n2408), .S(n4909), .Z(n3601) );
  OAI21_X1 U4215 ( .B1(n4334), .B2(n4830), .A(n3601), .ZN(U3529) );
  AND2_X1 U4216 ( .A1(n3668), .A2(n3667), .ZN(n3774) );
  XNOR2_X1 U4217 ( .A(n3602), .B(n3774), .ZN(n3614) );
  INV_X1 U4218 ( .A(n3603), .ZN(n3604) );
  AOI21_X1 U4219 ( .B1(n3606), .B2(n3605), .A(n3604), .ZN(n3608) );
  INV_X1 U4220 ( .A(n3774), .ZN(n3607) );
  XNOR2_X1 U4221 ( .A(n3608), .B(n3607), .ZN(n3612) );
  AOI22_X1 U4222 ( .A1(n4056), .A2(n4897), .B1(n3651), .B2(n4896), .ZN(n3609)
         );
  OAI21_X1 U4223 ( .B1(n3610), .B2(n4901), .A(n3609), .ZN(n3611) );
  AOI21_X1 U4224 ( .B1(n3612), .B2(n4891), .A(n3611), .ZN(n3613) );
  OAI21_X1 U4225 ( .B1(n3614), .B2(n4251), .A(n3613), .ZN(n4841) );
  INV_X1 U4226 ( .A(n4841), .ZN(n3621) );
  INV_X1 U4227 ( .A(n3614), .ZN(n4843) );
  OAI21_X1 U4228 ( .B1(n3616), .B2(n3615), .A(n3675), .ZN(n4840) );
  AOI22_X1 U4229 ( .A1(n4972), .A2(REG2_REG_13__SCAN_IN), .B1(n3617), .B2(
        n4917), .ZN(n3618) );
  OAI21_X1 U4230 ( .B1(n4840), .B2(n4259), .A(n3618), .ZN(n3619) );
  AOI21_X1 U4231 ( .B1(n4843), .B2(n4832), .A(n3619), .ZN(n3620) );
  OAI21_X1 U4232 ( .B1(n3621), .B2(n4972), .A(n3620), .ZN(U3277) );
  INV_X1 U4233 ( .A(n3622), .ZN(n3625) );
  OAI21_X1 U4234 ( .B1(n3625), .B2(n3624), .A(n3623), .ZN(n4815) );
  INV_X1 U4235 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3635) );
  NAND2_X1 U4236 ( .A1(n3807), .A2(n3808), .ZN(n3771) );
  XNOR2_X1 U4237 ( .A(n3626), .B(n3771), .ZN(n3630) );
  INV_X1 U4238 ( .A(n3630), .ZN(n4817) );
  XOR2_X1 U4239 ( .A(n3771), .B(n3627), .Z(n3633) );
  AOI22_X1 U4240 ( .A1(n4059), .A2(n4897), .B1(n3628), .B2(n4896), .ZN(n3629)
         );
  OAI21_X1 U4241 ( .B1(n4589), .B2(n4901), .A(n3629), .ZN(n3632) );
  NOR2_X1 U4242 ( .A1(n3630), .A2(n4251), .ZN(n3631) );
  AOI211_X1 U4243 ( .C1(n3633), .C2(n4891), .A(n3632), .B(n3631), .ZN(n4820)
         );
  INV_X1 U4244 ( .A(n4820), .ZN(n3634) );
  AOI21_X1 U4245 ( .B1(n4844), .B2(n4817), .A(n3634), .ZN(n3637) );
  MUX2_X1 U4246 ( .A(n3635), .B(n3637), .S(n4911), .Z(n3636) );
  OAI21_X1 U4247 ( .B1(n4815), .B2(n4334), .A(n3636), .ZN(U3528) );
  INV_X1 U4248 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3638) );
  MUX2_X1 U4249 ( .A(n3638), .B(n3637), .S(n4915), .Z(n3639) );
  OAI21_X1 U4250 ( .B1(n4815), .B2(n4374), .A(n3639), .ZN(U3487) );
  AOI21_X1 U4251 ( .B1(n3641), .B2(n4877), .A(n3640), .ZN(n3643) );
  MUX2_X1 U4252 ( .A(n4659), .B(n3643), .S(n4911), .Z(n3642) );
  OAI21_X1 U4253 ( .B1(n3646), .B2(n4334), .A(n3642), .ZN(U3530) );
  INV_X1 U4254 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3644) );
  MUX2_X1 U4255 ( .A(n3644), .B(n3643), .S(n4915), .Z(n3645) );
  OAI21_X1 U4256 ( .B1(n3646), .B2(n4374), .A(n3645), .ZN(U3491) );
  XNOR2_X1 U4257 ( .A(n3648), .B(n3647), .ZN(n3649) );
  XNOR2_X1 U4258 ( .A(n3650), .B(n3649), .ZN(n3656) );
  INV_X1 U4259 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4565) );
  NOR2_X1 U4260 ( .A1(STATE_REG_SCAN_IN), .A2(n4565), .ZN(n4677) );
  AOI21_X1 U4261 ( .B1(n4056), .B2(n4957), .A(n4677), .ZN(n3653) );
  AOI22_X1 U4262 ( .A1(n4862), .A2(n4948), .B1(n4960), .B2(n3651), .ZN(n3652)
         );
  OAI211_X1 U4263 ( .C1(n4966), .C2(n3654), .A(n3653), .B(n3652), .ZN(n3655)
         );
  AOI21_X1 U4264 ( .B1(n3656), .B2(n4961), .A(n3655), .ZN(n3657) );
  INV_X1 U4265 ( .A(n3657), .ZN(U3231) );
  INV_X1 U4266 ( .A(n4055), .ZN(n4859) );
  OAI22_X1 U4267 ( .A1(n4859), .A2(n4901), .B1(n4857), .B2(n4780), .ZN(n3662)
         );
  INV_X1 U4268 ( .A(n3658), .ZN(n3659) );
  AOI211_X1 U4269 ( .C1(n3660), .C2(n3788), .A(n4785), .B(n3659), .ZN(n3661)
         );
  AOI211_X1 U4270 ( .C1(n4897), .C2(n4862), .A(n3662), .B(n3661), .ZN(n4872)
         );
  INV_X1 U4271 ( .A(n3676), .ZN(n3663) );
  OAI21_X1 U4272 ( .B1(n3663), .B2(n4857), .A(n4890), .ZN(n4873) );
  INV_X1 U4273 ( .A(n4873), .ZN(n3666) );
  INV_X1 U4274 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3664) );
  OAI22_X1 U4275 ( .A1(n4825), .A2(n3664), .B1(n4871), .B2(n4827), .ZN(n3665)
         );
  AOI21_X1 U4276 ( .B1(n3666), .B2(n4968), .A(n3665), .ZN(n3674) );
  INV_X1 U4277 ( .A(n3667), .ZN(n3669) );
  OAI21_X1 U4278 ( .B1(n3602), .B2(n3669), .A(n3668), .ZN(n3680) );
  NAND2_X1 U4279 ( .A1(n3680), .A2(n3679), .ZN(n3678) );
  INV_X1 U4280 ( .A(n3670), .ZN(n3671) );
  NAND2_X1 U4281 ( .A1(n3678), .A2(n3671), .ZN(n3672) );
  XNOR2_X1 U4282 ( .A(n3672), .B(n3788), .ZN(n4876) );
  NAND2_X1 U4283 ( .A1(n4876), .A2(n4921), .ZN(n3673) );
  OAI211_X1 U4284 ( .C1(n4872), .C2(n4972), .A(n3674), .B(n3673), .ZN(U3275)
         );
  INV_X1 U4285 ( .A(n3675), .ZN(n3677) );
  OAI21_X1 U4286 ( .B1(n3677), .B2(n3683), .A(n3676), .ZN(n4851) );
  INV_X1 U4287 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3687) );
  OAI21_X1 U4288 ( .B1(n3680), .B2(n3679), .A(n3678), .ZN(n4853) );
  XNOR2_X1 U4289 ( .A(n3725), .B(n3780), .ZN(n3685) );
  NAND2_X1 U4290 ( .A1(n4898), .A2(n4274), .ZN(n3682) );
  NAND2_X1 U4291 ( .A1(n4591), .A2(n4897), .ZN(n3681) );
  OAI211_X1 U4292 ( .C1(n4780), .C2(n3683), .A(n3682), .B(n3681), .ZN(n3684)
         );
  AOI21_X1 U4293 ( .B1(n3685), .B2(n4891), .A(n3684), .ZN(n4856) );
  INV_X1 U4294 ( .A(n4856), .ZN(n3686) );
  AOI21_X1 U4295 ( .B1(n4853), .B2(n4877), .A(n3686), .ZN(n3689) );
  MUX2_X1 U4296 ( .A(n3687), .B(n3689), .S(n4915), .Z(n3688) );
  OAI21_X1 U4297 ( .B1(n4851), .B2(n4374), .A(n3688), .ZN(U3495) );
  INV_X1 U4298 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3690) );
  MUX2_X1 U4299 ( .A(n3690), .B(n3689), .S(n4911), .Z(n3691) );
  OAI21_X1 U4300 ( .B1(n4851), .B2(n4334), .A(n3691), .ZN(U3532) );
  NAND2_X1 U4301 ( .A1(n2303), .A2(n3693), .ZN(n3694) );
  XNOR2_X1 U4302 ( .A(n3692), .B(n3694), .ZN(n3700) );
  INV_X1 U4303 ( .A(n4850), .ZN(n3698) );
  NOR2_X1 U4304 ( .A1(n4536), .A2(STATE_REG_SCAN_IN), .ZN(n4684) );
  AOI21_X1 U4305 ( .B1(n4591), .B2(n4957), .A(n4684), .ZN(n3697) );
  AOI22_X1 U4306 ( .A1(n4898), .A2(n4948), .B1(n4960), .B2(n3695), .ZN(n3696)
         );
  OAI211_X1 U4307 ( .C1(n4966), .C2(n3698), .A(n3697), .B(n3696), .ZN(n3699)
         );
  AOI21_X1 U4308 ( .B1(n3700), .B2(n4961), .A(n3699), .ZN(n3701) );
  INV_X1 U4309 ( .A(n3701), .ZN(U3212) );
  NAND2_X1 U4310 ( .A1(n3895), .A2(n3894), .ZN(n3772) );
  XOR2_X1 U4311 ( .A(n3772), .B(n3702), .Z(n3713) );
  INV_X1 U4312 ( .A(n3713), .ZN(n3711) );
  XOR2_X1 U4313 ( .A(n3772), .B(n3897), .Z(n3705) );
  OAI22_X1 U4314 ( .A1(n3903), .A2(n4901), .B1(n3706), .B2(n4780), .ZN(n3703)
         );
  AOI21_X1 U4315 ( .B1(n4897), .B2(n4055), .A(n3703), .ZN(n3704) );
  OAI21_X1 U4316 ( .B1(n3705), .B2(n4785), .A(n3704), .ZN(n3712) );
  OAI21_X1 U4317 ( .B1(n4889), .B2(n3706), .A(n4264), .ZN(n3718) );
  NOR2_X1 U4318 ( .A1(n3718), .A2(n4259), .ZN(n3709) );
  INV_X1 U4319 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3707) );
  OAI22_X1 U4320 ( .A1(n4825), .A2(n3707), .B1(n4004), .B2(n4827), .ZN(n3708)
         );
  AOI211_X1 U4321 ( .C1(n3712), .C2(n4825), .A(n3709), .B(n3708), .ZN(n3710)
         );
  OAI21_X1 U4322 ( .B1(n3711), .B2(n4280), .A(n3710), .ZN(U3273) );
  AOI21_X1 U4323 ( .B1(n3713), .B2(n4877), .A(n3712), .ZN(n3715) );
  MUX2_X1 U4324 ( .A(n2620), .B(n3715), .S(n4911), .Z(n3714) );
  OAI21_X1 U4325 ( .B1(n4334), .B2(n3718), .A(n3714), .ZN(U3535) );
  INV_X1 U4326 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3716) );
  MUX2_X1 U4327 ( .A(n3716), .B(n3715), .S(n4915), .Z(n3717) );
  OAI21_X1 U4328 ( .B1(n3718), .B2(n4374), .A(n3717), .ZN(U3501) );
  NOR2_X1 U4329 ( .A1(n3738), .A2(n3719), .ZN(n4289) );
  NAND2_X1 U4330 ( .A1(n3720), .A2(n3723), .ZN(n3812) );
  AND2_X1 U4331 ( .A1(n3722), .A2(n3721), .ZN(n3844) );
  INV_X1 U4332 ( .A(n3844), .ZN(n3724) );
  NAND2_X1 U4333 ( .A1(n3724), .A2(n3723), .ZN(n3816) );
  OAI21_X1 U4334 ( .B1(n3725), .B2(n3812), .A(n3816), .ZN(n3727) );
  INV_X1 U4335 ( .A(n3854), .ZN(n3726) );
  INV_X1 U4336 ( .A(n3851), .ZN(n3785) );
  AOI211_X1 U4337 ( .C1(n3727), .C2(n3726), .A(n3848), .B(n3785), .ZN(n3731)
         );
  INV_X1 U4338 ( .A(n3728), .ZN(n3729) );
  OAI21_X1 U4339 ( .B1(n3729), .B2(n3784), .A(n3851), .ZN(n3856) );
  INV_X1 U4340 ( .A(n3856), .ZN(n3730) );
  AOI211_X1 U4341 ( .C1(n3852), .C2(n3731), .A(n3730), .B(n3858), .ZN(n3736)
         );
  INV_X1 U4342 ( .A(n3732), .ZN(n3735) );
  INV_X1 U4343 ( .A(n3733), .ZN(n3734) );
  NOR2_X1 U4344 ( .A1(n3734), .A2(n3766), .ZN(n3860) );
  OAI21_X1 U4345 ( .B1(n3736), .B2(n3735), .A(n3860), .ZN(n3743) );
  INV_X1 U4346 ( .A(n4125), .ZN(n4053) );
  INV_X1 U4347 ( .A(DATAI_31_), .ZN(n3737) );
  NOR2_X1 U4348 ( .A1(n3738), .A2(n3737), .ZN(n4115) );
  OR2_X1 U4349 ( .A1(n4114), .A2(n4115), .ZN(n3874) );
  NAND2_X1 U4350 ( .A1(n3753), .A2(n4289), .ZN(n3739) );
  AND2_X1 U4351 ( .A1(n3874), .A2(n3739), .ZN(n3759) );
  OAI21_X1 U4352 ( .B1(n4053), .B2(n3740), .A(n3759), .ZN(n3748) );
  NAND2_X1 U4353 ( .A1(n3742), .A2(n3741), .ZN(n3749) );
  AOI211_X1 U4354 ( .C1(n3863), .C2(n3743), .A(n3748), .B(n3749), .ZN(n3751)
         );
  INV_X1 U4355 ( .A(n3744), .ZN(n3865) );
  OR2_X1 U4356 ( .A1(n4125), .A2(n3745), .ZN(n3747) );
  AND2_X1 U4357 ( .A1(n3747), .A2(n3746), .ZN(n3868) );
  AOI21_X1 U4358 ( .B1(n3749), .B2(n3868), .A(n3748), .ZN(n3877) );
  NAND3_X1 U4359 ( .A1(n3761), .A2(n3868), .A3(n3867), .ZN(n3750) );
  AOI22_X1 U4360 ( .A1(n3751), .A2(n3865), .B1(n3877), .B2(n3750), .ZN(n3752)
         );
  AOI21_X1 U4361 ( .B1(n4114), .B2(n4289), .A(n3752), .ZN(n3758) );
  OR2_X1 U4362 ( .A1(n3753), .A2(n4289), .ZN(n3755) );
  NAND2_X1 U4363 ( .A1(n4114), .A2(n4115), .ZN(n3754) );
  NAND2_X1 U4364 ( .A1(n3755), .A2(n3754), .ZN(n3875) );
  INV_X1 U4365 ( .A(n3875), .ZN(n3760) );
  INV_X1 U4366 ( .A(n4115), .ZN(n4112) );
  NOR2_X1 U4367 ( .A1(n3760), .A2(n4112), .ZN(n3757) );
  NOR3_X1 U4368 ( .A1(n3758), .A2(n3757), .A3(n3756), .ZN(n3883) );
  XNOR2_X1 U4369 ( .A(n4944), .B(n3908), .ZN(n3902) );
  NAND4_X1 U4370 ( .A1(n3761), .A2(n4123), .A3(n3760), .A4(n3759), .ZN(n3762)
         );
  NOR3_X1 U4371 ( .A1(n4269), .A2(n3902), .A3(n3762), .ZN(n3799) );
  NAND2_X1 U4372 ( .A1(n3763), .A2(n3867), .ZN(n4153) );
  INV_X1 U4373 ( .A(n4153), .ZN(n3797) );
  XNOR2_X1 U4374 ( .A(n4232), .B(n4221), .ZN(n4212) );
  INV_X1 U4375 ( .A(n4725), .ZN(n3770) );
  INV_X1 U4376 ( .A(n3855), .ZN(n4209) );
  NAND2_X1 U4377 ( .A1(n4209), .A2(n4207), .ZN(n3922) );
  INV_X1 U4378 ( .A(n3922), .ZN(n3769) );
  NAND2_X1 U4379 ( .A1(n4151), .A2(n3764), .ZN(n4171) );
  INV_X1 U4380 ( .A(n3765), .ZN(n4169) );
  OR2_X1 U4381 ( .A1(n4169), .A2(n3766), .ZN(n4186) );
  NOR4_X1 U4382 ( .A1(n3767), .A2(n4230), .A3(n4171), .A4(n4186), .ZN(n3768)
         );
  NAND3_X1 U4383 ( .A1(n3770), .A2(n3769), .A3(n3768), .ZN(n3794) );
  NOR4_X1 U4384 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3792)
         );
  NOR4_X1 U4385 ( .A1(n3777), .A2(n4789), .A3(n3776), .A4(n3775), .ZN(n3791)
         );
  INV_X1 U4386 ( .A(n3778), .ZN(n3783) );
  INV_X1 U4387 ( .A(n3779), .ZN(n3782) );
  AND4_X1 U4388 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3790)
         );
  OR2_X1 U4389 ( .A1(n3785), .A2(n3784), .ZN(n4327) );
  NOR2_X1 U4390 ( .A1(n3786), .A2(n4732), .ZN(n3819) );
  INV_X1 U4391 ( .A(n3819), .ZN(n3787) );
  NAND2_X1 U4392 ( .A1(n3787), .A2(n4724), .ZN(n4714) );
  NOR4_X1 U4393 ( .A1(n4905), .A2(n3788), .A3(n4327), .A4(n4714), .ZN(n3789)
         );
  NAND4_X1 U4394 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3793)
         );
  NOR4_X1 U4395 ( .A1(n3795), .A2(n4212), .A3(n3794), .A4(n3793), .ZN(n3796)
         );
  NAND4_X1 U4396 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3801)
         );
  NOR3_X1 U4397 ( .A1(n3801), .A2(n3800), .A3(n2687), .ZN(n3882) );
  NAND3_X1 U4398 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3838) );
  NOR3_X1 U4399 ( .A1(n3838), .A2(n3806), .A3(n3805), .ZN(n3811) );
  INV_X1 U4400 ( .A(n3807), .ZN(n3810) );
  AND2_X1 U4401 ( .A1(n3809), .A2(n3808), .ZN(n3845) );
  OAI21_X1 U4402 ( .B1(n3811), .B2(n3810), .A(n3845), .ZN(n3815) );
  INV_X1 U4403 ( .A(n3812), .ZN(n3814) );
  NAND3_X1 U4404 ( .A1(n3815), .A2(n3814), .A3(n3813), .ZN(n3817) );
  NAND2_X1 U4405 ( .A1(n3817), .A2(n3816), .ZN(n3850) );
  OAI21_X1 U4406 ( .B1(n3819), .B2(n3818), .A(n4724), .ZN(n3825) );
  INV_X1 U4407 ( .A(n3820), .ZN(n3823) );
  INV_X1 U4408 ( .A(n3821), .ZN(n3822) );
  AOI211_X1 U4409 ( .C1(n3825), .C2(n3824), .A(n3823), .B(n3822), .ZN(n3830)
         );
  NAND2_X1 U4410 ( .A1(n3827), .A2(n3826), .ZN(n3829) );
  OAI21_X1 U4411 ( .B1(n3830), .B2(n3829), .A(n3828), .ZN(n3834) );
  NAND4_X1 U4412 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3840)
         );
  INV_X1 U4413 ( .A(n3835), .ZN(n3837) );
  NOR2_X1 U4414 ( .A1(n3837), .A2(n3836), .ZN(n3839) );
  AOI21_X1 U4415 ( .B1(n3840), .B2(n3839), .A(n3838), .ZN(n3847) );
  AOI21_X1 U4416 ( .B1(n3843), .B2(n3842), .A(n3841), .ZN(n3846) );
  OAI211_X1 U4417 ( .C1(n3847), .C2(n3846), .A(n3845), .B(n3844), .ZN(n3849)
         );
  AOI21_X1 U4418 ( .B1(n3850), .B2(n3849), .A(n3848), .ZN(n3853) );
  OAI211_X1 U4419 ( .C1(n3854), .C2(n3853), .A(n3852), .B(n3851), .ZN(n3857)
         );
  AOI21_X1 U4420 ( .B1(n3857), .B2(n3856), .A(n3855), .ZN(n3859) );
  NOR2_X1 U4421 ( .A1(n3859), .A2(n3858), .ZN(n3862) );
  OAI21_X1 U4422 ( .B1(n3862), .B2(n3861), .A(n3860), .ZN(n3864) );
  NAND2_X1 U4423 ( .A1(n3864), .A2(n3863), .ZN(n3866) );
  NAND2_X1 U4424 ( .A1(n3866), .A2(n3865), .ZN(n3873) );
  INV_X1 U4425 ( .A(n3867), .ZN(n3870) );
  INV_X1 U4426 ( .A(n3868), .ZN(n3869) );
  NOR4_X1 U4427 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3875), .ZN(n3872)
         );
  NAND2_X1 U4428 ( .A1(n3873), .A2(n3872), .ZN(n3880) );
  AND2_X1 U4429 ( .A1(n3875), .A2(n3874), .ZN(n3876) );
  OR2_X1 U4430 ( .A1(n3877), .A2(n3876), .ZN(n3879) );
  AOI21_X1 U4431 ( .B1(n3880), .B2(n3879), .A(n3878), .ZN(n3881) );
  NOR3_X1 U4432 ( .A1(n3883), .A2(n3882), .A3(n3881), .ZN(n3884) );
  INV_X1 U4433 ( .A(n3884), .ZN(n3885) );
  MUX2_X1 U4434 ( .A(n3885), .B(n3884), .S(n4787), .Z(n3892) );
  NOR4_X1 U4435 ( .A1(n2767), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n3891)
         );
  OAI21_X1 U4436 ( .B1(n4388), .B2(n3889), .A(B_REG_SCAN_IN), .ZN(n3890) );
  OAI22_X1 U4437 ( .A1(n3892), .A2(n4388), .B1(n3891), .B2(n3890), .ZN(U3239)
         );
  XNOR2_X1 U4438 ( .A(n3893), .B(n3902), .ZN(n3915) );
  INV_X1 U4439 ( .A(n3915), .ZN(n3913) );
  INV_X1 U4440 ( .A(n3894), .ZN(n3896) );
  OAI21_X1 U4441 ( .B1(n3897), .B2(n3896), .A(n3895), .ZN(n4270) );
  INV_X1 U4442 ( .A(n3898), .ZN(n3900) );
  OAI21_X1 U4443 ( .B1(n4270), .B2(n3900), .A(n3899), .ZN(n3901) );
  XOR2_X1 U4444 ( .A(n3902), .B(n3901), .Z(n3906) );
  OAI22_X1 U4445 ( .A1(n3903), .A2(n4268), .B1(n3908), .B2(n4780), .ZN(n3904)
         );
  AOI21_X1 U4446 ( .B1(n4274), .B2(n4958), .A(n3904), .ZN(n3905) );
  OAI21_X1 U4447 ( .B1(n3906), .B2(n4785), .A(n3905), .ZN(n3914) );
  INV_X1 U4448 ( .A(n4265), .ZN(n3909) );
  INV_X1 U4449 ( .A(n4254), .ZN(n3907) );
  OAI21_X1 U4450 ( .B1(n3909), .B2(n3908), .A(n3907), .ZN(n3920) );
  NOR2_X1 U4451 ( .A1(n3920), .A2(n4259), .ZN(n3911) );
  OAI22_X1 U4452 ( .A1(n4825), .A2(n2659), .B1(n4938), .B2(n4827), .ZN(n3910)
         );
  AOI211_X1 U4453 ( .C1(n3914), .C2(n4825), .A(n3911), .B(n3910), .ZN(n3912)
         );
  OAI21_X1 U4454 ( .B1(n3913), .B2(n4280), .A(n3912), .ZN(U3271) );
  INV_X1 U4455 ( .A(REG0_REG_19__SCAN_IN), .ZN(n3916) );
  AOI21_X1 U4456 ( .B1(n4877), .B2(n3915), .A(n3914), .ZN(n3918) );
  MUX2_X1 U4457 ( .A(n3916), .B(n3918), .S(n4915), .Z(n3917) );
  OAI21_X1 U4458 ( .B1(n3920), .B2(n4374), .A(n3917), .ZN(U3505) );
  MUX2_X1 U4459 ( .A(n2623), .B(n3918), .S(n4911), .Z(n3919) );
  OAI21_X1 U4460 ( .B1(n4334), .B2(n3920), .A(n3919), .ZN(U3537) );
  XNOR2_X1 U4461 ( .A(n3921), .B(n3922), .ZN(n4324) );
  INV_X1 U4462 ( .A(n4324), .ZN(n3932) );
  XNOR2_X1 U4463 ( .A(n4210), .B(n3922), .ZN(n3925) );
  OAI22_X1 U4464 ( .A1(n4214), .A2(n4901), .B1(n4780), .B2(n3926), .ZN(n3923)
         );
  AOI21_X1 U4465 ( .B1(n4897), .B2(n4958), .A(n3923), .ZN(n3924) );
  OAI21_X1 U4466 ( .B1(n3925), .B2(n4785), .A(n3924), .ZN(n4323) );
  OR2_X1 U4467 ( .A1(n4256), .A2(n3926), .ZN(n3927) );
  NAND2_X1 U4468 ( .A1(n2266), .A2(n3927), .ZN(n4370) );
  AOI22_X1 U4469 ( .A1(n4972), .A2(REG2_REG_21__SCAN_IN), .B1(n3928), .B2(
        n4917), .ZN(n3929) );
  OAI21_X1 U4470 ( .B1(n4370), .B2(n4259), .A(n3929), .ZN(n3930) );
  AOI21_X1 U4471 ( .B1(n4323), .B2(n4825), .A(n3930), .ZN(n3931) );
  OAI21_X1 U4472 ( .B1(n3932), .B2(n4280), .A(n3931), .ZN(U3269) );
  AND2_X1 U4473 ( .A1(n3933), .A2(n4067), .ZN(U3148) );
  NAND2_X1 U4474 ( .A1(n4068), .A2(n4386), .ZN(n3945) );
  OAI211_X1 U4475 ( .C1(n3936), .C2(n3935), .A(n4663), .B(n3934), .ZN(n3944)
         );
  AOI22_X1 U4476 ( .A1(n4697), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3943) );
  INV_X1 U4477 ( .A(n3937), .ZN(n3941) );
  NAND3_X1 U4478 ( .A1(n3939), .A2(n4069), .A3(n3938), .ZN(n3940) );
  NAND3_X1 U4479 ( .A1(n4698), .A2(n3941), .A3(n3940), .ZN(n3942) );
  NAND4_X1 U4480 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3946)
         );
  OR2_X1 U4481 ( .A1(n3947), .A2(n3946), .ZN(U3242) );
  XNOR2_X1 U4482 ( .A(n3949), .B(n3948), .ZN(n3954) );
  INV_X1 U4483 ( .A(n4141), .ZN(n3952) );
  AOI22_X1 U4484 ( .A1(n4137), .A2(n4948), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3951) );
  AOI22_X1 U4485 ( .A1(n4175), .A2(n4957), .B1(n4960), .B2(n4136), .ZN(n3950)
         );
  OAI211_X1 U4486 ( .C1(n4966), .C2(n3952), .A(n3951), .B(n3950), .ZN(n3953)
         );
  AOI21_X1 U4487 ( .B1(n3954), .B2(n4961), .A(n3953), .ZN(n3955) );
  INV_X1 U4488 ( .A(n3955), .ZN(U3211) );
  NAND3_X1 U4489 ( .A1(n3956), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3957) );
  OAI22_X1 U4490 ( .A1(n2671), .A2(n3957), .B1(STATE_REG_SCAN_IN), .B2(n3737), 
        .ZN(U3321) );
  INV_X1 U4491 ( .A(n3958), .ZN(n3960) );
  OAI211_X1 U4492 ( .C1(n3965), .C2(n3964), .A(n3963), .B(n4961), .ZN(n3970)
         );
  AOI21_X1 U4493 ( .B1(n4783), .B2(n4957), .A(n3966), .ZN(n3969) );
  AOI22_X1 U4494 ( .A1(n4060), .A2(n4948), .B1(n4960), .B2(n4774), .ZN(n3968)
         );
  OR2_X1 U4495 ( .A1(n4966), .A2(n4796), .ZN(n3967) );
  NAND4_X1 U4496 ( .A1(n3970), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(U3210)
         );
  AOI22_X1 U4497 ( .A1(n4216), .A2(n4948), .B1(n4960), .B2(n3971), .ZN(n3973)
         );
  NAND2_X1 U4498 ( .A1(U3149), .A2(REG3_REG_23__SCAN_IN), .ZN(n3972) );
  OAI211_X1 U4499 ( .C1(n4214), .C2(n4588), .A(n3973), .B(n3972), .ZN(n3979)
         );
  AOI211_X1 U4500 ( .C1(n3977), .C2(n3976), .A(n3975), .B(n3974), .ZN(n3978)
         );
  AOI211_X1 U4501 ( .C1(n4222), .C2(n4026), .A(n3979), .B(n3978), .ZN(n3980)
         );
  INV_X1 U4502 ( .A(n3980), .ZN(U3213) );
  INV_X1 U4503 ( .A(n3981), .ZN(n3982) );
  NOR2_X1 U4504 ( .A1(n3983), .A2(n3982), .ZN(n3991) );
  NAND2_X1 U4505 ( .A1(n3985), .A2(n3984), .ZN(n4009) );
  NAND2_X1 U4506 ( .A1(n4009), .A2(n3986), .ZN(n3989) );
  NAND2_X1 U4507 ( .A1(n3988), .A2(n3987), .ZN(n4008) );
  INV_X1 U4508 ( .A(n3992), .ZN(n4179) );
  AOI22_X1 U4509 ( .A1(n4216), .A2(n4957), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3995) );
  AOI22_X1 U4510 ( .A1(n4175), .A2(n4948), .B1(n4960), .B2(n3993), .ZN(n3994)
         );
  OAI211_X1 U4511 ( .C1(n4966), .C2(n4179), .A(n3995), .B(n3994), .ZN(n3996)
         );
  XNOR2_X1 U4512 ( .A(n3998), .B(n3997), .ZN(n3999) );
  XNOR2_X1 U4513 ( .A(n4000), .B(n3999), .ZN(n4006) );
  INV_X1 U4514 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4555) );
  NOR2_X1 U4515 ( .A1(STATE_REG_SCAN_IN), .A2(n4555), .ZN(n4098) );
  AOI21_X1 U4516 ( .B1(n4055), .B2(n4957), .A(n4098), .ZN(n4003) );
  AOI22_X1 U4517 ( .A1(n4927), .A2(n4948), .B1(n4960), .B2(n4001), .ZN(n4002)
         );
  OAI211_X1 U4518 ( .C1(n4966), .C2(n4004), .A(n4003), .B(n4002), .ZN(n4005)
         );
  AOI21_X1 U4519 ( .B1(n4006), .B2(n4961), .A(n4005), .ZN(n4007) );
  INV_X1 U4520 ( .A(n4007), .ZN(U3225) );
  NAND2_X1 U4521 ( .A1(n4009), .A2(n4008), .ZN(n4011) );
  XNOR2_X1 U4522 ( .A(n4011), .B(n4010), .ZN(n4017) );
  INV_X1 U4523 ( .A(n4196), .ZN(n4015) );
  AOI22_X1 U4524 ( .A1(n4232), .A2(n4957), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n4014) );
  AOI22_X1 U4525 ( .A1(n4190), .A2(n4948), .B1(n4960), .B2(n4012), .ZN(n4013)
         );
  OAI211_X1 U4526 ( .C1(n4966), .C2(n4015), .A(n4014), .B(n4013), .ZN(n4016)
         );
  AOI21_X1 U4527 ( .B1(n4017), .B2(n4961), .A(n4016), .ZN(n4018) );
  INV_X1 U4528 ( .A(n4018), .ZN(U3226) );
  OAI21_X1 U4529 ( .B1(n4021), .B2(n4020), .A(n4019), .ZN(n4022) );
  NAND2_X1 U4530 ( .A1(n4022), .A2(n4961), .ZN(n4028) );
  OAI22_X1 U4531 ( .A1(n4245), .A2(n4588), .B1(STATE_REG_SCAN_IN), .B2(n4023), 
        .ZN(n4025) );
  OAI22_X1 U4532 ( .A1(n4188), .A2(n4931), .B1(n4858), .B2(n4235), .ZN(n4024)
         );
  AOI211_X1 U4533 ( .C1(n4238), .C2(n4026), .A(n4025), .B(n4024), .ZN(n4027)
         );
  NAND2_X1 U4534 ( .A1(n4028), .A2(n4027), .ZN(U3232) );
  INV_X1 U4535 ( .A(n4029), .ZN(n4031) );
  NAND2_X1 U4536 ( .A1(n4031), .A2(n4030), .ZN(n4032) );
  XNOR2_X1 U4537 ( .A(n4033), .B(n4032), .ZN(n4040) );
  INV_X1 U4538 ( .A(n4034), .ZN(n4275) );
  NOR2_X1 U4539 ( .A1(STATE_REG_SCAN_IN), .A2(n4035), .ZN(n4105) );
  AOI21_X1 U4540 ( .B1(n4054), .B2(n4957), .A(n4105), .ZN(n4038) );
  AOI22_X1 U4541 ( .A1(n4944), .A2(n4948), .B1(n4960), .B2(n4036), .ZN(n4037)
         );
  OAI211_X1 U4542 ( .C1(n4966), .C2(n4275), .A(n4038), .B(n4037), .ZN(n4039)
         );
  AOI21_X1 U4543 ( .B1(n4040), .B2(n4961), .A(n4039), .ZN(n4041) );
  INV_X1 U4544 ( .A(n4041), .ZN(U3235) );
  NAND2_X1 U4545 ( .A1(n2297), .A2(n4042), .ZN(n4043) );
  XNOR2_X1 U4546 ( .A(n4044), .B(n4043), .ZN(n4051) );
  NOR2_X1 U4547 ( .A1(n4045), .A2(STATE_REG_SCAN_IN), .ZN(n4046) );
  AOI21_X1 U4548 ( .B1(n4156), .B2(n4948), .A(n4046), .ZN(n4048) );
  AOI22_X1 U4549 ( .A1(n4190), .A2(n4957), .B1(n4960), .B2(n4160), .ZN(n4047)
         );
  OAI211_X1 U4550 ( .C1(n4966), .C2(n4049), .A(n4048), .B(n4047), .ZN(n4050)
         );
  AOI21_X1 U4551 ( .B1(n4051), .B2(n4961), .A(n4050), .ZN(n4052) );
  INV_X1 U4552 ( .A(n4052), .ZN(U3237) );
  MUX2_X1 U4553 ( .A(DATAO_REG_29__SCAN_IN), .B(n4053), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4554 ( .A(n4137), .B(DATAO_REG_28__SCAN_IN), .S(n4067), .Z(U3578)
         );
  MUX2_X1 U4555 ( .A(n4156), .B(DATAO_REG_27__SCAN_IN), .S(n4067), .Z(U3577)
         );
  MUX2_X1 U4556 ( .A(n4175), .B(DATAO_REG_26__SCAN_IN), .S(n4067), .Z(U3576)
         );
  MUX2_X1 U4557 ( .A(n4190), .B(DATAO_REG_25__SCAN_IN), .S(n4067), .Z(U3575)
         );
  MUX2_X1 U4558 ( .A(n4216), .B(DATAO_REG_24__SCAN_IN), .S(n4067), .Z(U3574)
         );
  MUX2_X1 U4559 ( .A(n4232), .B(DATAO_REG_23__SCAN_IN), .S(n4067), .Z(U3573)
         );
  INV_X1 U4560 ( .A(n4214), .ZN(n4949) );
  MUX2_X1 U4561 ( .A(DATAO_REG_22__SCAN_IN), .B(n4949), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4562 ( .A(n4939), .B(DATAO_REG_21__SCAN_IN), .S(n4067), .Z(U3571)
         );
  MUX2_X1 U4563 ( .A(n4958), .B(DATAO_REG_20__SCAN_IN), .S(n4067), .Z(U3570)
         );
  MUX2_X1 U4564 ( .A(n4944), .B(DATAO_REG_19__SCAN_IN), .S(n4067), .Z(U3569)
         );
  MUX2_X1 U4565 ( .A(n4927), .B(DATAO_REG_18__SCAN_IN), .S(n4067), .Z(U3568)
         );
  MUX2_X1 U4566 ( .A(n4054), .B(DATAO_REG_17__SCAN_IN), .S(n4067), .Z(U3567)
         );
  MUX2_X1 U4567 ( .A(n4055), .B(DATAO_REG_16__SCAN_IN), .S(n4067), .Z(U3566)
         );
  MUX2_X1 U4568 ( .A(n4898), .B(DATAO_REG_15__SCAN_IN), .S(n4067), .Z(U3565)
         );
  MUX2_X1 U4569 ( .A(n4862), .B(DATAO_REG_14__SCAN_IN), .S(n4067), .Z(U3564)
         );
  MUX2_X1 U4570 ( .A(n4591), .B(DATAO_REG_13__SCAN_IN), .S(n4067), .Z(U3563)
         );
  MUX2_X1 U4571 ( .A(n4056), .B(DATAO_REG_12__SCAN_IN), .S(n4067), .Z(U3562)
         );
  MUX2_X1 U4572 ( .A(n4057), .B(DATAO_REG_11__SCAN_IN), .S(n4067), .Z(U3561)
         );
  MUX2_X1 U4573 ( .A(n4058), .B(DATAO_REG_10__SCAN_IN), .S(n4067), .Z(U3560)
         );
  MUX2_X1 U4574 ( .A(n4059), .B(DATAO_REG_9__SCAN_IN), .S(n4067), .Z(U3559) );
  MUX2_X1 U4575 ( .A(n4060), .B(DATAO_REG_8__SCAN_IN), .S(n4067), .Z(U3558) );
  MUX2_X1 U4576 ( .A(n4061), .B(DATAO_REG_7__SCAN_IN), .S(n4067), .Z(U3557) );
  MUX2_X1 U4577 ( .A(n4783), .B(DATAO_REG_6__SCAN_IN), .S(n4067), .Z(U3556) );
  MUX2_X1 U4578 ( .A(n4062), .B(DATAO_REG_5__SCAN_IN), .S(n4067), .Z(U3555) );
  MUX2_X1 U4579 ( .A(n4063), .B(DATAO_REG_4__SCAN_IN), .S(n4067), .Z(U3554) );
  MUX2_X1 U4580 ( .A(n4064), .B(DATAO_REG_3__SCAN_IN), .S(n4067), .Z(U3553) );
  MUX2_X1 U4581 ( .A(n4065), .B(DATAO_REG_2__SCAN_IN), .S(n4067), .Z(U3552) );
  MUX2_X1 U4582 ( .A(n4066), .B(DATAO_REG_1__SCAN_IN), .S(n4067), .Z(U3551) );
  MUX2_X1 U4583 ( .A(n4721), .B(DATAO_REG_0__SCAN_IN), .S(n4067), .Z(U3550) );
  NAND2_X1 U4584 ( .A1(n4068), .A2(n4387), .ZN(n4078) );
  OAI211_X1 U4585 ( .C1(n4071), .C2(n4070), .A(n4698), .B(n4069), .ZN(n4077)
         );
  OAI211_X1 U4586 ( .C1(n4074), .C2(n4073), .A(n4663), .B(n4072), .ZN(n4076)
         );
  AOI22_X1 U4587 ( .A1(n4697), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4075) );
  NAND4_X1 U4588 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(U3241)
         );
  OAI211_X1 U4589 ( .C1(n4081), .C2(n2617), .A(n4080), .B(n4698), .ZN(n4090)
         );
  AND2_X1 U4590 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4861) );
  INV_X1 U4591 ( .A(n4082), .ZN(n4083) );
  AOI211_X1 U4592 ( .C1(n2302), .C2(n4084), .A(n4083), .B(n4692), .ZN(n4085)
         );
  NOR2_X1 U4593 ( .A1(n4861), .A2(n4085), .ZN(n4089) );
  OR2_X1 U4594 ( .A1(n4703), .A2(n4086), .ZN(n4088) );
  NAND2_X1 U4595 ( .A1(n4697), .A2(ADDR_REG_15__SCAN_IN), .ZN(n4087) );
  NAND4_X1 U4596 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(U3255)
         );
  AOI21_X1 U4597 ( .B1(n4093), .B2(n4092), .A(n4091), .ZN(n4103) );
  AOI221_X1 U4598 ( .B1(n4096), .B2(n4095), .C1(n4094), .C2(n4095), .A(n4692), 
        .ZN(n4097) );
  OR2_X1 U4599 ( .A1(n4098), .A2(n4097), .ZN(n4099) );
  AOI21_X1 U4600 ( .B1(n4697), .B2(ADDR_REG_17__SCAN_IN), .A(n4099), .ZN(n4102) );
  OR2_X1 U4601 ( .A1(n4703), .A2(n4100), .ZN(n4101) );
  OAI211_X1 U4602 ( .C1(n4103), .C2(n4680), .A(n4102), .B(n4101), .ZN(U3257)
         );
  XNOR2_X1 U4603 ( .A(n4107), .B(n4106), .ZN(n4108) );
  NAND2_X1 U4604 ( .A1(n4698), .A2(n4108), .ZN(n4109) );
  OAI211_X1 U4605 ( .C1(n4111), .C2(n4703), .A(n4110), .B(n4109), .ZN(U3258)
         );
  XNOR2_X1 U4606 ( .A(n4287), .B(n4112), .ZN(n4341) );
  NOR2_X1 U4607 ( .A1(n4114), .A2(n4113), .ZN(n4291) );
  AOI21_X1 U4608 ( .B1(n4115), .B2(n4896), .A(n4291), .ZN(n4338) );
  NOR2_X1 U4609 ( .A1(n4338), .A2(n4972), .ZN(n4116) );
  AOI21_X1 U4610 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4972), .A(n4116), .ZN(n4117) );
  OAI21_X1 U4611 ( .B1(n4341), .B2(n4259), .A(n4117), .ZN(U3260) );
  XNOR2_X1 U4612 ( .A(n4118), .B(n4123), .ZN(n4297) );
  AOI22_X1 U4613 ( .A1(n4972), .A2(REG2_REG_28__SCAN_IN), .B1(n4119), .B2(
        n4917), .ZN(n4133) );
  INV_X1 U4614 ( .A(n4144), .ZN(n4122) );
  INV_X1 U4615 ( .A(n4120), .ZN(n4121) );
  OAI211_X1 U4616 ( .C1(n4122), .C2(n4126), .A(n4121), .B(n4908), .ZN(n4295)
         );
  XNOR2_X1 U4617 ( .A(n4124), .B(n4123), .ZN(n4130) );
  NOR2_X1 U4618 ( .A1(n4125), .A2(n4901), .ZN(n4129) );
  OAI22_X1 U4619 ( .A1(n4127), .A2(n4268), .B1(n4126), .B2(n4780), .ZN(n4128)
         );
  AOI211_X1 U4620 ( .C1(n4130), .C2(n4891), .A(n4129), .B(n4128), .ZN(n4296)
         );
  OAI21_X1 U4621 ( .B1(n4379), .B2(n4295), .A(n4296), .ZN(n4131) );
  NAND2_X1 U4622 ( .A1(n4131), .A2(n4825), .ZN(n4132) );
  OAI211_X1 U4623 ( .C1(n4297), .C2(n4280), .A(n4133), .B(n4132), .ZN(U3262)
         );
  XNOR2_X1 U4624 ( .A(n4134), .B(n4142), .ZN(n4135) );
  NAND2_X1 U4625 ( .A1(n4135), .A2(n4891), .ZN(n4139) );
  AOI22_X1 U4626 ( .A1(n4137), .A2(n4274), .B1(n4136), .B2(n4896), .ZN(n4138)
         );
  OAI211_X1 U4627 ( .C1(n4140), .C2(n4268), .A(n4139), .B(n4138), .ZN(n4298)
         );
  AOI21_X1 U4628 ( .B1(n4141), .B2(n4917), .A(n4298), .ZN(n4150) );
  XNOR2_X1 U4629 ( .A(n4143), .B(n4142), .ZN(n4299) );
  NAND2_X1 U4630 ( .A1(n4299), .A2(n4921), .ZN(n4149) );
  INV_X1 U4631 ( .A(n4162), .ZN(n4146) );
  OAI21_X1 U4632 ( .B1(n4146), .B2(n4145), .A(n4144), .ZN(n4349) );
  INV_X1 U4633 ( .A(n4349), .ZN(n4147) );
  AOI22_X1 U4634 ( .A1(n4147), .A2(n4968), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4972), .ZN(n4148) );
  OAI211_X1 U4635 ( .C1(n4972), .C2(n4150), .A(n4149), .B(n4148), .ZN(U3263)
         );
  XNOR2_X1 U4636 ( .A(n2272), .B(n4153), .ZN(n4303) );
  INV_X1 U4637 ( .A(n4303), .ZN(n4167) );
  INV_X1 U4638 ( .A(n4151), .ZN(n4152) );
  NOR2_X1 U4639 ( .A1(n2295), .A2(n4152), .ZN(n4154) );
  XNOR2_X1 U4640 ( .A(n4154), .B(n4153), .ZN(n4155) );
  NAND2_X1 U4641 ( .A1(n4155), .A2(n4891), .ZN(n4158) );
  AOI22_X1 U4642 ( .A1(n4156), .A2(n4274), .B1(n4896), .B2(n4160), .ZN(n4157)
         );
  OAI211_X1 U4643 ( .C1(n4159), .C2(n4268), .A(n4158), .B(n4157), .ZN(n4302)
         );
  NAND2_X1 U4644 ( .A1(n4178), .A2(n4160), .ZN(n4161) );
  NAND2_X1 U4645 ( .A1(n4162), .A2(n4161), .ZN(n4353) );
  AOI22_X1 U4646 ( .A1(n4972), .A2(REG2_REG_26__SCAN_IN), .B1(n4163), .B2(
        n4917), .ZN(n4164) );
  OAI21_X1 U4647 ( .B1(n4353), .B2(n4259), .A(n4164), .ZN(n4165) );
  AOI21_X1 U4648 ( .B1(n4302), .B2(n4825), .A(n4165), .ZN(n4166) );
  OAI21_X1 U4649 ( .B1(n4167), .B2(n4280), .A(n4166), .ZN(U3264) );
  XNOR2_X1 U4650 ( .A(n4168), .B(n4171), .ZN(n4307) );
  INV_X1 U4651 ( .A(n4307), .ZN(n4184) );
  NOR2_X1 U4652 ( .A1(n4170), .A2(n4169), .ZN(n4172) );
  XNOR2_X1 U4653 ( .A(n4172), .B(n4171), .ZN(n4177) );
  OAI22_X1 U4654 ( .A1(n4173), .A2(n4268), .B1(n4780), .B2(n3191), .ZN(n4174)
         );
  AOI21_X1 U4655 ( .B1(n4274), .B2(n4175), .A(n4174), .ZN(n4176) );
  OAI21_X1 U4656 ( .B1(n4177), .B2(n4785), .A(n4176), .ZN(n4306) );
  OAI21_X1 U4657 ( .B1(n4195), .B2(n3191), .A(n4178), .ZN(n4357) );
  NOR2_X1 U4658 ( .A1(n4357), .A2(n4259), .ZN(n4182) );
  INV_X1 U4659 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4180) );
  OAI22_X1 U4660 ( .A1(n4825), .A2(n4180), .B1(n4179), .B2(n4827), .ZN(n4181)
         );
  AOI211_X1 U4661 ( .C1(n4306), .C2(n4825), .A(n4182), .B(n4181), .ZN(n4183)
         );
  OAI21_X1 U4662 ( .B1(n4184), .B2(n4280), .A(n4183), .ZN(U3265) );
  XOR2_X1 U4663 ( .A(n4186), .B(n4185), .Z(n4311) );
  INV_X1 U4664 ( .A(n4311), .ZN(n4200) );
  XNOR2_X1 U4665 ( .A(n4187), .B(n4186), .ZN(n4192) );
  OAI22_X1 U4666 ( .A1(n4188), .A2(n4268), .B1(n4780), .B2(n4193), .ZN(n4189)
         );
  AOI21_X1 U4667 ( .B1(n4274), .B2(n4190), .A(n4189), .ZN(n4191) );
  OAI21_X1 U4668 ( .B1(n4192), .B2(n4785), .A(n4191), .ZN(n4310) );
  NOR2_X1 U4669 ( .A1(n4219), .A2(n4193), .ZN(n4194) );
  OR2_X1 U4670 ( .A1(n4195), .A2(n4194), .ZN(n4361) );
  AOI22_X1 U4671 ( .A1(n4972), .A2(REG2_REG_24__SCAN_IN), .B1(n4196), .B2(
        n4917), .ZN(n4197) );
  OAI21_X1 U4672 ( .B1(n4361), .B2(n4259), .A(n4197), .ZN(n4198) );
  AOI21_X1 U4673 ( .B1(n4310), .B2(n4825), .A(n4198), .ZN(n4199) );
  OAI21_X1 U4674 ( .B1(n4200), .B2(n4280), .A(n4199), .ZN(U3266) );
  OAI21_X1 U4675 ( .B1(n3921), .B2(n4202), .A(n4201), .ZN(n4229) );
  INV_X1 U4676 ( .A(n4229), .ZN(n4204) );
  NOR2_X1 U4677 ( .A1(n4204), .A2(n4203), .ZN(n4227) );
  NOR2_X1 U4678 ( .A1(n4227), .A2(n4205), .ZN(n4206) );
  XNOR2_X1 U4679 ( .A(n4206), .B(n4212), .ZN(n4315) );
  INV_X1 U4680 ( .A(n4315), .ZN(n4226) );
  INV_X1 U4681 ( .A(n4207), .ZN(n4208) );
  AOI21_X1 U4682 ( .B1(n4210), .B2(n4209), .A(n4208), .ZN(n4231) );
  OAI21_X1 U4683 ( .B1(n4231), .B2(n4230), .A(n4211), .ZN(n4213) );
  XNOR2_X1 U4684 ( .A(n4213), .B(n4212), .ZN(n4218) );
  OAI22_X1 U4685 ( .A1(n4214), .A2(n4268), .B1(n4221), .B2(n4780), .ZN(n4215)
         );
  AOI21_X1 U4686 ( .B1(n4274), .B2(n4216), .A(n4215), .ZN(n4217) );
  OAI21_X1 U4687 ( .B1(n4218), .B2(n4785), .A(n4217), .ZN(n4314) );
  INV_X1 U4688 ( .A(n4219), .ZN(n4220) );
  OAI21_X1 U4689 ( .B1(n2351), .B2(n4221), .A(n4220), .ZN(n4365) );
  AOI22_X1 U4690 ( .A1(n4972), .A2(REG2_REG_23__SCAN_IN), .B1(n4222), .B2(
        n4917), .ZN(n4223) );
  OAI21_X1 U4691 ( .B1(n4365), .B2(n4259), .A(n4223), .ZN(n4224) );
  AOI21_X1 U4692 ( .B1(n4314), .B2(n4825), .A(n4224), .ZN(n4225) );
  OAI21_X1 U4693 ( .B1(n4226), .B2(n4280), .A(n4225), .ZN(U3267) );
  INV_X1 U4694 ( .A(n4227), .ZN(n4228) );
  OAI21_X1 U4695 ( .B1(n4229), .B2(n4230), .A(n4228), .ZN(n4322) );
  XNOR2_X1 U4696 ( .A(n4231), .B(n4230), .ZN(n4237) );
  NAND2_X1 U4697 ( .A1(n4232), .A2(n4274), .ZN(n4234) );
  NAND2_X1 U4698 ( .A1(n4939), .A2(n4897), .ZN(n4233) );
  OAI211_X1 U4699 ( .C1(n4780), .C2(n4235), .A(n4234), .B(n4233), .ZN(n4236)
         );
  AOI21_X1 U4700 ( .B1(n4237), .B2(n4891), .A(n4236), .ZN(n4321) );
  AOI22_X1 U4701 ( .A1(n4972), .A2(REG2_REG_22__SCAN_IN), .B1(n4238), .B2(
        n4917), .ZN(n4241) );
  NAND2_X1 U4702 ( .A1(n2266), .A2(n4239), .ZN(n4318) );
  NAND3_X1 U4703 ( .A1(n4319), .A2(n4968), .A3(n4318), .ZN(n4240) );
  OAI211_X1 U4704 ( .C1(n4321), .C2(n4972), .A(n4241), .B(n4240), .ZN(n4242)
         );
  INV_X1 U4705 ( .A(n4242), .ZN(n4243) );
  OAI21_X1 U4706 ( .B1(n4322), .B2(n4280), .A(n4243), .ZN(U3268) );
  INV_X1 U4707 ( .A(n4244), .ZN(n4328) );
  NAND2_X1 U4708 ( .A1(n4328), .A2(n4327), .ZN(n4252) );
  OAI22_X1 U4709 ( .A1(n4245), .A2(n4901), .B1(n4780), .B2(n4253), .ZN(n4249)
         );
  XNOR2_X1 U4710 ( .A(n4246), .B(n4327), .ZN(n4247) );
  NOR2_X1 U4711 ( .A1(n4247), .A2(n4785), .ZN(n4248) );
  AOI211_X1 U4712 ( .C1(n4897), .C2(n4944), .A(n4249), .B(n4248), .ZN(n4250)
         );
  OAI21_X1 U4713 ( .B1(n4252), .B2(n4251), .A(n4250), .ZN(n4329) );
  INV_X1 U4714 ( .A(n4329), .ZN(n4263) );
  INV_X1 U4715 ( .A(n4252), .ZN(n4331) );
  NOR2_X1 U4716 ( .A1(n4254), .A2(n4253), .ZN(n4255) );
  OR2_X1 U4717 ( .A1(n4256), .A2(n4255), .ZN(n4375) );
  AOI22_X1 U4718 ( .A1(n4972), .A2(REG2_REG_20__SCAN_IN), .B1(n4257), .B2(
        n4917), .ZN(n4258) );
  OAI21_X1 U4719 ( .B1(n4375), .B2(n4259), .A(n4258), .ZN(n4261) );
  NOR3_X1 U4720 ( .A1(n4328), .A2(n4280), .A3(n4327), .ZN(n4260) );
  AOI211_X1 U4721 ( .C1(n4832), .C2(n4331), .A(n4261), .B(n4260), .ZN(n4262)
         );
  OAI21_X1 U4722 ( .B1(n4972), .B2(n4263), .A(n4262), .ZN(U3270) );
  INV_X1 U4723 ( .A(n4264), .ZN(n4266) );
  OAI211_X1 U4724 ( .C1(n4266), .C2(n4267), .A(n4908), .B(n4265), .ZN(n4335)
         );
  OAI22_X1 U4725 ( .A1(n4902), .A2(n4268), .B1(n4780), .B2(n4267), .ZN(n4273)
         );
  XNOR2_X1 U4726 ( .A(n4270), .B(n4269), .ZN(n4271) );
  NOR2_X1 U4727 ( .A1(n4271), .A2(n4785), .ZN(n4272) );
  AOI211_X1 U4728 ( .C1(n4274), .C2(n4944), .A(n4273), .B(n4272), .ZN(n4336)
         );
  OAI21_X1 U4729 ( .B1(n4379), .B2(n4335), .A(n4336), .ZN(n4283) );
  OAI22_X1 U4730 ( .A1(n4825), .A2(n2658), .B1(n4275), .B2(n4827), .ZN(n4282)
         );
  INV_X1 U4731 ( .A(n4276), .ZN(n4277) );
  AOI21_X1 U4732 ( .B1(n4279), .B2(n4278), .A(n4277), .ZN(n4337) );
  NOR2_X1 U4733 ( .A1(n4337), .A2(n4280), .ZN(n4281) );
  AOI211_X1 U4734 ( .C1(n4825), .C2(n4283), .A(n4282), .B(n4281), .ZN(n4284)
         );
  INV_X1 U4735 ( .A(n4284), .ZN(U3272) );
  NOR2_X1 U4736 ( .A1(n4338), .A2(n4909), .ZN(n4285) );
  AOI21_X1 U4737 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4909), .A(n4285), .ZN(n4286) );
  OAI21_X1 U4738 ( .B1(n4341), .B2(n4334), .A(n4286), .ZN(U3549) );
  INV_X1 U4739 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4294) );
  AOI21_X1 U4740 ( .B1(n4289), .B2(n4288), .A(n4287), .ZN(n4969) );
  NAND2_X1 U4741 ( .A1(n4969), .A2(n4743), .ZN(n4293) );
  AND2_X1 U4742 ( .A1(n4289), .A2(n4896), .ZN(n4290) );
  OR2_X1 U4743 ( .A1(n4291), .A2(n4290), .ZN(n4967) );
  NAND2_X1 U4744 ( .A1(n4967), .A2(n4911), .ZN(n4292) );
  OAI211_X1 U4745 ( .C1(n4911), .C2(n4294), .A(n4293), .B(n4292), .ZN(U3548)
         );
  OAI211_X1 U4746 ( .C1(n4297), .C2(n4906), .A(n4296), .B(n4295), .ZN(n4345)
         );
  MUX2_X1 U4747 ( .A(REG1_REG_28__SCAN_IN), .B(n4345), .S(n4911), .Z(U3546) );
  INV_X1 U4748 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4300) );
  AOI21_X1 U4749 ( .B1(n4299), .B2(n4877), .A(n4298), .ZN(n4346) );
  MUX2_X1 U4750 ( .A(n4300), .B(n4346), .S(n4911), .Z(n4301) );
  OAI21_X1 U4751 ( .B1(n4334), .B2(n4349), .A(n4301), .ZN(U3545) );
  INV_X1 U4752 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4304) );
  AOI21_X1 U4753 ( .B1(n4303), .B2(n4877), .A(n4302), .ZN(n4350) );
  MUX2_X1 U4754 ( .A(n4304), .B(n4350), .S(n4911), .Z(n4305) );
  OAI21_X1 U4755 ( .B1(n4334), .B2(n4353), .A(n4305), .ZN(U3544) );
  INV_X1 U4756 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4308) );
  AOI21_X1 U4757 ( .B1(n4307), .B2(n4877), .A(n4306), .ZN(n4354) );
  MUX2_X1 U4758 ( .A(n4308), .B(n4354), .S(n4911), .Z(n4309) );
  OAI21_X1 U4759 ( .B1(n4334), .B2(n4357), .A(n4309), .ZN(U3543) );
  INV_X1 U4760 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4312) );
  AOI21_X1 U4761 ( .B1(n4311), .B2(n4877), .A(n4310), .ZN(n4358) );
  MUX2_X1 U4762 ( .A(n4312), .B(n4358), .S(n4911), .Z(n4313) );
  OAI21_X1 U4763 ( .B1(n4334), .B2(n4361), .A(n4313), .ZN(U3542) );
  INV_X1 U4764 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4316) );
  AOI21_X1 U4765 ( .B1(n4315), .B2(n4877), .A(n4314), .ZN(n4362) );
  MUX2_X1 U4766 ( .A(n4316), .B(n4362), .S(n4911), .Z(n4317) );
  OAI21_X1 U4767 ( .B1(n4334), .B2(n4365), .A(n4317), .ZN(U3541) );
  NAND3_X1 U4768 ( .A1(n4319), .A2(n4908), .A3(n4318), .ZN(n4320) );
  OAI211_X1 U4769 ( .C1(n4322), .C2(n4906), .A(n4321), .B(n4320), .ZN(n4366)
         );
  MUX2_X1 U4770 ( .A(REG1_REG_22__SCAN_IN), .B(n4366), .S(n4911), .Z(U3540) );
  INV_X1 U4771 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4325) );
  AOI21_X1 U4772 ( .B1(n4324), .B2(n4877), .A(n4323), .ZN(n4367) );
  MUX2_X1 U4773 ( .A(n4325), .B(n4367), .S(n4911), .Z(n4326) );
  OAI21_X1 U4774 ( .B1(n4334), .B2(n4370), .A(n4326), .ZN(U3539) );
  INV_X1 U4775 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4332) );
  NOR3_X1 U4776 ( .A1(n4328), .A2(n4906), .A3(n4327), .ZN(n4330) );
  AOI211_X1 U4777 ( .C1(n4331), .C2(n4844), .A(n4330), .B(n4329), .ZN(n4371)
         );
  MUX2_X1 U4778 ( .A(n4332), .B(n4371), .S(n4911), .Z(n4333) );
  OAI21_X1 U4779 ( .B1(n4334), .B2(n4375), .A(n4333), .ZN(U3538) );
  OAI211_X1 U4780 ( .C1(n4337), .C2(n4906), .A(n4336), .B(n4335), .ZN(n4376)
         );
  MUX2_X1 U4781 ( .A(REG1_REG_18__SCAN_IN), .B(n4376), .S(n4911), .Z(U3536) );
  NOR2_X1 U4782 ( .A1(n4338), .A2(n4912), .ZN(n4339) );
  AOI21_X1 U4783 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4912), .A(n4339), .ZN(n4340) );
  OAI21_X1 U4784 ( .B1(n4341), .B2(n4374), .A(n4340), .ZN(U3517) );
  INV_X1 U4785 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4344) );
  NAND2_X1 U4786 ( .A1(n4969), .A2(n4745), .ZN(n4343) );
  NAND2_X1 U4787 ( .A1(n4967), .A2(n4915), .ZN(n4342) );
  OAI211_X1 U4788 ( .C1(n4915), .C2(n4344), .A(n4343), .B(n4342), .ZN(U3516)
         );
  MUX2_X1 U4789 ( .A(REG0_REG_28__SCAN_IN), .B(n4345), .S(n4915), .Z(U3514) );
  INV_X1 U4790 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4347) );
  MUX2_X1 U4791 ( .A(n4347), .B(n4346), .S(n4915), .Z(n4348) );
  OAI21_X1 U4792 ( .B1(n4349), .B2(n4374), .A(n4348), .ZN(U3513) );
  INV_X1 U4793 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4351) );
  MUX2_X1 U4794 ( .A(n4351), .B(n4350), .S(n4915), .Z(n4352) );
  OAI21_X1 U4795 ( .B1(n4353), .B2(n4374), .A(n4352), .ZN(U3512) );
  INV_X1 U4796 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4355) );
  MUX2_X1 U4797 ( .A(n4355), .B(n4354), .S(n4915), .Z(n4356) );
  OAI21_X1 U4798 ( .B1(n4357), .B2(n4374), .A(n4356), .ZN(U3511) );
  INV_X1 U4799 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4359) );
  MUX2_X1 U4800 ( .A(n4359), .B(n4358), .S(n4915), .Z(n4360) );
  OAI21_X1 U4801 ( .B1(n4361), .B2(n4374), .A(n4360), .ZN(U3510) );
  INV_X1 U4802 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4363) );
  MUX2_X1 U4803 ( .A(n4363), .B(n4362), .S(n4915), .Z(n4364) );
  OAI21_X1 U4804 ( .B1(n4365), .B2(n4374), .A(n4364), .ZN(U3509) );
  MUX2_X1 U4805 ( .A(REG0_REG_22__SCAN_IN), .B(n4366), .S(n4915), .Z(U3508) );
  INV_X1 U4806 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4368) );
  MUX2_X1 U4807 ( .A(n4368), .B(n4367), .S(n4915), .Z(n4369) );
  OAI21_X1 U4808 ( .B1(n4370), .B2(n4374), .A(n4369), .ZN(U3507) );
  INV_X1 U4809 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4372) );
  MUX2_X1 U4810 ( .A(n4372), .B(n4371), .S(n4915), .Z(n4373) );
  OAI21_X1 U4811 ( .B1(n4375), .B2(n4374), .A(n4373), .ZN(U3506) );
  MUX2_X1 U4812 ( .A(REG0_REG_18__SCAN_IN), .B(n4376), .S(n4915), .Z(U3503) );
  MUX2_X1 U4813 ( .A(n4377), .B(D_REG_1__SCAN_IN), .S(n4389), .Z(U3459) );
  MUX2_X1 U4814 ( .A(DATAI_27_), .B(n4599), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U4815 ( .A(n4378), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U4816 ( .A(DATAI_19_), .B(n4379), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4817 ( .A(n4380), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U4818 ( .A(n4381), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U4819 ( .A(DATAI_8_), .B(n4382), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4820 ( .A(n4383), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4821 ( .A(DATAI_4_), .B(n4384), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4822 ( .A(n4385), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4823 ( .A(n4386), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4824 ( .A(n4387), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  OAI21_X1 U4825 ( .B1(STATE_REG_SCAN_IN), .B2(n4419), .A(n4388), .ZN(U3329)
         );
  AND2_X1 U4826 ( .A1(D_REG_2__SCAN_IN), .A2(n4389), .ZN(U3320) );
  AND2_X1 U4827 ( .A1(D_REG_3__SCAN_IN), .A2(n4389), .ZN(U3319) );
  AND2_X1 U4828 ( .A1(D_REG_4__SCAN_IN), .A2(n4389), .ZN(U3318) );
  AND2_X1 U4829 ( .A1(D_REG_5__SCAN_IN), .A2(n4389), .ZN(U3317) );
  AND2_X1 U4830 ( .A1(D_REG_6__SCAN_IN), .A2(n4389), .ZN(U3316) );
  AND2_X1 U4831 ( .A1(D_REG_7__SCAN_IN), .A2(n4389), .ZN(U3315) );
  AND2_X1 U4832 ( .A1(D_REG_8__SCAN_IN), .A2(n4389), .ZN(U3314) );
  AND2_X1 U4833 ( .A1(D_REG_9__SCAN_IN), .A2(n4389), .ZN(U3313) );
  AND2_X1 U4834 ( .A1(D_REG_10__SCAN_IN), .A2(n4389), .ZN(U3312) );
  AND2_X1 U4835 ( .A1(D_REG_11__SCAN_IN), .A2(n4389), .ZN(U3311) );
  AND2_X1 U4836 ( .A1(D_REG_12__SCAN_IN), .A2(n4389), .ZN(U3310) );
  AND2_X1 U4837 ( .A1(D_REG_13__SCAN_IN), .A2(n4389), .ZN(U3309) );
  AND2_X1 U4838 ( .A1(D_REG_14__SCAN_IN), .A2(n4389), .ZN(U3308) );
  AND2_X1 U4839 ( .A1(D_REG_15__SCAN_IN), .A2(n4389), .ZN(U3307) );
  AND2_X1 U4840 ( .A1(D_REG_16__SCAN_IN), .A2(n4389), .ZN(U3306) );
  AND2_X1 U4841 ( .A1(D_REG_17__SCAN_IN), .A2(n4389), .ZN(U3305) );
  AND2_X1 U4842 ( .A1(D_REG_18__SCAN_IN), .A2(n4389), .ZN(U3304) );
  AND2_X1 U4843 ( .A1(D_REG_19__SCAN_IN), .A2(n4389), .ZN(U3303) );
  AND2_X1 U4844 ( .A1(D_REG_20__SCAN_IN), .A2(n4389), .ZN(U3302) );
  AND2_X1 U4845 ( .A1(D_REG_21__SCAN_IN), .A2(n4389), .ZN(U3301) );
  AND2_X1 U4846 ( .A1(D_REG_22__SCAN_IN), .A2(n4389), .ZN(U3300) );
  AND2_X1 U4847 ( .A1(D_REG_23__SCAN_IN), .A2(n4389), .ZN(U3299) );
  AND2_X1 U4848 ( .A1(D_REG_24__SCAN_IN), .A2(n4389), .ZN(U3298) );
  AND2_X1 U4849 ( .A1(D_REG_25__SCAN_IN), .A2(n4389), .ZN(U3297) );
  AND2_X1 U4850 ( .A1(D_REG_26__SCAN_IN), .A2(n4389), .ZN(U3296) );
  AND2_X1 U4851 ( .A1(D_REG_27__SCAN_IN), .A2(n4389), .ZN(U3295) );
  AND2_X1 U4852 ( .A1(D_REG_28__SCAN_IN), .A2(n4389), .ZN(U3294) );
  AND2_X1 U4853 ( .A1(D_REG_29__SCAN_IN), .A2(n4389), .ZN(U3293) );
  AND2_X1 U4854 ( .A1(D_REG_30__SCAN_IN), .A2(n4389), .ZN(U3292) );
  AND2_X1 U4855 ( .A1(D_REG_31__SCAN_IN), .A2(n4389), .ZN(U3291) );
  OAI22_X1 U4856 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_114), .B1(
        keyinput_115), .B2(REG3_REG_9__SCAN_IN), .ZN(n4390) );
  AOI221_X1 U4857 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_114), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_115), .A(n4390), .ZN(n4467) );
  INV_X1 U4858 ( .A(keyinput_113), .ZN(n4465) );
  INV_X1 U4859 ( .A(keyinput_112), .ZN(n4463) );
  OAI22_X1 U4860 ( .A1(n4483), .A2(keyinput_109), .B1(keyinput_108), .B2(
        REG3_REG_12__SCAN_IN), .ZN(n4391) );
  AOI221_X1 U4861 ( .B1(n4483), .B2(keyinput_109), .C1(REG3_REG_12__SCAN_IN), 
        .C2(keyinput_108), .A(n4391), .ZN(n4461) );
  OAI22_X1 U4862 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_111), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_110), .ZN(n4392) );
  AOI221_X1 U4863 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_111), .C1(
        keyinput_110), .C2(REG3_REG_16__SCAN_IN), .A(n4392), .ZN(n4460) );
  INV_X1 U4864 ( .A(keyinput_107), .ZN(n4458) );
  INV_X1 U4865 ( .A(keyinput_106), .ZN(n4456) );
  AOI22_X1 U4866 ( .A1(n4394), .A2(keyinput_100), .B1(n4486), .B2(keyinput_101), .ZN(n4393) );
  OAI221_X1 U4867 ( .B1(n4394), .B2(keyinput_100), .C1(n4486), .C2(
        keyinput_101), .A(n4393), .ZN(n4448) );
  INV_X1 U4868 ( .A(keyinput_99), .ZN(n4446) );
  AOI22_X1 U4869 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_97), .B1(U3149), 
        .B2(keyinput_96), .ZN(n4395) );
  OAI221_X1 U4870 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_97), .C1(U3149), 
        .C2(keyinput_96), .A(n4395), .ZN(n4443) );
  OAI22_X1 U4871 ( .A1(DATAI_3_), .A2(keyinput_92), .B1(DATAI_2_), .B2(
        keyinput_93), .ZN(n4396) );
  AOI221_X1 U4872 ( .B1(DATAI_3_), .B2(keyinput_92), .C1(keyinput_93), .C2(
        DATAI_2_), .A(n4396), .ZN(n4441) );
  INV_X1 U4873 ( .A(DATAI_4_), .ZN(n4525) );
  INV_X1 U4874 ( .A(keyinput_91), .ZN(n4437) );
  OAI22_X1 U4875 ( .A1(DATAI_7_), .A2(keyinput_88), .B1(keyinput_89), .B2(
        DATAI_6_), .ZN(n4397) );
  AOI221_X1 U4876 ( .B1(DATAI_7_), .B2(keyinput_88), .C1(DATAI_6_), .C2(
        keyinput_89), .A(n4397), .ZN(n4434) );
  INV_X1 U4877 ( .A(DATAI_15_), .ZN(n4423) );
  INV_X1 U4878 ( .A(DATAI_17_), .ZN(n4399) );
  OAI22_X1 U4879 ( .A1(n4400), .A2(keyinput_77), .B1(n4399), .B2(keyinput_78), 
        .ZN(n4398) );
  AOI221_X1 U4880 ( .B1(n4400), .B2(keyinput_77), .C1(keyinput_78), .C2(n4399), 
        .A(n4398), .ZN(n4406) );
  OAI22_X1 U4881 ( .A1(n2981), .A2(keyinput_75), .B1(keyinput_74), .B2(
        DATAI_21_), .ZN(n4401) );
  AOI221_X1 U4882 ( .B1(n2981), .B2(keyinput_75), .C1(DATAI_21_), .C2(
        keyinput_74), .A(n4401), .ZN(n4405) );
  OAI22_X1 U4883 ( .A1(n4490), .A2(keyinput_73), .B1(keyinput_76), .B2(
        DATAI_19_), .ZN(n4402) );
  AOI221_X1 U4884 ( .B1(n4490), .B2(keyinput_73), .C1(DATAI_19_), .C2(
        keyinput_76), .A(n4402), .ZN(n4404) );
  INV_X1 U4885 ( .A(DATAI_16_), .ZN(n4881) );
  XOR2_X1 U4886 ( .A(n4881), .B(keyinput_79), .Z(n4403) );
  NAND4_X1 U4887 ( .A1(n4406), .A2(n4405), .A3(n4404), .A4(n4403), .ZN(n4421)
         );
  AOI22_X1 U4888 ( .A1(DATAI_24_), .A2(keyinput_71), .B1(n4408), .B2(
        keyinput_70), .ZN(n4407) );
  OAI221_X1 U4889 ( .B1(DATAI_24_), .B2(keyinput_71), .C1(n4408), .C2(
        keyinput_70), .A(n4407), .ZN(n4417) );
  INV_X1 U4890 ( .A(keyinput_69), .ZN(n4415) );
  OAI22_X1 U4891 ( .A1(n3092), .A2(keyinput_67), .B1(keyinput_66), .B2(
        DATAI_29_), .ZN(n4409) );
  AOI221_X1 U4892 ( .B1(n3092), .B2(keyinput_67), .C1(DATAI_29_), .C2(
        keyinput_66), .A(n4409), .ZN(n4412) );
  AOI22_X1 U4893 ( .A1(DATAI_31_), .A2(keyinput_64), .B1(DATAI_30_), .B2(
        keyinput_65), .ZN(n4410) );
  OAI221_X1 U4894 ( .B1(DATAI_31_), .B2(keyinput_64), .C1(DATAI_30_), .C2(
        keyinput_65), .A(n4410), .ZN(n4411) );
  OAI211_X1 U4895 ( .C1(DATAI_27_), .C2(keyinput_68), .A(n4412), .B(n4411), 
        .ZN(n4413) );
  AOI21_X1 U4896 ( .B1(DATAI_27_), .B2(keyinput_68), .A(n4413), .ZN(n4414) );
  AOI221_X1 U4897 ( .B1(DATAI_26_), .B2(keyinput_69), .C1(n3063), .C2(n4415), 
        .A(n4414), .ZN(n4416) );
  OAI22_X1 U4898 ( .A1(keyinput_72), .A2(n4419), .B1(n4417), .B2(n4416), .ZN(
        n4418) );
  AOI21_X1 U4899 ( .B1(keyinput_72), .B2(n4419), .A(n4418), .ZN(n4420) );
  OAI22_X1 U4900 ( .A1(keyinput_80), .A2(n4423), .B1(n4421), .B2(n4420), .ZN(
        n4422) );
  AOI21_X1 U4901 ( .B1(keyinput_80), .B2(n4423), .A(n4422), .ZN(n4432) );
  INV_X1 U4902 ( .A(DATAI_10_), .ZN(n4812) );
  INV_X1 U4903 ( .A(DATAI_12_), .ZN(n4837) );
  AOI22_X1 U4904 ( .A1(n4812), .A2(keyinput_85), .B1(n4837), .B2(keyinput_83), 
        .ZN(n4424) );
  OAI221_X1 U4905 ( .B1(n4812), .B2(keyinput_85), .C1(n4837), .C2(keyinput_83), 
        .A(n4424), .ZN(n4427) );
  INV_X1 U4906 ( .A(DATAI_13_), .ZN(n4838) );
  AOI22_X1 U4907 ( .A1(DATAI_14_), .A2(keyinput_81), .B1(n4838), .B2(
        keyinput_82), .ZN(n4425) );
  OAI221_X1 U4908 ( .B1(DATAI_14_), .B2(keyinput_81), .C1(n4838), .C2(
        keyinput_82), .A(n4425), .ZN(n4426) );
  AOI211_X1 U4909 ( .C1(keyinput_84), .C2(DATAI_11_), .A(n4427), .B(n4426), 
        .ZN(n4428) );
  OAI21_X1 U4910 ( .B1(keyinput_84), .B2(DATAI_11_), .A(n4428), .ZN(n4431) );
  OAI22_X1 U4911 ( .A1(DATAI_9_), .A2(keyinput_86), .B1(DATAI_8_), .B2(
        keyinput_87), .ZN(n4429) );
  AOI221_X1 U4912 ( .B1(DATAI_9_), .B2(keyinput_86), .C1(keyinput_87), .C2(
        DATAI_8_), .A(n4429), .ZN(n4430) );
  OAI21_X1 U4913 ( .B1(n4432), .B2(n4431), .A(n4430), .ZN(n4433) );
  AOI22_X1 U4914 ( .A1(n4434), .A2(n4433), .B1(keyinput_90), .B2(DATAI_5_), 
        .ZN(n4435) );
  OAI21_X1 U4915 ( .B1(keyinput_90), .B2(DATAI_5_), .A(n4435), .ZN(n4436) );
  OAI221_X1 U4916 ( .B1(DATAI_4_), .B2(keyinput_91), .C1(n4525), .C2(n4437), 
        .A(n4436), .ZN(n4440) );
  AOI22_X1 U4917 ( .A1(DATAI_1_), .A2(keyinput_94), .B1(n2399), .B2(
        keyinput_95), .ZN(n4438) );
  OAI221_X1 U4918 ( .B1(DATAI_1_), .B2(keyinput_94), .C1(n2399), .C2(
        keyinput_95), .A(n4438), .ZN(n4439) );
  AOI21_X1 U4919 ( .B1(n4441), .B2(n4440), .A(n4439), .ZN(n4442) );
  OAI22_X1 U4920 ( .A1(n4443), .A2(n4442), .B1(keyinput_98), .B2(
        REG3_REG_27__SCAN_IN), .ZN(n4444) );
  AOI21_X1 U4921 ( .B1(keyinput_98), .B2(REG3_REG_27__SCAN_IN), .A(n4444), 
        .ZN(n4445) );
  AOI221_X1 U4922 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_99), .C1(n4536), 
        .C2(n4446), .A(n4445), .ZN(n4447) );
  OAI22_X1 U4923 ( .A1(n4448), .A2(n4447), .B1(keyinput_102), .B2(
        REG3_REG_3__SCAN_IN), .ZN(n4449) );
  AOI21_X1 U4924 ( .B1(keyinput_102), .B2(REG3_REG_3__SCAN_IN), .A(n4449), 
        .ZN(n4453) );
  AOI22_X1 U4925 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_103), .B1(n4451), 
        .B2(keyinput_105), .ZN(n4450) );
  OAI221_X1 U4926 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_103), .C1(n4451), 
        .C2(keyinput_105), .A(n4450), .ZN(n4452) );
  AOI211_X1 U4927 ( .C1(n3139), .C2(keyinput_104), .A(n4453), .B(n4452), .ZN(
        n4454) );
  OAI21_X1 U4928 ( .B1(n3139), .B2(keyinput_104), .A(n4454), .ZN(n4455) );
  OAI221_X1 U4929 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_106), .C1(n3336), 
        .C2(n4456), .A(n4455), .ZN(n4457) );
  OAI221_X1 U4930 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_107), .C1(n4548), 
        .C2(n4458), .A(n4457), .ZN(n4459) );
  NAND3_X1 U4931 ( .A1(n4461), .A2(n4460), .A3(n4459), .ZN(n4462) );
  OAI221_X1 U4932 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_112), .C1(n4555), 
        .C2(n4463), .A(n4462), .ZN(n4464) );
  OAI221_X1 U4933 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_113), .C1(n4557), 
        .C2(n4465), .A(n4464), .ZN(n4466) );
  AOI22_X1 U4934 ( .A1(n4467), .A2(n4466), .B1(keyinput_116), .B2(
        REG3_REG_0__SCAN_IN), .ZN(n4468) );
  OAI21_X1 U4935 ( .B1(keyinput_116), .B2(REG3_REG_0__SCAN_IN), .A(n4468), 
        .ZN(n4476) );
  OAI22_X1 U4936 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_118), .B1(
        REG3_REG_20__SCAN_IN), .B2(keyinput_117), .ZN(n4469) );
  AOI221_X1 U4937 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_118), .C1(
        keyinput_117), .C2(REG3_REG_20__SCAN_IN), .A(n4469), .ZN(n4475) );
  XNOR2_X1 U4938 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n4472) );
  XNOR2_X1 U4939 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_121), .ZN(n4471) );
  XNOR2_X1 U4940 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_120), .ZN(n4470) );
  NAND4_X1 U4941 ( .A1(n4473), .A2(n4472), .A3(n4471), .A4(n4470), .ZN(n4474)
         );
  AOI21_X1 U4942 ( .B1(n4476), .B2(n4475), .A(n4474), .ZN(n4479) );
  AOI22_X1 U4943 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_123), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput_125), .ZN(n4477) );
  OAI221_X1 U4944 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_123), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_125), .A(n4477), .ZN(n4478) );
  AOI211_X1 U4945 ( .C1(IR_REG_5__SCAN_IN), .C2(keyinput_124), .A(n4479), .B(
        n4478), .ZN(n4480) );
  OAI21_X1 U4946 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_124), .A(n4480), .ZN(
        n4582) );
  OAI22_X1 U4947 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_126), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput_127), .ZN(n4481) );
  AOI221_X1 U4948 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_126), .C1(
        keyinput_127), .C2(IR_REG_8__SCAN_IN), .A(n4481), .ZN(n4581) );
  INV_X1 U4949 ( .A(keyinput_49), .ZN(n4558) );
  INV_X1 U4950 ( .A(keyinput_48), .ZN(n4554) );
  OAI22_X1 U4951 ( .A1(n4483), .A2(keyinput_45), .B1(keyinput_46), .B2(
        REG3_REG_16__SCAN_IN), .ZN(n4482) );
  AOI221_X1 U4952 ( .B1(n4483), .B2(keyinput_45), .C1(REG3_REG_16__SCAN_IN), 
        .C2(keyinput_46), .A(n4482), .ZN(n4552) );
  OAI22_X1 U4953 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_47), .B1(keyinput_44), .B2(REG3_REG_12__SCAN_IN), .ZN(n4484) );
  AOI221_X1 U4954 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_47), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_44), .A(n4484), .ZN(n4551) );
  INV_X1 U4955 ( .A(keyinput_43), .ZN(n4549) );
  INV_X1 U4956 ( .A(keyinput_42), .ZN(n4546) );
  AOI22_X1 U4957 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_36), .B1(n4486), 
        .B2(keyinput_37), .ZN(n4485) );
  OAI221_X1 U4958 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_36), .C1(n4486), 
        .C2(keyinput_37), .A(n4485), .ZN(n4539) );
  INV_X1 U4959 ( .A(keyinput_35), .ZN(n4537) );
  INV_X1 U4960 ( .A(keyinput_27), .ZN(n4524) );
  OAI22_X1 U4961 ( .A1(DATAI_21_), .A2(keyinput_10), .B1(DATAI_17_), .B2(
        keyinput_14), .ZN(n4487) );
  AOI221_X1 U4962 ( .B1(DATAI_21_), .B2(keyinput_10), .C1(keyinput_14), .C2(
        DATAI_17_), .A(n4487), .ZN(n4495) );
  INV_X1 U4963 ( .A(DATAI_19_), .ZN(n4489) );
  OAI22_X1 U4964 ( .A1(n4490), .A2(keyinput_9), .B1(n4489), .B2(keyinput_12), 
        .ZN(n4488) );
  AOI221_X1 U4965 ( .B1(n4490), .B2(keyinput_9), .C1(keyinput_12), .C2(n4489), 
        .A(n4488), .ZN(n4494) );
  XOR2_X1 U4966 ( .A(keyinput_11), .B(DATAI_20_), .Z(n4493) );
  OAI22_X1 U4967 ( .A1(n4881), .A2(keyinput_15), .B1(keyinput_13), .B2(
        DATAI_18_), .ZN(n4491) );
  AOI221_X1 U4968 ( .B1(n4881), .B2(keyinput_15), .C1(DATAI_18_), .C2(
        keyinput_13), .A(n4491), .ZN(n4492) );
  NAND4_X1 U4969 ( .A1(n4495), .A2(n4494), .A3(n4493), .A4(n4492), .ZN(n4508)
         );
  AOI22_X1 U4970 ( .A1(DATAI_25_), .A2(keyinput_6), .B1(n3036), .B2(keyinput_7), .ZN(n4496) );
  OAI221_X1 U4971 ( .B1(DATAI_25_), .B2(keyinput_6), .C1(n3036), .C2(
        keyinput_7), .A(n4496), .ZN(n4505) );
  INV_X1 U4972 ( .A(keyinput_5), .ZN(n4503) );
  OAI22_X1 U4973 ( .A1(n3092), .A2(keyinput_3), .B1(keyinput_2), .B2(DATAI_29_), .ZN(n4497) );
  AOI221_X1 U4974 ( .B1(n3092), .B2(keyinput_3), .C1(DATAI_29_), .C2(
        keyinput_2), .A(n4497), .ZN(n4500) );
  AOI22_X1 U4975 ( .A1(DATAI_31_), .A2(keyinput_0), .B1(DATAI_30_), .B2(
        keyinput_1), .ZN(n4498) );
  OAI221_X1 U4976 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(DATAI_30_), .C2(
        keyinput_1), .A(n4498), .ZN(n4499) );
  OAI211_X1 U4977 ( .C1(DATAI_27_), .C2(keyinput_4), .A(n4500), .B(n4499), 
        .ZN(n4501) );
  AOI21_X1 U4978 ( .B1(DATAI_27_), .B2(keyinput_4), .A(n4501), .ZN(n4502) );
  AOI221_X1 U4979 ( .B1(DATAI_26_), .B2(n4503), .C1(n3063), .C2(keyinput_5), 
        .A(n4502), .ZN(n4504) );
  OAI22_X1 U4980 ( .A1(n4505), .A2(n4504), .B1(keyinput_8), .B2(DATAI_23_), 
        .ZN(n4506) );
  AOI21_X1 U4981 ( .B1(keyinput_8), .B2(DATAI_23_), .A(n4506), .ZN(n4507) );
  OAI22_X1 U4982 ( .A1(n4508), .A2(n4507), .B1(keyinput_16), .B2(DATAI_15_), 
        .ZN(n4509) );
  AOI21_X1 U4983 ( .B1(keyinput_16), .B2(DATAI_15_), .A(n4509), .ZN(n4518) );
  AOI22_X1 U4984 ( .A1(n4812), .A2(keyinput_21), .B1(n4838), .B2(keyinput_18), 
        .ZN(n4510) );
  OAI221_X1 U4985 ( .B1(n4812), .B2(keyinput_21), .C1(n4838), .C2(keyinput_18), 
        .A(n4510), .ZN(n4513) );
  INV_X1 U4986 ( .A(DATAI_11_), .ZN(n4821) );
  AOI22_X1 U4987 ( .A1(DATAI_14_), .A2(keyinput_17), .B1(n4821), .B2(
        keyinput_20), .ZN(n4511) );
  OAI221_X1 U4988 ( .B1(DATAI_14_), .B2(keyinput_17), .C1(n4821), .C2(
        keyinput_20), .A(n4511), .ZN(n4512) );
  AOI211_X1 U4989 ( .C1(keyinput_19), .C2(DATAI_12_), .A(n4513), .B(n4512), 
        .ZN(n4514) );
  OAI21_X1 U4990 ( .B1(keyinput_19), .B2(DATAI_12_), .A(n4514), .ZN(n4517) );
  INV_X1 U4991 ( .A(DATAI_9_), .ZN(n4810) );
  OAI22_X1 U4992 ( .A1(n4810), .A2(keyinput_22), .B1(keyinput_23), .B2(
        DATAI_8_), .ZN(n4515) );
  AOI221_X1 U4993 ( .B1(n4810), .B2(keyinput_22), .C1(DATAI_8_), .C2(
        keyinput_23), .A(n4515), .ZN(n4516) );
  OAI21_X1 U4994 ( .B1(n4518), .B2(n4517), .A(n4516), .ZN(n4522) );
  OAI22_X1 U4995 ( .A1(DATAI_7_), .A2(keyinput_24), .B1(keyinput_25), .B2(
        DATAI_6_), .ZN(n4519) );
  AOI221_X1 U4996 ( .B1(DATAI_7_), .B2(keyinput_24), .C1(DATAI_6_), .C2(
        keyinput_25), .A(n4519), .ZN(n4521) );
  INV_X1 U4997 ( .A(DATAI_5_), .ZN(n4763) );
  NOR2_X1 U4998 ( .A1(n4763), .A2(keyinput_26), .ZN(n4520) );
  AOI221_X1 U4999 ( .B1(n4522), .B2(n4521), .C1(keyinput_26), .C2(n4763), .A(
        n4520), .ZN(n4523) );
  AOI221_X1 U5000 ( .B1(DATAI_4_), .B2(keyinput_27), .C1(n4525), .C2(n4524), 
        .A(n4523), .ZN(n4530) );
  AOI22_X1 U5001 ( .A1(DATAI_2_), .A2(keyinput_29), .B1(DATAI_3_), .B2(
        keyinput_28), .ZN(n4526) );
  OAI221_X1 U5002 ( .B1(DATAI_2_), .B2(keyinput_29), .C1(DATAI_3_), .C2(
        keyinput_28), .A(n4526), .ZN(n4529) );
  XOR2_X1 U5003 ( .A(DATAI_0_), .B(keyinput_31), .Z(n4528) );
  XNOR2_X1 U5004 ( .A(DATAI_1_), .B(keyinput_30), .ZN(n4527) );
  OAI211_X1 U5005 ( .C1(n4530), .C2(n4529), .A(n4528), .B(n4527), .ZN(n4534)
         );
  OAI22_X1 U5006 ( .A1(U3149), .A2(keyinput_32), .B1(keyinput_33), .B2(
        REG3_REG_7__SCAN_IN), .ZN(n4531) );
  AOI221_X1 U5007 ( .B1(U3149), .B2(keyinput_32), .C1(REG3_REG_7__SCAN_IN), 
        .C2(keyinput_33), .A(n4531), .ZN(n4533) );
  NOR2_X1 U5008 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_34), .ZN(n4532) );
  AOI221_X1 U5009 ( .B1(n4534), .B2(n4533), .C1(keyinput_34), .C2(
        REG3_REG_27__SCAN_IN), .A(n4532), .ZN(n4535) );
  AOI221_X1 U5010 ( .B1(REG3_REG_14__SCAN_IN), .B2(n4537), .C1(n4536), .C2(
        keyinput_35), .A(n4535), .ZN(n4538) );
  OAI22_X1 U5011 ( .A1(n4539), .A2(n4538), .B1(keyinput_38), .B2(
        REG3_REG_3__SCAN_IN), .ZN(n4540) );
  AOI21_X1 U5012 ( .B1(keyinput_38), .B2(REG3_REG_3__SCAN_IN), .A(n4540), .ZN(
        n4543) );
  AOI22_X1 U5013 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_39), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput_41), .ZN(n4541) );
  OAI221_X1 U5014 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_39), .C1(
        REG3_REG_8__SCAN_IN), .C2(keyinput_41), .A(n4541), .ZN(n4542) );
  AOI211_X1 U5015 ( .C1(REG3_REG_28__SCAN_IN), .C2(keyinput_40), .A(n4543), 
        .B(n4542), .ZN(n4544) );
  OAI21_X1 U5016 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_40), .A(n4544), 
        .ZN(n4545) );
  OAI221_X1 U5017 ( .B1(REG3_REG_1__SCAN_IN), .B2(n4546), .C1(n3336), .C2(
        keyinput_42), .A(n4545), .ZN(n4547) );
  OAI221_X1 U5018 ( .B1(REG3_REG_21__SCAN_IN), .B2(n4549), .C1(n4548), .C2(
        keyinput_43), .A(n4547), .ZN(n4550) );
  NAND3_X1 U5019 ( .A1(n4552), .A2(n4551), .A3(n4550), .ZN(n4553) );
  OAI221_X1 U5020 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_48), .C1(n4555), 
        .C2(n4554), .A(n4553), .ZN(n4556) );
  OAI221_X1 U5021 ( .B1(REG3_REG_24__SCAN_IN), .B2(n4558), .C1(n4557), .C2(
        keyinput_49), .A(n4556), .ZN(n4563) );
  OAI22_X1 U5022 ( .A1(n2837), .A2(keyinput_51), .B1(REG3_REG_4__SCAN_IN), 
        .B2(keyinput_50), .ZN(n4559) );
  AOI221_X1 U5023 ( .B1(n2837), .B2(keyinput_51), .C1(keyinput_50), .C2(
        REG3_REG_4__SCAN_IN), .A(n4559), .ZN(n4562) );
  INV_X1 U5024 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4561) );
  NOR2_X1 U5025 ( .A1(n4561), .A2(keyinput_52), .ZN(n4560) );
  AOI221_X1 U5026 ( .B1(n4563), .B2(n4562), .C1(keyinput_52), .C2(n4561), .A(
        n4560), .ZN(n4571) );
  AOI22_X1 U5027 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_53), .B1(n4565), 
        .B2(keyinput_54), .ZN(n4564) );
  OAI221_X1 U5028 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_53), .C1(n4565), 
        .C2(keyinput_54), .A(n4564), .ZN(n4570) );
  OAI22_X1 U5029 ( .A1(n4704), .A2(keyinput_55), .B1(keyinput_56), .B2(
        IR_REG_1__SCAN_IN), .ZN(n4566) );
  AOI221_X1 U5030 ( .B1(n4704), .B2(keyinput_55), .C1(IR_REG_1__SCAN_IN), .C2(
        keyinput_56), .A(n4566), .ZN(n4569) );
  OAI22_X1 U5031 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_57), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput_58), .ZN(n4567) );
  AOI221_X1 U5032 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_57), .C1(keyinput_58), 
        .C2(IR_REG_3__SCAN_IN), .A(n4567), .ZN(n4568) );
  OAI211_X1 U5033 ( .C1(n4571), .C2(n4570), .A(n4569), .B(n4568), .ZN(n4576)
         );
  XOR2_X1 U5034 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .Z(n4575) );
  XNOR2_X1 U5035 ( .A(n4572), .B(keyinput_61), .ZN(n4574) );
  XNOR2_X1 U5036 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_59), .ZN(n4573) );
  NAND4_X1 U5037 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(n4579)
         );
  XNOR2_X1 U5038 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .ZN(n4578) );
  XNOR2_X1 U5039 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_62), .ZN(n4577) );
  NAND3_X1 U5040 ( .A1(n4579), .A2(n4578), .A3(n4577), .ZN(n4580) );
  AOI21_X1 U5041 ( .B1(n4582), .B2(n4581), .A(n4580), .ZN(n4597) );
  NAND2_X1 U5042 ( .A1(n2304), .A2(n4583), .ZN(n4584) );
  XNOR2_X1 U5043 ( .A(n4585), .B(n4584), .ZN(n4595) );
  INV_X1 U5044 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4586) );
  NOR2_X1 U5045 ( .A1(STATE_REG_SCAN_IN), .A2(n4586), .ZN(n4660) );
  OAI22_X1 U5046 ( .A1(n4589), .A2(n4588), .B1(n4858), .B2(n4587), .ZN(n4590)
         );
  AOI211_X1 U5047 ( .C1(n4948), .C2(n4591), .A(n4660), .B(n4590), .ZN(n4592)
         );
  OAI21_X1 U5048 ( .B1(n4966), .B2(n4593), .A(n4592), .ZN(n4594) );
  AOI21_X1 U5049 ( .B1(n4595), .B2(n4961), .A(n4594), .ZN(n4596) );
  XNOR2_X1 U5050 ( .A(n4597), .B(n4596), .ZN(U3221) );
  INV_X1 U5051 ( .A(n4600), .ZN(n4598) );
  OAI211_X1 U5052 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4599), .A(n4601), .B(n4598), 
        .ZN(n4604) );
  AOI22_X1 U5053 ( .A1(n4601), .A2(n4600), .B1(n4698), .B2(n4707), .ZN(n4603)
         );
  AOI22_X1 U5054 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4697), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4602) );
  AOI211_X1 U5055 ( .C1(n4607), .C2(n4606), .A(n4605), .B(n4692), .ZN(n4609)
         );
  AOI211_X1 U5056 ( .C1(n4697), .C2(ADDR_REG_5__SCAN_IN), .A(n4609), .B(n4608), 
        .ZN(n4614) );
  OAI211_X1 U5057 ( .C1(n4612), .C2(n4611), .A(n4698), .B(n4610), .ZN(n4613)
         );
  OAI211_X1 U5058 ( .C1(n4703), .C2(n4764), .A(n4614), .B(n4613), .ZN(U3245)
         );
  AOI211_X1 U5059 ( .C1(n4617), .C2(n4616), .A(n4615), .B(n4692), .ZN(n4619)
         );
  AOI211_X1 U5060 ( .C1(n4697), .C2(ADDR_REG_6__SCAN_IN), .A(n4619), .B(n4618), 
        .ZN(n4623) );
  OAI211_X1 U5061 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4621), .A(n4698), .B(n4620), 
        .ZN(n4622) );
  OAI211_X1 U5062 ( .C1(n4703), .C2(n4624), .A(n4623), .B(n4622), .ZN(U3246)
         );
  INV_X1 U5063 ( .A(n4625), .ZN(n4626) );
  NAND2_X1 U5064 ( .A1(n4627), .A2(n4626), .ZN(n4629) );
  OAI21_X1 U5065 ( .B1(n4630), .B2(n4629), .A(n4698), .ZN(n4628) );
  AOI21_X1 U5066 ( .B1(n4630), .B2(n4629), .A(n4628), .ZN(n4632) );
  AOI211_X1 U5067 ( .C1(n4697), .C2(ADDR_REG_9__SCAN_IN), .A(n4632), .B(n4631), 
        .ZN(n4637) );
  OAI211_X1 U5068 ( .C1(n4635), .C2(n4634), .A(n4663), .B(n4633), .ZN(n4636)
         );
  OAI211_X1 U5069 ( .C1(n4703), .C2(n4811), .A(n4637), .B(n4636), .ZN(U3249)
         );
  OAI211_X1 U5070 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4639), .A(n4663), .B(n4638), .ZN(n4642) );
  OAI211_X1 U5071 ( .C1(n4703), .C2(n4813), .A(n4642), .B(n4641), .ZN(n4643)
         );
  AOI211_X1 U5072 ( .C1(n4697), .C2(ADDR_REG_10__SCAN_IN), .A(n4644), .B(n4643), .ZN(n4645) );
  INV_X1 U5073 ( .A(n4645), .ZN(U3250) );
  AOI22_X1 U5074 ( .A1(n4646), .A2(REG1_REG_11__SCAN_IN), .B1(n2408), .B2(
        n4822), .ZN(n4649) );
  OAI21_X1 U5075 ( .B1(n4649), .B2(n4648), .A(n4698), .ZN(n4647) );
  AOI21_X1 U5076 ( .B1(n4649), .B2(n4648), .A(n4647), .ZN(n4651) );
  AOI211_X1 U5077 ( .C1(n4697), .C2(ADDR_REG_11__SCAN_IN), .A(n4651), .B(n4650), .ZN(n4656) );
  OAI211_X1 U5078 ( .C1(n4654), .C2(n4653), .A(n4663), .B(n4652), .ZN(n4655)
         );
  OAI211_X1 U5079 ( .C1(n4703), .C2(n4822), .A(n4656), .B(n4655), .ZN(U3251)
         );
  AOI211_X1 U5080 ( .C1(n4659), .C2(n4658), .A(n4657), .B(n4680), .ZN(n4661)
         );
  AOI211_X1 U5081 ( .C1(n4697), .C2(ADDR_REG_12__SCAN_IN), .A(n4661), .B(n4660), .ZN(n4666) );
  OAI211_X1 U5082 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4664), .A(n4663), .B(n4662), .ZN(n4665) );
  OAI211_X1 U5083 ( .C1(n4703), .C2(n2609), .A(n4666), .B(n4665), .ZN(U3252)
         );
  OAI21_X1 U5084 ( .B1(n4668), .B2(REG1_REG_13__SCAN_IN), .A(n4667), .ZN(n4670) );
  XNOR2_X1 U5085 ( .A(n4670), .B(n4669), .ZN(n4679) );
  AOI21_X1 U5086 ( .B1(n4839), .B2(n4672), .A(n4671), .ZN(n4674) );
  XNOR2_X1 U5087 ( .A(n4674), .B(n4673), .ZN(n4675) );
  OAI22_X1 U5088 ( .A1(n4839), .A2(n4703), .B1(n4692), .B2(n4675), .ZN(n4676)
         );
  AOI211_X1 U5089 ( .C1(n4697), .C2(ADDR_REG_13__SCAN_IN), .A(n4677), .B(n4676), .ZN(n4678) );
  OAI21_X1 U5090 ( .B1(n4680), .B2(n4679), .A(n4678), .ZN(U3253) );
  AOI211_X1 U5091 ( .C1(n4683), .C2(n4682), .A(n4681), .B(n4692), .ZN(n4685)
         );
  AOI211_X1 U5092 ( .C1(n4697), .C2(ADDR_REG_14__SCAN_IN), .A(n4685), .B(n4684), .ZN(n4689) );
  OAI211_X1 U5093 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4687), .A(n4698), .B(n4686), .ZN(n4688) );
  OAI211_X1 U5094 ( .C1(n4703), .C2(n4690), .A(n4689), .B(n4688), .ZN(U3254)
         );
  NOR2_X1 U5095 ( .A1(STATE_REG_SCAN_IN), .A2(n4691), .ZN(n4884) );
  AOI221_X1 U5096 ( .B1(n4695), .B2(n4694), .C1(n4693), .C2(n4694), .A(n4692), 
        .ZN(n4696) );
  AOI211_X1 U5097 ( .C1(n4697), .C2(ADDR_REG_16__SCAN_IN), .A(n4884), .B(n4696), .ZN(n4702) );
  OAI221_X1 U5098 ( .B1(n4700), .B2(REG1_REG_16__SCAN_IN), .C1(n4700), .C2(
        n4699), .A(n4698), .ZN(n4701) );
  OAI211_X1 U5099 ( .C1(n4703), .C2(n2315), .A(n4702), .B(n4701), .ZN(U3256)
         );
  AOI22_X1 U5100 ( .A1(STATE_REG_SCAN_IN), .A2(n4704), .B1(n2399), .B2(U3149), 
        .ZN(U3352) );
  AND2_X1 U5101 ( .A1(n4732), .A2(n4705), .ZN(n4713) );
  OAI21_X1 U5102 ( .B1(n4824), .B2(n4891), .A(n4714), .ZN(n4706) );
  OAI21_X1 U5103 ( .B1(n3156), .B2(n4901), .A(n4706), .ZN(n4711) );
  AOI211_X1 U5104 ( .C1(n4844), .C2(n4714), .A(n4713), .B(n4711), .ZN(n4709)
         );
  AOI22_X1 U5105 ( .A1(n4911), .A2(n4709), .B1(n4707), .B2(n4909), .ZN(U3518)
         );
  INV_X1 U5106 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4708) );
  AOI22_X1 U5107 ( .A1(n4915), .A2(n4709), .B1(n4708), .B2(n4912), .ZN(U3467)
         );
  INV_X1 U5108 ( .A(n4710), .ZN(n4712) );
  AOI21_X1 U5109 ( .B1(n4713), .B2(n4712), .A(n4711), .ZN(n4717) );
  AOI22_X1 U5110 ( .A1(n4714), .A2(n4832), .B1(REG3_REG_0__SCAN_IN), .B2(n4917), .ZN(n4715) );
  OAI221_X1 U5111 ( .B1(n4972), .B2(n4717), .C1(n4825), .C2(n4716), .A(n4715), 
        .ZN(U3290) );
  OAI21_X1 U5112 ( .B1(n4725), .B2(n4719), .A(n4718), .ZN(n4720) );
  INV_X1 U5113 ( .A(n4720), .ZN(n4737) );
  AOI22_X1 U5114 ( .A1(n4721), .A2(n4897), .B1(n4731), .B2(n4896), .ZN(n4722)
         );
  OAI21_X1 U5115 ( .B1(n4723), .B2(n4901), .A(n4722), .ZN(n4729) );
  NAND2_X1 U5116 ( .A1(n4725), .A2(n4724), .ZN(n4726) );
  AOI21_X1 U5117 ( .B1(n4727), .B2(n4726), .A(n4785), .ZN(n4728) );
  AOI211_X1 U5118 ( .C1(n4737), .C2(n4824), .A(n4729), .B(n4728), .ZN(n4740)
         );
  AOI21_X1 U5119 ( .B1(n4732), .B2(n4731), .A(n4730), .ZN(n4736) );
  AOI22_X1 U5120 ( .A1(n4737), .A2(n4844), .B1(n4908), .B2(n4736), .ZN(n4733)
         );
  AND2_X1 U5121 ( .A1(n4740), .A2(n4733), .ZN(n4735) );
  AOI22_X1 U5122 ( .A1(n4911), .A2(n4735), .B1(n2577), .B2(n4909), .ZN(U3519)
         );
  INV_X1 U5123 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5124 ( .A1(n4915), .A2(n4735), .B1(n4734), .B2(n4912), .ZN(U3469)
         );
  AOI22_X1 U5125 ( .A1(REG2_REG_1__SCAN_IN), .A2(n4972), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4917), .ZN(n4739) );
  AOI22_X1 U5126 ( .A1(n4737), .A2(n4832), .B1(n4968), .B2(n4736), .ZN(n4738)
         );
  OAI211_X1 U5127 ( .C1(n4972), .C2(n4740), .A(n4739), .B(n4738), .ZN(U3289)
         );
  AOI21_X1 U5128 ( .B1(n4844), .B2(n4742), .A(n4741), .ZN(n4748) );
  AOI22_X1 U5129 ( .A1(n4746), .A2(n4743), .B1(REG1_REG_2__SCAN_IN), .B2(n4909), .ZN(n4744) );
  OAI21_X1 U5130 ( .B1(n4748), .B2(n4909), .A(n4744), .ZN(U3520) );
  AOI22_X1 U5131 ( .A1(n4746), .A2(n4745), .B1(REG0_REG_2__SCAN_IN), .B2(n4912), .ZN(n4747) );
  OAI21_X1 U5132 ( .B1(n4748), .B2(n4912), .A(n4747), .ZN(U3471) );
  AOI22_X1 U5133 ( .A1(n4972), .A2(REG2_REG_3__SCAN_IN), .B1(n4917), .B2(n2757), .ZN(n4753) );
  INV_X1 U5134 ( .A(n4749), .ZN(n4750) );
  AOI22_X1 U5135 ( .A1(n4751), .A2(n4832), .B1(n4968), .B2(n4750), .ZN(n4752)
         );
  OAI211_X1 U5136 ( .C1(n4972), .C2(n4754), .A(n4753), .B(n4752), .ZN(U3287)
         );
  AND2_X1 U5137 ( .A1(n4755), .A2(n4844), .ZN(n4758) );
  INV_X1 U5138 ( .A(n4756), .ZN(n4757) );
  NOR3_X1 U5139 ( .A1(n4759), .A2(n4758), .A3(n4757), .ZN(n4762) );
  INV_X1 U5140 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4760) );
  AOI22_X1 U5141 ( .A1(n4911), .A2(n4762), .B1(n4760), .B2(n4909), .ZN(U3522)
         );
  INV_X1 U5142 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4761) );
  AOI22_X1 U5143 ( .A1(n4915), .A2(n4762), .B1(n4761), .B2(n4912), .ZN(U3475)
         );
  AOI22_X1 U5144 ( .A1(STATE_REG_SCAN_IN), .A2(n4764), .B1(n4763), .B2(U3149), 
        .ZN(U3347) );
  OAI22_X1 U5145 ( .A1(U3149), .A2(n4765), .B1(DATAI_6_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4766) );
  INV_X1 U5146 ( .A(n4766), .ZN(U3346) );
  AOI22_X1 U5147 ( .A1(n4767), .A2(n4917), .B1(REG2_REG_6__SCAN_IN), .B2(n4972), .ZN(n4772) );
  INV_X1 U5148 ( .A(n4768), .ZN(n4769) );
  AOI22_X1 U5149 ( .A1(n4770), .A2(n4832), .B1(n4968), .B2(n4769), .ZN(n4771)
         );
  OAI211_X1 U5150 ( .C1(n4972), .C2(n4773), .A(n4772), .B(n4771), .ZN(U3284)
         );
  AOI21_X1 U5151 ( .B1(n4775), .B2(n4774), .A(n4874), .ZN(n4777) );
  AND2_X1 U5152 ( .A1(n4777), .A2(n4776), .ZN(n4798) );
  XOR2_X1 U5153 ( .A(n4789), .B(n4778), .Z(n4786) );
  OAI22_X1 U5154 ( .A1(n4781), .A2(n4901), .B1(n4780), .B2(n4779), .ZN(n4782)
         );
  AOI21_X1 U5155 ( .B1(n4897), .B2(n4783), .A(n4782), .ZN(n4784) );
  OAI21_X1 U5156 ( .B1(n4786), .B2(n4785), .A(n4784), .ZN(n4797) );
  AOI211_X1 U5157 ( .C1(n4798), .C2(n4787), .A(n4972), .B(n4797), .ZN(n4793)
         );
  XOR2_X1 U5158 ( .A(n4790), .B(n4789), .Z(n4799) );
  NAND2_X1 U5159 ( .A1(n4799), .A2(n4791), .ZN(n4792) );
  NAND2_X1 U5160 ( .A1(n4793), .A2(n4792), .ZN(n4794) );
  OAI21_X1 U5161 ( .B1(REG2_REG_7__SCAN_IN), .B2(n4825), .A(n4794), .ZN(n4795)
         );
  OAI21_X1 U5162 ( .B1(n4796), .B2(n4827), .A(n4795), .ZN(U3283) );
  AOI211_X1 U5163 ( .C1(n4799), .C2(n4877), .A(n4798), .B(n4797), .ZN(n4802)
         );
  INV_X1 U5164 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4800) );
  AOI22_X1 U5165 ( .A1(n4911), .A2(n4802), .B1(n4800), .B2(n4909), .ZN(U3525)
         );
  INV_X1 U5166 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4801) );
  AOI22_X1 U5167 ( .A1(n4915), .A2(n4802), .B1(n4801), .B2(n4912), .ZN(U3481)
         );
  AOI22_X1 U5168 ( .A1(n4803), .A2(n4917), .B1(REG2_REG_8__SCAN_IN), .B2(n4972), .ZN(n4808) );
  INV_X1 U5169 ( .A(n4804), .ZN(n4805) );
  AOI22_X1 U5170 ( .A1(n4806), .A2(n4832), .B1(n4968), .B2(n4805), .ZN(n4807)
         );
  OAI211_X1 U5171 ( .C1(n4972), .C2(n4809), .A(n4808), .B(n4807), .ZN(U3282)
         );
  AOI22_X1 U5172 ( .A1(STATE_REG_SCAN_IN), .A2(n4811), .B1(n4810), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5173 ( .A1(STATE_REG_SCAN_IN), .A2(n4813), .B1(n4812), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5174 ( .A1(n4814), .A2(n4917), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4972), .ZN(n4819) );
  INV_X1 U5175 ( .A(n4815), .ZN(n4816) );
  AOI22_X1 U5176 ( .A1(n4817), .A2(n4832), .B1(n4968), .B2(n4816), .ZN(n4818)
         );
  OAI211_X1 U5177 ( .C1(n4972), .C2(n4820), .A(n4819), .B(n4818), .ZN(U3280)
         );
  AOI22_X1 U5178 ( .A1(STATE_REG_SCAN_IN), .A2(n4822), .B1(n4821), .B2(U3149), 
        .ZN(U3341) );
  AOI21_X1 U5179 ( .B1(n4824), .B2(n4833), .A(n4823), .ZN(n4836) );
  OAI22_X1 U5180 ( .A1(n4828), .A2(n4827), .B1(n4826), .B2(n4825), .ZN(n4829)
         );
  INV_X1 U5181 ( .A(n4829), .ZN(n4835) );
  INV_X1 U5182 ( .A(n4830), .ZN(n4831) );
  AOI22_X1 U5183 ( .A1(n4833), .A2(n4832), .B1(n4968), .B2(n4831), .ZN(n4834)
         );
  OAI211_X1 U5184 ( .C1(n4972), .C2(n4836), .A(n4835), .B(n4834), .ZN(U3279)
         );
  AOI22_X1 U5185 ( .A1(STATE_REG_SCAN_IN), .A2(n2609), .B1(n4837), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5186 ( .A1(STATE_REG_SCAN_IN), .A2(n4839), .B1(n4838), .B2(U3149), 
        .ZN(U3339) );
  NOR2_X1 U5187 ( .A1(n4840), .A2(n4874), .ZN(n4842) );
  AOI211_X1 U5188 ( .C1(n4844), .C2(n4843), .A(n4842), .B(n4841), .ZN(n4847)
         );
  AOI22_X1 U5189 ( .A1(n4911), .A2(n4847), .B1(n4845), .B2(n4909), .ZN(U3531)
         );
  INV_X1 U5190 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4846) );
  AOI22_X1 U5191 ( .A1(n4915), .A2(n4847), .B1(n4846), .B2(n4912), .ZN(U3493)
         );
  OAI22_X1 U5192 ( .A1(U3149), .A2(n4848), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4849) );
  INV_X1 U5193 ( .A(n4849), .ZN(U3338) );
  AOI22_X1 U5194 ( .A1(n4850), .A2(n4917), .B1(REG2_REG_14__SCAN_IN), .B2(
        n4972), .ZN(n4855) );
  INV_X1 U5195 ( .A(n4851), .ZN(n4852) );
  AOI22_X1 U5196 ( .A1(n4853), .A2(n4921), .B1(n4968), .B2(n4852), .ZN(n4854)
         );
  OAI211_X1 U5197 ( .C1(n4972), .C2(n4856), .A(n4855), .B(n4854), .ZN(U3276)
         );
  OAI22_X1 U5198 ( .A1(n4859), .A2(n4931), .B1(n4858), .B2(n4857), .ZN(n4860)
         );
  AOI211_X1 U5199 ( .C1(n4957), .C2(n4862), .A(n4861), .B(n4860), .ZN(n4870)
         );
  INV_X1 U5200 ( .A(n4863), .ZN(n4864) );
  NOR2_X1 U5201 ( .A1(n4865), .A2(n4864), .ZN(n4867) );
  XNOR2_X1 U5202 ( .A(n4867), .B(n4866), .ZN(n4868) );
  NAND2_X1 U5203 ( .A1(n4868), .A2(n4961), .ZN(n4869) );
  OAI211_X1 U5204 ( .C1(n4966), .C2(n4871), .A(n4870), .B(n4869), .ZN(U3238)
         );
  OAI21_X1 U5205 ( .B1(n4874), .B2(n4873), .A(n4872), .ZN(n4875) );
  AOI21_X1 U5206 ( .B1(n4877), .B2(n4876), .A(n4875), .ZN(n4880) );
  AOI22_X1 U5207 ( .A1(n4911), .A2(n4880), .B1(n4878), .B2(n4909), .ZN(U3533)
         );
  INV_X1 U5208 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4879) );
  AOI22_X1 U5209 ( .A1(n4915), .A2(n4880), .B1(n4879), .B2(n4912), .ZN(U3497)
         );
  AOI22_X1 U5210 ( .A1(STATE_REG_SCAN_IN), .A2(n2315), .B1(n4881), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5211 ( .A(n4918), .ZN(n4888) );
  AOI22_X1 U5212 ( .A1(n4898), .A2(n4957), .B1(n4960), .B2(n4895), .ZN(n4887)
         );
  XNOR2_X1 U5213 ( .A(n2301), .B(n4882), .ZN(n4885) );
  NOR2_X1 U5214 ( .A1(n4902), .A2(n4931), .ZN(n4883) );
  AOI211_X1 U5215 ( .C1(n4885), .C2(n4961), .A(n4884), .B(n4883), .ZN(n4886)
         );
  OAI211_X1 U5216 ( .C1(n4966), .C2(n4888), .A(n4887), .B(n4886), .ZN(U3223)
         );
  AOI21_X1 U5217 ( .B1(n4895), .B2(n4890), .A(n4889), .ZN(n4920) );
  OAI211_X1 U5218 ( .C1(n4894), .C2(n4893), .A(n4892), .B(n4891), .ZN(n4900)
         );
  AOI22_X1 U5219 ( .A1(n4898), .A2(n4897), .B1(n4896), .B2(n4895), .ZN(n4899)
         );
  OAI211_X1 U5220 ( .C1(n4902), .C2(n4901), .A(n4900), .B(n4899), .ZN(n4916)
         );
  OAI21_X1 U5221 ( .B1(n2491), .B2(n4905), .A(n4904), .ZN(n4919) );
  NOR2_X1 U5222 ( .A1(n4919), .A2(n4906), .ZN(n4907) );
  AOI211_X1 U5223 ( .C1(n4908), .C2(n4920), .A(n4916), .B(n4907), .ZN(n4914)
         );
  INV_X1 U5224 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4910) );
  AOI22_X1 U5225 ( .A1(n4911), .A2(n4914), .B1(n4910), .B2(n4909), .ZN(U3534)
         );
  INV_X1 U5226 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4913) );
  AOI22_X1 U5227 ( .A1(n4915), .A2(n4914), .B1(n4913), .B2(n4912), .ZN(U3499)
         );
  INV_X1 U5228 ( .A(n4916), .ZN(n4925) );
  AOI22_X1 U5229 ( .A1(n4918), .A2(n4917), .B1(REG2_REG_16__SCAN_IN), .B2(
        n4972), .ZN(n4924) );
  INV_X1 U5230 ( .A(n4919), .ZN(n4922) );
  AOI22_X1 U5231 ( .A1(n4922), .A2(n4921), .B1(n4968), .B2(n4920), .ZN(n4923)
         );
  OAI211_X1 U5232 ( .C1(n4972), .C2(n4925), .A(n4924), .B(n4923), .ZN(U3274)
         );
  AOI22_X1 U5233 ( .A1(n4927), .A2(n4957), .B1(n4960), .B2(n4926), .ZN(n4937)
         );
  OAI21_X1 U5234 ( .B1(n4930), .B2(n4929), .A(n4928), .ZN(n4935) );
  NOR2_X1 U5235 ( .A1(n4932), .A2(n4931), .ZN(n4934) );
  AOI211_X1 U5236 ( .C1(n4935), .C2(n4961), .A(n4934), .B(n4933), .ZN(n4936)
         );
  OAI211_X1 U5237 ( .C1(n4966), .C2(n4938), .A(n4937), .B(n4936), .ZN(U3216)
         );
  AOI22_X1 U5238 ( .A1(n4939), .A2(n4948), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n4946) );
  INV_X1 U5239 ( .A(n4952), .ZN(n4940) );
  NOR2_X1 U5240 ( .A1(n4940), .A2(n4953), .ZN(n4941) );
  XNOR2_X1 U5241 ( .A(n4954), .B(n4941), .ZN(n4943) );
  AOI222_X1 U5242 ( .A1(n4944), .A2(n4957), .B1(n4961), .B2(n4943), .C1(n4960), 
        .C2(n4942), .ZN(n4945) );
  OAI211_X1 U5243 ( .C1(n4966), .C2(n4947), .A(n4946), .B(n4945), .ZN(U3230)
         );
  AOI22_X1 U5244 ( .A1(n4949), .A2(n4948), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n4964) );
  NOR2_X1 U5245 ( .A1(n4951), .A2(n4950), .ZN(n4956) );
  OAI21_X1 U5246 ( .B1(n4954), .B2(n4953), .A(n4952), .ZN(n4955) );
  XOR2_X1 U5247 ( .A(n4956), .B(n4955), .Z(n4962) );
  AOI222_X1 U5248 ( .A1(n4962), .A2(n4961), .B1(n4960), .B2(n4959), .C1(n4958), 
        .C2(n4957), .ZN(n4963) );
  OAI211_X1 U5249 ( .C1(n4966), .C2(n4965), .A(n4964), .B(n4963), .ZN(U3220)
         );
  INV_X1 U5250 ( .A(n4967), .ZN(n4971) );
  AOI22_X1 U5251 ( .A1(n4969), .A2(n4968), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4972), .ZN(n4970) );
  OAI21_X1 U5252 ( .B1(n4972), .B2(n4971), .A(n4970), .ZN(U3261) );
  CLKBUF_X1 U2297 ( .A(n3078), .Z(n2261) );
  CLKBUF_X3 U2299 ( .A(n2756), .Z(n3081) );
endmodule

